
module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_63 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15;
    VMW_AOI21 U3 ( .A(A[5]), .B(n15), .C(A[6]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[2]), .B(A[3]), .C(A[4]), .Z(n15) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_62 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n16, n17;
    VMW_NOR2 U3 ( .A(A[6]), .B(n16), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n17) );
    VMW_AND3 U4 ( .A(A[5]), .B(n17), .C(A[4]), .Z(n16) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_61 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n18;
    VMW_NOR3 U3 ( .A(n18), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[4]), .C(A[2]), .Z(n18) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_60 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n19;
    VMW_AOI21 U3 ( .A(A[5]), .B(n19), .C(A[6]), .Z(LT_LE) );
    VMW_OR4 U4 ( .A(A[2]), .B(A[1]), .C(A[4]), .D(A[3]), .Z(n19) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_59 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI211 U3 ( .A(A[3]), .B(A[4]), .C(A[6]), .D(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_58 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI21 U3 ( .A(A[4]), .B(A[5]), .C(A[6]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_57 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n20, n21;
    VMW_AOI211 U3 ( .A(A[3]), .B(n20), .C(n21), .D(A[4]), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n20) );
    VMW_OR2 U4 ( .A(A[6]), .B(A[5]), .Z(n21) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_56 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n23, n24, n22;
    VMW_NOR2 U3 ( .A(A[6]), .B(n22), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[1]), .B(A[0]), .Z(n24) );
    VMW_AO21 U6 ( .A(A[2]), .B(n24), .C(A[3]), .Z(n23) );
    VMW_AND3 U4 ( .A(A[5]), .B(n23), .C(A[4]), .Z(n22) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_55 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n25, n26;
    VMW_NOR4 U3 ( .A(n25), .B(A[4]), .C(A[6]), .D(A[5]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n26), .Z(n25) );
    VMW_AOI211 U4 ( .A(A[0]), .B(A[1]), .C(A[3]), .D(A[2]), .Z(n26) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_54 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR4 U3 ( .A(A[6]), .B(A[5]), .C(A[4]), .D(A[3]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_53 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n27, n28;
    VMW_NOR2 U3 ( .A(A[6]), .B(n27), .Z(LT_LE) );
    VMW_OR4 U5 ( .A(A[1]), .B(A[0]), .C(A[3]), .D(A[2]), .Z(n28) );
    VMW_AND3 U4 ( .A(A[5]), .B(n28), .C(A[4]), .Z(n27) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_52 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n29, n30;
    VMW_NOR4 U3 ( .A(A[6]), .B(A[5]), .C(A[4]), .D(n29), .Z(LT_LE) );
    VMW_INV U5 ( .A(n30), .Z(n29) );
    VMW_OAI21 U4 ( .A(A[2]), .B(A[1]), .C(A[3]), .Z(n30) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_50 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n31, n32;
    VMW_NOR3 U3 ( .A(n31), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[1]), .B(A[0]), .Z(n32) );
    VMW_AND4 U4 ( .A(A[3]), .B(A[4]), .C(A[2]), .D(n32), .Z(n31) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_49 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n33, n34;
    VMW_NOR4 U3 ( .A(A[6]), .B(A[5]), .C(A[4]), .D(n33), .Z(LT_LE) );
    VMW_INV U5 ( .A(n34), .Z(n33) );
    VMW_OAI211 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(A[3]), .Z(n34) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_48 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR5 U3 ( .A(A[3]), .B(A[2]), .C(A[4]), .D(A[6]), .E(A[5]), .Z(LT_LE)
         );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_47 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n35, n36;
    VMW_NOR3 U3 ( .A(n35), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n36), .Z(n35) );
    VMW_OAI211 U4 ( .A(A[2]), .B(A[1]), .C(A[4]), .D(A[3]), .Z(n36) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_46 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n37;
    VMW_AOI21 U3 ( .A(A[5]), .B(n37), .C(A[6]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[4]), .B(A[3]), .C(A[2]), .Z(n37) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_45 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n40, n38, n39;
    VMW_NOR2 U3 ( .A(A[6]), .B(n38), .Z(LT_LE) );
    VMW_AND3 U5 ( .A(A[5]), .B(n40), .C(A[4]), .Z(n38) );
    VMW_INV U6 ( .A(n39), .Z(n40) );
    VMW_AOI211 U4 ( .A(A[0]), .B(A[1]), .C(A[3]), .D(A[2]), .Z(n39) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_44 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n41;
    VMW_NOR2 U3 ( .A(A[6]), .B(n41), .Z(LT_LE) );
    VMW_AND5 U4 ( .A(A[5]), .B(A[2]), .C(A[4]), .D(A[1]), .E(A[3]), .Z(n41) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_43 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n42, n43, n44;
    VMW_NOR2 U3 ( .A(n42), .B(A[6]), .Z(LT_LE) );
    VMW_OAI211 U5 ( .A(A[3]), .B(n43), .C(A[5]), .D(A[4]), .Z(n44) );
    VMW_INV U6 ( .A(n44), .Z(n42) );
    VMW_AND3 U4 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n43) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_42 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n46, n45;
    VMW_AOI21 U3 ( .A(A[5]), .B(n45), .C(A[6]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[4]), .B(n46), .Z(n45) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n46) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_41 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n47, n48;
    VMW_NOR2 U3 ( .A(A[6]), .B(n47), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n48) );
    VMW_AND4 U4 ( .A(A[5]), .B(A[3]), .C(A[4]), .D(n48), .Z(n47) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_40 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR2 U3 ( .A(A[6]), .B(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_39 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n49;
    VMW_AOI211 U3 ( .A(A[4]), .B(n49), .C(A[5]), .D(A[6]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[1]), .B(A[2]), .C(A[3]), .Z(n49) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_38 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n50;
    VMW_AOI211 U3 ( .A(A[1]), .B(A[2]), .C(n50), .D(A[3]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[6]), .B(A[5]), .C(A[4]), .Z(n50) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_37 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n51, n52;
    VMW_AOI211 U3 ( .A(A[3]), .B(n51), .C(n52), .D(A[4]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n51) );
    VMW_OR2 U4 ( .A(A[6]), .B(A[5]), .Z(n52) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_36 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n53;
    VMW_AOI211 U3 ( .A(A[4]), .B(n53), .C(A[6]), .D(A[5]), .Z(LT_LE) );
    VMW_OR4 U4 ( .A(A[1]), .B(A[0]), .C(A[3]), .D(A[2]), .Z(n53) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_35 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n54;
    VMW_NOR4 U3 ( .A(n54), .B(A[0]), .C(A[2]), .D(A[1]), .Z(LT_LE) );
    VMW_OR4 U4 ( .A(A[4]), .B(A[3]), .C(A[6]), .D(A[5]), .Z(n54) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_34 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55;
    VMW_NOR4 U3 ( .A(A[6]), .B(A[5]), .C(A[4]), .D(n55), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[1]), .B(A[3]), .C(A[0]), .D(A[2]), .Z(n55) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_33 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n56, n58, n57;
    VMW_AOI21 U3 ( .A(A[5]), .B(n56), .C(A[6]), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[4]), .B(n58), .C(A[3]), .Z(n56) );
    VMW_INV U6 ( .A(n57), .Z(n58) );
    VMW_OAI21 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .Z(n57) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_32 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n60, n59;
    VMW_AOI21 U3 ( .A(A[5]), .B(n59), .C(A[6]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[3]), .B(n60), .C(A[4]), .Z(n59) );
    VMW_OR2 U4 ( .A(A[2]), .B(A[1]), .Z(n60) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_31 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n61, n62;
    VMW_NOR2 U3 ( .A(A[6]), .B(n61), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[1]), .B(A[0]), .Z(n62) );
    VMW_AND5 U4 ( .A(A[2]), .B(n62), .C(A[4]), .D(A[5]), .E(A[3]), .Z(n61) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_30 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n63;
    VMW_NOR2 U3 ( .A(A[6]), .B(n63), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[4]), .B(A[5]), .C(A[3]), .Z(n63) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_29 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n66, n65;
    VMW_AOI21 U3 ( .A(A[5]), .B(n64), .C(A[6]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(n66), .B(A[4]), .Z(n64) );
    VMW_INV U6 ( .A(n65), .Z(n66) );
    VMW_OAI211 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(A[3]), .Z(n65) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_28 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n67;
    VMW_AND3 U3 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n67) );
    VMW_NOR5 U4 ( .A(A[3]), .B(n67), .C(A[4]), .D(A[6]), .E(A[5]), .Z(LT_LE)
         );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_27 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n68;
    VMW_AND5 U3 ( .A(A[1]), .B(A[2]), .C(A[4]), .D(A[0]), .E(A[3]), .Z(n68) );
    VMW_NOR3 U4 ( .A(n68), .B(A[6]), .C(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_26 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n69, n70;
    VMW_AOI21 U3 ( .A(A[5]), .B(n69), .C(A[6]), .Z(LT_LE) );
    VMW_OR4 U5 ( .A(A[2]), .B(n70), .C(A[4]), .D(A[3]), .Z(n69) );
    VMW_AND2 U4 ( .A(A[0]), .B(A[1]), .Z(n70) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_25 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n71, n72;
    VMW_NOR3 U3 ( .A(n71), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n72) );
    VMW_AND3 U4 ( .A(A[4]), .B(n72), .C(A[3]), .Z(n71) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_24 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n73, n74;
    VMW_NOR2 U3 ( .A(n73), .B(A[6]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n74), .Z(n73) );
    VMW_OAI211 U4 ( .A(A[3]), .B(A[2]), .C(A[5]), .D(A[4]), .Z(n74) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_23 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n75, n76;
    VMW_NOR3 U3 ( .A(n75), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n76) );
    VMW_AND3 U4 ( .A(A[4]), .B(n76), .C(A[3]), .Z(n75) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_22 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n77;
    VMW_NOR4 U3 ( .A(n77), .B(A[1]), .C(A[3]), .D(A[2]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[6]), .B(A[5]), .C(A[4]), .Z(n77) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_21 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR3 U3 ( .A(A[4]), .B(A[6]), .C(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_20 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n78, n79;
    VMW_AOI21 U3 ( .A(A[5]), .B(n78), .C(A[6]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[3]), .B(n79), .C(A[4]), .Z(n78) );
    VMW_OR3 U4 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n79) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_19 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n81, n80;
    VMW_AOI211 U3 ( .A(A[4]), .B(n80), .C(A[6]), .D(A[5]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[2]), .B(n81), .C(A[3]), .Z(n80) );
    VMW_OR2 U4 ( .A(A[1]), .B(A[0]), .Z(n81) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_18 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n82, n83;
    VMW_AOI211 U3 ( .A(A[2]), .B(n82), .C(n83), .D(A[3]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[1]), .B(A[0]), .Z(n82) );
    VMW_OR3 U4 ( .A(A[6]), .B(A[5]), .C(A[4]), .Z(n83) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_17 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n84;
    VMW_NOR3 U3 ( .A(n84), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[2]), .B(A[3]), .C(A[4]), .Z(n84) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_16 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n85, n86;
    VMW_AOI21 U3 ( .A(A[5]), .B(n85), .C(A[6]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[4]), .B(n86), .Z(n85) );
    VMW_AND4 U4 ( .A(A[1]), .B(A[3]), .C(A[0]), .D(A[2]), .Z(n86) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_15 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n87;
    VMW_NOR2 U3 ( .A(A[6]), .B(n87), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[2]), .B(A[3]), .C(A[4]), .D(A[5]), .Z(n87) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_14 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n88;
    VMW_AOI211 U3 ( .A(A[4]), .B(n88), .C(A[6]), .D(A[5]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n88) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_13 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n89;
    VMW_NOR3 U3 ( .A(n89), .B(A[6]), .C(A[5]), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[1]), .B(A[3]), .C(A[4]), .D(A[2]), .Z(n89) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_12 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n90, n91;
    VMW_NOR2 U3 ( .A(A[6]), .B(n90), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n91) );
    VMW_AND4 U4 ( .A(A[3]), .B(A[4]), .C(A[5]), .D(n91), .Z(n90) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_11 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n93, n92;
    VMW_NOR2 U3 ( .A(A[6]), .B(n92), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[1]), .B(A[2]), .C(A[3]), .Z(n93) );
    VMW_AND3 U4 ( .A(A[5]), .B(n93), .C(A[4]), .Z(n92) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_10 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n94, n95;
    VMW_NOR2 U3 ( .A(A[6]), .B(n94), .Z(LT_LE) );
    VMW_AND3 U5 ( .A(A[5]), .B(A[2]), .C(A[1]), .Z(n95) );
    VMW_AND4 U4 ( .A(A[3]), .B(A[4]), .C(A[0]), .D(n95), .Z(n94) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_9 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n97, n96;
    VMW_AOI21 U3 ( .A(A[5]), .B(n96), .C(A[6]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n97), .Z(n96) );
    VMW_AOI211 U4 ( .A(A[1]), .B(A[2]), .C(A[4]), .D(A[3]), .Z(n97) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_8 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n99, n98;
    VMW_AOI21 U3 ( .A(A[5]), .B(n98), .C(A[6]), .Z(LT_LE) );
    VMW_OR4 U5 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(n99), .Z(n98) );
    VMW_OR2 U4 ( .A(A[4]), .B(A[3]), .Z(n99) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_7 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n100, n101;
    VMW_AND3 U3 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n100) );
    VMW_OR2 U5 ( .A(n100), .B(A[3]), .Z(n101) );
    VMW_AOI211 U4 ( .A(A[4]), .B(n101), .C(A[6]), .D(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_6 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n103, n102;
    VMW_AOI21 U3 ( .A(A[5]), .B(n102), .C(A[6]), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[4]), .B(A[3]), .C(n103), .Z(n102) );
    VMW_AND3 U4 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n103) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_5 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n104;
    VMW_AOI21 U3 ( .A(A[5]), .B(n104), .C(A[6]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[4]), .B(A[3]), .Z(n104) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_4 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n105;
    VMW_AOI211 U3 ( .A(A[4]), .B(n105), .C(A[5]), .D(A[6]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[3]), .B(A[2]), .Z(n105) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_3 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n107, n106;
    VMW_NOR2 U3 ( .A(A[6]), .B(n106), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[2]), .B(A[1]), .Z(n107) );
    VMW_AND4 U4 ( .A(A[3]), .B(A[4]), .C(A[5]), .D(n107), .Z(n106) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_2 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n108;
    VMW_NOR4 U3 ( .A(A[6]), .B(A[5]), .C(A[4]), .D(n108), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n108) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n109, n110;
    VMW_AOI21 U3 ( .A(A[5]), .B(n109), .C(A[6]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[3]), .B(n110), .C(A[4]), .Z(n109) );
    VMW_AO21 U4 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n110) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_0 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [6:0] A;
input  [6:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n112, n111;
    VMW_AOI211 U3 ( .A(A[4]), .B(n111), .C(A[6]), .D(A[5]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n112), .Z(n111) );
    VMW_AOI211 U4 ( .A(A[0]), .B(A[1]), .C(A[3]), .D(A[2]), .Z(n112) );
endmodule


module NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, CallIn, ReturnIn, ColIn, PDiagIn, 
    NDiagIn, CallOut, ReturnOut, ColOut, PDiagOut, NDiagOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [6:0] Id;
input  [63:0] ColIn;
output [63:0] ColOut;
input  [6:0] ScanIn;
output [6:0] ScanOut;
input  [63:0] NDiagIn;
output [63:0] PDiagOut;
output [63:0] NDiagOut;
input  [63:0] PDiagIn;
input  Clk, Reset, RD, WR, ScanEnable, CallIn, ReturnIn;
output CallOut, ReturnOut;
    wire \NDiagOut[0] , n7456, n7824, n7888, n7918, n7766, n7471, n7741, n1526, 
        n7803, n7634, n1590, n7494, n7504, n7523, n7613, n7783, n7876, n7404, 
        n7423, n7438, n7683, n7698, n7708, n1574, n7713, n758, n7851, n7594, 
        n7734, n7608, n7798, n7538, n7893, n7903, n7571, ReturnOut1761, n7641, 
        n7666, n7556, n7924, n7478, n7818, n7748, n7881, n1638, n7911, n7563, 
        n7653, n7936, n7674, n7431, n7544, n7691, n7701, n934, n998, n7843, 
        n7864, n7586, n7397, n7416, n7726, n1350, Logic11, n7626, n7858, n7486, 
        n7516, n7531, n7601, n7791, n966, n7444, n7578, n7648, n7836, n7463, 
        n7774, n7753, n1302, n7811, n7878, n7443, n7464, n7668, n7558, n7816, 
        n7754, n7773, n7831, n1270, n7606, n7796, n7536, n7411, n7481, n7511, 
        n7621, n1446, n7721, n7581, n7863, n7436, n7844, n7696, n7458, n7706, 
        n7768, n7931, n7543, n694, n7654, n7673, n1414, n1222, n7886, n7916, 
        n7564, n7923, n7551, n7661, n7646, n7894, n7904, n7403, n7576, n7871, 
        n7733, n854, n7838, n7593, n7424, n7856, n7488, n7684, n7714, n7518, 
        n7628, n7493, n7524, n7614, n7784, n7503, n678, n7633, n806, n7399, 
        n7588, n7418, n7728, n7804, n1190, n7476, n7746, n7938, n7451, n7761, 
        n7823, n7459, n7769, n7930, n7542, n7887, \n1806[1] , n7672, n7655, 
        n7565, n7917, n7720, n7410, n7580, n7437, n7862, n7845, n7707, n7697, 
        n7879, n7607, n7797, n7537, n7480, n7510, n7620, n1238, n7442, n7465, 
        n7559, n7669, n7817, n7755, n7772, n7830, n7805, n7477, n7747, n7450, 
        n7760, n1286, n7822, \n1806[5] , n7615, n7785, n7492, n7525, n1174, 
        n7502, n7632, n7398, n7419, n7402, n7870, n7589, n7729, n7732, n7425, 
        n7592, n7857, n7489, n7685, n7715, n7629, n7519, n662, n7922, n1126, 
        n7550, n7660, n7647, n7895, n7905, n7892, n7577, n7570, n7839, n7902, 
        n7640, n7667, n7557, n7877, n7925, n7405, n7422, n7682, n7712, n7819, 
        n710, n7595, n7850, n7539, n7609, n7735, n7799, n7635, n7495, n7505, 
        n7522, n7612, n7782, n7439, n7457, n7699, n7709, n742, n7825, n7889, 
        n7767, n7740, n7470, n7802, n7919, n7445, n7579, n7649, n1622, n7837, 
        n7462, n7775, n7752, n7810, n1014, n7627, n982, n7859, n7487, n7517, 
        n7530, n7600, n7790, n7430, n7690, n7700, n7842, n1046, n7396, n7865, 
        n7417, n7587, n7727, n7479, n7749, n7880, n7910, n1318, n7937, 
        \n1806[3] , n7562, n7652, n7675, n7545, n7569, n7659, n950, n1398, 
        n7455, n7472, n7742, n7800, n1334, n7827, n7520, n7765, n7849, n7610, 
        n7780, n7637, n7497, n7507, n7875, n902, n7407, n7597, n7680, n7710, 
        n7737, n7420, n1366, n7852, n7890, n7927, n7469, \n1806[2] , n7665, 
        n7759, n7555, n1094, n7900, n7572, n7642, n7935, n7677, n7547, n7882, 
        n7912, n7560, n7394, n7650, n7809, n7415, n7432, n7585, n7725, n1542, 
        n7867, n7692, n7702, n7840, n7429, n7485, \n1806[6] , n7529, n7619, 
        n7789, n7532, n7602, n7792, n7625, n7515, n7689, n7719, n1078, n7447, 
        n7460, n7750, n7812, n7899, n7909, n1510, n7835, n7777, n7770, n790, 
        n7440, n7832, n7815, n7929, n7467, n7757, n7409, n7482, n7512, 
        \n1806[4] , n7605, n7622, n7795, n1254, n1462, n7535, n7599, n7739, 
        n7393, n7412, n7435, n7847, n7582, n7695, n7705, n7722, n7860, n1158, 
        n7499, n7509, n7639, n7657, n1430, n7885, n7915, n7932, n7567, n7540, 
        n7670, n1206, n7829, n7897, n7907, n7449, \n1806[0] , n7779, n870, 
        n7575, n7645, n7920, n7552, n7427, n7662, CallOut1768, n7855, n7687, 
        n7717, n7400, n7730, n7490, n7872, n7590, n822, n7869, n7500, n7630, 
        n7527, n7617, n7787, n7549, n7679, n7452, n7762, n7475, n7820, n7745, 
        n7807, n7656, n7884, n7914, n1110, n7933, n7566, n7413, n7434, n7541, 
        n7671, n7828, n7846, n7694, n7704, n7723, n7861, n7583, n7483, n7638, 
        n1478, n886, n7498, n7508, n7513, n7604, n7623, n7794, n7408, n1142, 
        n7534, n7598, n7738, n7441, n7771, n7833, n7814, n7466, n7756, n7928, 
        n7548, n7678, n7453, n7763, n1494, n7474, n7821, n7744, n7806, n7868, 
        n7491, n7501, n7631, n7786, n7616, n7526, n7426, n646, n7854, n7686, 
        n7716, n7401, n7591, n7731, n838, n7873, n7448, n7778, n7896, n7574, 
        n7644, n7906, n7921, n7553, n7663, n7468, n7664, n7758, n1382, n7891, 
        n7901, n7926, n7554, n7573, n7643, n7874, n7406, n7596, n7736, n7421, 
        n7681, n7711, n7853, n7521, n7848, n7611, n7781, n918, n7636, n7496, 
        n7506, n7658, n7568, n7454, n7473, n7743, n7801, n7826, n7461, n7751, 
        n7764, n1606, n7813, n7446, n1030, n7834, n7776, n7898, n7908, n7533, 
        n7603, n7793, n7428, n7484, n7514, n7624, n7688, n7718, n1558, n774, 
        n7395, n7414, n7584, n1062, n7866, n7433, n7724, n7693, n7703, n7841, 
        n7528, n7618, n7788, n7676, n7934, n7546, n7883, n7561, n7913, n7651, 
        n7808, n726;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 , UNCONNECTED_23 , UNCONNECTED_24 , 
	UNCONNECTED_25 , UNCONNECTED_26 , UNCONNECTED_27 , UNCONNECTED_28 , 
	UNCONNECTED_29 , UNCONNECTED_30 , UNCONNECTED_31 , UNCONNECTED_32 , 
	UNCONNECTED_33 , UNCONNECTED_34 , UNCONNECTED_35 , UNCONNECTED_36 , 
	UNCONNECTED_37 , UNCONNECTED_38 , UNCONNECTED_39 , UNCONNECTED_40 , 
	UNCONNECTED_41 , UNCONNECTED_42 , UNCONNECTED_43 , UNCONNECTED_44 , 
	UNCONNECTED_45 , UNCONNECTED_46 , UNCONNECTED_47 , UNCONNECTED_48 , 
	UNCONNECTED_49 , UNCONNECTED_50 , UNCONNECTED_51 , UNCONNECTED_52 , 
	UNCONNECTED_53 , UNCONNECTED_54 , UNCONNECTED_55 , UNCONNECTED_56 , 
	UNCONNECTED_57 ;
    assign PDiagOut[63] = \NDiagOut[0] ;
    assign NDiagOut[0] = \NDiagOut[0] ;
    VMW_PULLDOWN U1325 ( .Z(n7880) );
    VMW_PULLDOWN U1350 ( .Z(n7905) );
    VMW_PULLDOWN U1377 ( .Z(n7932) );
    VMW_NOR3 U1656 ( .A(n7677), .B(n7691), .C(n7679), .Z(n7690) );
    VMW_NAND4 U1828 ( .A(n7806), .B(n7506), .C(n7482), .D(n7458), .Z(n7740) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_12 gt_104_4 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7888), .TC(n7888), .LT_LE(
        n710) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_47 gt_104_37 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_1}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7923), .TC(n7923), 
        .LT_LE(n1238) );
    VMW_NOR2 U1884 ( .A(CallIn), .B(n758), .Z(n7828) );
    VMW_OR4 U1914 ( .A(n7847), .B(NDiagIn[33]), .C(ColIn[33]), .D(PDiagIn[33]), 
        .Z(n7673) );
    VMW_OR2 U1541 ( .A(NDiagIn[41]), .B(n7415), .Z(NDiagOut[42]) );
    VMW_OR2 U1566 ( .A(NDiagIn[16]), .B(n7448), .Z(NDiagOut[17]) );
    VMW_OAI211 U1933 ( .A(n7643), .B(n7646), .C(n7580), .D(n7860), .Z(n7859)
         );
    VMW_OR2 U1389 ( .A(n7396), .B(PDiagIn[60]), .Z(PDiagOut[59]) );
    VMW_OR2 U1392 ( .A(n7399), .B(PDiagIn[57]), .Z(PDiagOut[56]) );
    VMW_NAND2 U1434 ( .A(n7449), .B(n7450), .Z(PDiagOut[14]) );
    VMW_OR2 U1498 ( .A(ColIn[14]), .B(n7451), .Z(ColOut[14]) );
    VMW_OR2 U1508 ( .A(ColIn[4]), .B(n7466), .Z(ColOut[4]) );
    VMW_AND2 U1638 ( .A(n7621), .B(n7652), .Z(n7586) );
    VMW_NAND2 U1671 ( .A(ScanOut[4]), .B(ScanOut[3]), .Z(n7711) );
    VMW_INV U2050 ( .A(n7569), .Z(n7654) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_56 gt_104_10 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7931), .TC(n7931), .LT_LE(
        n806) );
    VMW_INV U2019 ( .A(n7677), .Z(n7802) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_48 gt_104_59 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_2, UNCONNECTED_3}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n7924), .TC(n7924), .LT_LE(n1590) );
    VMW_NOR2 U1846 ( .A(CallIn), .B(n1238), .Z(n7811) );
    VMW_AND2 U1583 ( .A(n7510), .B(n7511), .Z(ReturnOut1761) );
    VMW_NOR4 U1694 ( .A(n7735), .B(NDiagIn[10]), .C(ColIn[10]), .D(PDiagIn[10]
        ), .Z(n7614) );
    VMW_OR4 U1704 ( .A(n7745), .B(NDiagIn[36]), .C(ColIn[36]), .D(PDiagIn[36]), 
        .Z(n7680) );
    VMW_OAI211 U1723 ( .A(CallIn), .B(n1302), .C(n7633), .D(n7636), .Z(n7758)
         );
    VMW_NOR2 U1861 ( .A(CallIn), .B(n1014), .Z(n7818) );
    VMW_OR2 U1413 ( .A(n7420), .B(PDiagIn[36]), .Z(PDiagOut[35]) );
    VMW_AOI211 U1598 ( .A(n7548), .B(n7549), .C(n7545), .D(n7550), .Z(n7547)
         );
    VMW_OR2 U1408 ( .A(n7415), .B(PDiagIn[41]), .Z(PDiagOut[40]) );
    VMW_NAND2 U1483 ( .A(n7429), .B(n7472), .Z(ColOut[29]) );
    VMW_NAND2 U1513 ( .A(n7487), .B(n7488), .Z(\n1806[6] ) );
    VMW_AO21 U1738 ( .A(n7649), .B(n7774), .C(n7585), .Z(n7773) );
    VMW_INV U1961 ( .A(PDiagIn[13]), .Z(n7452) );
    VMW_OR4 U1604 ( .A(n7572), .B(n7566), .C(n7573), .D(n7574), .Z(n7571) );
    VMW_NOR2 U1623 ( .A(n7555), .B(n7614), .Z(n7552) );
    VMW_AND2 U1794 ( .A(n7790), .B(n7705), .Z(n7442) );
    VMW_INV U2002 ( .A(ReturnIn), .Z(n7703) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_19 gt_104_42 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7895), .TC(n7895), .LT_LE(
        n1318) );
    VMW_OAI211 U1946 ( .A(n7582), .B(n7635), .C(n7640), .D(n7637), .Z(n7865)
         );
    VMW_INV U2025 ( .A(n7512), .Z(n7511) );
    VMW_OR2 U1441 ( .A(n7460), .B(PDiagIn[8]), .Z(PDiagOut[7]) );
    VMW_OR2 U1534 ( .A(NDiagIn[48]), .B(n7408), .Z(NDiagOut[49]) );
    VMW_NOR2 U1771 ( .A(n7608), .B(n7611), .Z(n7413) );
    VMW_NOR2 U1928 ( .A(CallIn), .B(n1590), .Z(n7857) );
    VMW_NOR2 U1833 ( .A(CallIn), .B(n1494), .Z(n7735) );
    VMW_OR2 U1453 ( .A(ColIn[59]), .B(n7397), .Z(ColOut[59]) );
    VMW_OR2 U1466 ( .A(ColIn[46]), .B(n7410), .Z(ColOut[46]) );
    VMW_AND2 U1814 ( .A(n7705), .B(n7800), .Z(n7486) );
    VMW_INV U1984 ( .A(ScanOut[1]), .Z(n7610) );
    VMW_NOR2 U1756 ( .A(n7612), .B(n7715), .Z(n7398) );
    VMW_NOR2 U1763 ( .A(n7608), .B(n7720), .Z(n7405) );
    VMW_OR4 U1821 ( .A(PDiagIn[0]), .B(n7487), .C(ColIn[0]), .D(NDiagIn[0]), 
        .Z(n7697) );
    VMW_PULLDOWN U1322 ( .Z(n7877) );
    VMW_PULLDOWN U1330 ( .Z(n7885) );
    VMW_PULLDOWN U1337 ( .Z(n7892) );
    VMW_PULLDOWN U1359 ( .Z(n7914) );
    VMW_OR2 U1474 ( .A(ColIn[38]), .B(n7418), .Z(ColOut[38]) );
    VMW_OR2 U1678 ( .A(n7604), .B(n7717), .Z(n7718) );
    VMW_NAND2 U1744 ( .A(n7780), .B(n7680), .Z(n7779) );
    VMW_AND2 U1806 ( .A(n7796), .B(n7705), .Z(n7460) );
    VMW_INV U1996 ( .A(NDiagIn[11]), .Z(n7505) );
    VMW_INV U2059 ( .A(n7826), .Z(n7656) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_63 gt_104_19 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_4, UNCONNECTED_5}), .B({\NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n7938), .TC(n7938), .LT_LE(n950) );
    VMW_NAND2 U1491 ( .A(n7441), .B(n7476), .Z(ColOut[21]) );
    VMW_OR2 U1548 ( .A(NDiagIn[34]), .B(n7422), .Z(NDiagOut[35]) );
    VMW_NAND2 U1501 ( .A(n7456), .B(n7481), .Z(ColOut[11]) );
    VMW_OR2 U1526 ( .A(NDiagIn[56]), .B(n7400), .Z(NDiagOut[57]) );
    VMW_NAND2 U1616 ( .A(ScanOut[2]), .B(ScanOut[1]), .Z(n7604) );
    VMW_NAND3 U1631 ( .A(n7636), .B(n7637), .C(n7633), .Z(n7635) );
    VMW_INV U1973 ( .A(ColIn[19]), .Z(n7477) );
    VMW_INV U2010 ( .A(n7633), .Z(n7854) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_49 gt_104_50 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7925), .TC(n7925), .LT_LE(
        n1446) );
    VMW_AND2 U1786 ( .A(n7786), .B(n7705), .Z(n7430) );
    VMW_INV U2037 ( .A(n7721), .Z(n7798) );
    VMW_PULLDOWN U1342 ( .Z(n7897) );
    VMW_PULLDOWN U1365 ( .Z(n7920) );
    VMW_PULLDOWN U1380 ( .Z(n7935) );
    VMW_NAND2 U1426 ( .A(n7437), .B(n7438), .Z(PDiagOut[22]) );
    VMW_NOR2 U1868 ( .A(CallIn), .B(n918), .Z(n7737) );
    VMW_INV U1954 ( .A(PDiagIn[27]), .Z(n7431) );
    VMW_NOR2 U1686 ( .A(n7511), .B(n7727), .Z(n7726) );
    VMW_OR2 U1854 ( .A(CallIn), .B(n1190), .Z(n7644) );
    VMW_MUX2I U1716 ( .A(ScanOut[5]), .B(ScanIn[5]), .S(ScanEnable), .Z(n7489)
         );
    VMW_AO22 U1731 ( .A(n7727), .B(ScanOut[4]), .C(n7726), .D(ScanIn[4]), .Z(
        n7523) );
    VMW_OR2 U1401 ( .A(n7408), .B(PDiagIn[48]), .Z(PDiagOut[47]) );
    VMW_OR2 U1574 ( .A(NDiagIn[8]), .B(n7460), .Z(NDiagOut[9]) );
    VMW_AO21 U1591 ( .A(n7527), .B(n7528), .C(n7529), .Z(n7526) );
    VMW_NAND2 U1644 ( .A(n7664), .B(n7665), .Z(n7663) );
    VMW_NOR2 U1873 ( .A(CallIn), .B(n870), .Z(n7757) );
    VMW_INV U1968 ( .A(ColIn[29]), .Z(n7472) );
    VMW_INV U2065 ( .A(n7676), .Z(n7850) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_9 gt_104_25 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_6}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7885), .TC(
        n7885), .LT_LE(n1046) );
    VMW_OR4 U1896 ( .A(n7835), .B(NDiagIn[61]), .C(ColIn[61]), .D(PDiagIn[61]), 
        .Z(n7694) );
    VMW_OAI211 U1906 ( .A(n7542), .B(n7677), .C(n7780), .D(n7801), .Z(n7844)
         );
    VMW_PULLDOWN U1345 ( .Z(n7900) );
    VMW_OR2 U1448 ( .A(n7470), .B(PDiagIn[1]), .Z(PDiagOut[0]) );
    VMW_NAND2 U1553 ( .A(n7429), .B(n7496), .Z(NDiagOut[30]) );
    VMW_AO21 U1663 ( .A(n7703), .B(n7487), .C(Reset), .Z(n7512) );
    VMW_OAI211 U1921 ( .A(n7547), .B(n7641), .C(n7853), .D(n7639), .Z(n7782)
         );
    VMW_INV U2042 ( .A(n7730), .Z(n7630) );
    VMW_OR2 U1554 ( .A(NDiagIn[28]), .B(n7430), .Z(NDiagOut[29]) );
    VMW_NOR2 U1664 ( .A(ScanOut[6]), .B(ScanOut[5]), .Z(n7704) );
    VMW_NOR2 U1778 ( .A(n7612), .B(n7721), .Z(n7420) );
    VMW_OR2 U1926 ( .A(CallIn), .B(n1574), .Z(n7856) );
    VMW_INV U2045 ( .A(n7680), .Z(n7562) );
    VMW_PULLDOWN U1362 ( .Z(n7917) );
    VMW_OR4 U1891 ( .A(n7833), .B(NDiagIn[60]), .C(ColIn[60]), .D(PDiagIn[60]), 
        .Z(n7695) );
    VMW_AO21 U1901 ( .A(n7839), .B(n7657), .C(n7659), .Z(n7840) );
    VMW_OR2 U1387 ( .A(n7394), .B(PDiagIn[62]), .Z(PDiagOut[61]) );
    VMW_OR2 U1406 ( .A(n7413), .B(PDiagIn[43]), .Z(PDiagOut[42]) );
    VMW_OR2 U1468 ( .A(ColIn[44]), .B(n7412), .Z(ColOut[44]) );
    VMW_NAND2 U1573 ( .A(n7459), .B(n7506), .Z(NDiagOut[10]) );
    VMW_AND2 U1643 ( .A(n7662), .B(n7658), .Z(n7557) );
    VMW_INV U2062 ( .A(n7694), .Z(n7837) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_20 gt_104_22 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7896), .TC(n7896), 
        .LT_LE(n998) );
    VMW_AOI211 U1596 ( .A(n7543), .B(n7544), .C(n7539), .D(n7535), .Z(n7542)
         );
    VMW_NOR2 U1758 ( .A(n7612), .B(n7716), .Z(n7400) );
    VMW_NOR2 U1874 ( .A(CallIn), .B(n854), .Z(n7750) );
    VMW_OR2 U1421 ( .A(n7430), .B(PDiagIn[28]), .Z(PDiagOut[27]) );
    VMW_OR2 U1681 ( .A(n7709), .B(n7713), .Z(n7721) );
    VMW_NAND4 U1711 ( .A(n7753), .B(n7503), .C(n7479), .D(n7449), .Z(n7639) );
    VMW_OAI21 U1736 ( .A(n7556), .B(n7771), .C(n7772), .Z(n7565) );
    VMW_OR4 U1853 ( .A(n7814), .B(NDiagIn[28]), .C(ColIn[28]), .D(PDiagIn[28]), 
        .Z(n7815) );
    VMW_OAI211 U1948 ( .A(n7651), .B(n7584), .C(n7627), .D(n7628), .Z(n7866)
         );
    VMW_INV U1953 ( .A(PDiagIn[29]), .Z(n7428) );
    VMW_PULLDOWN U1379 ( .Z(n7934) );
    VMW_OR2 U1454 ( .A(ColIn[58]), .B(n7398), .Z(ColOut[58]) );
    VMW_OR2 U1473 ( .A(ColIn[39]), .B(n7417), .Z(ColOut[39]) );
    VMW_OR2 U1496 ( .A(ColIn[16]), .B(n7448), .Z(ColOut[16]) );
    VMW_NAND2 U1506 ( .A(n7463), .B(n7483), .Z(ColOut[6]) );
    VMW_OR2 U1521 ( .A(NDiagIn[61]), .B(n7395), .Z(NDiagOut[62]) );
    VMW_AND3 U1611 ( .A(n7594), .B(n7511), .C(n7595), .Z(n7522) );
    VMW_NOR2 U1781 ( .A(n7608), .B(n7725), .Z(n7423) );
    VMW_INV U2030 ( .A(n7712), .Z(n7785) );
    VMW_NOR2 U1636 ( .A(n7550), .B(n7641), .Z(n7649) );
    VMW_INV U2017 ( .A(n7663), .Z(n7693) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_38 gt_104_57 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_7}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7914), .TC(
        n7914), .LT_LE(n1558) );
    VMW_INV U1974 ( .A(ColIn[17]), .Z(n7478) );
    VMW_OR2 U1743 ( .A(n7688), .B(n7691), .Z(n7577) );
    VMW_NOR2 U1848 ( .A(CallIn), .B(n1254), .Z(n7812) );
    VMW_NAND2 U1801 ( .A(n7794), .B(n7708), .Z(n7453) );
    VMW_INV U1991 ( .A(NDiagIn[21]), .Z(n7500) );
    VMW_OR2 U1826 ( .A(CallIn), .B(n1606), .Z(n7755) );
    VMW_AND4 U1658 ( .A(n7666), .B(n7693), .C(n7694), .D(n7695), .Z(n7573) );
    VMW_NOR2 U1764 ( .A(n7612), .B(n7720), .Z(n7406) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_59 gt_104_39 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , UNCONNECTED_8, 
        UNCONNECTED_9, UNCONNECTED_10}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n7934), .TC(n7934), .LT_LE(n1270) );
    VMW_NAND2 U1428 ( .A(n7440), .B(n7441), .Z(PDiagOut[20]) );
    VMW_NAND2 U1446 ( .A(n7467), .B(n7468), .Z(PDiagOut[2]) );
    VMW_OR2 U1461 ( .A(ColIn[51]), .B(n7405), .Z(ColOut[51]) );
    VMW_OR2 U1568 ( .A(NDiagIn[14]), .B(n7451), .Z(NDiagOut[15]) );
    VMW_NOR2 U1751 ( .A(n7608), .B(n7712), .Z(n7393) );
    VMW_AO21 U1898 ( .A(n7664), .B(n7836), .C(n7831), .Z(n7534) );
    VMW_NOR2 U1908 ( .A(CallIn), .B(n1110), .Z(n7845) );
    VMW_AND2 U1813 ( .A(n7800), .B(n7708), .Z(n7470) );
    VMW_INV U1983 ( .A(ScanOut[4]), .Z(n7606) );
    VMW_NOR2 U1776 ( .A(n7612), .B(n7710), .Z(n7418) );
    VMW_OR2 U1834 ( .A(CallIn), .B(n1350), .Z(n7729) );
    VMW_OR2 U1533 ( .A(NDiagIn[49]), .B(n7407), .Z(NDiagOut[50]) );
    VMW_OR4 U1688 ( .A(n7728), .B(NDiagIn[18]), .C(ColIn[18]), .D(PDiagIn[18]), 
        .Z(n7632) );
    VMW_MUX2I U1718 ( .A(ScanOut[3]), .B(ScanIn[3]), .S(ScanEnable), .Z(n7491)
         );
    VMW_PULLDOWN U1331 ( .Z(n7886) );
    VMW_PULLDOWN U1339 ( .Z(n7894) );
    VMW_OR2 U1484 ( .A(ColIn[28]), .B(n7430), .Z(ColOut[28]) );
    VMW_NOR2 U1603 ( .A(CallIn), .B(n646), .Z(n7570) );
    VMW_NOR3 U1941 ( .A(n7574), .B(n7771), .C(n7699), .Z(n7762) );
    VMW_INV U2022 ( .A(n7687), .Z(n7543) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_35 gt_104_62 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7911), 
        .TC(n7911), .LT_LE(n1638) );
    VMW_NAND4 U1624 ( .A(n7616), .B(n7504), .C(n7480), .D(n7452), .Z(n7615) );
    VMW_NAND2 U1793 ( .A(n7790), .B(n7708), .Z(n7441) );
    VMW_INV U2005 ( .A(n7759), .Z(n7618) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_14 gt_104_45 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_11}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7890), 
        .TC(n7890), .LT_LE(n1366) );
    VMW_NAND2 U1514 ( .A(n7487), .B(n7489), .Z(\n1806[5] ) );
    VMW_OR2 U1528 ( .A(NDiagIn[54]), .B(n7402), .Z(NDiagOut[55]) );
    VMW_OR2 U1618 ( .A(n7604), .B(n7605), .Z(n7607) );
    VMW_INV U1966 ( .A(PDiagIn[3]), .Z(n7467) );
    VMW_AND2 U1788 ( .A(n7787), .B(n7705), .Z(n7433) );
    VMW_INV U2039 ( .A(n7723), .Z(n7794) );
    VMW_PULLDOWN U1357 ( .Z(n7912) );
    VMW_OR2 U1395 ( .A(n7402), .B(PDiagIn[54]), .Z(PDiagOut[53]) );
    VMW_OR2 U1414 ( .A(n7421), .B(PDiagIn[35]), .Z(PDiagOut[34]) );
    VMW_OR2 U1433 ( .A(n7448), .B(PDiagIn[16]), .Z(PDiagOut[15]) );
    VMW_NOR2 U1584 ( .A(n7512), .B(n7510), .Z(CallOut1768) );
    VMW_NAND4 U1693 ( .A(n7734), .B(n7505), .C(n7481), .D(n7455), .Z(n7622) );
    VMW_OAI211 U1724 ( .A(CallIn), .B(n1430), .C(n7759), .D(n7615), .Z(n7752)
         );
    VMW_NOR2 U1866 ( .A(CallIn), .B(n966), .Z(n7681) );
    VMW_NOR4 U1703 ( .A(n7744), .B(NDiagIn[39]), .C(ColIn[39]), .D(PDiagIn[39]
        ), .Z(n7691) );
    VMW_OR2 U1676 ( .A(n7711), .B(n7706), .Z(n7716) );
    VMW_NAND2 U1808 ( .A(n7705), .B(n7797), .Z(n7463) );
    VMW_OR4 U1841 ( .A(n7809), .B(NDiagIn[20]), .C(ColIn[20]), .D(PDiagIn[20]), 
        .Z(n7636) );
    VMW_INV U1998 ( .A(NDiagIn[6]), .Z(n7507) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_15 gt_104_3 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_12, UNCONNECTED_13}), .B({\NDiagOut[0] , Logic11, Logic11, 
        Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n7891), .TC(
        n7891), .LT_LE(n694) );
    VMW_INV U2057 ( .A(n7821), .Z(n7700) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_42 gt_104_17 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_14}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7918), .TC(n7918), .LT_LE(
        n918) );
    VMW_PULLDOWN U1370 ( .Z(n7925) );
    VMW_OR2 U1546 ( .A(NDiagIn[36]), .B(n7420), .Z(NDiagOut[37]) );
    VMW_NAND2 U1561 ( .A(n7441), .B(n7500), .Z(NDiagOut[22]) );
    VMW_OAI21 U1934 ( .A(n7561), .B(n7645), .C(n7859), .Z(n7774) );
    VMW_PULLDOWN U1378 ( .Z(n7933) );
    VMW_OR2 U1455 ( .A(ColIn[57]), .B(n7399), .Z(ColOut[57]) );
    VMW_OR2 U1472 ( .A(ColIn[40]), .B(n7416), .Z(ColOut[40]) );
    VMW_OR4 U1651 ( .A(n7681), .B(NDiagIn[43]), .C(ColIn[43]), .D(PDiagIn[43]), 
        .Z(n7536) );
    VMW_OR4 U1883 ( .A(n7827), .B(NDiagIn[55]), .C(ColIn[55]), .D(PDiagIn[55]), 
        .Z(n7661) );
    VMW_NOR2 U1913 ( .A(CallIn), .B(n1126), .Z(n7847) );
    VMW_AO21 U1742 ( .A(n7557), .B(n7558), .C(n7777), .Z(n7572) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_8 gt_104_30 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7884), .TC(n7884), 
        .LT_LE(n1126) );
    VMW_AND2 U1800 ( .A(n7705), .B(n7793), .Z(n7451) );
    VMW_INV U1990 ( .A(NDiagIn[23]), .Z(n7499) );
    VMW_OR2 U1827 ( .A(CallIn), .B(n1510), .Z(n7806) );
    VMW_NAND2 U1569 ( .A(n7453), .B(n7504), .Z(NDiagOut[14]) );
    VMW_AND4 U1659 ( .A(n7586), .B(n7696), .C(n7649), .D(n7548), .Z(n7592) );
    VMW_NOR2 U1765 ( .A(n7608), .B(n7722), .Z(n7407) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_25 gt_104_38 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7901), .TC(n7901), 
        .LT_LE(n1254) );
    VMW_OR2 U1520 ( .A(NDiagIn[62]), .B(n7394), .Z(NDiagOut[63]) );
    VMW_INV U1952 ( .A(PDiagIn[30]), .Z(n7426) );
    VMW_OR2 U1386 ( .A(n7393), .B(PDiagIn[63]), .Z(PDiagOut[62]) );
    VMW_NAND2 U1497 ( .A(n7450), .B(n7479), .Z(ColOut[15]) );
    VMW_AND4 U1610 ( .A(n7511), .B(n7591), .C(n7592), .D(n7593), .Z(n7524) );
    VMW_OR2 U1637 ( .A(n7651), .B(n7625), .Z(n7650) );
    VMW_NOR2 U1780 ( .A(n7612), .B(n7724), .Z(n7422) );
    VMW_INV U2031 ( .A(n7714), .Z(n7786) );
    VMW_INV U1975 ( .A(ColIn[15]), .Z(n7479) );
    VMW_INV U2016 ( .A(n7558), .Z(n7667) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_28 gt_104_56 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11, Logic11}), .LEQ(n7904), .TC(n7904), 
        .LT_LE(n1542) );
    VMW_NAND2 U1507 ( .A(n7465), .B(n7484), .Z(ColOut[5]) );
    VMW_NOR4 U1849 ( .A(n7812), .B(NDiagIn[25]), .C(ColIn[25]), .D(PDiagIn[25]
        ), .Z(n7529) );
    VMW_NOR2 U1875 ( .A(CallIn), .B(n838), .Z(n7751) );
    VMW_OR2 U1407 ( .A(n7414), .B(PDiagIn[42]), .Z(PDiagOut[41]) );
    VMW_AND2 U1597 ( .A(n7546), .B(n7526), .Z(n7545) );
    VMW_PULLDOWN U1323 ( .Z(n7878) );
    VMW_PULLDOWN U1338 ( .Z(n7893) );
    VMW_PULLDOWN U1344 ( .Z(n7899) );
    VMW_NAND2 U1420 ( .A(n7428), .B(n7429), .Z(PDiagOut[28]) );
    VMW_OR2 U1680 ( .A(n7609), .B(n7717), .Z(n7720) );
    VMW_AO21 U1737 ( .A(n7690), .B(n7689), .C(n7669), .Z(n7564) );
    VMW_NOR4 U1710 ( .A(PDiagIn[14]), .B(ColIn[14]), .C(NDiagIn[14]), .D(n7752
        ), .Z(n7619) );
    VMW_NOR2 U1852 ( .A(CallIn), .B(n1206), .Z(n7814) );
    VMW_AND2 U1665 ( .A(n7613), .B(n7704), .Z(n7705) );
    VMW_NAND3 U1949 ( .A(n7866), .B(n7626), .C(n7623), .Z(n7867) );
    VMW_INV U2044 ( .A(n7622), .Z(n7741) );
    VMW_FD CallOut_reg ( .D(CallOut1768), .CP(Clk), .Q(CallOut) );
    VMW_NAND4 U1927 ( .A(n7856), .B(n7508), .C(n7484), .D(n7464), .Z(n7626) );
    VMW_PULLDOWN U1356 ( .Z(n7911) );
    VMW_PULLDOWN U1363 ( .Z(n7918) );
    VMW_NAND2 U1555 ( .A(n7432), .B(n7497), .Z(NDiagOut[28]) );
    VMW_OR2 U1572 ( .A(NDiagIn[10]), .B(n7457), .Z(NDiagOut[11]) );
    VMW_NOR2 U1890 ( .A(CallIn), .B(n694), .Z(n7833) );
    VMW_AO21 U1900 ( .A(n7838), .B(n7660), .C(n7826), .Z(n7839) );
    VMW_FD \MyColumn_reg[5]  ( .D(n7870), .CP(Clk), .Q(ScanOut[5]) );
    VMW_OR2 U1469 ( .A(ColIn[43]), .B(n7413), .Z(ColOut[43]) );
    VMW_NAND2 U1642 ( .A(n7660), .B(n7661), .Z(n7558) );
    VMW_INV U2063 ( .A(n7780), .Z(n7678) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_5 gt_104_23 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , UNCONNECTED_15, 
        UNCONNECTED_16, UNCONNECTED_17}), .B({\NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n7881), .TC(n7881), .LT_LE(n1014) );
    VMW_OR2 U1547 ( .A(NDiagIn[35]), .B(n7421), .Z(NDiagOut[36]) );
    VMW_OR2 U1677 ( .A(n7606), .B(ScanOut[3]), .Z(n7717) );
    VMW_NOR2 U1759 ( .A(n7608), .B(n7718), .Z(n7401) );
    VMW_NAND2 U1809 ( .A(n7798), .B(n7708), .Z(n7465) );
    VMW_INV U1999 ( .A(NDiagIn[5]), .Z(n7508) );
    VMW_INV U2056 ( .A(n7536), .Z(n7683) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_31 gt_104_2 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, Logic11, 
        \NDiagOut[0] , Logic11}), .LEQ(n7907), .TC(n7907), .LT_LE(n678) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_16 gt_104_16 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        Logic11, Logic11, Logic11}), .LEQ(n7892), .TC(n7892), .LT_LE(n902) );
    VMW_PULLDOWN U1371 ( .Z(n7926) );
    VMW_OAI21 U1935 ( .A(n7773), .B(n7775), .C(n7586), .Z(n7861) );
    VMW_OR2 U1560 ( .A(NDiagIn[22]), .B(n7439), .Z(NDiagOut[23]) );
    VMW_NAND2 U1619 ( .A(ScanOut[0]), .B(n7602), .Z(n7608) );
    VMW_NAND2 U1650 ( .A(n7563), .B(n7680), .Z(n7679) );
    VMW_NOR2 U1882 ( .A(CallIn), .B(n774), .Z(n7827) );
    VMW_NOR4 U1912 ( .A(n7846), .B(NDiagIn[31]), .C(ColIn[31]), .D(PDiagIn[31]
        ), .Z(n7671) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_40 gt_104_31 ( .A({
        \n1806[6] , \n1806[5] , UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22}), .B({\NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] }), .LEQ(n7916), .TC(n7916), .LT_LE(n1142) );
    VMW_AND2 U1789 ( .A(n7788), .B(n7708), .Z(n7434) );
    VMW_INV U2038 ( .A(n7722), .Z(n7792) );
    VMW_OR2 U1394 ( .A(n7401), .B(PDiagIn[55]), .Z(PDiagOut[54]) );
    VMW_OR2 U1529 ( .A(NDiagIn[53]), .B(n7403), .Z(NDiagOut[54]) );
    VMW_OR3 U1585 ( .A(n7513), .B(n7514), .C(n7515), .Z(n7875) );
    VMW_OR2 U1415 ( .A(n7422), .B(PDiagIn[34]), .Z(PDiagOut[33]) );
    VMW_OR2 U1429 ( .A(n7442), .B(PDiagIn[20]), .Z(PDiagOut[19]) );
    VMW_NAND2 U1432 ( .A(n7446), .B(n7447), .Z(PDiagOut[16]) );
    VMW_AND2 U1692 ( .A(n7586), .B(n7639), .Z(n7595) );
    VMW_OR2 U1702 ( .A(n7648), .B(n7529), .Z(n7581) );
    VMW_AND4 U1725 ( .A(n7573), .B(n7739), .C(n7760), .D(n7530), .Z(n7702) );
    VMW_NOR2 U1867 ( .A(CallIn), .B(n902), .Z(n7736) );
    VMW_NOR2 U1840 ( .A(CallIn), .B(n1334), .Z(n7809) );
    VMW_NAND4 U1689 ( .A(n7729), .B(n7501), .C(n7477), .D(n7443), .Z(n7640) );
    VMW_MUX2I U1719 ( .A(ScanOut[2]), .B(ScanIn[2]), .S(ScanEnable), .Z(n7492)
         );
    VMW_PULLDOWN U1324 ( .Z(n7879) );
    VMW_OR2 U1388 ( .A(n7395), .B(PDiagIn[61]), .Z(PDiagOut[60]) );
    VMW_OR2 U1409 ( .A(n7416), .B(PDiagIn[40]), .Z(PDiagOut[39]) );
    VMW_NAND2 U1440 ( .A(n7458), .B(n7459), .Z(PDiagOut[8]) );
    VMW_OR2 U1447 ( .A(n7469), .B(PDiagIn[2]), .Z(PDiagOut[1]) );
    VMW_OR2 U1460 ( .A(ColIn[52]), .B(n7404), .Z(ColOut[52]) );
    VMW_NAND2 U1485 ( .A(n7432), .B(n7473), .Z(ColOut[27]) );
    VMW_NAND2 U1515 ( .A(n7487), .B(n7490), .Z(\n1806[4] ) );
    VMW_OR2 U1532 ( .A(NDiagIn[50]), .B(n7406), .Z(NDiagOut[51]) );
    VMW_NOR3 U1602 ( .A(n7567), .B(n7568), .C(n7569), .Z(n7566) );
    VMW_AND2 U1792 ( .A(n7789), .B(n7705), .Z(n7439) );
    VMW_NAND4 U1940 ( .A(n7740), .B(n7803), .C(n7639), .D(n7769), .Z(n7597) );
    VMW_FD \MyColumn_reg[1]  ( .D(n7874), .CP(Clk), .Q(ScanOut[1]) );
    VMW_OR3 U1625 ( .A(n7618), .B(n7619), .C(n7620), .Z(n7617) );
    VMW_INV U2023 ( .A(n7692), .Z(n7771) );
    VMW_INV U2004 ( .A(n7611), .Z(n7795) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_0 gt_104_44 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7876), .TC(n7876), .LT_LE(
        n1350) );
    VMW_AO22 U1750 ( .A(n7727), .B(ScanOut[0]), .C(n7726), .D(ScanIn[0]), .Z(
        n7515) );
    VMW_OAI21 U1899 ( .A(n7829), .B(n7532), .C(n7661), .Z(n7838) );
    VMW_INV U1967 ( .A(ColIn[30]), .Z(n7471) );
    VMW_OR4 U1909 ( .A(n7845), .B(NDiagIn[34]), .C(ColIn[34]), .D(PDiagIn[34]), 
        .Z(n7676) );
    VMW_AND2 U1812 ( .A(n7799), .B(n7705), .Z(n7469) );
    VMW_INV U1982 ( .A(ScanOut[6]), .Z(n7603) );
    VMW_NOR2 U1770 ( .A(n7612), .B(n7723), .Z(n7412) );
    VMW_NOR2 U1777 ( .A(n7608), .B(n7721), .Z(n7419) );
    VMW_NOR2 U1835 ( .A(CallIn), .B(n1398), .Z(n7808) );
    VMW_OR4 U1929 ( .A(n7857), .B(NDiagIn[4]), .C(ColIn[4]), .D(PDiagIn[4]), 
        .Z(n7624) );
    VMW_OR2 U1832 ( .A(CallIn), .B(n1478), .Z(n7734) );
    VMW_OR2 U1467 ( .A(ColIn[45]), .B(n7411), .Z(ColOut[45]) );
    VMW_AND2 U1815 ( .A(n7726), .B(CallIn), .Z(n7513) );
    VMW_INV U1985 ( .A(ScanOut[0]), .Z(n7613) );
    VMW_NOR2 U1757 ( .A(n7608), .B(n7716), .Z(n7399) );
    VMW_NAND2 U1482 ( .A(n7427), .B(n7471), .Z(ColOut[30]) );
    VMW_AOI211 U1599 ( .A(n7552), .B(n7553), .C(n7554), .D(n7555), .Z(n7551)
         );
    VMW_AO22 U1739 ( .A(n7550), .B(n7776), .C(n7638), .D(n7635), .Z(n7775) );
    VMW_INV U1960 ( .A(PDiagIn[15]), .Z(n7449) );
    VMW_FD \MyColumn_reg[3]  ( .D(n7872), .CP(Clk), .Q(ScanOut[3]) );
    VMW_OR2 U1512 ( .A(ColIn[0]), .B(n7486), .Z(ColOut[0]) );
    VMW_OR2 U1535 ( .A(NDiagIn[47]), .B(n7409), .Z(NDiagOut[48]) );
    VMW_AOI211 U1605 ( .A(n7543), .B(n7576), .C(n7577), .D(n7578), .Z(n7575)
         );
    VMW_NAND2 U1622 ( .A(n7602), .B(n7613), .Z(n7612) );
    VMW_INV U2003 ( .A(n7607), .Z(n7793) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_4 gt_104_43 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_23, UNCONNECTED_24}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n7880), .TC(n7880), .LT_LE(n1334) );
    VMW_INV U2024 ( .A(n7699), .Z(n7739) );
    VMW_NAND2 U1795 ( .A(n7791), .B(n7708), .Z(n7444) );
    VMW_AO21 U1947 ( .A(n7629), .B(n7865), .C(n7764), .Z(n7781) );
    VMW_PULLDOWN U1336 ( .Z(n7891) );
    VMW_PULLDOWN U1343 ( .Z(n7898) );
    VMW_PULLDOWN U1351 ( .Z(n7906) );
    VMW_PULLDOWN U1376 ( .Z(n7931) );
    VMW_OR2 U1393 ( .A(n7400), .B(PDiagIn[56]), .Z(PDiagOut[55]) );
    VMW_OR2 U1412 ( .A(n7419), .B(PDiagIn[37]), .Z(PDiagOut[36]) );
    VMW_OR2 U1435 ( .A(n7451), .B(PDiagIn[14]), .Z(PDiagOut[13]) );
    VMW_NAND2 U1499 ( .A(n7453), .B(n7480), .Z(ColOut[13]) );
    VMW_OR3 U1639 ( .A(n7567), .B(n7568), .C(n7654), .Z(n7653) );
    VMW_INV U2018 ( .A(n7669), .Z(n7593) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_18 gt_104_58 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7894), .TC(
        n7894), .LT_LE(n1574) );
    VMW_NAND2 U1509 ( .A(n7468), .B(n7485), .Z(ColOut[3]) );
    VMW_OR4 U1847 ( .A(n7811), .B(NDiagIn[26]), .C(ColIn[26]), .D(PDiagIn[26]), 
        .Z(n7528) );
    VMW_NOR4 U1695 ( .A(n7736), .B(NDiagIn[47]), .C(ColIn[47]), .D(PDiagIn[47]
        ), .Z(n7574) );
    VMW_NOR4 U1705 ( .A(PDiagIn[44]), .B(ColIn[44]), .C(NDiagIn[44]), .D(n7746
        ), .Z(n7689) );
    VMW_OAI211 U1722 ( .A(CallIn), .B(n950), .C(n7682), .D(n7684), .Z(n7746)
         );
    VMW_OR4 U1860 ( .A(n7817), .B(NDiagIn[37]), .C(ColIn[37]), .D(PDiagIn[37]), 
        .Z(n7780) );
    VMW_NAND2 U1567 ( .A(n7450), .B(n7503), .Z(NDiagOut[16]) );
    VMW_OR2 U1582 ( .A(n7486), .B(NDiagIn[0]), .Z(NDiagOut[1]) );
    VMW_AND2 U1657 ( .A(n7690), .B(n7543), .Z(n7692) );
    VMW_OR2 U1829 ( .A(CallIn), .B(n1446), .Z(n7616) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_3 gt_104_5 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_25}), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7879), .TC(n7879), 
        .LT_LE(n726) );
    VMW_NOR4 U1885 ( .A(n7828), .B(NDiagIn[56]), .C(ColIn[56]), .D(PDiagIn[56]
        ), .Z(n7829) );
    VMW_NOR2 U1915 ( .A(CallIn), .B(n1142), .Z(n7848) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_23 gt_104_36 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7899), .TC(n7899), .LT_LE(
        n1222) );
    VMW_AO21 U1932 ( .A(n7801), .B(n7802), .C(n7679), .Z(n7772) );
    VMW_PULLDOWN U1364 ( .Z(n7919) );
    VMW_OR2 U1540 ( .A(NDiagIn[42]), .B(n7414), .Z(NDiagOut[43]) );
    VMW_AND4 U1645 ( .A(n7557), .B(n7667), .C(n7533), .D(n7668), .Z(n7666) );
    VMW_OR2 U1670 ( .A(n7709), .B(n7604), .Z(n7710) );
    VMW_INV U2051 ( .A(n7740), .Z(n7555) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_24 gt_104_11 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_26, UNCONNECTED_27}), .B({\NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n7900), 
        .TC(n7900), .LT_LE(n822) );
    VMW_INV U2064 ( .A(n7844), .Z(n7852) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_6 gt_104_24 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11, Logic11}), .LEQ(n7882), .TC(n7882), .LT_LE(n1030) );
    VMW_NAND2 U1552 ( .A(n7427), .B(n7495), .Z(NDiagOut[31]) );
    VMW_OR2 U1575 ( .A(NDiagIn[7]), .B(n7461), .Z(NDiagOut[8]) );
    VMW_OAI21 U1897 ( .A(n7530), .B(n7837), .C(n7695), .Z(n7836) );
    VMW_NOR2 U1907 ( .A(CallIn), .B(n1078), .Z(n7745) );
    VMW_PULLDOWN U1381 ( .Z(n7936) );
    VMW_OR2 U1400 ( .A(n7407), .B(PDiagIn[49]), .Z(PDiagOut[48]) );
    VMW_OR2 U1427 ( .A(n7439), .B(PDiagIn[22]), .Z(PDiagOut[21]) );
    VMW_OR2 U1449 ( .A(n7393), .B(ColIn[63]), .Z(ColOut[63]) );
    VMW_AND4 U1662 ( .A(n7591), .B(n7592), .C(n7692), .D(n7702), .Z(n7510) );
    VMW_NAND3 U1920 ( .A(n7854), .B(n7636), .C(n7638), .Z(n7853) );
    VMW_INV U2043 ( .A(n7766), .Z(n7594) );
    VMW_NOR2 U1779 ( .A(n7608), .B(n7724), .Z(n7421) );
    VMW_OR3 U1590 ( .A(n7513), .B(n7524), .C(n7525), .Z(n7870) );
    VMW_NOR3 U1687 ( .A(ScanEnable), .B(CallIn), .C(n7511), .Z(n7727) );
    VMW_MUX2I U1717 ( .A(ScanOut[4]), .B(ScanIn[4]), .S(ScanEnable), .Z(n7490)
         );
    VMW_AO21 U1855 ( .A(n7815), .B(n7643), .C(n7743), .Z(n7527) );
    VMW_OAI211 U1730 ( .A(n7761), .B(n7765), .C(n7696), .D(n7591), .Z(n7766)
         );
    VMW_OR2 U1490 ( .A(ColIn[22]), .B(n7439), .Z(ColOut[22]) );
    VMW_OR2 U1500 ( .A(ColIn[12]), .B(n7454), .Z(ColOut[12]) );
    VMW_NOR4 U1872 ( .A(n7822), .B(NDiagIn[48]), .C(ColIn[48]), .D(PDiagIn[48]
        ), .Z(n7568) );
    VMW_INV U1969 ( .A(ColIn[27]), .Z(n7473) );
    VMW_NAND2 U1617 ( .A(ScanOut[3]), .B(n7606), .Z(n7605) );
    VMW_NAND4 U1630 ( .A(n7634), .B(n7500), .C(n7476), .D(n7440), .Z(n7633) );
    VMW_INV U1972 ( .A(ColIn[21]), .Z(n7476) );
    VMW_INV U2011 ( .A(n7641), .Z(n7776) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_17 gt_104_51 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_28, UNCONNECTED_29}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n7893), .TC(n7893), .LT_LE(n1462) );
    VMW_NAND2 U1787 ( .A(n7787), .B(n7708), .Z(n7432) );
    VMW_INV U2036 ( .A(n7720), .Z(n7791) );
    VMW_OR2 U1452 ( .A(ColIn[60]), .B(n7396), .Z(ColOut[60]) );
    VMW_OR2 U1527 ( .A(NDiagIn[55]), .B(n7401), .Z(NDiagOut[56]) );
    VMW_NOR2 U1762 ( .A(n7612), .B(n7719), .Z(n7404) );
    VMW_NOR2 U1869 ( .A(CallIn), .B(n934), .Z(n7820) );
    VMW_INV U1955 ( .A(PDiagIn[24]), .Z(n7435) );
    VMW_OR2 U1475 ( .A(ColIn[37]), .B(n7419), .Z(ColOut[37]) );
    VMW_NOR2 U1820 ( .A(n7538), .B(n7682), .Z(n7688) );
    VMW_AND2 U1807 ( .A(n7797), .B(n7708), .Z(n7461) );
    VMW_INV U1997 ( .A(NDiagIn[9]), .Z(n7506) );
    VMW_PULLDOWN U1321 ( .Z(n7876) );
    VMW_PULLDOWN U1326 ( .Z(n7881) );
    VMW_PULLDOWN U1353 ( .Z(n7908) );
    VMW_PULLDOWN U1358 ( .Z(n7913) );
    VMW_OR2 U1549 ( .A(NDiagIn[33]), .B(n7423), .Z(NDiagOut[34]) );
    VMW_OR2 U1679 ( .A(n7713), .B(n7717), .Z(n7719) );
    VMW_AO22 U1745 ( .A(n7619), .B(n7621), .C(n7595), .D(n7781), .Z(n7587) );
    VMW_INV U2058 ( .A(n7568), .Z(n7842) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_29 gt_104_18 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7905), .TC(n7905), .LT_LE(
        n934) );
    VMW_FD \MyColumn_reg[6]  ( .D(n7869), .CP(Clk), .Q(ScanOut[6]) );
    VMW_PULLDOWN U1374 ( .Z(n7929) );
    VMW_OR2 U1542 ( .A(NDiagIn[40]), .B(n7416), .Z(NDiagOut[41]) );
    VMW_NAND2 U1565 ( .A(n7447), .B(n7502), .Z(NDiagOut[18]) );
    VMW_OR4 U1655 ( .A(n7685), .B(n7541), .C(n7688), .D(n7689), .Z(n7687) );
    VMW_OR2 U1672 ( .A(n7711), .B(n7604), .Z(n7712) );
    VMW_NOR2 U1930 ( .A(CallIn), .B(n1526), .Z(n7858) );
    VMW_INV U2053 ( .A(n7528), .Z(n7647) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_62 gt_104_13 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_30}), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7937), .TC(n7937), 
        .LT_LE(n854) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_50 gt_104_34 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7926), .TC(n7926), .LT_LE(
        n1190) );
    VMW_OR2 U1391 ( .A(n7398), .B(PDiagIn[58]), .Z(PDiagOut[57]) );
    VMW_OR2 U1410 ( .A(n7417), .B(PDiagIn[39]), .Z(PDiagOut[38]) );
    VMW_OR2 U1459 ( .A(ColIn[53]), .B(n7403), .Z(ColOut[53]) );
    VMW_NOR4 U1887 ( .A(n7830), .B(NDiagIn[58]), .C(ColIn[58]), .D(PDiagIn[58]
        ), .Z(n7831) );
    VMW_OAI21 U1917 ( .A(n7850), .B(n7675), .C(n7673), .Z(n7849) );
    VMW_MUX2I U1720 ( .A(ScanOut[1]), .B(ScanIn[1]), .S(ScanEnable), .Z(n7493)
         );
    VMW_NOR2 U1769 ( .A(n7608), .B(n7723), .Z(n7411) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_30 gt_104_7 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , UNCONNECTED_31, 
        UNCONNECTED_32, UNCONNECTED_33}), .B({\NDiagOut[0] , Logic11, Logic11, 
        Logic11, \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n7906), 
        .TC(n7906), .LT_LE(n758) );
    VMW_OR2 U1437 ( .A(n7454), .B(PDiagIn[12]), .Z(PDiagOut[11]) );
    VMW_OR2 U1580 ( .A(NDiagIn[2]), .B(n7469), .Z(NDiagOut[3]) );
    VMW_NOR4 U1862 ( .A(n7818), .B(NDiagIn[40]), .C(ColIn[40]), .D(PDiagIn[40]
        ), .Z(n7541) );
    VMW_OR2 U1537 ( .A(NDiagIn[45]), .B(n7411), .Z(NDiagOut[46]) );
    VMW_AOI211 U1607 ( .A(n7548), .B(n7583), .C(n7579), .D(n7550), .Z(n7582)
         );
    VMW_AO21 U1697 ( .A(n7739), .B(n7574), .C(n7700), .Z(n7738) );
    VMW_NAND4 U1845 ( .A(n7810), .B(n7498), .C(n7474), .D(n7435), .Z(n7546) );
    VMW_OAI21 U1707 ( .A(n7749), .B(n7628), .C(n7626), .Z(n7748) );
    VMW_INV U1979 ( .A(ColIn[6]), .Z(n7483) );
    VMW_NAND2 U1797 ( .A(n7792), .B(n7708), .Z(n7447) );
    VMW_INV U2026 ( .A(n7625), .Z(n7596) );
    VMW_PULLDOWN U1328 ( .Z(n7883) );
    VMW_PULLDOWN U1334 ( .Z(n7889) );
    VMW_PULLDOWN U1348 ( .Z(n7903) );
    VMW_OR2 U1442 ( .A(n7461), .B(PDiagIn[7]), .Z(PDiagOut[6]) );
    VMW_OR2 U1465 ( .A(ColIn[47]), .B(n7409), .Z(ColOut[47]) );
    VMW_OR2 U1480 ( .A(ColIn[32]), .B(n7424), .Z(ColOut[32]) );
    VMW_AO21 U1945 ( .A(n7672), .B(n7864), .C(n7669), .Z(n7583) );
    VMW_OR2 U1510 ( .A(ColIn[2]), .B(n7469), .Z(ColOut[2]) );
    VMW_OR2 U1620 ( .A(n7610), .B(ScanOut[2]), .Z(n7609) );
    VMW_INV U1962 ( .A(PDiagIn[11]), .Z(n7455) );
    VMW_OR4 U1879 ( .A(n7824), .B(NDiagIn[54]), .C(ColIn[54]), .D(PDiagIn[54]), 
        .Z(n7660) );
    VMW_INV U2001 ( .A(CallIn), .Z(n7487) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_39 gt_104_41 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_34}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7915), .TC(
        n7915), .LT_LE(n1302) );
    VMW_NOR2 U1755 ( .A(n7608), .B(n7715), .Z(n7397) );
    VMW_NAND2 U1817 ( .A(n7802), .B(n7691), .Z(n7801) );
    VMW_INV U1987 ( .A(NDiagIn[29]), .Z(n7496) );
    VMW_NOR2 U1772 ( .A(n7611), .B(n7612), .Z(n7414) );
    VMW_OR2 U1669 ( .A(ScanOut[4]), .B(ScanOut[3]), .Z(n7709) );
    VMW_NOR2 U1830 ( .A(CallIn), .B(n1462), .Z(n7807) );
    VMW_INV U2048 ( .A(n7639), .Z(n7585) );
    VMW_OR2 U1398 ( .A(n7405), .B(PDiagIn[51]), .Z(PDiagOut[50]) );
    VMW_NAND2 U1419 ( .A(n7426), .B(n7427), .Z(PDiagOut[29]) );
    VMW_OR2 U1450 ( .A(ColIn[62]), .B(n7394), .Z(ColOut[62]) );
    VMW_OR2 U1477 ( .A(ColIn[35]), .B(n7421), .Z(ColOut[35]) );
    VMW_NAND2 U1559 ( .A(n7438), .B(n7499), .Z(NDiagOut[24]) );
    VMW_NAND2 U1805 ( .A(n7708), .B(n7796), .Z(n7459) );
    VMW_OR3 U1939 ( .A(n7645), .B(n7669), .C(n7767), .Z(n7770) );
    VMW_INV U1995 ( .A(NDiagIn[13]), .Z(n7504) );
    VMW_AO22 U1747 ( .A(n7586), .B(n7782), .C(n7595), .D(n7732), .Z(n7554) );
    VMW_NOR2 U1760 ( .A(n7612), .B(n7718), .Z(n7402) );
    VMW_NOR2 U1822 ( .A(CallIn), .B(n1638), .Z(n7804) );
    VMW_OR3 U1589 ( .A(n7513), .B(n7522), .C(n7523), .Z(n7871) );
    VMW_AND2 U1615 ( .A(n7603), .B(ScanOut[5]), .Z(n7602) );
    VMW_OR4 U1729 ( .A(n7732), .B(n7669), .C(n7645), .D(n7635), .Z(n7765) );
    VMW_NAND2 U1785 ( .A(n7786), .B(n7708), .Z(n7429) );
    VMW_INV U1957 ( .A(PDiagIn[21]), .Z(n7440) );
    VMW_INV U2034 ( .A(n7718), .Z(n7789) );
    VMW_PULLDOWN U1341 ( .Z(n7896) );
    VMW_PULLDOWN U1383 ( .Z(n7938) );
    VMW_OR2 U1402 ( .A(n7409), .B(PDiagIn[47]), .Z(PDiagOut[46]) );
    VMW_NAND2 U1489 ( .A(n7438), .B(n7475), .Z(ColOut[23]) );
    VMW_OR2 U1492 ( .A(ColIn[20]), .B(n7442), .Z(ColOut[20]) );
    VMW_OR2 U1502 ( .A(ColIn[10]), .B(n7457), .Z(ColOut[10]) );
    VMW_OR2 U1525 ( .A(NDiagIn[57]), .B(n7399), .Z(NDiagOut[58]) );
    VMW_INV U1970 ( .A(ColIn[24]), .Z(n7474) );
    VMW_NAND2 U1519 ( .A(n7487), .B(n7494), .Z(\n1806[0] ) );
    VMW_AND3 U1629 ( .A(n7630), .B(n7631), .C(n7632), .Z(n7629) );
    VMW_AND3 U1632 ( .A(n7639), .B(n7640), .C(n7629), .Z(n7638) );
    VMW_FD \MyColumn_reg[2]  ( .D(n7873), .CP(Clk), .Q(ScanOut[2]) );
    VMW_INV U2008 ( .A(n7640), .Z(n7733) );
    VMW_INV U2013 ( .A(n7650), .Z(n7696) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_52 gt_104_53 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_35}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7927), .TC(
        n7927), .LT_LE(n1494) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_34 gt_104_48 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        Logic11, Logic11, Logic11}), .LEQ(n7910), .TC(n7910), .LT_LE(n1414) );
    VMW_OR4 U1592 ( .A(n7531), .B(NDiagIn[62]), .C(ColIn[62]), .D(PDiagIn[62]), 
        .Z(n7530) );
    VMW_AO22 U1732 ( .A(n7690), .B(n7687), .C(n7692), .D(n7768), .Z(n7767) );
    VMW_OR4 U1870 ( .A(n7820), .B(NDiagIn[45]), .C(ColIn[45]), .D(PDiagIn[45]), 
        .Z(n7821) );
    VMW_NAND2 U1425 ( .A(n7435), .B(n7436), .Z(PDiagOut[23]) );
    VMW_AND4 U1857 ( .A(n7816), .B(n7495), .C(n7471), .D(n7426), .Z(n7670) );
    VMW_OR2 U1550 ( .A(NDiagIn[32]), .B(n7424), .Z(NDiagOut[33]) );
    VMW_OR2 U1685 ( .A(n7706), .B(n7709), .Z(n7725) );
    VMW_MUX2I U1715 ( .A(ScanOut[6]), .B(ScanIn[6]), .S(ScanEnable), .Z(n7488)
         );
    VMW_OR2 U1839 ( .A(CallIn), .B(n1414), .Z(n7753) );
    VMW_OAI21 U1922 ( .A(n7618), .B(n7615), .C(n7622), .Z(n7553) );
    VMW_PULLDOWN U1346 ( .Z(n7901) );
    VMW_PULLDOWN U1361 ( .Z(n7916) );
    VMW_PULLDOWN U1366 ( .Z(n7921) );
    VMW_AND2 U1647 ( .A(n7673), .B(n7674), .Z(n7672) );
    VMW_AND2 U1660 ( .A(n7697), .B(n7698), .Z(n7591) );
    VMW_INV U2041 ( .A(n7725), .Z(n7800) );
    VMW_INV U2066 ( .A(n7627), .Z(n7749) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_33 gt_104_26 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , Logic11}), .LEQ(n7909), .TC(n7909), .LT_LE(
        n1062) );
    VMW_NOR2 U1895 ( .A(CallIn), .B(n678), .Z(n7835) );
    VMW_NOR4 U1905 ( .A(n7843), .B(NDiagIn[38]), .C(ColIn[38]), .D(PDiagIn[38]
        ), .Z(n7578) );
    VMW_OR2 U1570 ( .A(NDiagIn[12]), .B(n7454), .Z(NDiagOut[13]) );
    VMW_NAND2 U1577 ( .A(n7465), .B(n7508), .Z(NDiagOut[6]) );
    VMW_NAND2 U1819 ( .A(n7617), .B(n7621), .Z(n7803) );
    VMW_INV U1989 ( .A(NDiagIn[24]), .Z(n7498) );
    VMW_NAND2 U1640 ( .A(n7656), .B(n7657), .Z(n7655) );
    VMW_NOR2 U1892 ( .A(CallIn), .B(n710), .Z(n7834) );
    VMW_AO22 U1902 ( .A(n7567), .B(n7842), .C(n7778), .D(n7840), .Z(n7841) );
    VMW_OR2 U1667 ( .A(n7605), .B(n7706), .Z(n7707) );
    VMW_INV U2061 ( .A(n7831), .Z(n7665) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_32 gt_104_21 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_36}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7908), .TC(n7908), 
        .LT_LE(n982) );
    VMW_INV U2046 ( .A(n7748), .Z(n7863) );
    VMW_OR2 U1539 ( .A(NDiagIn[43]), .B(n7413), .Z(NDiagOut[44]) );
    VMW_OR2 U1557 ( .A(NDiagIn[25]), .B(n7434), .Z(NDiagOut[26]) );
    VMW_AOI211 U1609 ( .A(n7511), .B(n7510), .C(n7590), .D(n7513), .Z(n7589)
         );
    VMW_NAND4 U1925 ( .A(n7855), .B(n7507), .C(n7483), .D(n7462), .Z(n7627) );
    VMW_NAND2 U1799 ( .A(n7708), .B(n7793), .Z(n7450) );
    VMW_INV U2028 ( .A(n7707), .Z(n7796) );
    VMW_PULLDOWN U1333 ( .Z(n7888) );
    VMW_PULLUP U1384 ( .Z(Logic11) );
    VMW_NAND2 U1422 ( .A(n7431), .B(n7432), .Z(PDiagOut[26]) );
    VMW_OR2 U1682 ( .A(n7706), .B(n7717), .Z(n7722) );
    VMW_AND4 U1712 ( .A(n7755), .B(n7509), .C(n7485), .D(n7467), .Z(n7754) );
    VMW_OR2 U1850 ( .A(CallIn), .B(n1222), .Z(n7813) );
    VMW_OR2 U1405 ( .A(n7412), .B(PDiagIn[44]), .Z(PDiagOut[43]) );
    VMW_OR2 U1439 ( .A(n7457), .B(PDiagIn[10]), .Z(PDiagOut[9]) );
    VMW_NOR2 U1595 ( .A(n7540), .B(n7541), .Z(n7539) );
    VMW_AO22 U1735 ( .A(n7693), .B(n7666), .C(n7655), .D(n7658), .Z(n7559) );
    VMW_OR4 U1877 ( .A(n7823), .B(NDiagIn[52]), .C(ColIn[52]), .D(PDiagIn[52]), 
        .Z(n7657) );
    VMW_NAND2 U1495 ( .A(n7447), .B(n7478), .Z(ColOut[17]) );
    VMW_OR4 U1635 ( .A(n7526), .B(n7646), .C(n7647), .D(n7648), .Z(n7645) );
    VMW_AO22 U1699 ( .A(n7614), .B(n7740), .C(n7741), .D(n7552), .Z(n7588) );
    VMW_NOR4 U1709 ( .A(n7751), .B(NDiagIn[51]), .C(ColIn[51]), .D(PDiagIn[51]
        ), .Z(n7659) );
    VMW_INV U2014 ( .A(n7653), .Z(n7778) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_57 gt_104_54 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7932), .TC(n7932), 
        .LT_LE(n1510) );
    VMW_OR2 U1505 ( .A(ColIn[7]), .B(n7461), .Z(ColOut[7]) );
    VMW_OR2 U1522 ( .A(NDiagIn[60]), .B(n7396), .Z(NDiagOut[61]) );
    VMW_INV U1977 ( .A(ColIn[11]), .Z(n7481) );
    VMW_FD \MyColumn_reg[0]  ( .D(n7875), .CP(Clk), .Q(ScanOut[0]) );
    VMW_PULLDOWN U1368 ( .Z(n7923) );
    VMW_OR2 U1445 ( .A(n7466), .B(PDiagIn[4]), .Z(PDiagOut[3]) );
    VMW_OR2 U1457 ( .A(ColIn[55]), .B(n7401), .Z(ColOut[55]) );
    VMW_AND4 U1612 ( .A(n7511), .B(n7591), .C(n7596), .D(n7597), .Z(n7520) );
    VMW_NAND3 U1950 ( .A(n7867), .B(n7599), .C(n7598), .Z(n7601) );
    VMW_INV U2033 ( .A(n7716), .Z(n7788) );
    VMW_NOR2 U1782 ( .A(n7612), .B(n7725), .Z(n7424) );
    VMW_OR4 U1889 ( .A(n7832), .B(NDiagIn[57]), .C(ColIn[57]), .D(PDiagIn[57]), 
        .Z(n7533) );
    VMW_OAI22 U1919 ( .A(n7679), .B(n7852), .C(n7851), .D(n7670), .Z(n7549) );
    VMW_OR2 U1470 ( .A(ColIn[42]), .B(n7414), .Z(ColOut[42]) );
    VMW_AO22 U1740 ( .A(n7727), .B(ScanOut[2]), .C(n7726), .D(ScanIn[2]), .Z(
        n7519) );
    VMW_NOR2 U1767 ( .A(n7607), .B(n7608), .Z(n7409) );
    VMW_OR4 U1825 ( .A(n7805), .B(NDiagIn[2]), .C(ColIn[2]), .D(PDiagIn[2]), 
        .Z(n7599) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_11 gt_104_9 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_37}), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7887), .TC(n7887), .LT_LE(
        n790) );
    VMW_AND2 U1802 ( .A(n7794), .B(n7705), .Z(n7454) );
    VMW_INV U1992 ( .A(NDiagIn[19]), .Z(n7501) );
    VMW_OR2 U1837 ( .A(CallIn), .B(n1382), .Z(n7731) );
    VMW_OR2 U1462 ( .A(ColIn[50]), .B(n7406), .Z(ColOut[50]) );
    VMW_NOR2 U1752 ( .A(n7612), .B(n7712), .Z(n7394) );
    VMW_NOR2 U1775 ( .A(n7608), .B(n7710), .Z(n7417) );
    VMW_AND2 U1810 ( .A(n7798), .B(n7705), .Z(n7466) );
    VMW_INV U1980 ( .A(ColIn[5]), .Z(n7484) );
    VMW_OR2 U1649 ( .A(n7678), .B(n7578), .Z(n7677) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_26 gt_104_28 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7902), .TC(n7902), .LT_LE(
        n1094) );
    VMW_OR2 U1487 ( .A(ColIn[25]), .B(n7434), .Z(ColOut[25]) );
    VMW_NAND2 U1517 ( .A(n7487), .B(n7492), .Z(\n1806[2] ) );
    VMW_NAND2 U1579 ( .A(n7468), .B(n7509), .Z(NDiagOut[4]) );
    VMW_AND3 U1627 ( .A(n7598), .B(n7599), .C(n7624), .Z(n7623) );
    VMW_INV U2006 ( .A(n7617), .Z(n7652) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_36 gt_104_46 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7912), .TC(n7912), 
        .LT_LE(n1382) );
    VMW_INV U1965 ( .A(PDiagIn[5]), .Z(n7464) );
    VMW_OR4 U1942 ( .A(NDiagIn[63]), .B(n7570), .C(ColIn[63]), .D(PDiagIn[63]), 
        .Z(n7760) );
    VMW_PULLDOWN U1327 ( .Z(n7882) );
    VMW_PULLDOWN U1329 ( .Z(n7884) );
    VMW_PULLDOWN U1332 ( .Z(n7887) );
    VMW_PULLDOWN U1354 ( .Z(n7909) );
    VMW_PULLDOWN U1373 ( .Z(n7928) );
    VMW_OR2 U1396 ( .A(n7403), .B(PDiagIn[53]), .Z(PDiagOut[52]) );
    VMW_NAND2 U1430 ( .A(n7443), .B(n7444), .Z(PDiagOut[18]) );
    VMW_OR2 U1530 ( .A(NDiagIn[52]), .B(n7404), .Z(NDiagOut[53]) );
    VMW_AOI211 U1600 ( .A(n7557), .B(n7558), .C(n7559), .D(n7560), .Z(n7556)
         );
    VMW_NAND2 U1790 ( .A(n7705), .B(n7788), .Z(n7436) );
    VMW_INV U2021 ( .A(n7540), .Z(n7685) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_22 gt_104_61 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_38}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7898), 
        .TC(n7898), .LT_LE(n1622) );
    VMW_AND4 U1690 ( .A(n7731), .B(n7502), .C(n7478), .D(n7446), .Z(n7730) );
    VMW_OR4 U1700 ( .A(n7742), .B(NDiagIn[7]), .C(ColIn[7]), .D(PDiagIn[7]), 
        .Z(n7628) );
    VMW_NOR2 U1859 ( .A(CallIn), .B(n1062), .Z(n7817) );
    VMW_OR2 U1842 ( .A(CallIn), .B(n1318), .Z(n7634) );
    VMW_OR3 U1587 ( .A(n7513), .B(n7518), .C(n7519), .Z(n7873) );
    VMW_NOR2 U1865 ( .A(CallIn), .B(n998), .Z(n7686) );
    VMW_OR2 U1417 ( .A(n7424), .B(PDiagIn[32]), .Z(PDiagOut[31]) );
    VMW_AO22 U1727 ( .A(n7727), .B(ScanOut[5]), .C(n7726), .D(ScanIn[5]), .Z(
        n7525) );
    VMW_NOR2 U1880 ( .A(CallIn), .B(n806), .Z(n7825) );
    VMW_INV U1959 ( .A(PDiagIn[17]), .Z(n7446) );
    VMW_NOR2 U1910 ( .A(CallIn), .B(n1094), .Z(n7756) );
    VMW_OR2 U1545 ( .A(NDiagIn[37]), .B(n7419), .Z(NDiagOut[38]) );
    VMW_OR2 U1562 ( .A(NDiagIn[20]), .B(n7442), .Z(NDiagOut[21]) );
    VMW_NOR2 U1652 ( .A(n7683), .B(n7537), .Z(n7682) );
    VMW_FD \MyColumn_reg[4]  ( .D(n7871), .CP(Clk), .Q(ScanOut[4]) );
    VMW_OR2 U1675 ( .A(n7609), .B(n7711), .Z(n7715) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_13 gt_104_33 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_39}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7889), .TC(n7889), .LT_LE(
        n1174) );
    VMW_NAND4 U1937 ( .A(n7863), .B(n7862), .C(n7624), .D(n7627), .Z(n7600) );
    VMW_INV U2054 ( .A(n7815), .Z(n7646) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_53 gt_104_14 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7928), .TC(n7928), 
        .LT_LE(n870) );
    VMW_NAND2 U1438 ( .A(n7455), .B(n7456), .Z(PDiagOut[10]) );
    VMW_OR2 U1456 ( .A(ColIn[56]), .B(n7400), .Z(ColOut[56]) );
    VMW_OR2 U1479 ( .A(ColIn[33]), .B(n7423), .Z(ColOut[33]) );
    VMW_AO22 U1749 ( .A(n7599), .B(n7754), .C(n7748), .D(n7623), .Z(n7784) );
    VMW_NOR2 U1888 ( .A(CallIn), .B(n742), .Z(n7832) );
    VMW_AOI21 U1918 ( .A(n7849), .B(n7674), .C(n7671), .Z(n7851) );
    VMW_OR2 U1471 ( .A(ColIn[41]), .B(n7415), .Z(ColOut[41]) );
    VMW_AO22 U1741 ( .A(n7663), .B(n7666), .C(n7778), .D(n7659), .Z(n7777) );
    VMW_NOR2 U1766 ( .A(n7612), .B(n7722), .Z(n7408) );
    VMW_NOR2 U1824 ( .A(CallIn), .B(n1622), .Z(n7805) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_43 gt_104_8 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        Logic11, Logic11, Logic11}), .LEQ(n7919), .TC(n7919), .LT_LE(n774) );
    VMW_NAND2 U1803 ( .A(n7708), .B(n7795), .Z(n7456) );
    VMW_INV U1993 ( .A(NDiagIn[17]), .Z(n7502) );
    VMW_OR2 U1494 ( .A(ColIn[18]), .B(n7445), .Z(ColOut[18]) );
    VMW_OR2 U1504 ( .A(ColIn[8]), .B(n7460), .Z(ColOut[8]) );
    VMW_AND4 U1634 ( .A(n7644), .B(n7496), .C(n7472), .D(n7428), .Z(n7643) );
    VMW_OR2 U1698 ( .A(n7738), .B(n7701), .Z(n7560) );
    VMW_OR4 U1708 ( .A(n7750), .B(NDiagIn[50]), .C(ColIn[50]), .D(PDiagIn[50]), 
        .Z(n7569) );
    VMW_INV U2015 ( .A(n7655), .Z(n7662) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_54 gt_104_55 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , UNCONNECTED_40, 
        UNCONNECTED_41, UNCONNECTED_42}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n7929), .TC(n7929), .LT_LE(n1526) );
    VMW_INV U1976 ( .A(ColIn[13]), .Z(n7480) );
    VMW_OR2 U1523 ( .A(NDiagIn[59]), .B(n7397), .Z(NDiagOut[60]) );
    VMW_AOI211 U1608 ( .A(n7585), .B(n7586), .C(n7587), .D(n7588), .Z(n7584)
         );
    VMW_AND5 U1613 ( .A(n7598), .B(n7599), .C(n7600), .D(n7511), .E(n7591), 
        .Z(n7518) );
    VMW_AND2 U1783 ( .A(n7785), .B(n7708), .Z(n7425) );
    VMW_OAI211 U1951 ( .A(n7783), .B(n7784), .C(n7697), .D(n7511), .Z(n7868)
         );
    VMW_AND2 U1798 ( .A(n7792), .B(n7705), .Z(n7448) );
    VMW_INV U2029 ( .A(n7710), .Z(n7797) );
    VMW_INV U2032 ( .A(n7715), .Z(n7787) );
    VMW_PULLDOWN U1347 ( .Z(n7902) );
    VMW_PULLDOWN U1360 ( .Z(n7915) );
    VMW_PULLDOWN U1385 ( .Z(\NDiagOut[0] ) );
    VMW_OR2 U1404 ( .A(n7411), .B(PDiagIn[45]), .Z(PDiagOut[44]) );
    VMW_OR2 U1423 ( .A(n7433), .B(PDiagIn[26]), .Z(PDiagOut[25]) );
    VMW_OR2 U1538 ( .A(NDiagIn[44]), .B(n7412), .Z(NDiagOut[45]) );
    VMW_OR2 U1683 ( .A(n7605), .B(n7713), .Z(n7723) );
    VMW_OR4 U1713 ( .A(n7756), .B(NDiagIn[35]), .C(ColIn[35]), .D(PDiagIn[35]), 
        .Z(n7675) );
    VMW_NOR3 U1594 ( .A(n7536), .B(n7537), .C(n7538), .Z(n7535) );
    VMW_AND4 U1851 ( .A(n7813), .B(n7497), .C(n7473), .D(n7431), .Z(n7743) );
    VMW_AO22 U1734 ( .A(n7727), .B(ScanOut[3]), .C(n7726), .D(ScanIn[3]), .Z(
        n7521) );
    VMW_NOR2 U1876 ( .A(CallIn), .B(n822), .Z(n7823) );
    VMW_OR4 U1818 ( .A(PDiagIn[22]), .B(ColIn[22]), .C(NDiagIn[22]), .D(n7758), 
        .Z(n7637) );
    VMW_INV U1988 ( .A(NDiagIn[27]), .Z(n7497) );
    VMW_OR2 U1556 ( .A(NDiagIn[26]), .B(n7433), .Z(NDiagOut[27]) );
    VMW_NAND2 U1571 ( .A(n7456), .B(n7505), .Z(NDiagOut[12]) );
    VMW_NOR3 U1641 ( .A(n7659), .B(n7574), .C(n7653), .Z(n7658) );
    VMW_OR4 U1893 ( .A(n7834), .B(NDiagIn[59]), .C(ColIn[59]), .D(PDiagIn[59]), 
        .Z(n7664) );
    VMW_AO21 U1903 ( .A(n7739), .B(n7841), .C(n7738), .Z(n7544) );
    VMW_INV U2060 ( .A(n7829), .Z(n7668) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_1 gt_104_20 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7877), .TC(n7877), .LT_LE(
        n966) );
    VMW_OR2 U1666 ( .A(ScanOut[2]), .B(ScanOut[1]), .Z(n7706) );
    VMW_INV U2047 ( .A(n7615), .Z(n7620) );
    VMW_PULLDOWN U1349 ( .Z(n7904) );
    VMW_PULLDOWN U1355 ( .Z(n7910) );
    VMW_PULLDOWN U1372 ( .Z(n7927) );
    VMW_NAND2 U1563 ( .A(n7444), .B(n7501), .Z(NDiagOut[20]) );
    VMW_NOR4 U1881 ( .A(n7825), .B(NDiagIn[53]), .C(ColIn[53]), .D(PDiagIn[53]
        ), .Z(n7826) );
    VMW_NOR2 U1911 ( .A(CallIn), .B(n1158), .Z(n7846) );
    VMW_OR2 U1924 ( .A(CallIn), .B(n1558), .Z(n7855) );
    VMW_NOR2 U1653 ( .A(n7541), .B(n7685), .Z(n7684) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_27 gt_104_32 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        Logic11, Logic11, Logic11}), .LEQ(n7903), .TC(n7903), .LT_LE(n1158) );
    VMW_OR2 U1674 ( .A(n7711), .B(n7713), .Z(n7714) );
    VMW_INV U2055 ( .A(n7581), .Z(n7860) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_58 gt_104_15 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , UNCONNECTED_43, UNCONNECTED_44, 
        UNCONNECTED_45, UNCONNECTED_46}), .B({\NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), .LEQ(
        n7933), .TC(n7933), .LT_LE(n886) );
    VMW_AO21 U1936 ( .A(n7803), .B(n7861), .C(n7651), .Z(n7862) );
    VMW_PULLDOWN U1369 ( .Z(n7924) );
    VMW_OR2 U1397 ( .A(n7404), .B(PDiagIn[52]), .Z(PDiagOut[51]) );
    VMW_OR2 U1416 ( .A(n7423), .B(PDiagIn[33]), .Z(PDiagOut[32]) );
    VMW_OR2 U1431 ( .A(n7445), .B(PDiagIn[18]), .Z(PDiagOut[17]) );
    VMW_OR2 U1478 ( .A(ColIn[34]), .B(n7422), .Z(ColOut[34]) );
    VMW_OR2 U1544 ( .A(NDiagIn[38]), .B(n7418), .Z(NDiagOut[39]) );
    VMW_AO22 U1691 ( .A(n7631), .B(n7730), .C(n7629), .D(n7733), .Z(n7732) );
    VMW_OAI21 U1748 ( .A(n7551), .B(n7650), .C(n7698), .Z(n7783) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_44 gt_104_1 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_47}), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7920), .TC(n7920), .LT_LE(
        n662) );
    VMW_NOR2 U1701 ( .A(n7743), .B(n7647), .Z(n7580) );
    VMW_OR2 U1843 ( .A(CallIn), .B(n1286), .Z(n7747) );
    VMW_NOR4 U1864 ( .A(n7819), .B(NDiagIn[42]), .C(ColIn[42]), .D(PDiagIn[42]
        ), .Z(n7537) );
    VMW_NAND2 U1444 ( .A(n7464), .B(n7465), .Z(PDiagOut[4]) );
    VMW_OR2 U1486 ( .A(ColIn[26]), .B(n7433), .Z(ColOut[26]) );
    VMW_OR3 U1586 ( .A(n7513), .B(n7516), .C(n7517), .Z(n7874) );
    VMW_AND2 U1626 ( .A(n7622), .B(n7552), .Z(n7621) );
    VMW_AO22 U1726 ( .A(n7727), .B(ScanOut[6]), .C(n7726), .D(ScanIn[6]), .Z(
        n7590) );
    VMW_INV U1958 ( .A(PDiagIn[19]), .Z(n7443) );
    VMW_INV U1964 ( .A(PDiagIn[6]), .Z(n7462) );
    VMW_INV U2007 ( .A(n7763), .Z(n7631) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_21 gt_104_47 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , UNCONNECTED_48, UNCONNECTED_49, 
        UNCONNECTED_50, UNCONNECTED_51}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n7897), .TC(n7897), .LT_LE(n1398) );
    VMW_NAND2 U1516 ( .A(n7487), .B(n7491), .Z(\n1806[3] ) );
    VMW_OR2 U1531 ( .A(NDiagIn[51]), .B(n7405), .Z(NDiagOut[52]) );
    VMW_AO22 U1943 ( .A(n7821), .B(n7701), .C(n7571), .D(n7739), .Z(n7576) );
    VMW_AOI211 U1601 ( .A(n7562), .B(n7563), .C(n7564), .D(n7565), .Z(n7561)
         );
    VMW_NAND2 U1791 ( .A(n7789), .B(n7708), .Z(n7438) );
    VMW_NOR4 U1836 ( .A(n7808), .B(NDiagIn[16]), .C(ColIn[16]), .D(PDiagIn[16]
        ), .Z(n7763) );
    VMW_NOR2 U1858 ( .A(CallIn), .B(n1030), .Z(n7744) );
    VMW_INV U2020 ( .A(n7684), .Z(n7538) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_55 gt_104_60 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7930), .TC(
        n7930), .LT_LE(n1606) );
    VMW_OR2 U1463 ( .A(ColIn[49]), .B(n7407), .Z(ColOut[49]) );
    VMW_NOR2 U1753 ( .A(n7608), .B(n7714), .Z(n7395) );
    VMW_NOR2 U1774 ( .A(n7612), .B(n7707), .Z(n7416) );
    VMW_NAND2 U1811 ( .A(n7799), .B(n7708), .Z(n7468) );
    VMW_INV U1981 ( .A(ColIn[3]), .Z(n7485) );
    VMW_OR2 U1578 ( .A(NDiagIn[4]), .B(n7466), .Z(NDiagOut[5]) );
    VMW_AND4 U1648 ( .A(n7672), .B(n7593), .C(n7675), .D(n7676), .Z(n7563) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_60 gt_104_29 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_52}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n7935), 
        .TC(n7935), .LT_LE(n1110) );
    VMW_NAND2 U1443 ( .A(n7462), .B(n7463), .Z(PDiagOut[5]) );
    VMW_OR2 U1464 ( .A(ColIn[48]), .B(n7408), .Z(ColOut[48]) );
    VMW_NOR2 U1754 ( .A(n7612), .B(n7714), .Z(n7396) );
    VMW_NOR3 U1816 ( .A(n7730), .B(n7763), .C(n7632), .Z(n7764) );
    VMW_INV U1986 ( .A(NDiagIn[30]), .Z(n7495) );
    VMW_NOR2 U1773 ( .A(n7608), .B(n7707), .Z(n7415) );
    VMW_NAND2 U1558 ( .A(n7436), .B(n7498), .Z(NDiagOut[25]) );
    VMW_AND2 U1668 ( .A(n7704), .B(ScanOut[0]), .Z(n7708) );
    VMW_OR4 U1831 ( .A(n7807), .B(NDiagIn[12]), .C(ColIn[12]), .D(PDiagIn[12]), 
        .Z(n7759) );
    VMW_INV U2049 ( .A(n7754), .Z(n7598) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_10 gt_104 ( .A({\n1806[6] , 
        \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , \n1806[0] 
        }), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, Logic11, Logic11, 
        Logic11}), .LEQ(n7886), .TC(n7886), .LT_LE(n646) );
    VMW_NOR2 U1606 ( .A(n7580), .B(n7581), .Z(n7579) );
    VMW_AND2 U1796 ( .A(n7791), .B(n7705), .Z(n7445) );
    VMW_INV U2027 ( .A(n7589), .Z(n7869) );
    VMW_PULLDOWN U1335 ( .Z(n7890) );
    VMW_PULLDOWN U1340 ( .Z(n7895) );
    VMW_PULLDOWN U1352 ( .Z(n7907) );
    VMW_OR2 U1390 ( .A(n7397), .B(PDiagIn[59]), .Z(PDiagOut[58]) );
    VMW_OR2 U1481 ( .A(ColIn[31]), .B(n7425), .Z(ColOut[31]) );
    VMW_OR2 U1511 ( .A(ColIn[1]), .B(n7470), .Z(ColOut[1]) );
    VMW_OR2 U1536 ( .A(NDiagIn[46]), .B(n7410), .Z(NDiagOut[47]) );
    VMW_OAI211 U1944 ( .A(n7575), .B(n7779), .C(n7675), .D(n7676), .Z(n7864)
         );
    VMW_OR2 U1581 ( .A(NDiagIn[1]), .B(n7470), .Z(NDiagOut[2]) );
    VMW_OR2 U1621 ( .A(n7605), .B(n7609), .Z(n7611) );
    VMW_INV U1963 ( .A(PDiagIn[9]), .Z(n7458) );
    VMW_INV U2000 ( .A(NDiagIn[3]), .Z(n7509) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_7 gt_104_40 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        Logic11, Logic11, Logic11}), .LEQ(n7883), .TC(n7883), .LT_LE(n1286) );
    VMW_MUX2I U1721 ( .A(ScanOut[0]), .B(ScanIn[0]), .S(ScanEnable), .Z(n7494)
         );
    VMW_NOR2 U1878 ( .A(CallIn), .B(n790), .Z(n7824) );
    VMW_FD ReturnOut_reg ( .D(ReturnOut1761), .CP(Clk), .Q(ReturnOut) );
    VMW_OR2 U1411 ( .A(n7418), .B(PDiagIn[38]), .Z(PDiagOut[37]) );
    VMW_NAND2 U1436 ( .A(n7452), .B(n7453), .Z(PDiagOut[12]) );
    VMW_NOR2 U1863 ( .A(CallIn), .B(n982), .Z(n7819) );
    VMW_OR2 U1543 ( .A(NDiagIn[39]), .B(n7417), .Z(NDiagOut[40]) );
    VMW_NOR4 U1696 ( .A(n7737), .B(NDiagIn[46]), .C(ColIn[46]), .D(PDiagIn[46]
        ), .Z(n7701) );
    VMW_AND4 U1706 ( .A(n7747), .B(n7499), .C(n7475), .D(n7437), .Z(n7550) );
    VMW_OR2 U1844 ( .A(CallIn), .B(n1270), .Z(n7810) );
    VMW_INV U1978 ( .A(ColIn[9]), .Z(n7482) );
    VMW_PULLDOWN U1375 ( .Z(n7930) );
    VMW_OR4 U1654 ( .A(n7686), .B(NDiagIn[41]), .C(ColIn[41]), .D(PDiagIn[41]), 
        .Z(n7540) );
    VMW_NAND2 U1673 ( .A(ScanOut[2]), .B(n7610), .Z(n7713) );
    VMW_NOR4 U1931 ( .A(n7858), .B(NDiagIn[8]), .C(ColIn[8]), .D(PDiagIn[8]), 
        .Z(n7651) );
    VMW_INV U2052 ( .A(n7546), .Z(n7648) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_45 gt_104_12 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7921), .TC(n7921), .LT_LE(
        n838) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_61 gt_104_35 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_53, UNCONNECTED_54}), .B({\NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n7936), 
        .TC(n7936), .LT_LE(n1206) );
    VMW_OR2 U1458 ( .A(ColIn[54]), .B(n7402), .Z(ColOut[54]) );
    VMW_OR2 U1564 ( .A(NDiagIn[18]), .B(n7445), .Z(NDiagOut[19]) );
    VMW_NOR2 U1886 ( .A(CallIn), .B(n726), .Z(n7830) );
    VMW_OR4 U1916 ( .A(n7848), .B(NDiagIn[32]), .C(ColIn[32]), .D(PDiagIn[32]), 
        .Z(n7674) );
    VMW_NOR2 U1768 ( .A(n7607), .B(n7612), .Z(n7410) );
    VMW_NOR2 U1838 ( .A(CallIn), .B(n1366), .Z(n7728) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_41 gt_104_6 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11}), .LEQ(n7917), .TC(n7917), 
        .LT_LE(n742) );
    VMW_NOR2 U1923 ( .A(CallIn), .B(n1542), .Z(n7742) );
    VMW_PULLDOWN U1367 ( .Z(n7922) );
    VMW_OR2 U1551 ( .A(NDiagIn[31]), .B(n7425), .Z(NDiagOut[32]) );
    VMW_NAND2 U1576 ( .A(n7463), .B(n7507), .Z(NDiagOut[7]) );
    VMW_OR2 U1646 ( .A(n7670), .B(n7671), .Z(n7669) );
    VMW_OR2 U1661 ( .A(n7700), .B(n7701), .Z(n7699) );
    VMW_INV U2040 ( .A(n7724), .Z(n7799) );
    VMW_NOR2 U1894 ( .A(CallIn), .B(n662), .Z(n7531) );
    VMW_NOR2 U1904 ( .A(CallIn), .B(n1046), .Z(n7843) );
    VMW_INV U2067 ( .A(n7868), .Z(n7514) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_46 gt_104_27 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , 
        UNCONNECTED_55, UNCONNECTED_56}), .B({\NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] }), 
        .LEQ(n7922), .TC(n7922), .LT_LE(n1078) );
    VMW_PULLDOWN U1382 ( .Z(n7937) );
    VMW_NAND2 U1488 ( .A(n7436), .B(n7474), .Z(ColOut[24]) );
    VMW_NAND4 U1628 ( .A(n7623), .B(n7626), .C(n7627), .D(n7628), .Z(n7625) );
    VMW_INV U2009 ( .A(n7635), .Z(n7642) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_2 gt_104_49 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        UNCONNECTED_57}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11, Logic11, \NDiagOut[0] }), .LEQ(n7878), .TC(n7878), 
        .LT_LE(n1430) );
    VMW_NAND2 U1518 ( .A(n7487), .B(n7493), .Z(\n1806[1] ) );
    VMW_AOI211 U1733 ( .A(n7649), .B(n7770), .C(n7588), .D(n7651), .Z(n7769)
         );
    VMW_NOR2 U1871 ( .A(CallIn), .B(n886), .Z(n7822) );
    VMW_OR2 U1399 ( .A(n7406), .B(PDiagIn[50]), .Z(PDiagOut[49]) );
    VMW_OR2 U1403 ( .A(n7410), .B(PDiagIn[46]), .Z(PDiagOut[45]) );
    VMW_OR2 U1424 ( .A(n7434), .B(PDiagIn[25]), .Z(PDiagOut[24]) );
    VMW_AND2 U1593 ( .A(n7533), .B(n7534), .Z(n7532) );
    VMW_OR2 U1856 ( .A(CallIn), .B(n1174), .Z(n7816) );
    VMW_OR2 U1684 ( .A(n7609), .B(n7709), .Z(n7724) );
    VMW_NOR4 U1714 ( .A(n7757), .B(NDiagIn[49]), .C(ColIn[49]), .D(PDiagIn[49]
        ), .Z(n7567) );
    VMW_OR2 U1418 ( .A(n7425), .B(PDiagIn[31]), .Z(PDiagOut[30]) );
    VMW_OR2 U1524 ( .A(NDiagIn[58]), .B(n7398), .Z(NDiagOut[59]) );
    VMW_OR3 U1588 ( .A(n7513), .B(n7520), .C(n7521), .Z(n7872) );
    VMW_AND3 U1614 ( .A(n7591), .B(n7601), .C(n7511), .Z(n7516) );
    VMW_OR4 U1728 ( .A(n7762), .B(n7550), .C(n7763), .D(n7764), .Z(n7761) );
    VMW_INV U2035 ( .A(n7719), .Z(n7790) );
    VMW_NAND2 U1784 ( .A(n7705), .B(n7785), .Z(n7427) );
    VMW_INV U1956 ( .A(PDiagIn[23]), .Z(n7437) );
    VMW_OR2 U1451 ( .A(ColIn[61]), .B(n7395), .Z(ColOut[61]) );
    VMW_OR2 U1476 ( .A(ColIn[36]), .B(n7420), .Z(ColOut[36]) );
    VMW_NAND2 U1493 ( .A(n7444), .B(n7477), .Z(ColOut[19]) );
    VMW_INV U1971 ( .A(ColIn[23]), .Z(n7475) );
    VMW_NAND2 U1503 ( .A(n7459), .B(n7482), .Z(ColOut[9]) );
    VMW_NAND2 U1633 ( .A(n7638), .B(n7642), .Z(n7641) );
    VMW_INV U2012 ( .A(n7645), .Z(n7548) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1_DW01_cmp2_7_37 gt_104_52 ( .A({
        \n1806[6] , \n1806[5] , \n1806[4] , \n1806[3] , \n1806[2] , \n1806[1] , 
        \n1806[0] }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, Logic11}), .LEQ(n7913), .TC(n7913), .LT_LE(
        n1478) );
    VMW_AND2 U1804 ( .A(n7705), .B(n7795), .Z(n7457) );
    VMW_AO21 U1938 ( .A(n7667), .B(n7557), .C(n7560), .Z(n7768) );
    VMW_INV U1994 ( .A(NDiagIn[15]), .Z(n7503) );
    VMW_AO22 U1746 ( .A(n7727), .B(ScanOut[1]), .C(n7726), .D(ScanIn[1]), .Z(
        n7517) );
    VMW_NOR2 U1761 ( .A(n7608), .B(n7719), .Z(n7403) );
    VMW_OR4 U1823 ( .A(n7804), .B(NDiagIn[1]), .C(ColIn[1]), .D(PDiagIn[1]), 
        .Z(n7698) );
endmodule


module NQueens_Control_IDWIDTH7_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, CallIn, ReturnIn, 
    CallOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [6:0] Id;
input  [6:0] ScanIn;
output [6:0] ScanOut;
input  [6:0] ScanId;
input  Clk, Reset, RD, WR, CallIn, ReturnIn;
output ScanEnable, CallOut;
    wire n421, n433, n387, n406, n395, n414, n446, n428, n441, n389, n408, 
        n413, n434, n392, n426, n401, n448, n453, n435, n393, n412, 
        \status[4] , n440, \ScanReg[2] , n388, n409, n449, n452, \status[0] , 
        n427, n400, \ScanReg[6] , n420, \ScanReg[4] , n386, n407, \status[2] , 
        n429, n447, \ScanReg[0] , n432, n415, n394, \status[6] , n439, 
        \ScanReg[1] , n422, n405, \status[7] , \ScanReg[5] , n417, n430, n396, 
        n445, \status[3] , \status[1] , n442, n437, n391, n402, n425, n410, 
        n450, \status[5] , n390, n398, \ScanReg[3] , n419, n436, n411, n443, 
        n418, n451, n399, n424, n403, n423, n385, n404, Logic01, n438, n444, 
        n416, n397, n431;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    assign ScanOut[6] = Logic01;
    assign ScanOut[5] = Logic01;
    assign ScanOut[4] = Logic01;
    assign ScanOut[3] = Logic01;
    assign ScanOut[2] = Logic01;
    assign ScanOut[1] = Logic01;
    assign ScanOut[0] = Logic01;
    VMW_PULLDOWN U96 ( .Z(n438) );
    VMW_AND4 U113 ( .A(n397), .B(n398), .C(n399), .D(n400), .Z(n387) );
    VMW_XNOR2 U134 ( .A(Addr[0]), .B(Id[0]), .Z(n411) );
    VMW_AND2 U108 ( .A(n387), .B(\status[7] ), .Z(n439) );
    VMW_INV U141 ( .A(n387), .Z(n385) );
    VMW_BUFIZ U166 ( .A(n431), .E(n418), .Z(\arr[30] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_PULLDOWN U83 ( .Z(n422) );
    VMW_PULLDOWN U84 ( .Z(n423) );
    VMW_INV U148 ( .A(n406), .Z(n389) );
    VMW_BUFIZ U153 ( .A(n417), .E(n418), .Z(\arr[9] ) );
    VMW_BUFIZ U174 ( .A(n439), .E(n418), .Z(\arr[7] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U101 ( .Z(Logic01) );
    VMW_AND2 U106 ( .A(\status[6] ), .B(n386), .Z(n447) );
    VMW_AO22 U121 ( .A(\status[4] ), .B(n387), .C(\ScanReg[4] ), .D(n385), .Z(
        n419) );
    VMW_AND4 U126 ( .A(n408), .B(n409), .C(n410), .D(n411), .Z(n400) );
    VMW_BUFIZ U168 ( .A(n433), .E(n418), .Z(\arr[20] ) );
    VMW_PULLDOWN U91 ( .Z(n432) );
    VMW_PULLDOWN U98 ( .Z(n442) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_NAND2 U128 ( .A(n387), .B(WR), .Z(n391) );
    VMW_BUFIZ U154 ( .A(n419), .E(n418), .Z(\arr[4] ) );
    VMW_BUFIZ U173 ( .A(n438), .E(n418), .Z(\arr[15] ) );
    VMW_INV U146 ( .A(n386), .Z(n393) );
    VMW_BUFIZ U161 ( .A(n426), .E(n418), .Z(\arr[31] ) );
    VMW_PULLDOWN U99 ( .Z(n443) );
    VMW_NOR5 U114 ( .A(\status[6] ), .B(\status[7] ), .C(\status[5] ), .D(
        \status[3] ), .E(\status[4] ), .Z(n401) );
    VMW_AO21 U133 ( .A(n389), .B(n391), .C(Reset), .Z(n396) );
    VMW_FD \status_reg[7]  ( .D(n446), .CP(Clk), .Q(\status[7] ) );
    VMW_BUFIZ U155 ( .A(n420), .E(n418), .Z(\arr[27] ) );
    VMW_BUFIZ U172 ( .A(n437), .E(n418), .Z(\arr[26] ) );
    VMW_PULLDOWN U82 ( .Z(n421) );
    VMW_BUFIZ U169 ( .A(n434), .E(n418), .Z(\arr[24] ) );
    VMW_PULLDOWN U85 ( .Z(n424) );
    VMW_PULLDOWN U90 ( .Z(n431) );
    VMW_AND2 U107 ( .A(\status[7] ), .B(n386), .Z(n446) );
    VMW_AO22 U120 ( .A(\status[5] ), .B(n387), .C(\ScanReg[5] ), .D(n385), .Z(
        n440) );
    VMW_AND4 U115 ( .A(\status[1] ), .B(n401), .C(n395), .D(n403), .Z(n402) );
    VMW_NAND3 U132 ( .A(n390), .B(n391), .C(n412), .Z(n394) );
    VMW_FD \status_reg[3]  ( .D(n450), .CP(Clk), .Q(\status[3] ) );
    VMW_PULLDOWN U97 ( .Z(n441) );
    VMW_OR2 U109 ( .A(n387), .B(RD), .Z(n418) );
    VMW_AND2 U129 ( .A(n402), .B(CallIn), .Z(n406) );
    VMW_INV U147 ( .A(n405), .Z(n412) );
    VMW_BUFIZ U160 ( .A(n425), .E(n418), .Z(\arr[6] ) );
    VMW_XNOR2 U140 ( .A(Addr[3]), .B(Id[3]), .Z(n399) );
    VMW_BUFIZ U167 ( .A(n432), .E(n418), .Z(\arr[29] ) );
    VMW_PULLDOWN U100 ( .Z(n445) );
    VMW_OAI21 U112 ( .A(n395), .B(n393), .C(n396), .Z(n453) );
    VMW_XNOR2 U135 ( .A(Addr[1]), .B(Id[1]), .Z(n410) );
    VMW_FD \status_reg[1]  ( .D(n452), .CP(Clk), .Q(\status[1] ) );
    VMW_AND2 U127 ( .A(n403), .B(n404), .Z(CallOut) );
    VMW_BUFIZ U149 ( .A(n413), .E(n418), .Z(\arr[19] ) );
    VMW_BUFIZ U152 ( .A(n416), .E(n418), .Z(\arr[10] ) );
    VMW_BUFIZ U175 ( .A(n440), .E(n418), .Z(\arr[5] ) );
    VMW_FD \status_reg[5]  ( .D(n448), .CP(Clk), .Q(\status[5] ) );
    VMW_PULLDOWN U77 ( .Z(n413) );
    VMW_PULLDOWN U79 ( .Z(n416) );
    VMW_PULLDOWN U95 ( .Z(n437) );
    VMW_AND4 U110 ( .A(n388), .B(n389), .C(n390), .D(n391), .Z(n451) );
    VMW_XNOR2 U137 ( .A(Addr[6]), .B(Id[6]), .Z(n408) );
    VMW_BUFIZ U159 ( .A(n424), .E(n418), .Z(\arr[12] ) );
    VMW_AO22 U119 ( .A(\status[6] ), .B(n387), .C(\ScanReg[6] ), .D(n385), .Z(
        n425) );
    VMW_INV U142 ( .A(\status[2] ), .Z(n403) );
    VMW_FD \status_reg[4]  ( .D(n449), .CP(Clk), .Q(\status[4] ) );
    VMW_BUFIZ U165 ( .A(n430), .E(n418), .Z(\arr[13] ) );
    VMW_BUFIZ U180 ( .A(n445), .E(n418), .Z(\arr[8] ) );
    VMW_PULLDOWN U80 ( .Z(n417) );
    VMW_PULLDOWN U87 ( .Z(n427) );
    VMW_BUFIZ U150 ( .A(n414), .E(n418), .Z(\arr[0] ) );
    VMW_BUFIZ U177 ( .A(n442), .E(n418), .Z(\arr[18] ) );
    VMW_AND2 U102 ( .A(RD), .B(n385), .Z(ScanEnable) );
    VMW_AO22 U125 ( .A(\status[0] ), .B(n387), .C(\ScanReg[0] ), .D(n385), .Z(
        n414) );
    VMW_AND2 U105 ( .A(\status[5] ), .B(n386), .Z(n448) );
    VMW_FD \status_reg[0]  ( .D(n453), .CP(Clk), .Q(\status[0] ) );
    VMW_AO22 U122 ( .A(\status[3] ), .B(n387), .C(\ScanReg[3] ), .D(n385), .Z(
        n436) );
    VMW_FD \status_reg[2]  ( .D(n451), .CP(Clk), .Q(\status[2] ) );
    VMW_PULLDOWN U89 ( .Z(n430) );
    VMW_XNOR2 U139 ( .A(Addr[5]), .B(Id[5]), .Z(n397) );
    VMW_BUFIZ U157 ( .A(n422), .E(n418), .Z(\arr[25] ) );
    VMW_BUFIZ U170 ( .A(n435), .E(n418), .Z(\arr[17] ) );
    VMW_PULLDOWN U92 ( .Z(n433) );
    VMW_INV U145 ( .A(Reset), .Z(n390) );
    VMW_BUFIZ U162 ( .A(n427), .E(n418), .Z(\arr[21] ) );
    VMW_FD \status_reg[6]  ( .D(n447), .CP(Clk), .Q(\status[6] ) );
    VMW_BUFIZ U179 ( .A(n444), .E(n418), .Z(\arr[1] ) );
    VMW_NOR2 U117 ( .A(n406), .B(CallOut), .Z(n405) );
    VMW_PULLDOWN U78 ( .Z(n415) );
    VMW_PULLDOWN U81 ( .Z(n420) );
    VMW_NAND2 U130 ( .A(ReturnIn), .B(n402), .Z(n407) );
    VMW_XNOR2 U138 ( .A(Addr[2]), .B(Id[2]), .Z(n398) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_BUFIZ U156 ( .A(n421), .E(n418), .Z(\arr[14] ) );
    VMW_BUFIZ U171 ( .A(n436), .E(n418), .Z(\arr[3] ) );
    VMW_PULLDOWN U86 ( .Z(n426) );
    VMW_PULLDOWN U88 ( .Z(n428) );
    VMW_PULLDOWN U93 ( .Z(n434) );
    VMW_AND2 U104 ( .A(\status[4] ), .B(n386), .Z(n449) );
    VMW_AND3 U116 ( .A(n401), .B(n392), .C(\status[0] ), .Z(n404) );
    VMW_AO22 U123 ( .A(\status[2] ), .B(n387), .C(\ScanReg[2] ), .D(n385), .Z(
        n429) );
    VMW_OAI21 U131 ( .A(n404), .B(n386), .C(n403), .Z(n388) );
    VMW_BUFIZ U178 ( .A(n443), .E(n418), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_PULLDOWN U94 ( .Z(n435) );
    VMW_INV U143 ( .A(\status[1] ), .Z(n392) );
    VMW_INV U144 ( .A(\status[0] ), .Z(n395) );
    VMW_BUFIZ U163 ( .A(n428), .E(n418), .Z(\arr[28] ) );
    VMW_BUFIZ U158 ( .A(n423), .E(n418), .Z(\arr[16] ) );
    VMW_BUFIZ U164 ( .A(n429), .E(n418), .Z(\arr[2] ) );
    VMW_AND2 U103 ( .A(\status[3] ), .B(n386), .Z(n450) );
    VMW_OAI21 U111 ( .A(n392), .B(n393), .C(n394), .Z(n452) );
    VMW_XNOR2 U136 ( .A(Addr[4]), .B(Id[4]), .Z(n409) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AO22 U124 ( .A(\status[1] ), .B(n387), .C(\ScanReg[1] ), .D(n385), .Z(
        n444) );
    VMW_AND4 U118 ( .A(n405), .B(n407), .C(n390), .D(n391), .Z(n386) );
    VMW_BUFIZ U151 ( .A(n415), .E(n418), .Z(\arr[23] ) );
    VMW_BUFIZ U176 ( .A(n441), .E(n418), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wColumn_13[27] , \wNDiag_29[0] , \wColumn_30[16] , \wColumn_45[26] , 
        \wColumn_33[3] , \wColumn_50[12] , \wPDiag_61[2] , \wColumn_6[31] , 
        \wPDiag_6[53] , \wPDiag_12[18] , \wColumn_25[22] , \wNDiag_25[57] , 
        \wNDiag_38[35] , \wPDiag_51[34] , \wNDiag_58[31] , \wNDiag_58[28] , 
        \wPDiag_59[62] , \wNDiag_30[63] , \wPDiag_44[19] , \wNDiag_45[53] , 
        \wPDiag_31[30] , \wPDiag_31[29] , \wNDiag_13[52] , \wColumn_30[0] , 
        \wColumn_38[59] , \wColumn_38[40] , \wColumn_58[44] , \wPDiag_59[51] , 
        \wPDiag_62[1] , \wColumn_6[28] , \wPDiag_59[48] , \wPDiag_8[4] , 
        \wPDiag_18[9] , \wPDiag_39[55] , \wColumn_25[11] , \wColumn_50[38] , 
        \wColumn_50[21] , \wScan_0[6] , \wColumn_1[43] , \wPDiag_1[38] , 
        \wNDiag_3[60] , \wNDiag_3[53] , \wPDiag_5[23] , \wPDiag_6[60] , 
        \wNDiag_8[46] , \wColumn_30[25] , \wColumn_13[14] , \wColumn_45[15] , 
        \wCall_63[0] , \wColumn_57[7] , \wNDiag_10[22] , \wPDiag_12[32] , 
        \wColumn_54[4] , \wNDiag_13[61] , \wNDiag_30[50] , \wNDiag_45[60] , 
        \wNDiag_53[8] , \wPDiag_24[37] , \wNDiag_30[49] , \wPDiag_44[33] , 
        \wNDiag_26[27] , \wNDiag_50[54] , \wNDiag_53[17] , \wPDiag_52[44] , 
        \wPDiag_32[59] , \wPDiag_32[40] , \wNDiag_33[13] , \wNDiag_46[23] , 
        \wNDiag_32[1] , \wColumn_18[18] , \wColumn_10[57] , \wColumn_28[2] , 
        \wColumn_18[32] , \wScan_19[0] , \wPDiag_19[27] , \wColumn_26[52] , 
        \wNDiag_31[2] , \wColumn_46[56] , \wColumn_53[62] , \wColumn_5[58] , 
        \wPDiag_5[10] , \wNDiag_56[5] , \wNDiag_10[11] , \wNDiag_33[39] , 
        \wPDiag_11[42] , \wNDiag_33[20] , \wPDiag_47[43] , \wNDiag_26[14] , 
        \wNDiag_46[10] , \wPDiag_27[47] , \wColumn_51[9] , \wNDiag_53[24] , 
        \wNDiag_48[9] , \wColumn_5[41] , \wNDiag_7[51] , \wNDiag_7[48] , 
        \wColumn_14[55] , \wNDiag_18[47] , \wPDiag_19[14] , \wColumn_22[50] , 
        \wColumn_26[61] , \wNDiag_55[6] , \wColumn_33[55] , \wReturn_39[0] , 
        \wColumn_53[51] , \wColumn_53[48] , \wPDiag_39[2] , \wColumn_57[60] , 
        \wScan_59[2] , \wColumn_22[49] , \wColumn_42[54] , \wPDiag_1[21] , 
        \wColumn_9[26] , \wNDiag_14[39] , \wNDiag_14[20] , \wNDiag_42[38] , 
        \wNDiag_61[10] , \wPDiag_36[42] , \wNDiag_42[21] , \wPDiag_60[43] , 
        \wNDiag_22[25] , \wNDiag_37[11] , \wNDiag_57[15] , \wPDiag_56[46] , 
        \wPDiag_9[44] , \wNDiag_15[4] , \wColumn_37[57] , \wColumn_61[56] , 
        \wColumn_22[63] , \wColumn_57[53] , \wColumn_12[8] , \wPDiag_40[9] , 
        \wPDiag_1[12] , \wColumn_3[4] , \wColumn_9[15] , \wNDiag_22[16] , 
        \wPDiag_23[45] , \wNDiag_57[26] , \wNDiag_14[13] , \wPDiag_15[59] , 
        \wPDiag_15[40] , \wNDiag_37[22] , \wPDiag_43[41] , \wNDiag_61[23] , 
        \wNDiag_42[12] , \wPDiag_43[58] , \wColumn_2[33] , \wColumn_2[19] , 
        \wPDiag_2[51] , \wNDiag_4[38] , \wNDiag_4[21] , \wNDiag_7[62] , 
        \wNDiag_16[7] , \wPDiag_22[3] , \wPDiag_2[48] , \wNDiag_17[50] , 
        \wNDiag_17[49] , \wNDiag_34[61] , \wNDiag_41[51] , \wPDiag_63[33] , 
        \wPDiag_35[32] , \wNDiag_41[48] , \wNDiag_62[60] , \wNDiag_21[55] , 
        \wScan_42[3] , \wPDiag_55[36] , \wPDiag_28[50] , \wPDiag_28[49] , 
        \wPDiag_2[62] , \wColumn_6[9] , \wColumn_17[25] , \wColumn_21[39] , 
        \wScan_41[0] , \wPDiag_48[54] , \wColumn_21[20] , \wPDiag_21[0] , 
        \wColumn_54[10] , \wColumn_34[14] , \wColumn_41[24] , \wColumn_62[15] , 
        \wPDiag_20[35] , \wPDiag_16[30] , \wNDiag_54[56] , \wPDiag_16[29] , 
        \wNDiag_17[63] , \wNDiag_34[52] , \wPDiag_35[18] , \wPDiag_40[28] , 
        \wNDiag_41[62] , \wPDiag_40[31] , \wNDiag_62[53] , \wPDiag_63[19] , 
        \wNDiag_4[12] , \wColumn_14[6] , \wPDiag_46[7] , \wColumn_29[45] , 
        \wNDiag_9[4] , \wColumn_17[16] , \wColumn_34[27] , \wColumn_49[58] , 
        \wColumn_49[41] , \wColumn_41[17] , \wColumn_17[5] , \wPDiag_45[4] , 
        \wColumn_21[13] , \wColumn_62[26] , \wNDiag_49[34] , \wColumn_54[23] , 
        \wReturn_61[0] , \wNDiag_10[9] , \wScan_3[5] , \wColumn_3[39] , 
        \wColumn_3[20] , \wNDiag_6[42] , \wColumn_8[35] , \wPDiag_8[57] , 
        \wPDiag_14[53] , \wPDiag_22[56] , \wScan_25[4] , \wPDiag_28[63] , 
        \wNDiag_29[29] , \wNDiag_29[30] , \wScan_33[0] , \wNDiag_56[35] , 
        \wNDiag_36[28] , \wPDiag_53[0] , \wPDiag_37[62] , \wPDiag_42[52] , 
        \wNDiag_43[18] , \wNDiag_60[30] , \wNDiag_15[19] , \wNDiag_18[1] , 
        \wNDiag_36[31] , \wPDiag_50[3] , \wNDiag_60[29] , \wPDiag_61[63] , 
        \wColumn_36[44] , \wColumn_60[45] , \wColumn_56[40] , \wReturn_13[0] , 
        \wPDiag_14[60] , \wNDiag_15[33] , \wScan_30[3] , \wColumn_56[59] , 
        \wPDiag_37[51] , \wPDiag_42[61] , \wPDiag_61[49] , \wPDiag_37[4] , 
        \wPDiag_37[48] , \wNDiag_43[32] , \wPDiag_61[50] , \wNDiag_23[36] , 
        \wPDiag_57[55] , \wColumn_15[46] , \wColumn_23[43] , \wScan_57[4] , 
        \wNDiag_62[9] , \wPDiag_29[8] , \wPDiag_34[7] , \wColumn_43[47] , 
        \wPDiag_48[1] , \wNDiag_48[27] , \wColumn_3[13] , \wNDiag_4[1] , 
        \wNDiag_28[23] , \wColumn_35[34] , \wNDiag_5[18] , \wNDiag_7[2] , 
        \wColumn_20[19] , \wColumn_63[35] , \wScan_28[1] , \wColumn_55[29] , 
        \wColumn_55[30] , \wColumn_28[56] , \wColumn_48[52] , \wColumn_16[36] , 
        \wPDiag_17[23] , \wColumn_19[3] , \wPDiag_21[26] , \wPDiag_54[16] , 
        \wNDiag_55[45] , \wNDiag_35[41] , \wColumn_20[33] , \wPDiag_34[12] , 
        \wNDiag_35[58] , \wPDiag_62[13] , \wNDiag_63[59] , \wPDiag_41[22] , 
        \wNDiag_63[40] , \wColumn_40[37] , \wPDiag_29[43] , \wPDiag_3[42] , 
        \wNDiag_5[32] , \wNDiag_16[43] , \wPDiag_17[10] , \wNDiag_28[10] , 
        \wNDiag_40[42] , \wNDiag_48[14] , \wCall_49[0] , \wPDiag_49[47] , 
        \wPDiag_62[20] , \wPDiag_34[38] , \wPDiag_41[11] , \wPDiag_62[39] , 
        \wNDiag_20[46] , \wPDiag_21[15] , \wPDiag_34[21] , \wPDiag_54[25] , 
        \wPDiag_32[9] , \wColumn_48[61] , \wColumn_60[8] , \wPDiag_6[2] , 
        \wNDiag_31[43] , \wNDiag_43[2] , \wPDiag_13[38] , \wPDiag_13[21] , 
        \wPDiag_30[10] , \wPDiag_45[39] , \wPDiag_25[24] , \wPDiag_45[20] , 
        \wColumn_39[60] , \wPDiag_50[14] , \wNDiag_51[47] , \wColumn_59[1] , 
        \wNDiag_1[30] , \wPDiag_5[1] , \wColumn_7[22] , \wNDiag_9[55] , 
        \wColumn_31[36] , \wColumn_51[32] , \wPDiag_58[42] , \wNDiag_59[11] , 
        \wPDiag_7[59] , \wPDiag_7[40] , \wPDiag_38[46] , \wNDiag_39[15] , 
        \wNDiag_40[1] , \wColumn_39[53] , \wColumn_59[57] , \wNDiag_1[29] , 
        \wColumn_4[61] , \wColumn_4[52] , \wColumn_7[11] , \wNDiag_12[58] , 
        \wNDiag_24[44] , \wPDiag_25[17] , \wPDiag_50[27] , \wNDiag_27[6] , 
        \wNDiag_44[40] , \wNDiag_12[41] , \wPDiag_13[12] , \wNDiag_44[59] , 
        \wPDiag_45[13] , \wNDiag_24[5] , \wPDiag_30[23] , \wNDiag_39[26] , 
        \wColumn_12[34] , \wColumn_44[35] , \wNDiag_59[22] , \wColumn_23[9] , 
        \wColumn_24[31] , \wColumn_24[28] , \wColumn_51[18] , \wColumn_32[46] , 
        \wColumn_52[42] , \wNDiag_58[3] , \wPDiag_10[51] , \wPDiag_10[48] , 
        \wPDiag_10[1] , \wNDiag_19[54] , \wColumn_42[0] , \wPDiag_33[60] , 
        \wPDiag_46[50] , \wPDiag_13[2] , \wPDiag_26[54] , \wNDiag_32[33] , 
        \wPDiag_46[49] , \wNDiag_52[37] , \wPDiag_18[34] , \wColumn_19[38] , 
        \wColumn_19[21] , \wColumn_41[3] , \wColumn_26[4] , \wColumn_11[44] , 
        \wScan_14[5] , \wNDiag_21[8] , \wNDiag_1[39] , \wNDiag_1[5] , 
        \wNDiag_2[59] , \wPDiag_4[30] , \wPDiag_4[29] , \wColumn_27[58] , 
        \wColumn_27[41] , \wColumn_47[45] , \wScan_17[6] , \wColumn_19[12] , 
        \wNDiag_2[40] , \wColumn_38[8] , \wNDiag_2[6] , \wColumn_3[30] , 
        \wColumn_3[29] , \wPDiag_3[52] , \wPDiag_10[62] , \wCall_11[0] , 
        \wNDiag_27[34] , \wPDiag_53[57] , \wNDiag_11[31] , \wColumn_25[7] , 
        \wPDiag_33[53] , \wPDiag_46[63] , \wNDiag_47[29] , \wNDiag_32[19] , 
        \wNDiag_11[28] , \wNDiag_47[30] , \wColumn_16[26] , \wColumn_63[16] , 
        \wNDiag_16[53] , \wColumn_20[23] , \wColumn_35[17] , \wColumn_40[27] , 
        \wColumn_55[13] , \wNDiag_20[56] , \wNDiag_28[19] , \wPDiag_31[3] , 
        \wColumn_63[2] , \wPDiag_49[57] , \wScan_51[3] , \wPDiag_29[53] , 
        \wPDiag_34[31] , \wScan_52[0] , \wPDiag_54[35] , \wPDiag_62[29] , 
        \wNDiag_63[63] , \wPDiag_17[19] , \wPDiag_34[28] , \wNDiag_40[52] , 
        \wPDiag_62[30] , \wPDiag_41[18] , \wNDiag_35[62] , \wNDiag_5[22] , 
        \wPDiag_32[0] , \wColumn_60[1] , \wNDiag_28[33] , \wPDiag_3[61] , 
        \wNDiag_4[8] , \wColumn_8[6] , \wColumn_16[15] , \wColumn_20[10] , 
        \wPDiag_29[60] , \wPDiag_48[8] , \wNDiag_48[37] , \wColumn_55[39] , 
        \wColumn_55[20] , \wPDiag_55[7] , \wColumn_63[25] , \wColumn_35[24] , 
        \wNDiag_5[11] , \wColumn_40[14] , \wColumn_28[46] , \wColumn_48[42] , 
        \wNDiag_6[61] , \wNDiag_6[52] , \wColumn_8[25] , \wNDiag_16[60] , 
        \wPDiag_56[4] , \wPDiag_17[33] , \wNDiag_35[48] , \wScan_36[4] , 
        \wPDiag_41[32] , \wNDiag_63[50] , \wPDiag_21[36] , \wNDiag_35[51] , 
        \wNDiag_40[61] , \wNDiag_55[55] , \wNDiag_63[49] , \wPDiag_57[45] , 
        \wNDiag_15[23] , \wNDiag_23[26] , \wNDiag_56[16] , \wNDiag_36[12] , 
        \wPDiag_37[58] , \wNDiag_43[22] , \wPDiag_61[40] , \wNDiag_60[13] , 
        \wPDiag_61[59] , \wPDiag_37[41] , \wNDiag_62[0] , \wColumn_15[56] , 
        \wColumn_43[57] , \wNDiag_61[3] , \wColumn_23[53] , \wPDiag_29[1] , 
        \wColumn_56[63] , \wScan_49[1] , \wPDiag_14[43] , \wCall_28[0] , 
        \wNDiag_36[21] , \wNDiag_15[10] , \wNDiag_36[38] , \wNDiag_43[11] , 
        \wNDiag_60[39] , \wPDiag_22[46] , \wPDiag_42[42] , \wNDiag_60[20] , 
        \wColumn_8[16] , \wNDiag_18[8] , \wNDiag_23[15] , \wPDiag_53[9] , 
        \wNDiag_56[25] , \wNDiag_2[63] , \wNDiag_2[50] , \wPDiag_8[47] , 
        \wColumn_11[54] , \wPDiag_18[24] , \wColumn_23[60] , \wColumn_56[49] , 
        \wColumn_36[54] , \wColumn_56[50] , \wColumn_60[55] , \wNDiag_21[1] , 
        \wColumn_27[51] , \wColumn_27[48] , \wColumn_52[61] , \wColumn_47[55] , 
        \wNDiag_2[49] , \wColumn_38[1] , \wColumn_4[42] , \wPDiag_4[39] , 
        \wPDiag_4[20] , \wPDiag_10[8] , \wNDiag_11[38] , \wNDiag_22[2] , 
        \wNDiag_47[20] , \wNDiag_11[21] , \wNDiag_32[10] , \wNDiag_47[39] , 
        \wPDiag_18[17] , \wColumn_27[62] , \wNDiag_27[24] , \wPDiag_33[43] , 
        \wNDiag_52[14] , \wPDiag_53[47] , \wColumn_32[56] , \wColumn_42[9] , 
        \wNDiag_45[5] , \wColumn_52[52] , \wNDiag_19[44] , \wPDiag_4[13] , 
        \wScan_5[2] , \wScan_6[1] , \wPDiag_10[58] , \wPDiag_10[41] , 
        \wPDiag_26[44] , \wNDiag_27[17] , \wNDiag_32[23] , \wNDiag_52[27] , 
        \wPDiag_46[59] , \wNDiag_47[13] , \wNDiag_11[12] , \wPDiag_46[40] , 
        \wPDiag_3[6] , \wColumn_19[31] , \wColumn_19[28] , \wNDiag_46[6] , 
        \wNDiag_1[20] , \wColumn_20[3] , \wColumn_39[43] , \wNDiag_1[13] , 
        \wColumn_7[18] , \wPDiag_7[50] , \wPDiag_7[49] , \wColumn_59[47] , 
        \wScan_12[2] , \wNDiag_12[51] , \wPDiag_30[33] , \wNDiag_44[49] , 
        \wNDiag_12[48] , \wNDiag_31[60] , \wNDiag_44[50] , \wNDiag_24[54] , 
        \wPDiag_50[37] , \wNDiag_59[32] , \wPDiag_7[63] , \wScan_11[1] , 
        \wPDiag_58[61] , \wColumn_12[24] , \wColumn_23[0] , \wColumn_24[38] , 
        \wColumn_24[21] , \wNDiag_39[36] , \wColumn_51[11] , \wNDiag_39[3] , 
        \wNDiag_12[62] , \wPDiag_13[28] , \wPDiag_25[34] , \wColumn_31[15] , 
        \wColumn_44[25] , \wNDiag_51[57] , \wColumn_59[8] , \wPDiag_13[31] , 
        \wPDiag_45[30] , \wPDiag_30[19] , \wNDiag_31[53] , \wNDiag_44[63] , 
        \wPDiag_45[29] , \wPDiag_16[6] , \wColumn_44[7] , \wColumn_2[23] , 
        \wNDiag_3[43] , \wColumn_5[51] , \wPDiag_5[19] , \wPDiag_5[8] , 
        \wNDiag_9[45] , \wColumn_12[17] , \wPDiag_15[5] , \wColumn_31[26] , 
        \wColumn_47[4] , \wColumn_24[12] , \wColumn_44[16] , \wPDiag_38[56] , 
        \wColumn_51[22] , \wColumn_7[32] , \wPDiag_58[52] , \wNDiag_59[18] , 
        \wNDiag_40[8] , \wNDiag_10[18] , \wColumn_18[22] , \wScan_63[1] , 
        \wPDiag_27[57] , \wColumn_51[0] , \wNDiag_53[34] , \wPDiag_11[52] , 
        \wNDiag_18[57] , \wPDiag_32[63] , \wNDiag_33[30] , \wNDiag_33[29] , 
        \wNDiag_46[19] , \wPDiag_47[53] , \wNDiag_48[0] , \wColumn_52[3] , 
        \wColumn_5[48] , \wNDiag_10[32] , \wPDiag_11[61] , \wPDiag_32[49] , 
        \wColumn_33[45] , \wNDiag_46[33] , \wColumn_53[58] , \wColumn_53[41] , 
        \wScan_60[2] , \wPDiag_32[50] , \wPDiag_47[60] , \wColumn_35[4] , 
        \wNDiag_26[37] , \wPDiag_52[54] , \wColumn_5[62] , \wPDiag_5[33] , 
        \wColumn_18[11] , \wNDiag_32[8] , \wColumn_10[47] , \wColumn_26[42] , 
        \wColumn_46[46] , \wColumn_36[7] , \wColumn_6[38] , \wPDiag_18[0] , 
        \wPDiag_19[37] , \wPDiag_39[45] , \wNDiag_38[16] , \wNDiag_50[2] , 
        \wNDiag_58[12] , \wPDiag_59[58] , \wColumn_6[21] , \wPDiag_59[41] , 
        \wColumn_6[12] , \wNDiag_8[56] , \wColumn_30[35] , \wPDiag_12[22] , 
        \wPDiag_24[27] , \wColumn_25[18] , \wColumn_50[31] , \wColumn_38[63] , 
        \wColumn_50[28] , \wColumn_49[2] , \wNDiag_50[44] , \wNDiag_30[59] , 
        \wPDiag_31[13] , \wPDiag_51[17] , \wNDiag_30[40] , \wPDiag_44[23] , 
        \wNDiag_53[1] , \wColumn_13[37] , \wColumn_25[32] , \wNDiag_29[9] , 
        \wColumn_45[36] , \wNDiag_58[38] , \wNDiag_58[21] , \wColumn_6[0] , 
        \wPDiag_6[43] , \wPDiag_12[11] , \wNDiag_13[42] , \wNDiag_34[6] , 
        \wReturn_58[0] , \wNDiag_38[25] , \wPDiag_44[10] , \wPDiag_31[20] , 
        \wNDiag_45[43] , \wPDiag_24[14] , \wNDiag_25[47] , \wPDiag_31[39] , 
        \wNDiag_37[5] , \wPDiag_51[24] , \wColumn_30[9] , \wColumn_38[50] , 
        \wColumn_38[49] , \wPDiag_62[8] , \wColumn_58[54] , \wNDiag_13[3] , 
        \wPDiag_16[39] , \wPDiag_35[11] , \wPDiag_40[21] , \wNDiag_62[43] , 
        \wPDiag_16[20] , \wNDiag_34[42] , \wPDiag_40[38] , \wPDiag_63[10] , 
        \wNDiag_54[46] , \wNDiag_10[0] , \wPDiag_20[25] , \wColumn_29[55] , 
        \wColumn_49[51] , \wColumn_49[48] , \wPDiag_55[15] , \wColumn_34[37] , 
        \wScan_38[2] , \wColumn_54[33] , \wColumn_62[36] , \wNDiag_29[20] , 
        \wPDiag_2[58] , \wColumn_5[3] , \wCall_6[0] , \wNDiag_29[39] , 
        \wNDiag_49[24] , \wPDiag_58[2] , \wPDiag_2[41] , \wNDiag_4[31] , 
        \wNDiag_4[28] , \wNDiag_21[45] , \wColumn_49[62] , \wColumn_1[60] , 
        \wColumn_1[53] , \wColumn_2[10] , \wPDiag_16[13] , \wNDiag_17[40] , 
        \wPDiag_20[16] , \wPDiag_55[26] , \wPDiag_40[12] , \wNDiag_41[58] , 
        \wPDiag_35[22] , \wNDiag_41[41] , \wPDiag_63[23] , \wNDiag_17[59] , 
        \wPDiag_28[59] , \wPDiag_48[44] , \wNDiag_49[17] , \wPDiag_28[40] , 
        \wNDiag_29[13] , \wPDiag_9[54] , \wColumn_17[35] , \wColumn_21[30] , 
        \wColumn_41[34] , \wColumn_21[29] , \wPDiag_21[9] , \wColumn_54[19] , 
        \wScan_20[0] , \wColumn_37[47] , \wColumn_57[43] , \wColumn_61[46] , 
        \wColumn_11[2] , \wColumn_12[1] , \wPDiag_40[0] , \wPDiag_15[50] , 
        \wPDiag_15[49] , \wNDiag_37[32] , \wPDiag_43[48] , \wPDiag_60[60] , 
        \wPDiag_23[55] , \wPDiag_36[61] , \wPDiag_43[51] , \wNDiag_61[33] , 
        \wPDiag_43[3] , \wScan_23[3] , \wNDiag_57[36] , \wPDiag_24[4] , 
        \wPDiag_1[31] , \wColumn_14[45] , \wColumn_42[44] , \wScan_44[4] , 
        \wColumn_22[59] , \wColumn_22[40] , \wPDiag_1[28] , \wNDiag_2[44] , 
        \wColumn_4[56] , \wNDiag_7[58] , \wNDiag_7[41] , \wColumn_9[36] , 
        \wPDiag_56[56] , \wPDiag_10[55] , \wPDiag_13[6] , \wNDiag_14[30] , 
        \wNDiag_14[29] , \wPDiag_15[63] , \wNDiag_22[35] , \wNDiag_42[31] , 
        \wPDiag_60[53] , \wNDiag_61[19] , \wPDiag_27[7] , \wPDiag_36[52] , 
        \wNDiag_37[18] , \wNDiag_42[28] , \wPDiag_43[62] , \wColumn_19[25] , 
        \wPDiag_26[50] , \wPDiag_26[49] , \wColumn_41[7] , \wPDiag_53[60] , 
        \wNDiag_52[33] , \wPDiag_10[5] , \wNDiag_19[50] , \wNDiag_19[49] , 
        \wNDiag_32[37] , \wPDiag_46[54] , \wColumn_42[4] , \wNDiag_58[7] , 
        \wNDiag_11[35] , \wColumn_25[3] , \wColumn_32[42] , \wPDiag_33[57] , 
        \wNDiag_45[8] , \wNDiag_47[34] , \wColumn_52[46] , \wPDiag_26[63] , 
        \wNDiag_27[29] , \wNDiag_52[19] , \wPDiag_53[53] , \wNDiag_27[30] , 
        \wPDiag_4[34] , \wColumn_19[16] , \wScan_17[2] , \wColumn_27[45] , 
        \wScan_0[2] , \wColumn_11[59] , \wColumn_47[41] , \wColumn_11[40] , 
        \wScan_14[1] , \wColumn_47[58] , \wPDiag_18[30] , \wColumn_26[0] , 
        \wPDiag_18[29] , \wNDiag_19[63] , \wPDiag_5[5] , \wPDiag_38[42] , 
        \wNDiag_39[11] , \wNDiag_59[15] , \wColumn_7[26] , \wNDiag_40[5] , 
        \wPDiag_58[46] , \wNDiag_9[51] , \wNDiag_9[48] , \wColumn_31[32] , 
        \wColumn_47[9] , \wPDiag_15[8] , \wColumn_51[36] , \wColumn_1[47] , 
        \wPDiag_1[25] , \wNDiag_1[34] , \wScan_3[1] , \wColumn_59[60] , 
        \wPDiag_6[6] , \wPDiag_25[39] , \wPDiag_25[20] , \wNDiag_51[43] , 
        \wColumn_59[5] , \wPDiag_30[14] , \wPDiag_50[10] , \wNDiag_31[47] , 
        \wNDiag_43[6] , \wPDiag_45[24] , \wColumn_7[15] , \wNDiag_9[62] , 
        \wColumn_12[30] , \wPDiag_13[25] , \wColumn_24[35] , \wColumn_31[18] , 
        \wColumn_44[28] , \wColumn_12[29] , \wColumn_44[31] , \wNDiag_59[26] , 
        \wNDiag_12[45] , \wNDiag_24[1] , \wNDiag_39[22] , \wPDiag_45[17] , 
        \wPDiag_13[16] , \wPDiag_30[27] , \wNDiag_44[44] , \wNDiag_24[59] , 
        \wNDiag_24[40] , \wNDiag_27[2] , \wPDiag_50[23] , \wPDiag_25[13] , 
        \wColumn_39[57] , \wNDiag_1[8] , \wColumn_3[24] , \wNDiag_4[5] , 
        \wPDiag_7[44] , \wColumn_59[53] , \wNDiag_7[6] , \wPDiag_17[27] , 
        \wPDiag_34[16] , \wNDiag_35[45] , \wPDiag_41[26] , \wNDiag_63[44] , 
        \wColumn_19[7] , \wNDiag_55[41] , \wPDiag_62[17] , \wPDiag_21[22] , 
        \wColumn_28[52] , \wColumn_48[56] , \wPDiag_54[12] , \wNDiag_55[58] , 
        \wPDiag_56[9] , \wScan_28[5] , \wColumn_55[34] , \wColumn_16[18] , 
        \wColumn_35[29] , \wColumn_40[19] , \wColumn_63[31] , \wNDiag_28[27] , 
        \wColumn_35[30] , \wColumn_63[28] , \wColumn_3[17] , \wPDiag_3[46] , 
        \wColumn_28[61] , \wPDiag_48[5] , \wNDiag_48[23] , \wNDiag_5[36] , 
        \wNDiag_16[47] , \wNDiag_20[42] , \wPDiag_54[38] , \wPDiag_21[11] , 
        \wPDiag_54[21] , \wPDiag_41[15] , \wPDiag_17[14] , \wPDiag_34[25] , 
        \wNDiag_40[46] , \wPDiag_62[24] , \wNDiag_28[14] , \wNDiag_48[10] , 
        \wPDiag_49[43] , \wPDiag_29[47] , \wPDiag_8[53] , \wColumn_16[32] , 
        \wColumn_20[37] , \wColumn_40[33] , \wNDiag_18[5] , \wColumn_36[59] , 
        \wColumn_36[40] , \wColumn_56[44] , \wColumn_60[58] , \wColumn_60[41] , 
        \wColumn_2[37] , \wPDiag_2[55] , \wNDiag_6[46] , \wPDiag_8[60] , 
        \wPDiag_14[57] , \wPDiag_50[7] , \wColumn_15[42] , \wPDiag_22[52] , 
        \wNDiag_36[35] , \wPDiag_42[56] , \wNDiag_60[34] , \wNDiag_23[18] , 
        \wScan_33[4] , \wPDiag_53[4] , \wNDiag_56[31] , \wNDiag_56[28] , 
        \wPDiag_57[62] , \wPDiag_34[3] , \wColumn_43[43] , \wScan_54[3] , 
        \wColumn_23[47] , \wScan_57[0] , \wColumn_8[31] , \wPDiag_57[51] , 
        \wColumn_8[28] , \wPDiag_22[61] , \wPDiag_57[48] , \wNDiag_15[37] , 
        \wNDiag_23[32] , \wPDiag_37[55] , \wNDiag_43[36] , \wPDiag_61[54] , 
        \wPDiag_37[0] , \wColumn_17[38] , \wColumn_17[21] , \wColumn_41[39] , 
        \wColumn_62[11] , \wColumn_41[20] , \wNDiag_17[54] , \wColumn_21[24] , 
        \wColumn_34[10] , \wColumn_54[14] , \wPDiag_21[4] , \wNDiag_21[51] , 
        \wPDiag_28[54] , \wScan_41[4] , \wPDiag_48[50] , \wPDiag_48[49] , 
        \wNDiag_54[61] , \wNDiag_21[48] , \wPDiag_55[32] , \wPDiag_35[36] , 
        \wNDiag_41[55] , \wPDiag_63[37] , \wNDiag_4[25] , \wPDiag_22[7] , 
        \wNDiag_29[34] , \wNDiag_4[16] , \wNDiag_9[0] , \wScan_25[0] , 
        \wPDiag_48[63] , \wNDiag_49[29] , \wColumn_17[12] , \wColumn_21[17] , 
        \wNDiag_49[30] , \wColumn_54[27] , \wColumn_17[1] , \wPDiag_45[0] , 
        \wColumn_34[23] , \wColumn_62[22] , \wColumn_41[13] , \wColumn_9[22] , 
        \wColumn_14[2] , \wColumn_29[58] , \wColumn_29[41] , \wColumn_49[45] , 
        \wPDiag_46[3] , \wPDiag_16[34] , \wScan_26[3] , \wPDiag_40[35] , 
        \wNDiag_62[57] , \wPDiag_20[31] , \wPDiag_20[28] , \wNDiag_21[62] , 
        \wNDiag_34[56] , \wNDiag_54[52] , \wPDiag_55[18] , \wPDiag_56[42] , 
        \wNDiag_14[24] , \wNDiag_22[38] , \wNDiag_22[21] , \wNDiag_57[11] , 
        \wNDiag_37[15] , \wNDiag_42[25] , \wPDiag_60[47] , \wNDiag_61[14] , 
        \wPDiag_36[46] , \wPDiag_1[16] , \wColumn_3[0] , \wNDiag_7[55] , 
        \wColumn_14[51] , \wColumn_14[48] , \wColumn_37[60] , \wColumn_42[50] , 
        \wColumn_42[49] , \wColumn_61[61] , \wNDiag_16[3] , \wColumn_22[54] , 
        \wPDiag_39[6] , \wPDiag_24[9] , \wScan_59[6] , \wColumn_9[11] , 
        \wNDiag_14[17] , \wPDiag_15[44] , \wNDiag_37[26] , \wNDiag_42[16] , 
        \wPDiag_23[41] , \wPDiag_43[45] , \wNDiag_61[27] , \wNDiag_22[12] , 
        \wPDiag_23[58] , \wNDiag_57[22] , \wCall_3[0] , \wPDiag_9[59] , 
        \wPDiag_9[40] , \wNDiag_15[0] , \wColumn_14[62] , \wColumn_37[53] , 
        \wColumn_57[57] , \wColumn_42[63] , \wNDiag_3[57] , \wColumn_10[53] , 
        \wScan_19[4] , \wPDiag_19[23] , \wColumn_61[52] , \wColumn_26[56] , 
        \wNDiag_31[6] , \wColumn_46[52] , \wColumn_33[62] , \wColumn_5[45] , 
        \wPDiag_5[27] , \wColumn_28[6] , \wColumn_10[60] , \wNDiag_10[26] , 
        \wNDiag_32[5] , \wNDiag_33[17] , \wColumn_35[9] , \wNDiag_46[27] , 
        \wNDiag_26[23] , \wPDiag_32[44] , \wPDiag_52[59] , \wPDiag_52[40] , 
        \wNDiag_53[13] , \wColumn_33[51] , \wColumn_46[61] , \wNDiag_18[43] , 
        \wPDiag_19[10] , \wColumn_33[48] , \wColumn_53[55] , \wNDiag_55[2] , 
        \wPDiag_5[14] , \wNDiag_10[15] , \wPDiag_11[46] , \wNDiag_26[10] , 
        \wPDiag_27[43] , \wNDiag_53[39] , \wNDiag_33[24] , \wNDiag_53[20] , 
        \wNDiag_46[14] , \wPDiag_47[47] , \wPDiag_6[57] , \wColumn_18[36] , 
        \wNDiag_56[1] , \wColumn_30[4] , \wColumn_38[44] , \wPDiag_62[5] , 
        \wColumn_58[40] , \wNDiag_13[56] , \wPDiag_31[34] , \wColumn_58[59] , 
        \wPDiag_24[19] , \wNDiag_45[57] , \wNDiag_50[63] , \wPDiag_51[29] , 
        \wNDiag_25[53] , \wNDiag_37[8] , \wPDiag_51[30] , \wNDiag_38[31] , 
        \wNDiag_38[28] , \wNDiag_58[35] , \wPDiag_39[62] , \wColumn_50[16] , 
        \wNDiag_8[42] , \wPDiag_12[36] , \wColumn_13[23] , \wColumn_25[26] , 
        \wNDiag_29[4] , \wColumn_33[7] , \wPDiag_61[6] , \wPDiag_24[33] , 
        \wNDiag_25[60] , \wColumn_30[12] , \wColumn_45[22] , \wNDiag_50[50] , 
        \wPDiag_44[37] , \wNDiag_50[49] , \wColumn_13[10] , \wColumn_30[38] , 
        \wNDiag_30[54] , \wColumn_54[0] , \wColumn_30[21] , \wColumn_57[3] , 
        \wColumn_25[15] , \wColumn_45[11] , \wColumn_50[25] , \wColumn_1[57] , 
        \wColumn_3[9] , \wColumn_6[35] , \wPDiag_8[0] , \wPDiag_39[51] , 
        \wPDiag_39[48] , \wPDiag_59[55] , \wColumn_9[18] , \wPDiag_23[48] , 
        \wNDiag_57[32] , \wColumn_11[6] , \wPDiag_23[51] , \wPDiag_43[7] , 
        \wPDiag_56[61] , \wColumn_12[5] , \wPDiag_15[54] , \wPDiag_43[55] , 
        \wNDiag_61[37] , \wNDiag_37[36] , \wPDiag_40[4] , \wPDiag_1[35] , 
        \wNDiag_7[45] , \wColumn_9[32] , \wPDiag_9[50] , \wPDiag_9[49] , 
        \wColumn_37[43] , \wColumn_61[42] , \wColumn_57[47] , \wNDiag_14[34] , 
        \wNDiag_15[9] , \wScan_20[4] , \wPDiag_27[3] , \wPDiag_36[56] , 
        \wNDiag_22[31] , \wNDiag_42[35] , \wPDiag_60[57] , \wPDiag_56[52] , 
        \wNDiag_57[18] , \wNDiag_22[28] , \wPDiag_23[62] , \wColumn_2[27] , 
        \wColumn_5[7] , \wPDiag_9[63] , \wColumn_22[44] , \wScan_47[3] , 
        \wColumn_14[58] , \wColumn_14[41] , \wColumn_42[59] , \wScan_44[0] , 
        \wColumn_42[40] , \wPDiag_24[0] , \wNDiag_49[20] , \wPDiag_58[6] , 
        \wNDiag_9[9] , \wNDiag_49[39] , \wColumn_2[14] , \wColumn_6[4] , 
        \wNDiag_10[4] , \wColumn_17[8] , \wNDiag_29[24] , \wColumn_34[33] , 
        \wColumn_29[51] , \wColumn_29[48] , \wScan_38[6] , \wPDiag_45[9] , 
        \wColumn_62[32] , \wColumn_54[37] , \wColumn_49[55] , \wNDiag_13[7] , 
        \wPDiag_20[38] , \wPDiag_20[21] , \wPDiag_55[11] , \wNDiag_54[42] , 
        \wPDiag_16[24] , \wNDiag_34[46] , \wColumn_17[31] , \wColumn_17[28] , 
        \wColumn_21[34] , \wPDiag_35[15] , \wPDiag_63[14] , \wPDiag_40[25] , 
        \wNDiag_62[47] , \wColumn_41[30] , \wColumn_62[18] , \wColumn_34[19] , 
        \wColumn_41[29] , \wPDiag_28[44] , \wPDiag_2[45] , \wNDiag_4[35] , 
        \wPDiag_16[17] , \wNDiag_29[17] , \wNDiag_41[45] , \wPDiag_48[59] , 
        \wPDiag_48[40] , \wNDiag_49[13] , \wPDiag_63[27] , \wNDiag_17[44] , 
        \wPDiag_40[16] , \wPDiag_20[12] , \wPDiag_35[26] , \wPDiag_55[22] , 
        \wNDiag_21[58] , \wNDiag_21[41] , \wPDiag_12[26] , \wColumn_29[62] , 
        \wNDiag_30[44] , \wNDiag_53[5] , \wPDiag_24[23] , \wPDiag_31[17] , 
        \wPDiag_44[27] , \wColumn_49[6] , \wNDiag_50[59] , \wPDiag_51[13] , 
        \wNDiag_50[40] , \wColumn_54[9] , \wColumn_58[63] , \wNDiag_1[24] , 
        \wNDiag_3[47] , \wColumn_5[55] , \wColumn_6[25] , \wPDiag_8[9] , 
        \wNDiag_8[52] , \wColumn_13[19] , \wColumn_50[35] , \wColumn_30[31] , 
        \wColumn_30[28] , \wColumn_45[18] , \wPDiag_59[45] , \wColumn_6[16] , 
        \wPDiag_6[47] , \wPDiag_18[4] , \wNDiag_50[6] , \wNDiag_58[16] , 
        \wNDiag_38[12] , \wPDiag_39[58] , \wPDiag_39[41] , \wPDiag_12[15] , 
        \wPDiag_24[10] , \wColumn_38[54] , \wColumn_58[50] , \wColumn_58[49] , 
        \wPDiag_51[20] , \wNDiag_25[43] , \wNDiag_37[1] , \wPDiag_51[39] , 
        \wNDiag_45[47] , \wNDiag_13[46] , \wPDiag_44[14] , \wPDiag_31[24] , 
        \wNDiag_34[2] , \wNDiag_38[38] , \wNDiag_38[21] , \wScan_8[3] , 
        \wNDiag_8[61] , \wNDiag_58[25] , \wColumn_13[33] , \wColumn_45[32] , 
        \wColumn_25[36] , \wColumn_53[45] , \wColumn_33[58] , \wScan_60[6] , 
        \wColumn_33[41] , \wNDiag_48[4] , \wPDiag_5[37] , \wColumn_10[43] , 
        \wPDiag_11[56] , \wNDiag_18[53] , \wPDiag_19[19] , \wPDiag_47[57] , 
        \wColumn_52[7] , \wColumn_18[26] , \wNDiag_26[19] , \wNDiag_33[34] , 
        \wNDiag_53[30] , \wPDiag_27[53] , \wColumn_51[4] , \wPDiag_52[63] , 
        \wNDiag_53[29] , \wNDiag_56[8] , \wScan_63[5] , \wNDiag_18[60] , 
        \wPDiag_19[33] , \wColumn_36[3] , \wColumn_26[46] , \wColumn_46[42] , 
        \wColumn_18[15] , \wPDiag_7[54] , \wNDiag_10[36] , \wNDiag_26[33] , 
        \wPDiag_52[49] , \wPDiag_27[60] , \wPDiag_52[50] , \wPDiag_32[54] , 
        \wColumn_35[0] , \wScan_11[5] , \wColumn_12[39] , \wColumn_44[21] , 
        \wNDiag_46[37] , \wColumn_12[20] , \wColumn_31[11] , \wNDiag_39[7] , 
        \wColumn_44[38] , \wColumn_23[4] , \wColumn_24[25] , \wColumn_51[15] , 
        \wNDiag_24[8] , \wNDiag_39[32] , \wPDiag_38[61] , \wScan_12[6] , 
        \wNDiag_24[49] , \wPDiag_50[33] , \wNDiag_59[36] , \wNDiag_12[55] , 
        \wNDiag_24[50] , \wNDiag_51[60] , \wPDiag_30[37] , \wNDiag_44[54] , 
        \wColumn_39[47] , \wColumn_59[43] , \wNDiag_1[17] , \wColumn_7[36] , 
        \wCall_14[0] , \wColumn_20[7] , \wPDiag_58[56] , \wNDiag_9[58] , 
        \wNDiag_9[41] , \wColumn_24[16] , \wPDiag_38[52] , \wNDiag_39[18] , 
        \wColumn_31[22] , \wColumn_51[26] , \wColumn_12[13] , \wColumn_44[12] , 
        \wPDiag_15[1] , \wColumn_47[0] , \wNDiag_2[54] , \wPDiag_4[24] , 
        \wNDiag_11[25] , \wPDiag_13[35] , \wPDiag_16[2] , \wColumn_44[3] , 
        \wNDiag_24[63] , \wPDiag_25[30] , \wNDiag_31[57] , \wPDiag_45[34] , 
        \wPDiag_25[29] , \wNDiag_27[39] , \wNDiag_27[20] , \wPDiag_50[19] , 
        \wNDiag_51[53] , \wNDiag_52[10] , \wPDiag_53[43] , \wNDiag_22[6] , 
        \wNDiag_32[14] , \wPDiag_33[47] , \wNDiag_47[24] , \wColumn_38[5] , 
        \wColumn_1[55] , \wNDiag_1[26] , \wNDiag_1[1] , \wPDiag_3[2] , 
        \wColumn_11[50] , \wColumn_47[48] , \wColumn_11[49] , \wNDiag_21[5] , 
        \wColumn_47[51] , \wColumn_32[61] , \wPDiag_18[39] , \wColumn_27[55] , 
        \wPDiag_18[20] , \wColumn_19[35] , \wColumn_26[9] , \wColumn_4[46] , 
        \wPDiag_4[17] , \wNDiag_46[2] , \wScan_6[5] , \wNDiag_11[16] , 
        \wPDiag_10[45] , \wNDiag_32[27] , \wPDiag_46[44] , \wPDiag_26[59] , 
        \wNDiag_47[17] , \wPDiag_26[40] , \wNDiag_27[13] , \wNDiag_52[23] , 
        \wScan_5[6] , \wNDiag_6[56] , \wColumn_11[63] , \wPDiag_18[13] , 
        \wNDiag_19[40] , \wNDiag_19[59] , \wNDiag_45[1] , \wColumn_52[56] , 
        \wColumn_15[52] , \wColumn_23[57] , \wPDiag_29[5] , \wColumn_32[52] , 
        \wColumn_47[62] , \wScan_49[5] , \wColumn_60[62] , \wColumn_36[63] , 
        \wColumn_43[53] , \wNDiag_61[7] , \wColumn_8[38] , \wNDiag_15[27] , 
        \wNDiag_60[17] , \wNDiag_62[4] , \wNDiag_36[16] , \wPDiag_37[45] , 
        \wPDiag_37[9] , \wNDiag_43[26] , \wPDiag_61[44] , \wNDiag_56[12] , 
        \wPDiag_57[58] , \wColumn_8[21] , \wNDiag_23[22] , \wPDiag_57[41] , 
        \wPDiag_8[43] , \wColumn_15[61] , \wColumn_36[50] , \wColumn_36[49] , 
        \wColumn_60[51] , \wColumn_43[60] , \wColumn_56[54] , \wColumn_60[48] , 
        \wNDiag_2[2] , \wPDiag_22[42] , \wNDiag_23[11] , \wNDiag_56[21] , 
        \wColumn_3[34] , \wPDiag_3[56] , \wNDiag_5[26] , \wColumn_8[12] , 
        \wNDiag_56[38] , \wPDiag_14[47] , \wNDiag_15[14] , \wNDiag_36[25] , 
        \wPDiag_42[46] , \wNDiag_60[24] , \wNDiag_43[15] , \wPDiag_32[4] , 
        \wColumn_60[5] , \wNDiag_5[15] , \wReturn_16[0] , \wColumn_16[22] , 
        \wNDiag_16[57] , \wPDiag_34[35] , \wNDiag_40[56] , \wPDiag_62[34] , 
        \wColumn_20[27] , \wNDiag_20[52] , \wScan_52[4] , \wPDiag_54[31] , 
        \wPDiag_54[28] , \wNDiag_55[62] , \wPDiag_21[18] , \wPDiag_29[57] , 
        \wPDiag_31[7] , \wNDiag_48[19] , \wPDiag_49[53] , \wColumn_63[6] , 
        \wColumn_55[17] , \wColumn_35[13] , \wColumn_40[23] , \wColumn_63[12] , 
        \wPDiag_17[37] , \wNDiag_20[61] , \wPDiag_21[32] , \wNDiag_55[48] , 
        \wNDiag_55[51] , \wColumn_28[42] , \wNDiag_35[55] , \wScan_36[0] , 
        \wPDiag_41[36] , \wPDiag_56[0] , \wNDiag_63[54] , \wColumn_8[2] , 
        \wColumn_35[20] , \wColumn_48[46] , \wColumn_16[11] , \wColumn_35[39] , 
        \wColumn_40[10] , \wColumn_63[38] , \wColumn_20[14] , \wPDiag_55[3] , 
        \wColumn_63[21] , \wNDiag_48[33] , \wColumn_55[24] , \wPDiag_49[60] , 
        \wNDiag_28[37] , \wScan_35[3] , \wNDiag_1[15] , \wPDiag_7[56] , 
        \wColumn_20[5] , \wColumn_39[45] , \wColumn_59[58] , \wScan_12[4] , 
        \wNDiag_12[57] , \wNDiag_44[56] , \wReturn_56[0] , \wColumn_59[41] , 
        \wPDiag_30[35] , \wColumn_12[22] , \wColumn_23[6] , \wNDiag_24[52] , 
        \wNDiag_27[9] , \wPDiag_50[31] , \wPDiag_25[18] , \wPDiag_38[63] , 
        \wNDiag_39[30] , \wPDiag_50[28] , \wNDiag_51[62] , \wNDiag_59[34] , 
        \wNDiag_39[29] , \wColumn_24[27] , \wColumn_31[13] , \wColumn_51[17] , 
        \wColumn_44[23] , \wPDiag_13[37] , \wNDiag_24[61] , \wPDiag_25[32] , 
        \wNDiag_39[5] , \wNDiag_51[48] , \wNDiag_51[51] , \wNDiag_31[55] , 
        \wPDiag_16[0] , \wColumn_44[1] , \wPDiag_45[36] , \wNDiag_1[3] , 
        \wNDiag_2[56] , \wColumn_7[34] , \wNDiag_9[43] , \wColumn_12[11] , 
        \wPDiag_15[3] , \wColumn_31[20] , \wColumn_44[10] , \wColumn_47[2] , 
        \wColumn_24[14] , \wColumn_31[39] , \wColumn_51[24] , \wPDiag_38[50] , 
        \wPDiag_38[49] , \wPDiag_58[54] , \wColumn_11[52] , \wPDiag_18[22] , 
        \wColumn_27[57] , \wNDiag_21[7] , \wColumn_32[63] , \wColumn_47[53] , 
        \wNDiag_2[0] , \wPDiag_3[0] , \wColumn_4[44] , \wPDiag_4[26] , 
        \wNDiag_22[4] , \wColumn_38[7] , \wScan_5[4] , \wColumn_11[61] , 
        \wNDiag_11[27] , \wPDiag_33[45] , \wColumn_25[8] , \wNDiag_27[22] , 
        \wNDiag_32[16] , \wNDiag_47[26] , \wColumn_32[49] , \wNDiag_52[12] , 
        \wPDiag_53[58] , \wPDiag_53[41] , \wPDiag_18[11] , \wNDiag_19[42] , 
        \wColumn_32[50] , \wColumn_47[60] , \wNDiag_45[3] , \wColumn_52[54] , 
        \wPDiag_4[15] , \wPDiag_10[47] , \wNDiag_11[14] , \wPDiag_26[42] , 
        \wNDiag_27[11] , \wNDiag_52[21] , \wNDiag_52[38] , \wPDiag_46[46] , 
        \wNDiag_47[15] , \wNDiag_32[25] , \wColumn_19[37] , \wNDiag_6[54] , 
        \wColumn_8[23] , \wNDiag_23[39] , \wNDiag_23[20] , \wNDiag_46[0] , 
        \wNDiag_56[10] , \wPDiag_57[43] , \wNDiag_15[25] , \wPDiag_37[47] , 
        \wNDiag_36[14] , \wNDiag_60[15] , \wNDiag_43[24] , \wPDiag_61[46] , 
        \wNDiag_62[6] , \wColumn_8[10] , \wPDiag_14[45] , \wColumn_15[50] , 
        \wColumn_15[49] , \wColumn_43[48] , \wColumn_60[60] , \wNDiag_15[16] , 
        \wColumn_23[55] , \wColumn_36[61] , \wColumn_43[51] , \wNDiag_61[5] , 
        \wPDiag_29[7] , \wPDiag_34[8] , \wPDiag_42[44] , \wNDiag_60[26] , 
        \wNDiag_43[17] , \wPDiag_22[59] , \wNDiag_36[27] , \wNDiag_56[23] , 
        \wNDiag_23[13] , \wPDiag_22[40] , \wColumn_3[36] , \wPDiag_3[54] , 
        \wPDiag_8[58] , \wColumn_56[56] , \wPDiag_8[41] , \wColumn_15[63] , 
        \wColumn_60[53] , \wColumn_16[39] , \wColumn_35[11] , \wColumn_36[52] , 
        \wColumn_43[62] , \wColumn_16[20] , \wColumn_40[21] , \wNDiag_16[55] , 
        \wColumn_20[25] , \wPDiag_31[5] , \wColumn_40[38] , \wColumn_63[10] , 
        \wColumn_63[4] , \wNDiag_20[50] , \wNDiag_20[49] , \wPDiag_29[55] , 
        \wPDiag_49[51] , \wPDiag_49[48] , \wColumn_55[15] , \wScan_51[5] , 
        \wScan_52[6] , \wPDiag_54[33] , \wNDiag_40[54] , \wNDiag_55[60] , 
        \wPDiag_62[36] , \wPDiag_34[37] , \wNDiag_5[24] , \wPDiag_32[6] , 
        \wScan_35[1] , \wCall_54[0] , \wColumn_60[7] , \wNDiag_5[17] , 
        \wColumn_8[0] , \wColumn_20[16] , \wNDiag_28[35] , \wNDiag_48[31] , 
        \wNDiag_48[28] , \wPDiag_49[62] , \wColumn_55[26] , \wColumn_40[12] , 
        \wColumn_16[13] , \wColumn_35[22] , \wPDiag_55[1] , \wColumn_63[23] , 
        \wCall_8[0] , \wColumn_28[59] , \wColumn_48[44] , \wColumn_28[40] , 
        \wPDiag_56[2] , \wPDiag_9[52] , \wPDiag_17[35] , \wNDiag_35[57] , 
        \wScan_20[6] , \wNDiag_20[63] , \wPDiag_21[30] , \wScan_36[2] , 
        \wNDiag_63[56] , \wPDiag_41[34] , \wPDiag_21[29] , \wPDiag_54[19] , 
        \wNDiag_55[53] , \wColumn_57[45] , \wColumn_37[58] , \wColumn_61[40] , 
        \wColumn_37[41] , \wColumn_61[59] , \wPDiag_1[37] , \wPDiag_9[61] , 
        \wColumn_11[4] , \wColumn_12[7] , \wPDiag_15[56] , \wCall_26[0] , 
        \wPDiag_40[6] , \wNDiag_37[34] , \wPDiag_43[57] , \wNDiag_61[35] , 
        \wNDiag_57[30] , \wColumn_14[43] , \wNDiag_16[8] , \wNDiag_22[19] , 
        \wPDiag_43[5] , \wPDiag_56[63] , \wNDiag_57[29] , \wScan_23[5] , 
        \wPDiag_23[53] , \wPDiag_24[2] , \wScan_44[2] , \wColumn_22[46] , 
        \wColumn_42[42] , \wScan_47[1] , \wColumn_2[25] , \wColumn_6[6] , 
        \wNDiag_7[47] , \wColumn_9[30] , \wColumn_9[29] , \wNDiag_22[33] , 
        \wPDiag_56[49] , \wPDiag_23[60] , \wPDiag_56[50] , \wNDiag_13[5] , 
        \wNDiag_14[36] , \wPDiag_27[1] , \wPDiag_36[54] , \wNDiag_42[37] , 
        \wPDiag_60[55] , \wPDiag_63[16] , \wPDiag_16[26] , \wPDiag_20[23] , 
        \wNDiag_34[44] , \wPDiag_35[17] , \wPDiag_40[27] , \wNDiag_62[45] , 
        \wNDiag_54[59] , \wPDiag_55[13] , \wColumn_14[9] , \wColumn_29[53] , 
        \wColumn_49[57] , \wNDiag_54[40] , \wPDiag_46[8] , \wColumn_17[19] , 
        \wColumn_34[31] , \wScan_38[4] , \wColumn_54[35] , \wColumn_62[29] , 
        \wColumn_34[28] , \wColumn_41[18] , \wColumn_62[30] , \wColumn_2[16] , 
        \wPDiag_2[47] , \wColumn_5[5] , \wNDiag_10[6] , \wNDiag_29[26] , 
        \wNDiag_49[22] , \wPDiag_58[4] , \wNDiag_4[37] , \wColumn_29[60] , 
        \wPDiag_16[15] , \wPDiag_20[10] , \wNDiag_21[43] , \wPDiag_55[20] , 
        \wPDiag_55[39] , \wNDiag_17[46] , \wPDiag_35[24] , \wNDiag_41[47] , 
        \wPDiag_63[25] , \wPDiag_40[14] , \wPDiag_48[42] , \wNDiag_49[11] , 
        \wColumn_6[27] , \wColumn_17[33] , \wPDiag_28[46] , \wNDiag_29[15] , 
        \wColumn_41[32] , \wPDiag_18[6] , \wColumn_21[36] , \wNDiag_38[10] , 
        \wPDiag_39[43] , \wPDiag_59[47] , \wNDiag_8[50] , \wNDiag_50[4] , 
        \wNDiag_58[14] , \wColumn_57[8] , \wNDiag_8[49] , \wColumn_30[33] , 
        \wPDiag_12[24] , \wPDiag_24[38] , \wPDiag_24[21] , \wColumn_50[37] , 
        \wPDiag_51[11] , \wColumn_58[61] , \wColumn_49[4] , \wNDiag_50[42] , 
        \wNDiag_53[7] , \wNDiag_30[46] , \wPDiag_31[15] , \wPDiag_44[25] , 
        \wColumn_25[34] , \wReturn_0[0] , \wColumn_1[45] , \wPDiag_1[27] , 
        \wColumn_2[35] , \wPDiag_2[57] , \wNDiag_3[45] , \wColumn_5[57] , 
        \wColumn_6[14] , \wNDiag_8[63] , \wColumn_13[28] , \wColumn_13[31] , 
        \wColumn_45[30] , \wColumn_30[19] , \wColumn_45[29] , \wPDiag_6[45] , 
        \wPDiag_12[17] , \wNDiag_34[0] , \wNDiag_58[27] , \wNDiag_38[23] , 
        \wNDiag_13[44] , \wPDiag_31[26] , \wNDiag_45[45] , \wPDiag_24[12] , 
        \wPDiag_44[16] , \wNDiag_25[58] , \wNDiag_25[41] , \wPDiag_51[22] , 
        \wNDiag_37[3] , \wColumn_38[56] , \wPDiag_11[54] , \wColumn_18[24] , 
        \wColumn_58[52] , \wPDiag_27[51] , \wPDiag_27[48] , \wNDiag_53[32] , 
        \wColumn_51[6] , \wPDiag_52[61] , \wNDiag_33[36] , \wPDiag_47[55] , 
        \wNDiag_18[51] , \wColumn_52[5] , \wNDiag_18[48] , \wReturn_24[0] , 
        \wNDiag_48[6] , \wScan_8[1] , \wColumn_33[43] , \wColumn_53[47] , 
        \wNDiag_10[34] , \wNDiag_55[9] , \wScan_60[4] , \wColumn_18[17] , 
        \wNDiag_26[31] , \wPDiag_32[56] , \wColumn_35[2] , \wNDiag_46[35] , 
        \wNDiag_26[28] , \wPDiag_27[62] , \wPDiag_52[52] , \wNDiag_53[18] , 
        \wNDiag_4[27] , \wPDiag_5[35] , \wColumn_10[58] , \wColumn_10[41] , 
        \wColumn_26[44] , \wColumn_46[59] , \wNDiag_18[62] , \wPDiag_19[28] , 
        \wColumn_36[1] , \wColumn_46[40] , \wPDiag_19[31] , \wPDiag_22[5] , 
        \wNDiag_4[14] , \wColumn_14[0] , \wPDiag_16[36] , \wColumn_17[23] , 
        \wNDiag_17[56] , \wPDiag_20[19] , \wPDiag_35[34] , \wNDiag_41[57] , 
        \wPDiag_63[35] , \wColumn_21[26] , \wNDiag_21[53] , \wPDiag_28[56] , 
        \wScan_42[5] , \wNDiag_54[63] , \wPDiag_55[29] , \wPDiag_55[30] , 
        \wScan_41[6] , \wPDiag_48[52] , \wNDiag_49[18] , \wPDiag_21[6] , 
        \wColumn_54[16] , \wCall_47[0] , \wPDiag_20[33] , \wNDiag_21[60] , 
        \wColumn_34[12] , \wColumn_62[13] , \wColumn_41[22] , \wNDiag_54[50] , 
        \wNDiag_54[49] , \wScan_26[1] , \wPDiag_40[37] , \wNDiag_62[55] , 
        \wNDiag_34[54] , \wColumn_29[43] , \wPDiag_46[1] , \wNDiag_9[2] , 
        \wColumn_17[10] , \wColumn_17[3] , \wColumn_49[47] , \wPDiag_45[2] , 
        \wColumn_62[20] , \wColumn_21[15] , \wColumn_34[38] , \wColumn_34[21] , 
        \wColumn_41[11] , \wColumn_62[39] , \wColumn_54[25] , \wPDiag_48[61] , 
        \wNDiag_49[32] , \wScan_25[2] , \wNDiag_29[36] , \wNDiag_7[57] , 
        \wColumn_14[53] , \wColumn_22[56] , \wScan_59[4] , \wColumn_37[62] , 
        \wPDiag_39[4] , \wColumn_42[52] , \wColumn_61[63] , \wColumn_9[39] , 
        \wColumn_9[20] , \wNDiag_14[26] , \wPDiag_27[8] , \wNDiag_37[17] , 
        \wPDiag_36[44] , \wNDiag_42[27] , \wPDiag_60[45] , \wPDiag_56[40] , 
        \wNDiag_61[16] , \wNDiag_22[23] , \wPDiag_56[59] , \wNDiag_57[13] , 
        \wPDiag_9[42] , \wColumn_14[60] , \wColumn_37[51] , \wColumn_42[61] , 
        \wColumn_61[49] , \wColumn_37[48] , \wColumn_61[50] , \wNDiag_15[2] , 
        \wColumn_57[55] , \wPDiag_1[14] , \wColumn_9[13] , \wNDiag_57[39] , 
        \wNDiag_14[15] , \wPDiag_15[46] , \wNDiag_22[10] , \wPDiag_23[43] , 
        \wNDiag_57[20] , \wNDiag_42[14] , \wNDiag_37[24] , \wPDiag_43[47] , 
        \wNDiag_61[25] , \wColumn_3[2] , \wNDiag_3[55] , \wPDiag_5[25] , 
        \wNDiag_10[24] , \wNDiag_16[1] , \wNDiag_26[38] , \wNDiag_26[21] , 
        \wPDiag_52[42] , \wPDiag_32[46] , \wNDiag_33[15] , \wNDiag_53[11] , 
        \wNDiag_46[25] , \wNDiag_32[7] , \wPDiag_5[16] , \wColumn_10[51] , 
        \wColumn_10[48] , \wColumn_28[4] , \wNDiag_31[4] , \wColumn_33[60] , 
        \wColumn_46[50] , \wColumn_18[34] , \wScan_19[6] , \wColumn_26[54] , 
        \wColumn_46[49] , \wPDiag_19[38] , \wPDiag_19[21] , \wColumn_36[8] , 
        \wNDiag_56[3] , \wNDiag_10[17] , \wPDiag_11[44] , \wNDiag_46[16] , 
        \wNDiag_33[26] , \wPDiag_47[45] , \wNDiag_26[12] , \wPDiag_27[41] , 
        \wNDiag_53[22] , \wPDiag_27[58] , \wColumn_5[47] , \wColumn_10[62] , 
        \wNDiag_18[58] , \wNDiag_18[41] , \wPDiag_19[12] , \wColumn_33[53] , 
        \wColumn_46[63] , \wColumn_53[57] , \wNDiag_55[0] , \wColumn_13[38] , 
        \wColumn_13[21] , \wNDiag_29[6] , \wColumn_30[10] , \wColumn_45[39] , 
        \wColumn_25[24] , \wReturn_45[0] , \wColumn_45[20] , \wColumn_50[14] , 
        \wColumn_6[37] , \wPDiag_6[55] , \wNDiag_13[54] , \wNDiag_25[51] , 
        \wColumn_33[5] , \wPDiag_61[4] , \wNDiag_34[9] , \wNDiag_38[33] , 
        \wPDiag_39[60] , \wNDiag_58[37] , \wNDiag_25[48] , \wNDiag_50[61] , 
        \wPDiag_51[32] , \wPDiag_31[36] , \wNDiag_45[55] , \wColumn_58[42] , 
        \wColumn_30[6] , \wPDiag_62[7] , \wColumn_38[46] , \wPDiag_59[57] , 
        \wNDiag_38[19] , \wPDiag_39[53] , \wColumn_50[27] , \wPDiag_3[9] , 
        \wColumn_4[54] , \wPDiag_8[2] , \wColumn_25[17] , \wNDiag_8[59] , 
        \wColumn_57[1] , \wNDiag_8[40] , \wColumn_13[12] , \wPDiag_12[34] , 
        \wColumn_30[23] , \wColumn_45[13] , \wNDiag_30[56] , \wPDiag_44[35] , 
        \wColumn_54[2] , \wPDiag_24[31] , \wPDiag_24[28] , \wNDiag_25[62] , 
        \wNDiag_50[52] , \wPDiag_51[18] , \wColumn_32[59] , \wColumn_32[40] , 
        \wColumn_52[44] , \wNDiag_58[5] , \wPDiag_10[57] , \wPDiag_10[7] , 
        \wPDiag_18[18] , \wColumn_42[6] , \wNDiag_19[52] , \wNDiag_32[35] , 
        \wReturn_37[0] , \wPDiag_13[4] , \wColumn_41[5] , \wPDiag_46[56] , 
        \wNDiag_52[28] , \wPDiag_53[62] , \wColumn_19[27] , \wPDiag_26[52] , 
        \wNDiag_27[18] , \wNDiag_52[31] , \wPDiag_18[32] , \wNDiag_46[9] , 
        \wNDiag_19[61] , \wColumn_26[2] , \wScan_0[0] , \wNDiag_2[46] , 
        \wPDiag_4[36] , \wColumn_11[42] , \wScan_14[3] , \wColumn_47[43] , 
        \wScan_17[0] , \wColumn_27[47] , \wScan_3[3] , \wPDiag_6[4] , 
        \wNDiag_11[37] , \wColumn_19[14] , \wPDiag_26[61] , \wNDiag_27[32] , 
        \wPDiag_53[51] , \wNDiag_47[36] , \wPDiag_53[48] , \wPDiag_13[27] , 
        \wColumn_25[1] , \wPDiag_30[16] , \wPDiag_33[55] , \wPDiag_45[26] , 
        \wNDiag_43[4] , \wPDiag_25[22] , \wNDiag_31[45] , \wPDiag_50[12] , 
        \wNDiag_51[58] , \wNDiag_51[41] , \wColumn_59[7] , \wPDiag_16[9] , 
        \wColumn_44[8] , \wColumn_51[34] , \wColumn_59[62] , \wNDiag_1[36] , 
        \wPDiag_5[7] , \wNDiag_9[53] , \wColumn_31[29] , \wColumn_44[19] , 
        \wColumn_12[18] , \wColumn_31[30] , \wColumn_7[24] , \wNDiag_40[7] , 
        \wNDiag_59[17] , \wPDiag_58[44] , \wPDiag_7[46] , \wPDiag_38[59] , 
        \wPDiag_38[40] , \wNDiag_39[13] , \wColumn_59[51] , \wColumn_59[48] , 
        \wColumn_2[38] , \wNDiag_2[9] , \wColumn_3[26] , \wColumn_7[17] , 
        \wNDiag_12[47] , \wNDiag_24[42] , \wColumn_39[55] , \wPDiag_25[11] , 
        \wNDiag_27[0] , \wPDiag_50[38] , \wPDiag_30[25] , \wPDiag_50[21] , 
        \wPDiag_13[14] , \wPDiag_45[15] , \wNDiag_24[3] , \wNDiag_39[39] , 
        \wNDiag_44[46] , \wNDiag_39[20] , \wNDiag_59[24] , \wNDiag_9[60] , 
        \wColumn_12[32] , \wColumn_24[37] , \wColumn_44[33] , \wNDiag_28[25] , 
        \wPDiag_48[7] , \wNDiag_48[38] , \wNDiag_48[21] , \wColumn_3[15] , 
        \wNDiag_4[7] , \wColumn_8[9] , \wColumn_63[33] , \wNDiag_7[4] , 
        \wColumn_28[50] , \wColumn_35[32] , \wPDiag_55[8] , \wColumn_55[36] , 
        \wColumn_28[49] , \wColumn_16[30] , \wPDiag_17[25] , \wColumn_19[5] , 
        \wColumn_48[54] , \wNDiag_55[43] , \wPDiag_21[39] , \wPDiag_21[20] , 
        \wPDiag_54[10] , \wPDiag_34[14] , \wPDiag_41[24] , \wNDiag_63[46] , 
        \wPDiag_62[15] , \wColumn_20[35] , \wNDiag_35[47] , \wColumn_16[29] , 
        \wColumn_35[18] , \wColumn_40[28] , \wNDiag_28[16] , \wColumn_40[31] , 
        \wColumn_63[19] , \wPDiag_3[44] , \wNDiag_5[34] , \wNDiag_16[45] , 
        \wPDiag_29[45] , \wPDiag_34[27] , \wNDiag_48[12] , \wPDiag_49[41] , 
        \wPDiag_49[58] , \wPDiag_17[16] , \wPDiag_41[17] , \wNDiag_20[59] , 
        \wNDiag_20[40] , \wNDiag_40[44] , \wPDiag_62[26] , \wPDiag_21[13] , 
        \wPDiag_54[23] , \wColumn_28[63] , \wColumn_8[19] , \wPDiag_22[50] , 
        \wScan_33[6] , \wCall_35[0] , \wPDiag_53[6] , \wPDiag_57[60] , 
        \wNDiag_56[33] , \wPDiag_22[49] , \wNDiag_3[58] , \wNDiag_3[41] , 
        \wColumn_5[60] , \wColumn_5[53] , \wNDiag_6[44] , \wColumn_8[33] , 
        \wPDiag_8[51] , \wPDiag_14[55] , \wNDiag_36[37] , \wNDiag_18[7] , 
        \wPDiag_42[54] , \wNDiag_60[36] , \wPDiag_50[5] , \wScan_30[5] , 
        \wColumn_36[42] , \wColumn_60[43] , \wPDiag_8[48] , \wColumn_56[46] , 
        \wNDiag_15[35] , \wNDiag_43[34] , \wPDiag_61[56] , \wPDiag_22[63] , 
        \wNDiag_23[29] , \wPDiag_37[57] , \wPDiag_37[2] , \wNDiag_56[19] , 
        \wPDiag_57[53] , \wNDiag_23[30] , \wScan_8[5] , \wPDiag_8[62] , 
        \wScan_57[2] , \wColumn_15[59] , \wColumn_23[45] , \wColumn_15[40] , 
        \wColumn_43[41] , \wScan_54[1] , \wPDiag_34[1] , \wColumn_43[58] , 
        \wColumn_53[43] , \wScan_60[0] , \wColumn_33[47] , \wNDiag_48[2] , 
        \wPDiag_11[50] , \wNDiag_18[55] , \wColumn_52[1] , \wNDiag_33[32] , 
        \wPDiag_47[48] , \wPDiag_11[49] , \wPDiag_32[61] , \wPDiag_47[51] , 
        \wColumn_18[39] , \wPDiag_27[55] , \wColumn_51[2] , \wNDiag_53[36] , 
        \wColumn_18[20] , \wScan_63[3] , \wPDiag_19[35] , \wColumn_36[5] , 
        \wReturn_40[0] , \wPDiag_5[31] , \wColumn_10[45] , \wColumn_46[44] , 
        \wColumn_26[59] , \wNDiag_31[9] , \wColumn_26[40] , \wPDiag_5[28] , 
        \wReturn_5[0] , \wNDiag_10[30] , \wNDiag_10[29] , \wPDiag_11[63] , 
        \wColumn_18[13] , \wColumn_28[9] , \wNDiag_26[35] , \wPDiag_52[56] , 
        \wNDiag_46[31] , \wPDiag_12[39] , \wPDiag_32[52] , \wNDiag_33[18] , 
        \wColumn_35[6] , \wPDiag_44[21] , \wNDiag_46[28] , \wPDiag_47[62] , 
        \wPDiag_12[20] , \wPDiag_31[11] , \wPDiag_44[38] , \wNDiag_53[3] , 
        \wPDiag_24[25] , \wNDiag_30[42] , \wColumn_49[0] , \wNDiag_50[46] , 
        \wPDiag_51[15] , \wColumn_38[61] , \wColumn_50[33] , \wColumn_5[1] , 
        \wColumn_6[23] , \wNDiag_8[54] , \wColumn_30[37] , \wNDiag_50[0] , 
        \wNDiag_58[10] , \wPDiag_59[43] , \wColumn_6[10] , \wPDiag_6[58] , 
        \wPDiag_18[2] , \wPDiag_39[47] , \wNDiag_38[14] , \wColumn_58[56] , 
        \wPDiag_6[41] , \wPDiag_12[13] , \wNDiag_13[40] , \wPDiag_24[16] , 
        \wNDiag_25[45] , \wColumn_38[52] , \wNDiag_37[7] , \wPDiag_31[22] , 
        \wPDiag_51[26] , \wPDiag_44[12] , \wNDiag_45[58] , \wNDiag_13[59] , 
        \wNDiag_34[4] , \wNDiag_45[41] , \wNDiag_38[27] , \wNDiag_58[23] , 
        \wColumn_13[35] , \wColumn_25[30] , \wColumn_45[34] , \wColumn_25[29] , 
        \wColumn_33[8] , \wPDiag_61[9] , \wColumn_50[19] , \wNDiag_10[2] , 
        \wNDiag_29[22] , \wNDiag_49[26] , \wPDiag_58[0] , \wColumn_2[21] , 
        \wColumn_2[12] , \wNDiag_4[19] , \wColumn_21[18] , \wColumn_34[35] , 
        \wColumn_62[34] , \wScan_38[0] , \wColumn_54[31] , \wColumn_54[28] , 
        \wColumn_29[57] , \wColumn_6[2] , \wPDiag_20[27] , \wColumn_49[53] , 
        \wNDiag_54[44] , \wPDiag_55[17] , \wNDiag_13[1] , \wNDiag_34[59] , 
        \wPDiag_35[13] , \wPDiag_40[23] , \wNDiag_62[41] , \wNDiag_62[58] , 
        \wPDiag_63[12] , \wPDiag_16[22] , \wColumn_17[37] , \wColumn_21[32] , 
        \wNDiag_34[40] , \wNDiag_29[11] , \wColumn_41[36] , \wPDiag_16[11] , 
        \wNDiag_17[42] , \wReturn_18[0] , \wPDiag_28[42] , \wPDiag_48[46] , 
        \wPDiag_35[20] , \wNDiag_49[15] , \wPDiag_35[39] , \wPDiag_40[10] , 
        \wPDiag_63[38] , \wNDiag_21[47] , \wNDiag_41[43] , \wPDiag_63[21] , 
        \wScan_0[4] , \wColumn_1[62] , \wColumn_1[51] , \wPDiag_1[19] , 
        \wPDiag_2[43] , \wNDiag_4[33] , \wPDiag_20[14] , \wPDiag_55[24] , 
        \wPDiag_22[8] , \wColumn_49[60] , \wColumn_11[0] , \wScan_23[1] , 
        \wColumn_12[3] , \wNDiag_14[18] , \wPDiag_23[57] , \wPDiag_43[1] , 
        \wNDiag_37[30] , \wNDiag_57[34] , \wPDiag_60[62] , \wNDiag_61[28] , 
        \wPDiag_15[52] , \wPDiag_36[63] , \wNDiag_42[19] , \wNDiag_61[31] , 
        \wPDiag_43[53] , \wNDiag_37[29] , \wPDiag_40[2] , \wColumn_1[48] , 
        \wPDiag_1[33] , \wNDiag_7[43] , \wColumn_9[34] , \wPDiag_9[56] , 
        \wScan_20[2] , \wColumn_37[45] , \wColumn_57[58] , \wColumn_61[44] , 
        \wNDiag_14[32] , \wPDiag_15[61] , \wColumn_57[41] , \wPDiag_36[49] , 
        \wNDiag_42[33] , \wPDiag_60[51] , \wPDiag_27[5] , \wPDiag_36[50] , 
        \wPDiag_43[60] , \wPDiag_56[54] , \wPDiag_60[48] , \wNDiag_22[37] , 
        \wScan_47[5] , \wColumn_14[47] , \wColumn_22[42] , \wPDiag_39[9] , 
        \wColumn_42[46] , \wScan_44[6] , \wPDiag_24[6] , \wNDiag_1[22] , 
        \wNDiag_1[7] , \wColumn_3[32] , \wColumn_3[18] , \wPDiag_3[50] , 
        \wPDiag_3[49] , \wNDiag_5[39] , \wPDiag_32[2] , \wCall_42[0] , 
        \wNDiag_5[20] , \wColumn_60[3] , \wNDiag_16[51] , \wNDiag_16[48] , 
        \wPDiag_34[33] , \wNDiag_40[49] , \wNDiag_63[61] , \wNDiag_20[54] , 
        \wNDiag_35[60] , \wNDiag_40[50] , \wPDiag_62[32] , \wScan_52[2] , 
        \wPDiag_54[37] , \wPDiag_3[63] , \wNDiag_7[9] , \wColumn_16[24] , 
        \wColumn_20[38] , \wColumn_20[21] , \wPDiag_29[51] , \wPDiag_29[48] , 
        \wPDiag_49[55] , \wScan_51[1] , \wColumn_55[11] , \wPDiag_31[1] , 
        \wColumn_63[0] , \wNDiag_16[62] , \wPDiag_17[28] , \wColumn_19[8] , 
        \wColumn_35[15] , \wColumn_63[14] , \wColumn_40[25] , \wNDiag_55[57] , 
        \wPDiag_21[34] , \wScan_36[6] , \wPDiag_62[18] , \wNDiag_63[52] , 
        \wPDiag_41[30] , \wPDiag_17[31] , \wPDiag_34[19] , \wNDiag_35[53] , 
        \wNDiag_40[63] , \wPDiag_41[29] , \wColumn_28[44] , \wNDiag_5[13] , 
        \wCall_30[0] , \wPDiag_56[6] , \wColumn_48[59] , \wColumn_8[4] , 
        \wColumn_16[17] , \wColumn_48[40] , \wPDiag_55[5] , \wColumn_63[27] , 
        \wColumn_35[26] , \wColumn_40[16] , \wColumn_20[12] , \wColumn_55[22] , 
        \wNDiag_28[31] , \wNDiag_48[35] , \wNDiag_28[28] , \wPDiag_29[62] , 
        \wScan_35[5] , \wNDiag_6[50] , \wColumn_15[54] , \wColumn_23[51] , 
        \wColumn_23[48] , \wScan_49[3] , \wPDiag_29[3] , \wColumn_43[55] , 
        \wColumn_56[61] , \wNDiag_61[1] , \wNDiag_6[49] , \wColumn_8[27] , 
        \wNDiag_15[38] , \wNDiag_36[10] , \wNDiag_62[2] , \wNDiag_15[21] , 
        \wPDiag_37[43] , \wNDiag_43[20] , \wPDiag_61[42] , \wNDiag_43[39] , 
        \wNDiag_60[11] , \wPDiag_57[47] , \wPDiag_8[45] , \wNDiag_23[24] , 
        \wColumn_36[56] , \wNDiag_56[14] , \wColumn_60[57] , \wColumn_23[62] , 
        \wColumn_56[52] , \wPDiag_50[8] , \wNDiag_2[61] , \wNDiag_2[52] , 
        \wNDiag_2[4] , \wColumn_8[14] , \wPDiag_22[44] , \wPDiag_4[22] , 
        \wNDiag_6[63] , \wPDiag_14[58] , \wPDiag_14[41] , \wNDiag_23[17] , 
        \wNDiag_56[27] , \wPDiag_42[59] , \wNDiag_43[13] , \wNDiag_36[23] , 
        \wPDiag_42[40] , \wNDiag_60[22] , \wNDiag_15[12] , \wNDiag_11[23] , 
        \wNDiag_27[26] , \wPDiag_53[45] , \wNDiag_32[12] , \wPDiag_33[58] , 
        \wNDiag_52[16] , \wPDiag_33[41] , \wNDiag_47[22] , \wNDiag_22[0] , 
        \wPDiag_3[4] , \wColumn_11[56] , \wColumn_19[19] , \wColumn_38[3] , 
        \wNDiag_21[3] , \wColumn_47[57] , \wPDiag_18[26] , \wColumn_27[53] , 
        \wColumn_52[63] , \wColumn_4[59] , \wColumn_4[40] , \wPDiag_4[11] , 
        \wColumn_19[33] , \wNDiag_46[4] , \wScan_5[0] , \wScan_6[3] , 
        \wPDiag_10[43] , \wNDiag_47[11] , \wNDiag_32[21] , \wNDiag_11[10] , 
        \wPDiag_46[42] , \wPDiag_13[9] , \wPDiag_26[46] , \wNDiag_32[38] , 
        \wNDiag_27[15] , \wColumn_41[8] , \wNDiag_52[25] , \wNDiag_58[8] , 
        \wPDiag_7[52] , \wScan_11[3] , \wColumn_12[26] , \wPDiag_18[15] , 
        \wNDiag_19[46] , \wColumn_27[60] , \wNDiag_45[7] , \wColumn_52[50] , 
        \wColumn_52[49] , \wColumn_32[54] , \wColumn_23[2] , \wColumn_24[23] , 
        \wColumn_31[17] , \wNDiag_39[1] , \wColumn_44[27] , \wColumn_51[13] , 
        \wScan_12[0] , \wNDiag_24[56] , \wNDiag_39[34] , \wPDiag_58[63] , 
        \wNDiag_59[30] , \wNDiag_59[29] , \wNDiag_12[53] , \wPDiag_50[35] , 
        \wPDiag_13[19] , \wPDiag_30[31] , \wPDiag_30[28] , \wNDiag_31[62] , 
        \wNDiag_44[52] , \wPDiag_45[18] , \wColumn_59[45] , \wColumn_20[1] , 
        \wColumn_39[58] , \wNDiag_1[11] , \wColumn_7[30] , \wColumn_7[29] , 
        \wColumn_39[41] , \wPDiag_58[49] , \wPDiag_58[50] , \wNDiag_9[47] , 
        \wColumn_12[15] , \wPDiag_15[7] , \wColumn_24[10] , \wPDiag_38[54] , 
        \wColumn_51[20] , \wColumn_47[6] , \wColumn_51[39] , \wColumn_31[24] , 
        \wColumn_44[14] , \wReturn_32[0] , \wColumn_3[22] , \wNDiag_4[3] , 
        \wPDiag_6[9] , \wPDiag_7[61] , \wPDiag_16[4] , \wColumn_44[5] , 
        \wNDiag_31[48] , \wNDiag_43[9] , \wPDiag_45[32] , \wNDiag_6[59] , 
        \wPDiag_8[55] , \wNDiag_12[60] , \wPDiag_13[33] , \wNDiag_31[51] , 
        \wNDiag_44[61] , \wPDiag_25[36] , \wNDiag_51[55] , \wScan_30[1] , 
        \wColumn_56[42] , \wPDiag_14[51] , \wPDiag_14[48] , \wNDiag_18[3] , 
        \wColumn_36[46] , \wColumn_60[47] , \wPDiag_37[60] , \wPDiag_42[50] , 
        \wPDiag_50[1] , \wNDiag_60[32] , \wNDiag_36[33] , \wPDiag_42[49] , 
        \wPDiag_61[61] , \wColumn_15[44] , \wPDiag_22[54] , \wPDiag_53[2] , 
        \wNDiag_56[37] , \wScan_33[2] , \wPDiag_34[5] , \wScan_54[5] , 
        \wColumn_23[58] , \wColumn_23[41] , \wColumn_43[45] , \wNDiag_61[8] , 
        \wScan_57[6] , \wNDiag_6[40] , \wNDiag_7[0] , \wColumn_8[37] , 
        \wNDiag_23[34] , \wPDiag_57[57] , \wPDiag_14[62] , \wNDiag_15[31] , 
        \wNDiag_15[28] , \wNDiag_36[19] , \wPDiag_37[53] , \wPDiag_37[6] , 
        \wPDiag_42[63] , \wNDiag_43[29] , \wCall_51[0] , \wPDiag_17[38] , 
        \wPDiag_17[21] , \wPDiag_41[39] , \wNDiag_43[30] , \wNDiag_60[18] , 
        \wPDiag_61[52] , \wPDiag_62[11] , \wNDiag_35[43] , \wPDiag_41[20] , 
        \wNDiag_63[42] , \wColumn_19[1] , \wPDiag_21[24] , \wPDiag_34[10] , 
        \wPDiag_54[14] , \wNDiag_55[47] , \wColumn_48[50] , \wColumn_48[49] , 
        \wScan_28[3] , \wColumn_28[54] , \wColumn_55[32] , \wColumn_35[36] , 
        \wColumn_63[37] , \wNDiag_28[38] , \wColumn_3[11] , \wPDiag_3[59] , 
        \wPDiag_3[40] , \wNDiag_28[21] , \wPDiag_48[3] , \wNDiag_48[25] , 
        \wNDiag_5[30] , \wNDiag_5[29] , \wColumn_48[63] , \wNDiag_16[58] , 
        \wNDiag_20[44] , \wPDiag_21[17] , \wPDiag_54[27] , \wNDiag_16[41] , 
        \wPDiag_17[12] , \wPDiag_34[23] , \wNDiag_40[40] , \wPDiag_62[22] , 
        \wNDiag_40[59] , \wPDiag_41[13] , \wNDiag_48[16] , \wPDiag_49[45] , 
        \wPDiag_5[3] , \wColumn_7[20] , \wColumn_16[34] , \wNDiag_28[12] , 
        \wPDiag_29[41] , \wPDiag_29[58] , \wColumn_40[35] , \wColumn_20[31] , 
        \wColumn_20[28] , \wColumn_55[18] , \wPDiag_31[8] , \wColumn_63[9] , 
        \wPDiag_38[44] , \wNDiag_39[17] , \wPDiag_58[40] , \wColumn_7[39] , 
        \wPDiag_58[59] , \wNDiag_59[13] , \wNDiag_9[57] , \wNDiag_40[3] , 
        \wColumn_31[34] , \wNDiag_1[32] , \wNDiag_1[18] , \wColumn_24[19] , 
        \wColumn_51[29] , \wColumn_39[62] , \wColumn_51[30] , \wPDiag_6[0] , 
        \wPDiag_13[23] , \wPDiag_25[26] , \wPDiag_50[16] , \wNDiag_43[0] , 
        \wNDiag_51[45] , \wColumn_59[3] , \wColumn_7[13] , \wColumn_12[36] , 
        \wColumn_24[33] , \wPDiag_30[12] , \wNDiag_31[58] , \wNDiag_31[41] , 
        \wPDiag_45[22] , \wNDiag_39[8] , \wColumn_44[37] , \wNDiag_59[39] , 
        \wNDiag_12[43] , \wPDiag_13[10] , \wNDiag_24[7] , \wNDiag_59[20] , 
        \wPDiag_30[38] , \wNDiag_39[24] , \wPDiag_30[21] , \wNDiag_44[42] , 
        \wNDiag_24[46] , \wPDiag_25[15] , \wPDiag_45[11] , \wPDiag_50[25] , 
        \wNDiag_27[4] , \wNDiag_2[42] , \wColumn_4[50] , \wColumn_4[49] , 
        \wPDiag_4[18] , \wPDiag_7[42] , \wColumn_20[8] , \wColumn_39[51] , 
        \wColumn_39[48] , \wColumn_59[55] , \wPDiag_10[53] , \wPDiag_13[0] , 
        \wColumn_19[23] , \wColumn_41[1] , \wNDiag_52[35] , \wPDiag_26[56] , 
        \wNDiag_32[31] , \wNDiag_32[28] , \wPDiag_46[52] , \wNDiag_47[18] , 
        \wPDiag_33[62] , \wPDiag_10[3] , \wNDiag_11[19] , \wNDiag_19[56] , 
        \wColumn_42[2] , \wNDiag_58[1] , \wPDiag_10[60] , \wNDiag_11[33] , 
        \wColumn_32[44] , \wColumn_52[59] , \wColumn_52[40] , \wColumn_25[5] , 
        \wPDiag_33[51] , \wPDiag_46[61] , \wColumn_19[10] , \wNDiag_27[36] , 
        \wPDiag_33[48] , \wNDiag_47[32] , \wReturn_53[0] , \wPDiag_53[55] , 
        \wPDiag_4[32] , \wScan_17[4] , \wColumn_11[46] , \wNDiag_22[9] , 
        \wColumn_27[43] , \wColumn_4[63] , \wColumn_26[6] , \wColumn_47[47] , 
        \wColumn_6[19] , \wPDiag_6[51] , \wPDiag_18[36] , \wColumn_30[2] , 
        \wColumn_38[42] , \wPDiag_62[3] , \wPDiag_6[48] , \wColumn_58[46] , 
        \wNDiag_13[50] , \wNDiag_13[49] , \wNDiag_30[61] , \wNDiag_45[51] , 
        \wNDiag_25[55] , \wPDiag_31[32] , \wNDiag_45[48] , \wPDiag_51[36] , 
        \wNDiag_58[33] , \wPDiag_59[60] , \wColumn_25[39] , \wNDiag_38[37] , 
        \wColumn_25[20] , \wColumn_33[1] , \wPDiag_61[0] , \wColumn_50[10] , 
        \wPDiag_6[62] , \wPDiag_12[30] , \wColumn_13[25] , \wColumn_30[14] , 
        \wColumn_45[24] , \wPDiag_24[35] , \wNDiag_29[2] , \wColumn_49[9] , 
        \wNDiag_30[52] , \wPDiag_31[18] , \wPDiag_44[28] , \wNDiag_45[62] , 
        \wNDiag_50[56] , \wPDiag_12[29] , \wNDiag_13[63] , \wPDiag_44[31] , 
        \wPDiag_8[6] , \wNDiag_8[44] , \wColumn_54[6] , \wColumn_13[16] , 
        \wColumn_30[27] , \wColumn_45[17] , \wColumn_57[5] , \wColumn_50[23] , 
        \wColumn_1[58] , \wPDiag_1[23] , \wNDiag_3[62] , \wNDiag_3[51] , 
        \wNDiag_3[48] , \wColumn_6[33] , \wReturn_21[0] , \wColumn_25[13] , 
        \wPDiag_39[57] , \wNDiag_50[9] , \wNDiag_58[19] , \wPDiag_59[53] , 
        \wColumn_10[55] , \wScan_19[2] , \wPDiag_19[25] , \wColumn_26[50] , 
        \wColumn_26[49] , \wColumn_53[60] , \wNDiag_31[0] , \wColumn_46[54] , 
        \wColumn_5[43] , \wPDiag_5[38] , \wColumn_28[0] , \wNDiag_32[3] , 
        \wPDiag_5[21] , \wNDiag_10[39] , \wNDiag_10[20] , \wPDiag_32[42] , 
        \wNDiag_33[11] , \wNDiag_46[38] , \wNDiag_18[45] , \wColumn_26[63] , 
        \wNDiag_26[25] , \wNDiag_46[21] , \wColumn_33[57] , \wPDiag_52[46] , 
        \wNDiag_53[15] , \wColumn_53[53] , \wNDiag_55[4] , \wPDiag_19[16] , 
        \wColumn_52[8] , \wPDiag_5[12] , \wNDiag_10[13] , \wNDiag_26[16] , 
        \wNDiag_53[26] , \wPDiag_27[45] , \wPDiag_47[41] , \wPDiag_11[59] , 
        \wPDiag_11[40] , \wNDiag_46[12] , \wPDiag_47[58] , \wNDiag_33[22] , 
        \wColumn_18[30] , \wColumn_18[29] , \wColumn_9[24] , \wNDiag_22[27] , 
        \wNDiag_56[7] , \wPDiag_56[44] , \wNDiag_57[17] , \wNDiag_14[22] , 
        \wPDiag_36[40] , \wPDiag_36[59] , \wNDiag_37[13] , \wPDiag_60[58] , 
        \wNDiag_61[12] , \wNDiag_42[23] , \wPDiag_60[41] , \wPDiag_1[10] , 
        \wNDiag_7[60] , \wNDiag_7[53] , \wColumn_14[57] , \wColumn_22[52] , 
        \wColumn_42[56] , \wPDiag_39[0] , \wColumn_57[62] , \wScan_59[0] , 
        \wNDiag_16[5] , \wColumn_3[6] , \wColumn_9[17] , \wColumn_11[9] , 
        \wNDiag_14[11] , \wPDiag_43[43] , \wNDiag_61[21] , \wPDiag_15[42] , 
        \wNDiag_37[39] , \wNDiag_42[10] , \wNDiag_61[38] , \wNDiag_37[20] , 
        \wPDiag_43[8] , \wNDiag_57[24] , \wNDiag_22[14] , \wPDiag_23[47] , 
        \wColumn_1[41] , \wColumn_1[8] , \wColumn_2[31] , \wPDiag_2[53] , 
        \wPDiag_9[46] , \wNDiag_15[6] , \wColumn_22[61] , \wColumn_57[51] , 
        \wColumn_57[48] , \wPDiag_16[18] , \wColumn_17[27] , \wColumn_34[16] , 
        \wColumn_37[55] , \wColumn_61[54] , \wColumn_41[26] , \wColumn_21[22] , 
        \wPDiag_21[2] , \wColumn_62[17] , \wNDiag_21[57] , \wPDiag_28[52] , 
        \wScan_41[2] , \wPDiag_48[56] , \wColumn_54[12] , \wNDiag_29[18] , 
        \wScan_42[1] , \wPDiag_55[34] , \wNDiag_34[63] , \wPDiag_35[29] , 
        \wPDiag_40[19] , \wNDiag_41[53] , \wPDiag_63[31] , \wNDiag_17[52] , 
        \wPDiag_35[30] , \wNDiag_62[62] , \wPDiag_63[28] , \wNDiag_4[23] , 
        \wPDiag_22[1] , \wScan_25[6] , \wPDiag_28[61] , \wColumn_2[28] , 
        \wNDiag_29[32] , \wPDiag_2[60] , \wNDiag_4[10] , \wColumn_5[8] , 
        \wNDiag_9[6] , \wColumn_17[14] , \wColumn_17[7] , \wColumn_21[11] , 
        \wNDiag_49[36] , \wColumn_54[38] , \wPDiag_58[9] , \wColumn_54[21] , 
        \wColumn_34[25] , \wColumn_41[15] , \wCall_23[0] , \wPDiag_45[6] , 
        \wColumn_62[24] , \wColumn_49[43] , \wNDiag_2[27] , \wNDiag_2[14] , 
        \wPDiag_10[36] , \wNDiag_13[8] , \wColumn_14[4] , \wPDiag_16[32] , 
        \wColumn_29[47] , \wPDiag_46[5] , \wNDiag_34[50] , \wNDiag_41[60] , 
        \wNDiag_62[48] , \wScan_26[5] , \wPDiag_40[33] , \wNDiag_62[51] , 
        \wNDiag_17[61] , \wNDiag_34[49] , \wPDiag_20[37] , \wNDiag_54[54] , 
        \wPDiag_26[33] , \wNDiag_32[54] , \wScan_46[1] , \wPDiag_46[37] , 
        \wNDiag_52[49] , \wNDiag_27[60] , \wNDiag_52[50] , \wColumn_4[35] , 
        \wColumn_11[10] , \wColumn_19[46] , \wPDiag_25[2] , \wPDiag_26[1] , 
        \wColumn_27[15] , \wColumn_52[25] , \wColumn_32[21] , \wColumn_47[11] , 
        \wColumn_32[38] , \wScan_45[2] , \wPDiag_4[57] , \wPDiag_18[60] , 
        \wNDiag_19[33] , \wColumn_10[4] , \wNDiag_11[56] , \wNDiag_17[8] , 
        \wScan_22[5] , \wPDiag_42[5] , \wPDiag_26[19] , \wPDiag_53[30] , 
        \wNDiag_27[53] , \wPDiag_33[34] , \wNDiag_47[57] , \wNDiag_52[63] , 
        \wPDiag_53[29] , \wPDiag_18[53] , \wNDiag_19[19] , \wScan_21[6] , 
        \wNDiag_1[57] , \wColumn_4[5] , \wColumn_7[45] , \wNDiag_9[32] , 
        \wColumn_11[23] , \wColumn_32[12] , \wColumn_47[22] , \wColumn_12[60] , 
        \wColumn_13[7] , \wCall_27[0] , \wPDiag_41[6] , \wColumn_27[26] , 
        \wColumn_51[55] , \wColumn_52[16] , \wColumn_31[48] , \wColumn_44[61] , 
        \wColumn_31[51] , \wPDiag_7[14] , \wNDiag_12[15] , \wPDiag_38[38] , 
        \wPDiag_38[21] , \wPDiag_58[25] , \wPDiag_45[47] , \wPDiag_13[46] , 
        \wNDiag_31[24] , \wNDiag_44[14] , \wNDiag_24[10] , \wNDiag_51[20] , 
        \wPDiag_25[43] , \wNDiag_51[39] , \wNDiag_9[18] , \wColumn_12[53] , 
        \wPDiag_38[12] , \wNDiag_39[58] , \wScan_39[4] , \wNDiag_39[41] , 
        \wPDiag_58[16] , \wNDiag_59[45] , \wNDiag_11[6] , \wColumn_31[62] , 
        \wColumn_44[52] , \wColumn_24[56] , \wPDiag_59[4] , \wColumn_7[6] , 
        \wPDiag_7[27] , \wNDiag_12[5] , \wColumn_59[30] , \wColumn_59[29] , 
        \wColumn_3[47] , \wPDiag_3[16] , \wNDiag_12[26] , \wNDiag_24[23] , 
        \wColumn_39[34] , \wPDiag_50[59] , \wNDiag_51[13] , \wPDiag_50[40] , 
        \wColumn_15[9] , \wPDiag_30[44] , \wNDiag_31[17] , \wPDiag_47[8] , 
        \wColumn_28[31] , \wNDiag_44[27] , \wColumn_28[28] , \wNDiag_16[17] , 
        \wNDiag_20[12] , \wNDiag_36[3] , \wColumn_48[35] , \wNDiag_55[22] , 
        \wPDiag_21[58] , \wPDiag_21[41] , \wPDiag_41[45] , \wNDiag_63[27] , 
        \wPDiag_17[44] , \wNDiag_35[26] , \wNDiag_40[16] , \wNDiag_28[44] , 
        \wNDiag_48[59] , \wNDiag_48[40] , \wPDiag_49[13] , \wPDiag_29[17] , 
        \wPDiag_3[25] , \wNDiag_5[55] , \wColumn_16[62] , \wColumn_63[52] , 
        \wNDiag_16[24] , \wColumn_35[53] , \wColumn_40[63] , \wNDiag_35[0] , 
        \wColumn_55[57] , \wNDiag_20[38] , \wNDiag_20[21] , \wPDiag_34[46] , 
        \wNDiag_35[15] , \wNDiag_63[14] , \wNDiag_40[25] , \wPDiag_62[47] , 
        \wNDiag_55[11] , \wColumn_48[4] , \wPDiag_54[42] , \wNDiag_52[7] , 
        \wNDiag_6[16] , \wPDiag_8[30] , \wColumn_15[12] , \wColumn_16[51] , 
        \wPDiag_19[6] , \wColumn_20[54] , \wColumn_16[48] , \wColumn_35[60] , 
        \wColumn_40[49] , \wColumn_63[61] , \wPDiag_29[24] , \wColumn_40[50] , 
        \wNDiag_51[4] , \wColumn_56[8] , \wColumn_36[23] , \wColumn_43[13] , 
        \wPDiag_49[39] , \wPDiag_49[20] , \wColumn_37[1] , \wColumn_60[22] , 
        \wPDiag_8[29] , \wColumn_56[27] , \wColumn_23[17] , \wColumn_34[2] , 
        \wColumn_8[61] , \wScan_9[1] , \wPDiag_14[34] , \wPDiag_22[31] , 
        \wPDiag_22[28] , \wNDiag_23[62] , \wNDiag_56[52] , \wPDiag_57[18] , 
        \wColumn_15[38] , \wColumn_23[24] , \wNDiag_36[56] , \wPDiag_42[35] , 
        \wColumn_53[5] , \wNDiag_60[57] , \wColumn_56[14] , \wColumn_15[21] , 
        \wReturn_25[0] , \wColumn_36[10] , \wColumn_43[20] , \wColumn_43[39] , 
        \wNDiag_49[6] , \wColumn_60[11] , \wScan_61[4] , \wColumn_1[17] , 
        \wPDiag_1[46] , \wColumn_2[54] , \wPDiag_2[36] , \wNDiag_4[46] , 
        \wNDiag_6[25] , \wColumn_8[52] , \wNDiag_15[54] , \wPDiag_37[36] , 
        \wNDiag_43[55] , \wNDiag_54[9] , \wPDiag_61[37] , \wNDiag_23[48] , 
        \wNDiag_23[51] , \wPDiag_57[32] , \wNDiag_56[61] , \wPDiag_14[3] , 
        \wColumn_46[2] , \wColumn_50[6] , \wColumn_17[42] , \wColumn_21[47] , 
        \wPDiag_28[37] , \wPDiag_48[33] , \wNDiag_49[60] , \wColumn_41[43] , 
        \wColumn_49[15] , \wColumn_29[11] , \wPDiag_17[0] , \wPDiag_35[55] , 
        \wColumn_45[1] , \wNDiag_17[37] , \wPDiag_20[61] , \wNDiag_21[32] , 
        \wNDiag_41[36] , \wPDiag_63[54] , \wPDiag_55[48] , \wColumn_22[6] , 
        \wColumn_34[59] , \wPDiag_55[51] , \wColumn_62[41] , \wColumn_34[40] , 
        \wColumn_62[58] , \wColumn_54[44] , \wNDiag_29[57] , \wPDiag_48[19] , 
        \wNDiag_49[53] , \wNDiag_7[36] , \wScan_13[4] , \wPDiag_16[57] , 
        \wPDiag_20[52] , \wColumn_21[5] , \wNDiag_38[5] , \wNDiag_54[31] , 
        \wNDiag_54[28] , \wPDiag_55[62] , \wNDiag_21[18] , \wPDiag_40[56] , 
        \wNDiag_62[34] , \wColumn_29[22] , \wNDiag_34[35] , \wReturn_57[0] , 
        \wNDiag_26[9] , \wColumn_49[26] , \wPDiag_2[0] , \wColumn_9[58] , 
        \wColumn_9[41] , \wNDiag_14[47] , \wPDiag_15[14] , \wNDiag_42[46] , 
        \wPDiag_60[24] , \wPDiag_23[11] , \wPDiag_36[25] , \wPDiag_43[15] , 
        \wNDiag_22[42] , \wPDiag_56[21] , \wNDiag_47[0] , \wPDiag_56[38] , 
        \wPDiag_1[3] , \wScan_4[4] , \wPDiag_9[10] , \wNDiag_44[3] , 
        \wColumn_22[37] , \wColumn_42[33] , \wColumn_14[32] , \wPDiag_15[27] , 
        \wPDiag_23[22] , \wPDiag_56[12] , \wNDiag_57[58] , \wNDiag_37[45] , 
        \wColumn_39[7] , \wNDiag_57[41] , \wPDiag_60[17] , \wNDiag_23[4] , 
        \wColumn_24[8] , \wPDiag_36[16] , \wPDiag_43[26] , \wNDiag_61[44] , 
        \wColumn_1[24] , \wPDiag_9[23] , \wColumn_14[18] , \wColumn_61[28] , 
        \wColumn_37[30] , \wColumn_37[29] , \wColumn_42[19] , \wColumn_61[31] , 
        \wColumn_57[34] , \wColumn_10[30] , \wColumn_10[29] , \wNDiag_20[7] , 
        \wColumn_33[18] , \wColumn_46[31] , \wColumn_26[35] , \wColumn_46[28] , 
        \wNDiag_3[34] , \wColumn_5[15] , \wNDiag_18[13] , \wPDiag_19[40] , 
        \wPDiag_19[59] , \wPDiag_5[44] , \wNDiag_10[45] , \wPDiag_11[16] , 
        \wNDiag_26[59] , \wNDiag_26[40] , \wPDiag_27[13] , \wPDiag_52[23] , 
        \wNDiag_46[44] , \wPDiag_32[27] , \wPDiag_47[17] , \wNDiag_3[0] , 
        \wColumn_5[26] , \wNDiag_18[39] , \wNDiag_60[5] , \wNDiag_18[20] , 
        \wPDiag_28[7] , \wScan_1[0] , \wColumn_1[34] , \wColumn_6[56] , 
        \wPDiag_6[34] , \wCall_9[0] , \wPDiag_11[25] , \wColumn_18[55] , 
        \wColumn_33[32] , \wPDiag_35[8] , \wColumn_53[36] , \wNDiag_33[47] , 
        \wNDiag_13[35] , \wPDiag_24[63] , \wNDiag_25[30] , \wPDiag_27[39] , 
        \wPDiag_27[20] , \wPDiag_32[14] , \wPDiag_47[24] , \wNDiag_63[6] , 
        \wPDiag_52[10] , \wNDiag_53[43] , \wNDiag_25[29] , \wPDiag_31[57] , 
        \wNDiag_50[19] , \wPDiag_51[53] , \wPDiag_57[2] , \wScan_37[2] , 
        \wNDiag_45[34] , \wColumn_58[23] , \wNDiag_8[12] , \wColumn_13[59] , 
        \wColumn_13[40] , \wColumn_38[27] , \wScan_34[1] , \wColumn_45[58] , 
        \wColumn_45[41] , \wColumn_9[0] , \wColumn_25[45] , \wNDiag_38[52] , 
        \wPDiag_39[18] , \wNDiag_58[56] , \wPDiag_12[55] , \wColumn_38[14] , 
        \wScan_53[6] , \wPDiag_54[1] , \wPDiag_44[54] , \wColumn_58[10] , 
        \wPDiag_24[50] , \wPDiag_24[49] , \wNDiag_30[37] , \wNDiag_50[33] , 
        \wPDiag_33[6] , \wPDiag_51[60] , \wColumn_61[7] , \wCall_55[0] , 
        \wNDiag_7[15] , \wNDiag_8[38] , \wPDiag_30[5] , \wPDiag_59[36] , 
        \wNDiag_38[61] , \wPDiag_39[32] , \wColumn_62[4] , \wScan_50[5] , 
        \wColumn_50[46] , \wNDiag_8[21] , \wColumn_9[62] , \wPDiag_15[37] , 
        \wScan_16[0] , \wColumn_30[42] , \wPDiag_43[36] , \wNDiag_61[54] , 
        \wNDiag_22[61] , \wNDiag_37[55] , \wNDiag_57[51] , \wPDiag_23[32] , 
        \wNDiag_57[48] , \wPDiag_9[33] , \wColumn_22[14] , \wColumn_24[1] , 
        \wColumn_57[24] , \wColumn_14[11] , \wColumn_27[2] , \wColumn_61[21] , 
        \wColumn_37[39] , \wScan_15[3] , \wColumn_37[20] , \wColumn_42[10] , 
        \wColumn_61[38] , \wPDiag_1[56] , \wReturn_36[0] , \wColumn_2[44] , 
        \wPDiag_2[9] , \wNDiag_7[26] , \wPDiag_12[4] , \wColumn_40[5] , 
        \wColumn_9[51] , \wColumn_9[48] , \wNDiag_22[52] , \wPDiag_23[18] , 
        \wNDiag_47[9] , \wPDiag_56[28] , \wNDiag_57[62] , \wPDiag_56[31] , 
        \wPDiag_9[19] , \wColumn_14[22] , \wNDiag_14[57] , \wPDiag_36[35] , 
        \wNDiag_42[56] , \wPDiag_60[34] , \wColumn_22[27] , \wColumn_37[13] , 
        \wNDiag_59[5] , \wColumn_61[12] , \wColumn_42[23] , \wPDiag_11[7] , 
        \wColumn_43[6] , \wColumn_57[17] , \wColumn_17[61] , \wNDiag_25[3] , 
        \wColumn_54[54] , \wColumn_34[50] , \wColumn_41[60] , \wColumn_62[48] , 
        \wColumn_62[51] , \wPDiag_28[14] , \wColumn_34[49] , \wPDiag_2[15] , 
        \wPDiag_16[47] , \wNDiag_29[47] , \wNDiag_34[25] , \wNDiag_41[15] , 
        \wPDiag_48[10] , \wNDiag_49[43] , \wNDiag_17[14] , \wPDiag_40[46] , 
        \wNDiag_62[24] , \wPDiag_20[42] , \wNDiag_54[38] , \wNDiag_21[11] , 
        \wNDiag_54[21] , \wNDiag_26[0] , \wColumn_49[36] , \wColumn_29[32] , 
        \wPDiag_48[23] , \wScan_2[3] , \wPDiag_2[26] , \wPDiag_4[7] , 
        \wPDiag_28[27] , \wColumn_34[63] , \wColumn_41[53] , \wNDiag_41[7] , 
        \wColumn_17[52] , \wColumn_21[57] , \wColumn_62[62] , \wNDiag_4[56] , 
        \wPDiag_7[4] , \wColumn_29[18] , \wNDiag_42[4] , \wColumn_58[7] , 
        \wColumn_5[36] , \wNDiag_5[7] , \wColumn_6[46] , \wPDiag_6[17] , 
        \wPDiag_17[9] , \wNDiag_21[22] , \wPDiag_55[41] , \wNDiag_54[12] , 
        \wPDiag_55[58] , \wNDiag_17[27] , \wNDiag_34[16] , \wColumn_45[8] , 
        \wNDiag_41[26] , \wPDiag_63[44] , \wPDiag_35[45] , \wNDiag_62[17] , 
        \wPDiag_12[45] , \wPDiag_24[59] , \wPDiag_24[40] , \wColumn_58[19] , 
        \wNDiag_50[23] , \wNDiag_25[13] , \wNDiag_30[27] , \wNDiag_45[17] , 
        \wNDiag_13[16] , \wPDiag_44[44] , \wPDiag_39[22] , \wPDiag_6[24] , 
        \wNDiag_6[4] , \wNDiag_8[31] , \wColumn_45[62] , \wPDiag_59[26] , 
        \wNDiag_8[28] , \wColumn_30[52] , \wColumn_13[63] , \wNDiag_13[25] , 
        \wNDiag_30[14] , \wColumn_50[56] , \wNDiag_45[24] , \wPDiag_31[47] , 
        \wColumn_18[5] , \wNDiag_25[39] , \wNDiag_25[20] , \wPDiag_51[43] , 
        \wNDiag_50[10] , \wColumn_38[37] , \wColumn_9[9] , \wColumn_13[50] , 
        \wColumn_13[49] , \wColumn_25[55] , \wColumn_58[33] , \wColumn_30[61] , 
        \wPDiag_49[7] , \wColumn_45[51] , \wColumn_45[48] , \wPDiag_59[15] , 
        \wNDiag_18[30] , \wNDiag_38[42] , \wPDiag_54[8] , \wNDiag_58[46] , 
        \wPDiag_39[11] , \wNDiag_18[29] , \wPDiag_19[63] , \wScan_55[1] , 
        \wColumn_10[13] , \wPDiag_35[1] , \wColumn_26[16] , \wColumn_33[22] , 
        \wColumn_46[12] , \wColumn_53[26] , \wNDiag_3[17] , \wColumn_18[45] , 
        \wPDiag_36[2] , \wColumn_10[39] , \wColumn_10[20] , \wPDiag_11[35] , 
        \wNDiag_26[63] , \wPDiag_27[29] , \wPDiag_52[19] , \wNDiag_53[53] , 
        \wPDiag_27[30] , \wPDiag_47[34] , \wScan_56[2] , \wColumn_26[25] , 
        \wNDiag_33[57] , \wPDiag_51[5] , \wColumn_53[15] , \wNDiag_19[7] , 
        \wColumn_46[38] , \wNDiag_10[55] , \wPDiag_19[50] , \wPDiag_19[49] , 
        \wScan_31[5] , \wColumn_33[11] , \wColumn_46[21] , \wPDiag_32[37] , 
        \wReturn_1[0] , \wColumn_1[1] , \wNDiag_1[47] , \wNDiag_3[24] , 
        \wNDiag_26[50] , \wNDiag_46[54] , \wNDiag_26[49] , \wNDiag_53[60] , 
        \wScan_32[6] , \wCall_34[0] , \wPDiag_52[33] , \wPDiag_52[6] , 
        \wNDiag_3[9] , \wPDiag_5[54] , \wNDiag_8[2] , \wColumn_16[3] , 
        \wColumn_24[46] , \wNDiag_39[51] , \wPDiag_44[2] , \wNDiag_59[55] , 
        \wNDiag_39[48] , \wNDiag_9[11] , \wColumn_44[42] , \wColumn_12[43] , 
        \wScan_24[2] , \wColumn_2[2] , \wNDiag_2[37] , \wColumn_7[55] , 
        \wPDiag_7[37] , \wScan_27[1] , \wColumn_39[24] , \wColumn_59[39] , 
        \wNDiag_9[22] , \wNDiag_12[36] , \wColumn_15[0] , \wPDiag_30[54] , 
        \wNDiag_44[37] , \wColumn_59[20] , \wNDiag_24[33] , \wPDiag_25[60] , 
        \wPDiag_47[1] , \wPDiag_50[50] , \wPDiag_50[49] , \wPDiag_20[6] , 
        \wColumn_31[58] , \wColumn_31[41] , \wPDiag_38[28] , \wScan_40[6] , 
        \wColumn_51[45] , \wNDiag_39[62] , \wPDiag_38[31] , \wCall_46[0] , 
        \wPDiag_13[56] , \wPDiag_23[5] , \wPDiag_58[35] , \wNDiag_24[19] , 
        \wPDiag_50[63] , \wNDiag_51[29] , \wPDiag_25[53] , \wNDiag_51[30] , 
        \wNDiag_31[34] , \wColumn_39[17] , \wPDiag_45[57] , \wColumn_59[13] , 
        \wScan_43[5] , \wPDiag_4[47] , \wNDiag_11[46] , \wPDiag_33[24] , 
        \wPDiag_46[14] , \wColumn_4[16] , \wPDiag_10[15] , \wNDiag_17[1] , 
        \wNDiag_27[43] , \wNDiag_47[47] , \wPDiag_26[10] , \wPDiag_53[39] , 
        \wPDiag_53[20] , \wColumn_4[25] , \wPDiag_10[26] , \wColumn_11[33] , 
        \wNDiag_14[2] , \wPDiag_18[43] , \wNDiag_19[10] , \wColumn_27[36] , 
        \wPDiag_26[23] , \wColumn_47[32] , \wNDiag_52[59] , \wNDiag_52[40] , 
        \wPDiag_53[13] , \wNDiag_32[44] , \wPDiag_33[17] , \wPDiag_46[27] , 
        \wColumn_11[19] , \wColumn_19[56] , \wPDiag_26[8] , \wColumn_32[28] , 
        \wColumn_47[18] , \wNDiag_19[23] , \wColumn_32[31] , \wColumn_52[35] , 
        \wScan_58[4] , \wPDiag_38[4] , \wColumn_15[31] , \wColumn_36[19] , 
        \wColumn_3[57] , \wPDiag_3[35] , \wNDiag_6[35] , \wColumn_8[42] , 
        \wPDiag_8[13] , \wColumn_15[28] , \wColumn_43[29] , \wColumn_23[34] , 
        \wColumn_43[30] , \wColumn_60[18] , \wPDiag_22[12] , \wNDiag_23[41] , 
        \wNDiag_54[0] , \wNDiag_57[3] , \wNDiag_23[58] , \wPDiag_14[17] , 
        \wNDiag_15[44] , \wPDiag_57[22] , \wPDiag_37[26] , \wPDiag_42[16] , 
        \wNDiag_43[45] , \wPDiag_61[27] , \wPDiag_8[39] , \wScan_18[6] , 
        \wNDiag_30[4] , \wColumn_56[37] , \wPDiag_8[20] , \wPDiag_14[24] , 
        \wColumn_36[33] , \wColumn_37[8] , \wColumn_60[32] , \wNDiag_36[46] , 
        \wPDiag_37[15] , \wPDiag_42[25] , \wNDiag_60[47] , \wPDiag_61[14] , 
        \wNDiag_16[34] , \wNDiag_20[31] , \wNDiag_20[28] , \wPDiag_21[62] , 
        \wPDiag_22[38] , \wColumn_29[4] , \wNDiag_33[7] , \wNDiag_56[42] , 
        \wPDiag_22[21] , \wPDiag_57[11] , \wPDiag_54[52] , \wNDiag_55[18] , 
        \wPDiag_34[56] , \wNDiag_40[35] , \wPDiag_62[57] , \wColumn_55[2] , 
        \wNDiag_5[45] , \wColumn_28[12] , \wColumn_48[16] , \wPDiag_9[2] , 
        \wColumn_16[58] , \wColumn_16[41] , \wColumn_40[40] , \wColumn_20[44] , 
        \wColumn_40[59] , \wScan_64[0] , \wNDiag_48[63] , \wPDiag_49[29] , 
        \wPDiag_49[30] , \wPDiag_17[54] , \wColumn_28[38] , \wPDiag_29[34] , 
        \wColumn_56[1] , \wColumn_48[25] , \wColumn_28[21] , \wPDiag_21[51] , 
        \wColumn_31[6] , \wNDiag_35[36] , \wPDiag_41[55] , \wPDiag_63[7] , 
        \wNDiag_63[37] , \wPDiag_54[61] , \wPDiag_21[48] , \wNDiag_55[32] , 
        \wNDiag_3[30] , \wNDiag_3[29] , \wColumn_6[61] , \wNDiag_28[54] , 
        \wNDiag_28[6] , \wColumn_32[5] , \wReturn_44[0] , \wNDiag_48[50] , 
        \wPDiag_60[4] , \wColumn_35[43] , \wNDiag_35[9] , \wNDiag_48[49] , 
        \wColumn_55[47] , \wColumn_63[42] , \wColumn_6[52] , \wPDiag_6[30] , 
        \wNDiag_8[16] , \wColumn_9[4] , \wPDiag_54[5] , \wNDiag_58[52] , 
        \wPDiag_59[18] , \wColumn_25[58] , \wNDiag_38[56] , \wColumn_25[41] , 
        \wColumn_45[45] , \wColumn_13[44] , \wColumn_18[8] , \wScan_34[5] , 
        \wColumn_38[23] , \wScan_37[6] , \wPDiag_6[29] , \wColumn_58[27] , 
        \wNDiag_6[9] , \wPDiag_12[62] , \wNDiag_13[28] , \wNDiag_45[30] , 
        \wNDiag_8[25] , \wNDiag_13[31] , \wNDiag_30[19] , \wPDiag_31[53] , 
        \wNDiag_25[34] , \wCall_31[0] , \wPDiag_57[6] , \wPDiag_44[63] , 
        \wNDiag_45[29] , \wPDiag_51[57] , \wColumn_30[46] , \wPDiag_30[1] , 
        \wScan_50[1] , \wColumn_50[42] , \wPDiag_39[36] , \wColumn_62[0] , 
        \wPDiag_12[51] , \wPDiag_24[54] , \wPDiag_33[2] , \wNDiag_58[61] , 
        \wPDiag_59[32] , \wColumn_61[3] , \wPDiag_44[49] , \wNDiag_50[37] , 
        \wPDiag_12[48] , \wNDiag_30[33] , \wPDiag_44[50] , \wPDiag_31[60] , 
        \wColumn_38[10] , \wColumn_58[14] , \wScan_53[2] , \wNDiag_3[4] , 
        \wColumn_18[62] , \wColumn_5[11] , \wPDiag_5[59] , \wPDiag_5[40] , 
        \wNDiag_10[58] , \wNDiag_10[41] , \wPDiag_32[23] , \wNDiag_46[59] , 
        \wPDiag_47[13] , \wPDiag_11[12] , \wNDiag_26[44] , \wNDiag_46[40] , 
        \wPDiag_27[17] , \wPDiag_52[27] , \wNDiag_18[17] , \wPDiag_19[44] , 
        \wColumn_26[31] , \wPDiag_51[8] , \wColumn_10[34] , \wColumn_26[28] , 
        \wColumn_53[18] , \wPDiag_11[38] , \wPDiag_27[24] , \wColumn_46[35] , 
        \wPDiag_52[14] , \wNDiag_53[47] , \wPDiag_32[10] , \wPDiag_47[20] , 
        \wPDiag_11[21] , \wNDiag_33[43] , \wPDiag_47[39] , \wColumn_18[51] , 
        \wNDiag_63[2] , \wColumn_18[48] , \wColumn_33[36] , \wScan_48[3] , 
        \wColumn_1[39] , \wColumn_1[13] , \wPDiag_1[7] , \wScan_4[0] , 
        \wColumn_5[22] , \wNDiag_18[24] , \wColumn_53[32] , \wPDiag_28[3] , 
        \wNDiag_60[1] , \wPDiag_9[14] , \wColumn_14[36] , \wColumn_22[33] , 
        \wColumn_42[37] , \wNDiag_59[8] , \wNDiag_44[7] , \wPDiag_1[42] , 
        \wPDiag_2[4] , \wNDiag_22[46] , \wNDiag_47[4] , \wScan_7[3] , 
        \wColumn_9[45] , \wPDiag_23[15] , \wNDiag_14[43] , \wPDiag_56[25] , 
        \wPDiag_15[10] , \wPDiag_36[21] , \wPDiag_43[11] , \wPDiag_60[39] , 
        \wPDiag_36[38] , \wNDiag_42[42] , \wPDiag_60[20] , \wNDiag_7[32] , 
        \wPDiag_12[9] , \wColumn_40[8] , \wColumn_1[20] , \wNDiag_20[3] , 
        \wColumn_2[63] , \wPDiag_2[32] , \wPDiag_7[9] , \wNDiag_7[18] , 
        \wPDiag_9[27] , \wColumn_22[19] , \wColumn_57[30] , \wColumn_57[29] , 
        \wColumn_37[34] , \wColumn_61[35] , \wPDiag_15[23] , \wPDiag_36[12] , 
        \wNDiag_37[58] , \wPDiag_43[22] , \wNDiag_61[40] , \wNDiag_37[41] , 
        \wPDiag_60[13] , \wNDiag_61[59] , \wPDiag_16[60] , \wNDiag_21[36] , 
        \wPDiag_23[26] , \wNDiag_23[0] , \wColumn_39[3] , \wPDiag_56[16] , 
        \wNDiag_57[45] , \wPDiag_55[55] , \wReturn_33[0] , \wPDiag_35[48] , 
        \wPDiag_17[4] , \wPDiag_35[51] , \wNDiag_41[32] , \wPDiag_63[50] , 
        \wColumn_45[5] , \wNDiag_17[33] , \wPDiag_40[61] , \wPDiag_63[49] , 
        \wNDiag_42[9] , \wNDiag_4[42] , \wColumn_29[15] , \wColumn_49[11] , 
        \wColumn_17[46] , \wColumn_41[47] , \wColumn_21[43] , \wPDiag_48[37] , 
        \wColumn_2[50] , \wPDiag_2[18] , \wScan_13[0] , \wPDiag_14[7] , 
        \wColumn_46[6] , \wPDiag_28[33] , \wNDiag_29[60] , \wColumn_49[22] , 
        \wPDiag_16[53] , \wColumn_29[26] , \wNDiag_62[29] , \wPDiag_63[63] , 
        \wNDiag_17[19] , \wPDiag_20[56] , \wColumn_21[1] , \wNDiag_34[31] , 
        \wNDiag_34[28] , \wPDiag_40[52] , \wNDiag_41[18] , \wNDiag_62[30] , 
        \wPDiag_35[62] , \wNDiag_54[35] , \wColumn_2[49] , \wPDiag_28[19] , 
        \wNDiag_38[1] , \wNDiag_29[53] , \wNDiag_6[38] , \wNDiag_6[12] , 
        \wScan_10[3] , \wColumn_22[2] , \wNDiag_49[57] , \wPDiag_14[30] , 
        \wPDiag_14[29] , \wNDiag_15[63] , \wColumn_34[44] , \wColumn_54[59] , 
        \wColumn_54[40] , \wPDiag_42[31] , \wColumn_62[45] , \wNDiag_60[53] , 
        \wPDiag_61[19] , \wPDiag_42[28] , \wNDiag_43[62] , \wPDiag_22[35] , 
        \wColumn_29[9] , \wNDiag_36[52] , \wPDiag_37[18] , \wNDiag_56[56] , 
        \wPDiag_8[34] , \wColumn_23[13] , \wColumn_34[6] , \wReturn_41[0] , 
        \wColumn_56[23] , \wColumn_15[16] , \wColumn_37[5] , \wColumn_60[26] , 
        \wNDiag_30[9] , \wColumn_36[27] , \wColumn_43[17] , \wColumn_50[2] , 
        \wNDiag_6[21] , \wColumn_8[56] , \wNDiag_23[55] , \wScan_62[3] , 
        \wNDiag_15[50] , \wPDiag_37[32] , \wPDiag_57[36] , \wNDiag_15[49] , 
        \wNDiag_36[61] , \wNDiag_43[48] , \wNDiag_60[60] , \wNDiag_43[51] , 
        \wPDiag_61[33] , \wScan_61[0] , \wColumn_1[5] , \wNDiag_1[60] , 
        \wColumn_3[43] , \wScan_9[5] , \wColumn_15[25] , \wColumn_20[63] , 
        \wColumn_23[39] , \wColumn_23[20] , \wColumn_36[14] , \wNDiag_49[2] , 
        \wColumn_60[15] , \wColumn_43[24] , \wColumn_53[1] , \wColumn_56[10] , 
        \wColumn_55[53] , \wNDiag_28[59] , \wColumn_35[57] , \wNDiag_35[4] , 
        \wColumn_63[56] , \wPDiag_29[13] , \wPDiag_3[38] , \wPDiag_3[21] , 
        \wPDiag_3[12] , \wNDiag_5[62] , \wNDiag_16[13] , \wPDiag_17[40] , 
        \wNDiag_28[40] , \wColumn_32[8] , \wNDiag_35[22] , \wNDiag_40[12] , 
        \wNDiag_48[44] , \wPDiag_60[9] , \wPDiag_49[17] , \wPDiag_41[58] , 
        \wPDiag_41[41] , \wNDiag_63[23] , \wPDiag_17[59] , \wNDiag_20[16] , 
        \wPDiag_21[45] , \wNDiag_55[26] , \wNDiag_36[7] , \wColumn_48[31] , 
        \wColumn_48[28] , \wReturn_4[0] , \wColumn_28[35] , \wPDiag_49[24] , 
        \wColumn_16[55] , \wPDiag_29[39] , \wPDiag_29[20] , \wColumn_40[54] , 
        \wNDiag_51[0] , \wPDiag_19[2] , \wColumn_20[49] , \wColumn_20[50] , 
        \wColumn_55[60] , \wNDiag_5[51] , \wColumn_48[0] , \wNDiag_52[3] , 
        \wNDiag_5[48] , \wPDiag_7[10] , \wNDiag_16[39] , \wNDiag_20[25] , 
        \wPDiag_54[46] , \wNDiag_55[15] , \wNDiag_16[20] , \wNDiag_35[11] , 
        \wNDiag_40[21] , \wPDiag_62[43] , \wPDiag_34[42] , \wNDiag_40[38] , 
        \wNDiag_63[10] , \wNDiag_1[53] , \wColumn_7[58] , \wColumn_7[41] , 
        \wNDiag_12[11] , \wPDiag_13[42] , \wPDiag_23[8] , \wPDiag_25[47] , 
        \wNDiag_51[24] , \wNDiag_24[14] , \wNDiag_31[20] , \wNDiag_44[10] , 
        \wNDiag_31[39] , \wPDiag_45[43] , \wPDiag_38[25] , \wPDiag_58[21] , 
        \wNDiag_9[36] , \wPDiag_58[38] , \wNDiag_12[22] , \wReturn_19[0] , 
        \wColumn_31[55] , \wColumn_51[48] , \wColumn_24[61] , \wColumn_51[51] , 
        \wPDiag_30[59] , \wNDiag_31[13] , \wNDiag_44[23] , \wNDiag_24[27] , 
        \wPDiag_30[40] , \wPDiag_50[44] , \wNDiag_51[17] , \wNDiag_2[23] , 
        \wNDiag_2[10] , \wColumn_4[31] , \wColumn_4[28] , \wColumn_4[1] , 
        \wColumn_7[2] , \wColumn_39[30] , \wColumn_39[29] , \wPDiag_7[23] , 
        \wNDiag_12[1] , \wColumn_59[34] , \wNDiag_11[2] , \wColumn_24[52] , 
        \wColumn_44[56] , \wColumn_51[62] , \wPDiag_59[0] , \wColumn_12[57] , 
        \wNDiag_19[37] , \wPDiag_38[16] , \wScan_39[0] , \wPDiag_58[12] , 
        \wNDiag_59[58] , \wNDiag_59[41] , \wNDiag_39[45] , \wPDiag_38[9] , 
        \wScan_45[6] , \wPDiag_4[60] , \wColumn_11[14] , \wPDiag_25[6] , 
        \wPDiag_26[5] , \wColumn_27[11] , \wColumn_32[25] , \wCall_43[0] , 
        \wColumn_47[15] , \wColumn_52[21] , \wColumn_52[38] , \wColumn_19[42] , 
        \wColumn_10[0] , \wPDiag_10[32] , \wNDiag_11[61] , \wPDiag_26[37] , 
        \wNDiag_52[54] , \wScan_46[5] , \wPDiag_46[33] , \wNDiag_32[49] , 
        \wNDiag_47[60] , \wPDiag_10[18] , \wColumn_11[27] , \wColumn_13[3] , 
        \wColumn_27[22] , \wNDiag_32[50] , \wColumn_52[12] , \wPDiag_41[2] , 
        \wPDiag_18[57] , \wScan_21[2] , \wColumn_32[16] , \wColumn_47[26] , 
        \wPDiag_33[30] , \wNDiag_11[52] , \wScan_22[1] , \wNDiag_27[57] , 
        \wNDiag_32[63] , \wPDiag_33[29] , \wPDiag_46[19] , \wNDiag_47[53] , 
        \wPDiag_53[34] , \wPDiag_42[1] , \wColumn_3[60] , \wPDiag_4[53] , 
        \wNDiag_28[63] , \wPDiag_29[29] , \wColumn_3[53] , \wPDiag_3[31] , 
        \wPDiag_3[28] , \wNDiag_5[58] , \wPDiag_9[6] , \wPDiag_29[30] , 
        \wColumn_56[5] , \wPDiag_49[34] , \wColumn_16[45] , \wReturn_20[0] , 
        \wColumn_20[59] , \wColumn_20[40] , \wColumn_40[44] , \wNDiag_51[9] , 
        \wScan_64[4] , \wColumn_48[9] , \wNDiag_5[41] , \wColumn_48[12] , 
        \wColumn_28[16] , \wNDiag_16[30] , \wPDiag_34[52] , \wNDiag_35[18] , 
        \wColumn_55[6] , \wNDiag_16[29] , \wPDiag_17[63] , \wNDiag_40[28] , 
        \wPDiag_41[62] , \wNDiag_20[35] , \wNDiag_40[31] , \wPDiag_62[53] , 
        \wNDiag_63[19] , \wNDiag_28[50] , \wColumn_32[1] , \wColumn_35[47] , 
        \wPDiag_54[56] , \wColumn_63[46] , \wColumn_55[43] , \wPDiag_60[0] , 
        \wNDiag_48[54] , \wNDiag_28[49] , \wColumn_4[12] , \wNDiag_6[31] , 
        \wPDiag_17[50] , \wPDiag_17[49] , \wPDiag_21[55] , \wNDiag_28[2] , 
        \wColumn_31[2] , \wNDiag_55[36] , \wPDiag_63[3] , \wPDiag_41[51] , 
        \wNDiag_63[33] , \wPDiag_34[61] , \wPDiag_41[48] , \wPDiag_62[60] , 
        \wColumn_28[25] , \wNDiag_35[32] , \wColumn_48[38] , \wColumn_48[21] , 
        \wNDiag_6[28] , \wColumn_8[46] , \wPDiag_14[13] , \wNDiag_15[59] , 
        \wNDiag_15[40] , \wNDiag_43[41] , \wPDiag_61[23] , \wPDiag_22[16] , 
        \wPDiag_37[22] , \wPDiag_42[12] , \wNDiag_43[58] , \wPDiag_8[24] , 
        \wPDiag_8[17] , \wNDiag_23[45] , \wPDiag_57[26] , \wNDiag_54[4] , 
        \wNDiag_57[7] , \wPDiag_14[39] , \wPDiag_14[20] , \wColumn_15[35] , 
        \wColumn_23[30] , \wColumn_23[29] , \wColumn_53[8] , \wColumn_56[19] , 
        \wColumn_43[34] , \wPDiag_22[25] , \wPDiag_57[15] , \wColumn_29[0] , 
        \wNDiag_36[42] , \wPDiag_42[38] , \wNDiag_56[46] , \wPDiag_61[10] , 
        \wNDiag_33[3] , \wPDiag_37[11] , \wPDiag_42[21] , \wNDiag_60[43] , 
        \wColumn_36[37] , \wColumn_60[36] , \wColumn_11[37] , \wScan_18[2] , 
        \wNDiag_30[0] , \wColumn_56[33] , \wColumn_47[36] , \wNDiag_14[6] , 
        \wPDiag_18[47] , \wColumn_27[32] , \wNDiag_19[14] , \wNDiag_1[43] , 
        \wColumn_2[6] , \wPDiag_10[11] , \wNDiag_17[5] , \wPDiag_26[14] , 
        \wNDiag_27[47] , \wPDiag_53[24] , \wNDiag_11[42] , \wPDiag_33[39] , 
        \wNDiag_47[43] , \wPDiag_33[20] , \wPDiag_46[10] , \wNDiag_2[33] , 
        \wPDiag_4[43] , \wColumn_10[9] , \wPDiag_42[8] , \wNDiag_2[19] , 
        \wColumn_4[38] , \wColumn_4[21] , \wColumn_19[61] , \wColumn_19[52] , 
        \wNDiag_19[27] , \wPDiag_38[0] , \wColumn_27[18] , \wColumn_52[28] , 
        \wColumn_32[35] , \wColumn_52[31] , \wScan_58[0] , \wPDiag_7[33] , 
        \wPDiag_10[22] , \wNDiag_32[40] , \wNDiag_12[32] , \wColumn_15[4] , 
        \wNDiag_24[37] , \wPDiag_26[27] , \wNDiag_32[59] , \wPDiag_33[13] , 
        \wPDiag_46[23] , \wPDiag_53[17] , \wNDiag_52[44] , \wPDiag_30[50] , 
        \wPDiag_50[54] , \wNDiag_12[8] , \wPDiag_13[61] , \wPDiag_30[49] , 
        \wPDiag_45[60] , \wPDiag_47[5] , \wScan_27[5] , \wNDiag_44[33] , 
        \wColumn_59[24] , \wColumn_39[39] , \wNDiag_3[39] , \wNDiag_3[20] , 
        \wNDiag_3[13] , \wColumn_4[8] , \wNDiag_9[15] , \wColumn_12[47] , 
        \wColumn_39[20] , \wScan_24[6] , \wColumn_44[46] , \wColumn_24[42] , 
        \wColumn_7[62] , \wNDiag_8[6] , \wNDiag_39[55] , \wPDiag_59[9] , 
        \wNDiag_59[51] , \wColumn_7[51] , \wColumn_7[48] , \wPDiag_7[19] , 
        \wColumn_16[7] , \wNDiag_59[48] , \wCall_22[0] , \wPDiag_44[6] , 
        \wColumn_39[13] , \wScan_43[1] , \wNDiag_12[18] , \wPDiag_30[63] , 
        \wNDiag_44[19] , \wColumn_59[17] , \wPDiag_45[53] , \wNDiag_31[29] , 
        \wPDiag_13[52] , \wPDiag_23[1] , \wNDiag_31[30] , \wNDiag_51[34] , 
        \wPDiag_25[57] , \wPDiag_58[28] , \wNDiag_59[62] , \wNDiag_9[26] , 
        \wPDiag_20[2] , \wPDiag_58[31] , \wPDiag_38[35] , \wScan_40[2] , 
        \wColumn_51[41] , \wColumn_51[58] , \wNDiag_10[62] , \wPDiag_11[31] , 
        \wColumn_31[45] , \wNDiag_46[63] , \wPDiag_47[29] , \wPDiag_11[28] , 
        \wPDiag_32[19] , \wNDiag_33[53] , \wPDiag_47[30] , \wScan_56[6] , 
        \wColumn_18[58] , \wPDiag_27[34] , \wNDiag_53[57] , \wColumn_5[32] , 
        \wPDiag_5[63] , \wColumn_18[41] , \wPDiag_36[6] , \wColumn_10[17] , 
        \wColumn_26[12] , \wCall_50[0] , \wColumn_53[22] , \wColumn_33[26] , 
        \wColumn_46[16] , \wPDiag_35[5] , \wScan_55[5] , \wPDiag_5[50] , 
        \wNDiag_18[34] , \wNDiag_60[8] , \wPDiag_5[49] , \wNDiag_26[54] , 
        \wScan_32[2] , \wPDiag_52[2] , \wPDiag_52[37] , \wNDiag_33[60] , 
        \wPDiag_2[11] , \wColumn_5[18] , \wNDiag_10[51] , \wNDiag_10[48] , 
        \wPDiag_32[33] , \wNDiag_46[50] , \wPDiag_19[54] , \wNDiag_46[49] , 
        \wScan_31[1] , \wNDiag_5[3] , \wColumn_6[42] , \wNDiag_8[35] , 
        \wColumn_10[24] , \wColumn_33[15] , \wColumn_46[25] , \wNDiag_19[3] , 
        \wColumn_25[62] , \wColumn_26[38] , \wPDiag_51[1] , \wColumn_26[21] , 
        \wColumn_50[52] , \wColumn_53[11] , \wColumn_30[56] , \wPDiag_6[13] , 
        \wPDiag_12[58] , \wPDiag_30[8] , \wPDiag_39[26] , \wPDiag_59[22] , 
        \wColumn_62[9] , \wPDiag_44[40] , \wPDiag_12[41] , \wNDiag_13[12] , 
        \wNDiag_30[23] , \wPDiag_44[59] , \wNDiag_45[13] , \wPDiag_24[44] , 
        \wNDiag_25[17] , \wNDiag_50[27] , \wColumn_38[19] , \wScan_29[3] , 
        \wPDiag_39[15] , \wNDiag_38[46] , \wNDiag_58[42] , \wPDiag_59[11] , 
        \wPDiag_6[39] , \wColumn_13[54] , \wColumn_25[51] , \wColumn_45[55] , 
        \wColumn_25[48] , \wPDiag_49[3] , \wColumn_50[61] , \wColumn_58[37] , 
        \wPDiag_6[20] , \wNDiag_6[0] , \wNDiag_13[21] , \wColumn_18[1] , 
        \wNDiag_25[24] , \wColumn_38[33] , \wNDiag_50[14] , \wPDiag_51[47] , 
        \wPDiag_31[43] , \wNDiag_45[39] , \wNDiag_13[38] , \wColumn_29[36] , 
        \wNDiag_30[10] , \wNDiag_45[20] , \wNDiag_4[61] , \wNDiag_26[4] , 
        \wColumn_49[32] , \wColumn_21[8] , \wNDiag_21[15] , \wNDiag_54[25] , 
        \wScan_1[4] , \wColumn_2[59] , \wPDiag_16[43] , \wNDiag_17[10] , 
        \wPDiag_20[46] , \wNDiag_34[38] , \wPDiag_40[42] , \wNDiag_62[20] , 
        \wNDiag_34[21] , \wNDiag_41[11] , \wNDiag_62[39] , \wNDiag_29[43] , 
        \wPDiag_48[14] , \wNDiag_49[47] , \wColumn_2[40] , \wPDiag_28[10] , 
        \wNDiag_38[8] , \wPDiag_2[22] , \wNDiag_4[52] , \wNDiag_17[23] , 
        \wColumn_21[60] , \wNDiag_25[7] , \wColumn_34[54] , \wColumn_62[55] , 
        \wColumn_54[50] , \wColumn_54[49] , \wNDiag_21[26] , \wNDiag_34[12] , 
        \wPDiag_35[58] , \wPDiag_35[41] , \wNDiag_62[13] , \wPDiag_63[59] , 
        \wNDiag_41[22] , \wPDiag_63[40] , \wColumn_49[18] , \wNDiag_54[16] , 
        \wPDiag_55[45] , \wColumn_58[3] , \wPDiag_7[0] , \wNDiag_42[0] , 
        \wPDiag_4[3] , \wColumn_17[56] , \wColumn_21[53] , \wColumn_54[63] , 
        \wColumn_41[57] , \wNDiag_41[3] , \wPDiag_28[23] , \wPDiag_48[27] , 
        \wColumn_1[30] , \wColumn_1[29] , \wPDiag_1[61] , \wPDiag_9[37] , 
        \wColumn_14[15] , \wColumn_27[6] , \wColumn_37[24] , \wColumn_42[14] , 
        \wColumn_61[25] , \wColumn_57[39] , \wColumn_22[10] , \wColumn_57[20] , 
        \wColumn_24[5] , \wPDiag_1[52] , \wNDiag_7[22] , \wNDiag_7[11] , 
        \wReturn_52[0] , \wColumn_9[55] , \wPDiag_11[3] , \wNDiag_14[60] , 
        \wPDiag_15[33] , \wPDiag_23[36] , \wNDiag_42[61] , \wNDiag_57[55] , 
        \wNDiag_61[49] , \wScan_16[4] , \wNDiag_37[51] , \wPDiag_43[32] , 
        \wNDiag_61[50] , \wNDiag_23[9] , \wNDiag_37[48] , \wColumn_43[2] , 
        \wColumn_14[26] , \wColumn_22[23] , \wColumn_37[17] , \wColumn_57[13] , 
        \wColumn_42[27] , \wNDiag_14[53] , \wPDiag_36[31] , \wPDiag_36[28] , 
        \wNDiag_59[1] , \wColumn_61[16] , \wNDiag_37[62] , \wNDiag_42[52] , 
        \wPDiag_60[30] , \wPDiag_43[18] , \wPDiag_15[19] , \wPDiag_60[29] , 
        \wNDiag_61[63] , \wNDiag_22[56] , \wPDiag_56[35] , \wPDiag_12[0] , 
        \wColumn_40[1] , \wNDiag_3[11] , \wColumn_5[30] , \wNDiag_18[36] , 
        \wPDiag_28[8] , \wColumn_5[29] , \wPDiag_5[61] , \wColumn_10[15] , 
        \wColumn_33[24] , \wColumn_46[14] , \wColumn_26[10] , \wPDiag_35[7] , 
        \wColumn_53[39] , \wPDiag_36[4] , \wColumn_53[20] , \wReturn_12[0] , 
        \wColumn_10[26] , \wNDiag_10[60] , \wPDiag_11[33] , \wColumn_18[43] , 
        \wPDiag_27[36] , \wNDiag_33[51] , \wNDiag_53[55] , \wNDiag_33[48] , 
        \wNDiag_46[61] , \wNDiag_19[1] , \wColumn_26[23] , \wPDiag_47[32] , 
        \wNDiag_63[9] , \wPDiag_51[3] , \wScan_56[4] , \wColumn_53[13] , 
        \wColumn_33[17] , \wColumn_46[27] , \wPDiag_19[56] , \wScan_31[3] , 
        \wNDiag_46[52] , \wPDiag_47[18] , \wScan_1[6] , \wColumn_2[42] , 
        \wNDiag_3[22] , \wNDiag_10[53] , \wPDiag_32[28] , \wNDiag_33[62] , 
        \wPDiag_11[19] , \wNDiag_26[56] , \wScan_32[0] , \wPDiag_32[31] , 
        \wPDiag_52[35] , \wPDiag_5[52] , \wPDiag_52[0] , \wNDiag_5[1] , 
        \wColumn_6[59] , \wPDiag_6[11] , \wCall_48[0] , \wPDiag_12[43] , 
        \wNDiag_13[10] , \wPDiag_24[46] , \wNDiag_25[15] , \wPDiag_33[9] , 
        \wNDiag_50[25] , \wColumn_61[8] , \wNDiag_30[38] , \wPDiag_44[42] , 
        \wNDiag_30[21] , \wPDiag_39[24] , \wNDiag_45[11] , \wColumn_6[40] , 
        \wPDiag_59[39] , \wPDiag_6[22] , \wNDiag_6[2] , \wNDiag_8[37] , 
        \wColumn_30[54] , \wPDiag_59[20] , \wColumn_25[60] , \wColumn_50[50] , 
        \wColumn_50[49] , \wNDiag_13[23] , \wPDiag_31[41] , \wColumn_18[3] , 
        \wNDiag_25[26] , \wNDiag_30[12] , \wPDiag_31[58] , \wNDiag_45[22] , 
        \wNDiag_50[16] , \wColumn_38[31] , \wColumn_38[28] , \wPDiag_51[45] , 
        \wColumn_58[35] , \wColumn_13[56] , \wColumn_25[53] , \wPDiag_49[1] , 
        \wColumn_50[63] , \wColumn_45[57] , \wNDiag_58[40] , \wColumn_21[62] , 
        \wScan_29[1] , \wNDiag_38[44] , \wPDiag_39[17] , \wNDiag_58[59] , 
        \wPDiag_59[13] , \wNDiag_25[5] , \wNDiag_29[41] , \wColumn_34[56] , 
        \wColumn_54[52] , \wColumn_62[57] , \wPDiag_2[13] , \wNDiag_4[63] , 
        \wPDiag_16[58] , \wColumn_22[9] , \wPDiag_28[12] , \wNDiag_29[58] , 
        \wPDiag_48[16] , \wNDiag_49[45] , \wPDiag_16[41] , \wNDiag_17[12] , 
        \wPDiag_40[40] , \wNDiag_62[22] , \wPDiag_20[44] , \wNDiag_21[17] , 
        \wNDiag_34[23] , \wPDiag_40[59] , \wNDiag_41[13] , \wNDiag_54[27] , 
        \wNDiag_26[6] , \wColumn_49[29] , \wColumn_49[30] , \wColumn_29[34] , 
        \wPDiag_48[25] , \wColumn_1[32] , \wPDiag_1[63] , \wScan_2[5] , 
        \wPDiag_2[39] , \wPDiag_4[1] , \wColumn_17[54] , \wPDiag_28[38] , 
        \wPDiag_28[21] , \wColumn_41[55] , \wNDiag_41[1] , \wPDiag_7[2] , 
        \wColumn_21[51] , \wColumn_54[61] , \wColumn_21[48] , \wNDiag_42[2] , 
        \wPDiag_2[20] , \wNDiag_4[50] , \wNDiag_4[49] , \wColumn_58[1] , 
        \wNDiag_21[24] , \wNDiag_54[14] , \wPDiag_55[47] , \wNDiag_7[13] , 
        \wNDiag_14[62] , \wPDiag_15[31] , \wNDiag_17[38] , \wNDiag_17[21] , 
        \wPDiag_35[43] , \wNDiag_41[39] , \wNDiag_62[11] , \wNDiag_34[10] , 
        \wNDiag_41[20] , \wPDiag_63[42] , \wPDiag_36[19] , \wNDiag_37[53] , 
        \wPDiag_15[28] , \wNDiag_42[63] , \wPDiag_43[29] , \wScan_16[6] , 
        \wPDiag_43[30] , \wPDiag_60[18] , \wNDiag_61[52] , \wPDiag_23[34] , 
        \wColumn_39[8] , \wNDiag_57[57] , \wCall_10[0] , \wColumn_24[7] , 
        \wPDiag_9[35] , \wColumn_14[17] , \wColumn_22[12] , \wColumn_37[26] , 
        \wColumn_57[22] , \wColumn_42[16] , \wColumn_27[4] , \wColumn_61[27] , 
        \wColumn_1[18] , \wPDiag_1[50] , \wScan_15[5] , \wNDiag_20[8] , 
        \wPDiag_1[49] , \wNDiag_7[39] , \wNDiag_7[20] , \wPDiag_12[2] , 
        \wColumn_9[57] , \wColumn_40[3] , \wNDiag_14[51] , \wNDiag_14[48] , 
        \wNDiag_22[54] , \wPDiag_56[37] , \wNDiag_42[50] , \wPDiag_60[32] , 
        \wNDiag_37[60] , \wNDiag_42[49] , \wNDiag_61[61] , \wPDiag_36[33] , 
        \wColumn_3[62] , \wPDiag_3[33] , \wPDiag_11[1] , \wColumn_14[24] , 
        \wColumn_37[15] , \wColumn_42[25] , \wNDiag_59[3] , \wColumn_61[14] , 
        \wNDiag_16[32] , \wNDiag_20[37] , \wColumn_22[38] , \wColumn_43[0] , 
        \wColumn_22[21] , \wColumn_57[11] , \wPDiag_41[60] , \wPDiag_54[54] , 
        \wPDiag_62[48] , \wPDiag_17[61] , \wPDiag_34[50] , \wNDiag_40[33] , 
        \wColumn_55[4] , \wPDiag_62[51] , \wColumn_28[14] , \wPDiag_34[49] , 
        \wNDiag_5[43] , \wColumn_48[10] , \wNDiag_52[8] , \wPDiag_9[4] , 
        \wColumn_16[47] , \wPDiag_19[9] , \wColumn_20[42] , \wColumn_40[46] , 
        \wScan_64[6] , \wNDiag_28[61] , \wPDiag_49[36] , \wPDiag_29[32] , 
        \wCall_62[0] , \wColumn_3[51] , \wColumn_3[48] , \wPDiag_3[19] , 
        \wColumn_28[27] , \wColumn_48[23] , \wColumn_56[7] , \wNDiag_16[18] , 
        \wPDiag_34[63] , \wNDiag_35[30] , \wNDiag_35[29] , \wNDiag_40[19] , 
        \wNDiag_63[31] , \wPDiag_41[53] , \wPDiag_17[52] , \wPDiag_21[57] , 
        \wNDiag_55[34] , \wPDiag_62[62] , \wNDiag_63[28] , \wColumn_31[0] , 
        \wPDiag_63[1] , \wNDiag_28[52] , \wPDiag_29[18] , \wPDiag_8[15] , 
        \wColumn_15[37] , \wNDiag_28[0] , \wColumn_32[3] , \wColumn_35[45] , 
        \wNDiag_48[56] , \wPDiag_60[2] , \wColumn_55[58] , \wColumn_55[41] , 
        \wColumn_63[44] , \wColumn_43[36] , \wNDiag_49[9] , \wColumn_23[32] , 
        \wColumn_1[7] , \wColumn_2[4] , \wNDiag_2[31] , \wNDiag_6[33] , 
        \wColumn_8[44] , \wReturn_38[0] , \wNDiag_54[6] , \wPDiag_14[11] , 
        \wPDiag_22[14] , \wPDiag_57[24] , \wNDiag_23[47] , \wNDiag_57[5] , 
        \wPDiag_37[39] , \wNDiag_43[43] , \wPDiag_61[21] , \wNDiag_15[42] , 
        \wPDiag_37[20] , \wPDiag_42[10] , \wPDiag_61[38] , \wColumn_50[9] , 
        \wNDiag_6[19] , \wPDiag_8[26] , \wNDiag_30[2] , \wScan_18[0] , 
        \wColumn_23[18] , \wColumn_56[31] , \wColumn_56[28] , \wColumn_36[35] , 
        \wColumn_60[34] , \wPDiag_14[22] , \wPDiag_22[27] , \wNDiag_33[1] , 
        \wNDiag_36[40] , \wNDiag_36[59] , \wPDiag_37[13] , \wNDiag_60[58] , 
        \wPDiag_61[12] , \wPDiag_42[23] , \wNDiag_60[41] , \wColumn_29[2] , 
        \wPDiag_57[17] , \wNDiag_56[44] , \wNDiag_2[28] , \wColumn_19[63] , 
        \wPDiag_4[58] , \wPDiag_4[41] , \wPDiag_10[13] , \wNDiag_47[41] , 
        \wNDiag_11[59] , \wNDiag_11[40] , \wPDiag_33[22] , \wPDiag_46[12] , 
        \wNDiag_47[58] , \wNDiag_17[7] , \wPDiag_26[16] , \wPDiag_53[26] , 
        \wNDiag_27[45] , \wNDiag_1[58] , \wColumn_4[23] , \wColumn_4[10] , 
        \wPDiag_10[39] , \wPDiag_10[20] , \wColumn_11[35] , \wColumn_13[8] , 
        \wNDiag_14[4] , \wPDiag_18[45] , \wNDiag_19[16] , \wColumn_27[29] , 
        \wColumn_52[19] , \wColumn_27[30] , \wPDiag_41[9] , \wColumn_47[34] , 
        \wPDiag_26[25] , \wNDiag_52[46] , \wPDiag_53[15] , \wNDiag_32[42] , 
        \wPDiag_46[38] , \wColumn_19[50] , \wColumn_19[49] , \wPDiag_33[11] , 
        \wPDiag_46[21] , \wNDiag_19[25] , \wColumn_32[37] , \wPDiag_38[2] , 
        \wColumn_52[33] , \wScan_58[2] , \wColumn_7[60] , \wPDiag_58[19] , 
        \wNDiag_59[53] , \wNDiag_8[4] , \wColumn_16[5] , \wPDiag_44[4] , 
        \wNDiag_39[57] , \wReturn_60[0] , \wNDiag_9[17] , \wNDiag_11[9] , 
        \wColumn_24[59] , \wColumn_24[40] , \wColumn_12[45] , \wScan_24[4] , 
        \wColumn_44[44] , \wNDiag_1[41] , \wColumn_7[9] , \wColumn_39[22] , 
        \wNDiag_6[10] , \wColumn_7[53] , \wPDiag_7[31] , \wPDiag_7[28] , 
        \wColumn_59[26] , \wNDiag_9[24] , \wNDiag_12[30] , \wNDiag_44[28] , 
        \wPDiag_45[62] , \wPDiag_47[7] , \wNDiag_12[29] , \wPDiag_13[63] , 
        \wColumn_15[6] , \wNDiag_31[18] , \wPDiag_30[52] , \wNDiag_44[31] , 
        \wNDiag_24[35] , \wColumn_31[47] , \wPDiag_50[56] , \wPDiag_20[0] , 
        \wPDiag_38[37] , \wScan_40[0] , \wColumn_51[43] , \wNDiag_59[60] , 
        \wPDiag_8[36] , \wPDiag_13[50] , \wPDiag_13[49] , \wPDiag_23[3] , 
        \wPDiag_25[55] , \wNDiag_51[36] , \wPDiag_58[33] , \wPDiag_30[61] , 
        \wNDiag_31[32] , \wPDiag_45[51] , \wColumn_15[14] , \wColumn_39[11] , 
        \wScan_43[3] , \wPDiag_45[48] , \wColumn_59[15] , \wColumn_23[11] , 
        \wColumn_36[25] , \wColumn_37[7] , \wColumn_60[24] , \wColumn_43[15] , 
        \wColumn_56[21] , \wColumn_34[4] , \wColumn_56[38] , \wPDiag_14[32] , 
        \wNDiag_15[61] , \wPDiag_22[37] , \wNDiag_56[54] , \wNDiag_36[49] , 
        \wNDiag_33[8] , \wNDiag_36[50] , \wPDiag_42[33] , \wNDiag_60[51] , 
        \wColumn_15[27] , \wColumn_23[22] , \wNDiag_43[60] , \wNDiag_60[48] , 
        \wColumn_56[12] , \wNDiag_49[0] , \wColumn_53[3] , \wColumn_60[17] , 
        \wColumn_36[16] , \wColumn_43[26] , \wColumn_3[58] , \wColumn_3[41] , 
        \wPDiag_3[10] , \wNDiag_6[23] , \wColumn_8[54] , \wPDiag_14[18] , 
        \wNDiag_60[62] , \wScan_61[2] , \wPDiag_61[28] , \wNDiag_15[52] , 
        \wNDiag_23[57] , \wNDiag_36[63] , \wPDiag_37[30] , \wPDiag_42[19] , 
        \wNDiag_43[53] , \wPDiag_61[31] , \wPDiag_37[29] , \wColumn_50[0] , 
        \wPDiag_57[34] , \wScan_62[1] , \wNDiag_5[60] , \wColumn_28[37] , 
        \wNDiag_36[5] , \wColumn_48[33] , \wNDiag_16[11] , \wPDiag_17[42] , 
        \wNDiag_20[14] , \wPDiag_21[47] , \wColumn_31[9] , \wNDiag_55[24] , 
        \wPDiag_63[8] , \wNDiag_35[20] , \wNDiag_40[10] , \wNDiag_63[38] , 
        \wNDiag_35[39] , \wPDiag_41[43] , \wNDiag_48[46] , \wNDiag_63[21] , 
        \wPDiag_49[15] , \wPDiag_29[11] , \wNDiag_16[22] , \wColumn_20[61] , 
        \wNDiag_28[42] , \wNDiag_28[9] , \wColumn_35[55] , \wNDiag_35[6] , 
        \wColumn_55[48] , \wReturn_59[0] , \wColumn_63[54] , \wPDiag_34[59] , 
        \wNDiag_35[13] , \wNDiag_40[23] , \wColumn_55[51] , \wPDiag_62[41] , 
        \wPDiag_34[40] , \wPDiag_62[58] , \wNDiag_63[12] , \wScanEnable[0] , 
        \wNDiag_1[62] , \wPDiag_3[23] , \wNDiag_5[53] , \wNDiag_20[27] , 
        \wPDiag_54[44] , \wNDiag_55[17] , \wColumn_48[2] , \wColumn_48[19] , 
        \wColumn_7[43] , \wNDiag_9[34] , \wColumn_16[57] , \wPDiag_19[0] , 
        \wColumn_20[52] , \wNDiag_52[1] , \wColumn_55[62] , \wColumn_40[56] , 
        \wNDiag_51[2] , \wColumn_24[63] , \wPDiag_29[22] , \wPDiag_49[26] , 
        \wColumn_31[57] , \wColumn_51[53] , \wNDiag_12[13] , \wPDiag_13[40] , 
        \wPDiag_20[9] , \wPDiag_58[23] , \wPDiag_38[27] , \wNDiag_31[22] , 
        \wNDiag_44[12] , \wPDiag_45[58] , \wPDiag_13[59] , \wNDiag_24[16] , 
        \wPDiag_25[45] , \wPDiag_45[41] , \wNDiag_51[26] , \wNDiag_1[51] , 
        \wColumn_4[3] , \wPDiag_7[12] , \wColumn_39[18] , \wNDiag_11[0] , 
        \wPDiag_38[14] , \wScan_39[2] , \wNDiag_39[47] , \wPDiag_58[10] , 
        \wNDiag_59[43] , \wColumn_12[55] , \wColumn_44[54] , \wCall_7[0] , 
        \wPDiag_7[38] , \wPDiag_7[21] , \wColumn_24[50] , \wColumn_24[49] , 
        \wColumn_51[60] , \wPDiag_59[2] , \wNDiag_12[3] , \wColumn_39[32] , 
        \wColumn_59[36] , \wNDiag_1[48] , \wColumn_7[0] , \wNDiag_2[38] , 
        \wNDiag_2[12] , \wPDiag_10[30] , \wPDiag_10[29] , \wNDiag_11[63] , 
        \wNDiag_12[39] , \wNDiag_24[25] , \wPDiag_50[46] , \wNDiag_51[15] , 
        \wNDiag_31[11] , \wNDiag_44[21] , \wNDiag_12[20] , \wPDiag_30[42] , 
        \wNDiag_44[38] , \wNDiag_32[52] , \wPDiag_33[18] , \wPDiag_46[31] , 
        \wColumn_19[40] , \wPDiag_26[35] , \wPDiag_46[28] , \wNDiag_47[62] , 
        \wNDiag_52[56] , \wColumn_4[33] , \wPDiag_4[62] , \wColumn_19[59] , 
        \wPDiag_26[7] , \wColumn_11[16] , \wColumn_27[13] , \wColumn_52[23] , 
        \wPDiag_25[4] , \wColumn_32[27] , \wColumn_47[17] , \wPDiag_4[51] , 
        \wPDiag_4[48] , \wNDiag_19[35] , \wScan_45[4] , \wColumn_10[2] , 
        \wPDiag_42[3] , \wNDiag_2[21] , \wColumn_4[19] , \wNDiag_11[50] , 
        \wScan_22[3] , \wNDiag_27[55] , \wPDiag_53[36] , \wNDiag_47[48] , 
        \wNDiag_11[49] , \wPDiag_33[32] , \wNDiag_47[51] , \wPDiag_18[55] , 
        \wScan_21[0] , \wNDiag_32[61] , \wNDiag_5[8] , \wColumn_6[63] , 
        \wPDiag_6[32] , \wColumn_11[25] , \wPDiag_12[60] , \wColumn_13[1] , 
        \wColumn_27[20] , \wColumn_32[14] , \wColumn_47[24] , \wColumn_52[10] , 
        \wPDiag_41[0] , \wNDiag_25[36] , \wColumn_27[39] , \wPDiag_51[55] , 
        \wNDiag_45[32] , \wNDiag_13[33] , \wPDiag_31[48] , \wPDiag_44[61] , 
        \wPDiag_57[4] , \wPDiag_31[51] , \wNDiag_8[14] , \wScan_37[4] , 
        \wColumn_38[38] , \wColumn_38[21] , \wColumn_58[25] , \wColumn_45[47] , 
        \wColumn_13[46] , \wColumn_25[43] , \wPDiag_49[8] , \wNDiag_38[54] , 
        \wColumn_9[6] , \wPDiag_54[7] , \wNDiag_58[49] , \wColumn_6[50] , 
        \wPDiag_6[18] , \wColumn_38[12] , \wNDiag_58[50] , \wScan_53[0] , 
        \wColumn_58[16] , \wPDiag_12[53] , \wNDiag_30[31] , \wNDiag_13[19] , 
        \wPDiag_24[56] , \wNDiag_30[28] , \wPDiag_31[62] , \wPDiag_44[52] , 
        \wNDiag_45[18] , \wPDiag_33[0] , \wColumn_61[1] , \wNDiag_50[35] , 
        \wColumn_6[49] , \wPDiag_59[30] , \wNDiag_8[27] , \wColumn_30[44] , 
        \wPDiag_30[3] , \wPDiag_39[34] , \wNDiag_58[63] , \wPDiag_59[29] , 
        \wColumn_62[2] , \wScan_50[3] , \wColumn_50[59] , \wColumn_50[40] , 
        \wColumn_10[36] , \wNDiag_19[8] , \wColumn_46[37] , \wNDiag_3[32] , 
        \wNDiag_3[6] , \wColumn_5[13] , \wNDiag_18[15] , \wColumn_26[33] , 
        \wPDiag_19[46] , \wPDiag_5[42] , \wNDiag_10[43] , \wNDiag_26[46] , 
        \wPDiag_27[15] , \wPDiag_52[25] , \wPDiag_32[21] , \wPDiag_47[11] , 
        \wPDiag_11[10] , \wCall_29[0] , \wNDiag_46[42] , \wPDiag_32[38] , 
        \wColumn_18[60] , \wColumn_5[39] , \wPDiag_52[9] , \wColumn_5[20] , 
        \wNDiag_60[3] , \wNDiag_18[26] , \wPDiag_28[1] , \wScan_48[1] , 
        \wColumn_53[30] , \wScan_1[2] , \wColumn_1[36] , \wColumn_1[22] , 
        \wColumn_1[11] , \wPDiag_1[59] , \wNDiag_3[18] , \wColumn_26[19] , 
        \wColumn_33[34] , \wColumn_53[29] , \wNDiag_7[30] , \wNDiag_7[29] , 
        \wPDiag_11[23] , \wColumn_18[53] , \wPDiag_32[12] , \wNDiag_33[58] , 
        \wPDiag_47[22] , \wPDiag_27[26] , \wNDiag_33[41] , \wNDiag_53[45] , 
        \wNDiag_63[0] , \wPDiag_52[16] , \wPDiag_1[40] , \wPDiag_2[6] , 
        \wScan_7[1] , \wNDiag_14[58] , \wNDiag_14[41] , \wPDiag_36[23] , 
        \wNDiag_42[59] , \wPDiag_43[13] , \wNDiag_42[40] , \wPDiag_60[22] , 
        \wPDiag_15[12] , \wNDiag_47[6] , \wColumn_9[47] , \wNDiag_22[44] , 
        \wPDiag_23[17] , \wPDiag_56[27] , \wPDiag_1[5] , \wScan_4[2] , 
        \wPDiag_9[16] , \wPDiag_11[8] , \wColumn_43[9] , \wNDiag_44[5] , 
        \wColumn_22[31] , \wColumn_22[28] , \wColumn_57[18] , \wColumn_14[34] , 
        \wPDiag_9[25] , \wPDiag_15[38] , \wPDiag_23[24] , \wColumn_39[1] , 
        \wColumn_42[35] , \wNDiag_57[47] , \wPDiag_56[14] , \wPDiag_15[21] , 
        \wPDiag_36[10] , \wPDiag_43[20] , \wNDiag_61[42] , \wNDiag_23[2] , 
        \wNDiag_37[43] , \wColumn_37[36] , \wPDiag_43[39] , \wPDiag_60[11] , 
        \wColumn_61[37] , \wColumn_57[32] , \wNDiag_20[1] , \wColumn_1[3] , 
        \wNDiag_1[45] , \wColumn_2[61] , \wPDiag_28[31] , \wColumn_2[52] , 
        \wPDiag_2[30] , \wPDiag_4[8] , \wPDiag_14[5] , \wColumn_21[58] , 
        \wPDiag_28[28] , \wNDiag_29[62] , \wColumn_46[4] , \wPDiag_48[35] , 
        \wColumn_21[41] , \wColumn_41[45] , \wNDiag_41[8] , \wNDiag_4[59] , 
        \wNDiag_4[40] , \wColumn_17[44] , \wColumn_49[13] , \wColumn_58[8] , 
        \wPDiag_2[29] , \wScan_10[1] , \wPDiag_16[62] , \wNDiag_17[28] , 
        \wColumn_29[17] , \wNDiag_41[30] , \wNDiag_62[18] , \wPDiag_63[52] , 
        \wPDiag_17[6] , \wNDiag_17[31] , \wPDiag_40[63] , \wNDiag_41[29] , 
        \wNDiag_21[34] , \wNDiag_34[19] , \wPDiag_35[53] , \wColumn_45[7] , 
        \wPDiag_55[57] , \wColumn_34[46] , \wColumn_62[47] , \wColumn_22[0] , 
        \wNDiag_49[55] , \wColumn_54[42] , \wPDiag_7[35] , \wNDiag_12[34] , 
        \wScan_13[2] , \wPDiag_16[51] , \wPDiag_20[54] , \wNDiag_29[51] , 
        \wNDiag_29[48] , \wNDiag_38[3] , \wColumn_21[3] , \wNDiag_34[33] , 
        \wNDiag_54[37] , \wPDiag_16[48] , \wPDiag_35[60] , \wPDiag_40[49] , 
        \wPDiag_63[61] , \wColumn_29[24] , \wPDiag_40[50] , \wNDiag_62[32] , 
        \wColumn_49[39] , \wColumn_49[20] , \wNDiag_24[31] , \wNDiag_24[28] , 
        \wPDiag_25[62] , \wPDiag_50[52] , \wNDiag_51[18] , \wNDiag_44[35] , 
        \wPDiag_47[3] , \wColumn_15[2] , \wPDiag_30[56] , \wScan_27[3] , 
        \wColumn_39[26] , \wColumn_59[22] , \wCall_2[0] , \wColumn_7[57] , 
        \wNDiag_8[0] , \wNDiag_9[13] , \wColumn_44[40] , \wColumn_12[58] , 
        \wColumn_12[41] , \wColumn_44[59] , \wScan_24[0] , \wPDiag_13[54] , 
        \wColumn_16[1] , \wColumn_24[44] , \wPDiag_38[19] , \wNDiag_39[53] , 
        \wPDiag_44[0] , \wNDiag_31[36] , \wColumn_39[15] , \wNDiag_59[57] , 
        \wColumn_59[11] , \wPDiag_23[7] , \wPDiag_25[51] , \wPDiag_45[55] , 
        \wPDiag_50[61] , \wPDiag_25[48] , \wNDiag_51[32] , \wNDiag_9[39] , 
        \wNDiag_9[20] , \wPDiag_20[4] , \wPDiag_38[33] , \wNDiag_39[60] , 
        \wPDiag_58[37] , \wColumn_31[43] , \wScan_40[4] , \wColumn_51[47] , 
        \wColumn_11[31] , \wColumn_47[29] , \wColumn_11[28] , \wColumn_32[19] , 
        \wColumn_47[30] , \wNDiag_14[0] , \wPDiag_18[58] , \wColumn_27[34] , 
        \wPDiag_18[41] , \wNDiag_19[12] , \wColumn_2[0] , \wColumn_4[14] , 
        \wNDiag_17[3] , \wPDiag_26[12] , \wNDiag_27[41] , \wPDiag_53[22] , 
        \wNDiag_27[58] , \wNDiag_2[35] , \wPDiag_4[45] , \wPDiag_10[17] , 
        \wNDiag_11[44] , \wPDiag_33[26] , \wPDiag_46[16] , \wNDiag_47[45] , 
        \wColumn_3[55] , \wPDiag_3[37] , \wColumn_4[27] , \wNDiag_5[47] , 
        \wNDiag_6[37] , \wPDiag_10[24] , \wColumn_19[54] , \wNDiag_19[38] , 
        \wNDiag_19[21] , \wPDiag_25[9] , \wColumn_32[33] , \wPDiag_38[6] , 
        \wColumn_52[37] , \wScan_58[6] , \wPDiag_33[15] , \wPDiag_46[25] , 
        \wPDiag_26[38] , \wNDiag_32[46] , \wPDiag_26[21] , \wNDiag_52[42] , 
        \wPDiag_53[11] , \wColumn_8[59] , \wPDiag_14[15] , \wNDiag_15[46] , 
        \wPDiag_37[24] , \wPDiag_42[14] , \wNDiag_43[47] , \wPDiag_61[25] , 
        \wNDiag_57[1] , \wColumn_8[40] , \wNDiag_23[43] , \wPDiag_57[39] , 
        \wPDiag_8[22] , \wPDiag_8[11] , \wPDiag_22[10] , \wPDiag_57[20] , 
        \wColumn_23[36] , \wNDiag_54[2] , \wPDiag_14[26] , \wColumn_15[33] , 
        \wPDiag_22[23] , \wColumn_29[6] , \wColumn_43[32] , \wNDiag_56[40] , 
        \wPDiag_37[17] , \wNDiag_56[59] , \wPDiag_57[13] , \wPDiag_42[27] , 
        \wNDiag_60[45] , \wColumn_15[19] , \wNDiag_33[5] , \wNDiag_36[44] , 
        \wColumn_34[9] , \wPDiag_61[16] , \wColumn_36[31] , \wColumn_36[28] , 
        \wColumn_43[18] , \wColumn_60[30] , \wScan_18[4] , \wColumn_56[35] , 
        \wColumn_60[29] , \wPDiag_9[0] , \wPDiag_29[36] , \wNDiag_30[6] , 
        \wNDiag_48[61] , \wColumn_56[3] , \wColumn_16[43] , \wColumn_20[46] , 
        \wPDiag_49[32] , \wColumn_40[42] , \wColumn_48[14] , \wScan_64[2] , 
        \wNDiag_16[36] , \wColumn_28[10] , \wNDiag_40[37] , \wPDiag_62[55] , 
        \wNDiag_20[33] , \wPDiag_21[60] , \wPDiag_34[54] , \wPDiag_54[50] , 
        \wColumn_55[0] , \wPDiag_54[49] , \wColumn_32[7] , \wColumn_35[58] , 
        \wColumn_35[41] , \wColumn_63[59] , \wNDiag_48[52] , \wColumn_55[45] , 
        \wColumn_63[40] , \wPDiag_49[18] , \wPDiag_60[6] , \wPDiag_17[56] , 
        \wNDiag_20[19] , \wNDiag_28[56] , \wNDiag_28[4] , \wPDiag_21[53] , 
        \wColumn_31[4] , \wPDiag_54[63] , \wNDiag_35[34] , \wNDiag_55[30] , 
        \wNDiag_55[29] , \wPDiag_63[5] , \wColumn_28[23] , \wPDiag_41[57] , 
        \wNDiag_63[35] , \wNDiag_36[8] , \wColumn_48[27] , \wPDiag_1[54] , 
        \wPDiag_1[8] , \wNDiag_7[17] , \wPDiag_9[31] , \wPDiag_9[28] , 
        \wColumn_14[13] , \wScan_15[1] , \wColumn_22[16] , \wColumn_27[0] , 
        \wColumn_61[23] , \wColumn_37[22] , \wColumn_42[12] , \wColumn_57[26] , 
        \wColumn_24[3] , \wColumn_9[60] , \wNDiag_22[63] , \wPDiag_23[29] , 
        \wPDiag_23[30] , \wPDiag_56[19] , \wNDiag_57[53] , \wPDiag_11[5] , 
        \wPDiag_15[35] , \wScan_16[2] , \wPDiag_43[34] , \wNDiag_61[56] , 
        \wNDiag_37[57] , \wColumn_22[25] , \wColumn_57[15] , \wColumn_14[39] , 
        \wColumn_14[20] , \wColumn_42[38] , \wColumn_43[4] , \wColumn_61[10] , 
        \wNDiag_59[7] , \wColumn_37[11] , \wColumn_42[21] , \wNDiag_7[24] , 
        \wColumn_9[53] , \wNDiag_14[55] , \wNDiag_44[8] , \wNDiag_22[50] , 
        \wPDiag_36[37] , \wNDiag_42[54] , \wNDiag_57[60] , \wPDiag_60[36] , 
        \wPDiag_12[6] , \wNDiag_22[49] , \wPDiag_56[33] , \wColumn_40[7] , 
        \wScan_2[1] , \wColumn_2[46] , \wPDiag_2[17] , \wPDiag_16[45] , 
        \wPDiag_20[59] , \wPDiag_20[40] , \wNDiag_26[2] , \wColumn_29[30] , 
        \wColumn_29[29] , \wColumn_49[34] , \wNDiag_21[13] , \wNDiag_54[23] , 
        \wNDiag_17[16] , \wNDiag_34[27] , \wNDiag_41[17] , \wPDiag_40[44] , 
        \wPDiag_48[12] , \wNDiag_49[41] , \wNDiag_62[26] , \wNDiag_49[58] , 
        \wColumn_17[63] , \wPDiag_28[16] , \wNDiag_29[45] , \wColumn_34[52] , 
        \wColumn_41[62] , \wNDiag_17[25] , \wNDiag_25[1] , \wColumn_62[53] , 
        \wNDiag_34[14] , \wNDiag_41[24] , \wColumn_54[56] , \wPDiag_63[46] , 
        \wPDiag_35[47] , \wNDiag_62[15] , \wPDiag_55[43] , \wPDiag_2[24] , 
        \wNDiag_4[54] , \wNDiag_21[39] , \wNDiag_21[20] , \wNDiag_54[10] , 
        \wColumn_58[5] , \wPDiag_4[5] , \wPDiag_7[6] , \wColumn_21[55] , 
        \wNDiag_42[6] , \wColumn_41[51] , \wNDiag_41[5] , \wPDiag_14[8] , 
        \wColumn_17[50] , \wColumn_17[49] , \wColumn_34[61] , \wColumn_41[48] , 
        \wColumn_62[60] , \wPDiag_28[25] , \wColumn_46[9] , \wPDiag_48[38] , 
        \wPDiag_48[21] , \wNDiag_3[26] , \wNDiag_3[15] , \wNDiag_5[5] , 
        \wColumn_6[44] , \wNDiag_8[33] , \wColumn_30[50] , \wColumn_50[54] , 
        \wColumn_45[60] , \wColumn_13[61] , \wColumn_30[49] , \wPDiag_6[15] , 
        \wPDiag_12[47] , \wPDiag_39[39] , \wPDiag_59[24] , \wPDiag_39[20] , 
        \wNDiag_13[14] , \wNDiag_30[25] , \wNDiag_45[15] , \wPDiag_24[42] , 
        \wPDiag_44[46] , \wNDiag_25[11] , \wNDiag_50[38] , \wNDiag_50[21] , 
        \wScan_29[5] , \wNDiag_38[40] , \wNDiag_38[59] , \wPDiag_39[13] , 
        \wPDiag_6[26] , \wNDiag_8[19] , \wColumn_30[63] , \wColumn_45[53] , 
        \wNDiag_58[44] , \wPDiag_59[17] , \wColumn_13[52] , \wColumn_25[57] , 
        \wPDiag_49[5] , \wNDiag_6[6] , \wColumn_18[7] , \wColumn_38[35] , 
        \wColumn_58[31] , \wColumn_58[28] , \wNDiag_25[22] , \wNDiag_50[12] , 
        \wPDiag_51[58] , \wPDiag_51[41] , \wNDiag_30[16] , \wNDiag_45[26] , 
        \wPDiag_57[9] , \wPDiag_11[37] , \wNDiag_13[27] , \wPDiag_31[45] , 
        \wNDiag_33[55] , \wPDiag_47[36] , \wScan_56[0] , \wColumn_18[47] , 
        \wNDiag_26[61] , \wPDiag_27[32] , \wNDiag_53[51] , \wNDiag_53[48] , 
        \wColumn_5[34] , \wColumn_10[11] , \wColumn_26[14] , \wPDiag_36[0] , 
        \wColumn_53[24] , \wColumn_33[39] , \wColumn_33[20] , \wPDiag_35[3] , 
        \wColumn_46[10] , \wPDiag_5[56] , \wNDiag_18[32] , \wScan_55[3] , 
        \wPDiag_19[61] , \wPDiag_52[4] , \wNDiag_10[57] , \wNDiag_26[52] , 
        \wPDiag_52[28] , \wNDiag_53[62] , \wPDiag_27[18] , \wScan_32[4] , 
        \wPDiag_52[31] , \wPDiag_32[35] , \wNDiag_46[56] , \wColumn_10[22] , 
        \wNDiag_18[18] , \wPDiag_19[52] , \wNDiag_19[5] , \wColumn_33[13] , 
        \wColumn_46[23] , \wColumn_53[17] , \wColumn_26[27] , \wColumn_1[26] , 
        \wColumn_1[15] , \wPDiag_1[1] , \wColumn_2[56] , \wPDiag_2[34] , 
        \wPDiag_17[2] , \wNDiag_17[35] , \wPDiag_20[63] , \wNDiag_21[30] , 
        \wPDiag_51[7] , \wNDiag_21[29] , \wNDiag_54[19] , \wPDiag_55[53] , 
        \wColumn_29[13] , \wPDiag_35[57] , \wNDiag_41[34] , \wColumn_45[3] , 
        \wPDiag_63[56] , \wNDiag_4[44] , \wColumn_49[17] , \wScan_13[6] , 
        \wPDiag_14[1] , \wColumn_17[59] , \wColumn_17[40] , \wColumn_41[58] , 
        \wColumn_41[41] , \wColumn_21[45] , \wPDiag_28[35] , \wPDiag_48[31] , 
        \wPDiag_48[28] , \wNDiag_49[62] , \wColumn_46[0] , \wCall_15[0] , 
        \wPDiag_16[55] , \wColumn_29[39] , \wColumn_29[20] , \wColumn_49[24] , 
        \wNDiag_34[37] , \wPDiag_40[54] , \wNDiag_62[36] , \wPDiag_20[49] , 
        \wNDiag_54[33] , \wPDiag_20[50] , \wColumn_21[7] , \wNDiag_29[55] , 
        \wPDiag_55[60] , \wScan_4[6] , \wScan_10[5] , \wColumn_22[4] , 
        \wNDiag_38[7] , \wNDiag_49[48] , \wNDiag_25[8] , \wNDiag_49[51] , 
        \wColumn_54[46] , \wColumn_14[30] , \wColumn_14[29] , \wColumn_34[42] , 
        \wColumn_62[43] , \wColumn_42[31] , \wColumn_61[19] , \wColumn_42[28] , 
        \wColumn_37[18] , \wPDiag_9[12] , \wColumn_22[35] , \wNDiag_44[1] , 
        \wPDiag_1[44] , \wPDiag_2[2] , \wColumn_9[43] , \wNDiag_22[59] , 
        \wPDiag_56[23] , \wPDiag_23[13] , \wNDiag_47[2] , \wNDiag_14[45] , 
        \wPDiag_15[16] , \wNDiag_22[40] , \wNDiag_42[44] , \wPDiag_60[26] , 
        \wPDiag_36[27] , \wPDiag_43[17] , \wScan_7[5] , \wNDiag_7[34] , 
        \wNDiag_3[36] , \wPDiag_9[38] , \wPDiag_9[21] , \wNDiag_20[5] , 
        \wPDiag_15[25] , \wColumn_27[9] , \wColumn_37[32] , \wColumn_57[36] , 
        \wColumn_61[33] , \wPDiag_23[39] , \wPDiag_23[20] , \wNDiag_23[6] , 
        \wNDiag_37[47] , \wPDiag_36[14] , \wPDiag_60[15] , \wPDiag_43[24] , 
        \wNDiag_61[46] , \wPDiag_56[10] , \wColumn_39[5] , \wNDiag_57[43] , 
        \wNDiag_3[2] , \wPDiag_5[46] , \wPDiag_11[14] , \wNDiag_46[46] , 
        \wPDiag_47[15] , \wColumn_5[17] , \wNDiag_10[47] , \wPDiag_32[25] , 
        \wNDiag_26[42] , \wPDiag_27[11] , \wPDiag_52[21] , \wPDiag_52[38] , 
        \wNDiag_18[11] , \wPDiag_19[42] , \wColumn_10[32] , \wColumn_26[37] , 
        \wColumn_46[33] , \wColumn_10[18] , \wPDiag_11[27] , \wPDiag_27[22] , 
        \wPDiag_52[12] , \wNDiag_53[58] , \wNDiag_53[41] , \wColumn_18[57] , 
        \wPDiag_32[16] , \wNDiag_33[45] , \wNDiag_63[4] , \wPDiag_36[9] , 
        \wPDiag_47[26] , \wColumn_33[30] , \wColumn_33[29] , \wColumn_46[19] , 
        \wScan_48[5] , \wColumn_53[34] , \wNDiag_1[55] , \wColumn_2[9] , 
        \wNDiag_2[16] , \wColumn_4[37] , \wColumn_5[24] , \wNDiag_18[22] , 
        \wPDiag_28[5] , \wColumn_6[54] , \wPDiag_6[36] , \wNDiag_8[10] , 
        \wColumn_9[2] , \wNDiag_60[7] , \wColumn_13[42] , \wColumn_25[47] , 
        \wNDiag_38[50] , \wNDiag_38[49] , \wPDiag_54[3] , \wNDiag_58[54] , 
        \wScan_34[3] , \wColumn_45[43] , \wColumn_38[25] , \wColumn_58[21] , 
        \wNDiag_8[23] , \wNDiag_13[37] , \wScan_37[0] , \wPDiag_57[0] , 
        \wColumn_58[38] , \wPDiag_24[61] , \wNDiag_25[32] , \wPDiag_31[55] , 
        \wNDiag_45[36] , \wPDiag_51[48] , \wPDiag_51[51] , \wColumn_30[59] , 
        \wColumn_30[40] , \wPDiag_30[7] , \wPDiag_39[30] , \wColumn_50[44] , 
        \wColumn_62[6] , \wNDiag_38[63] , \wPDiag_39[29] , \wPDiag_12[57] , 
        \wReturn_17[0] , \wPDiag_24[52] , \wNDiag_50[31] , \wPDiag_59[34] , 
        \wNDiag_25[18] , \wPDiag_33[4] , \wNDiag_50[28] , \wPDiag_51[62] , 
        \wColumn_61[5] , \wPDiag_44[56] , \wNDiag_30[35] , \wPDiag_18[62] , 
        \wNDiag_19[28] , \wColumn_38[16] , \wScan_53[4] , \wColumn_58[12] , 
        \wNDiag_19[31] , \wColumn_11[12] , \wColumn_32[23] , \wScan_45[0] , 
        \wColumn_47[13] , \wPDiag_25[0] , \wPDiag_26[3] , \wColumn_27[17] , 
        \wColumn_52[27] , \wPDiag_10[34] , \wColumn_19[44] , \wPDiag_26[31] , 
        \wPDiag_26[28] , \wNDiag_27[62] , \wNDiag_32[56] , \wNDiag_52[52] , 
        \wPDiag_53[18] , \wColumn_11[38] , \wColumn_13[5] , \wPDiag_41[4] , 
        \wScan_46[3] , \wPDiag_46[35] , \wColumn_27[24] , \wColumn_52[14] , 
        \wColumn_32[10] , \wColumn_47[20] , \wColumn_11[21] , \wColumn_47[39] , 
        \wNDiag_14[9] , \wPDiag_18[51] , \wPDiag_18[48] , \wScan_21[4] , 
        \wNDiag_47[55] , \wNDiag_2[25] , \wNDiag_11[54] , \wNDiag_27[51] , 
        \wNDiag_27[48] , \wPDiag_33[36] , \wPDiag_53[32] , \wNDiag_52[61] , 
        \wPDiag_4[55] , \wColumn_10[6] , \wPDiag_42[7] , \wColumn_7[47] , 
        \wPDiag_7[16] , \wColumn_59[18] , \wNDiag_12[17] , \wNDiag_24[12] , 
        \wPDiag_25[58] , \wPDiag_25[41] , \wNDiag_51[22] , \wPDiag_13[44] , 
        \wPDiag_45[45] , \wNDiag_31[26] , \wPDiag_38[23] , \wNDiag_44[16] , 
        \wColumn_7[4] , \wNDiag_9[30] , \wNDiag_9[29] , \wColumn_12[62] , 
        \wPDiag_58[27] , \wColumn_31[53] , \wColumn_44[63] , \wNDiag_12[24] , 
        \wPDiag_30[46] , \wColumn_51[57] , \wNDiag_24[38] , \wNDiag_24[21] , 
        \wNDiag_31[15] , \wNDiag_44[25] , \wNDiag_51[11] , \wPDiag_50[42] , 
        \wColumn_39[36] , \wColumn_3[45] , \wColumn_4[7] , \wPDiag_7[25] , 
        \wNDiag_12[7] , \wColumn_59[32] , \wColumn_24[54] , \wPDiag_59[6] , 
        \wNDiag_8[9] , \wNDiag_11[4] , \wColumn_12[51] , \wColumn_44[49] , 
        \wColumn_12[48] , \wColumn_44[50] , \wColumn_16[60] , \wColumn_16[8] , 
        \wColumn_31[60] , \wNDiag_59[47] , \wColumn_35[48] , \wNDiag_35[2] , 
        \wPDiag_38[10] , \wPDiag_44[9] , \wPDiag_58[14] , \wScan_39[6] , 
        \wNDiag_39[43] , \wColumn_55[55] , \wNDiag_28[46] , \wColumn_35[51] , 
        \wColumn_63[50] , \wColumn_40[61] , \wColumn_63[49] , \wPDiag_3[27] , 
        \wPDiag_3[14] , \wNDiag_16[15] , \wPDiag_29[15] , \wNDiag_48[42] , 
        \wPDiag_49[11] , \wPDiag_17[46] , \wPDiag_41[47] , \wNDiag_63[25] , 
        \wNDiag_20[10] , \wNDiag_35[24] , \wNDiag_40[14] , \wPDiag_21[43] , 
        \wNDiag_55[20] , \wColumn_28[33] , \wNDiag_36[1] , \wNDiag_55[39] , 
        \wColumn_48[37] , \wPDiag_9[9] , \wPDiag_49[22] , \wColumn_16[53] , 
        \wPDiag_29[26] , \wColumn_63[63] , \wPDiag_19[4] , \wColumn_20[56] , 
        \wColumn_35[62] , \wColumn_40[52] , \wNDiag_51[6] , \wColumn_28[19] , 
        \wNDiag_52[5] , \wNDiag_5[57] , \wColumn_48[6] , \wNDiag_6[27] , 
        \wNDiag_6[14] , \wColumn_8[63] , \wPDiag_14[36] , \wNDiag_16[26] , 
        \wNDiag_20[23] , \wPDiag_54[59] , \wNDiag_55[13] , \wPDiag_34[44] , 
        \wPDiag_54[40] , \wNDiag_63[16] , \wNDiag_35[17] , \wNDiag_40[27] , 
        \wPDiag_62[45] , \wColumn_55[9] , \wNDiag_36[54] , \wPDiag_22[33] , 
        \wPDiag_42[37] , \wNDiag_60[55] , \wNDiag_23[60] , \wNDiag_56[49] , 
        \wNDiag_56[50] , \wPDiag_8[32] , \wColumn_34[0] , \wColumn_15[10] , 
        \wColumn_23[15] , \wColumn_36[21] , \wColumn_56[25] , \wColumn_43[11] , 
        \wColumn_60[39] , \wColumn_36[38] , \wColumn_37[3] , \wColumn_60[20] , 
        \wColumn_8[50] , \wColumn_50[4] , \wNDiag_57[8] , \wColumn_8[49] , 
        \wPDiag_57[30] , \wScan_62[5] , \wScan_9[3] , \wNDiag_15[56] , 
        \wPDiag_22[19] , \wNDiag_56[63] , \wPDiag_57[29] , \wNDiag_23[53] , 
        \wNDiag_43[57] , \wPDiag_61[35] , \wPDiag_37[34] , \wScan_1[3] , 
        \wColumn_1[2] , \wColumn_2[1] , \wPDiag_8[18] , \wColumn_15[23] , 
        \wColumn_36[12] , \wColumn_43[22] , \wScan_61[6] , \wNDiag_49[4] , 
        \wColumn_60[13] , \wColumn_53[7] , \wColumn_56[16] , \wPDiag_10[16] , 
        \wColumn_23[26] , \wNDiag_47[44] , \wNDiag_2[34] , \wNDiag_11[45] , 
        \wPDiag_33[27] , \wPDiag_46[17] , \wNDiag_17[2] , \wPDiag_26[13] , 
        \wNDiag_27[59] , \wPDiag_53[23] , \wNDiag_27[40] , \wPDiag_4[44] , 
        \wColumn_11[30] , \wColumn_11[29] , \wColumn_27[35] , \wColumn_47[31] , 
        \wColumn_47[28] , \wColumn_32[18] , \wNDiag_1[44] , \wColumn_4[26] , 
        \wColumn_4[15] , \wPDiag_10[25] , \wNDiag_14[1] , \wPDiag_18[59] , 
        \wPDiag_18[40] , \wNDiag_19[13] , \wColumn_19[55] , \wPDiag_26[39] , 
        \wPDiag_26[20] , \wPDiag_53[10] , \wNDiag_52[43] , \wNDiag_19[39] , 
        \wNDiag_32[47] , \wPDiag_33[14] , \wPDiag_38[7] , \wPDiag_46[24] , 
        \wNDiag_19[20] , \wNDiag_8[1] , \wPDiag_25[8] , \wColumn_32[32] , 
        \wColumn_52[36] , \wNDiag_9[12] , \wColumn_12[40] , \wScan_24[1] , 
        \wColumn_24[45] , \wColumn_44[58] , \wColumn_12[59] , \wColumn_44[41] , 
        \wNDiag_12[35] , \wColumn_16[0] , \wPDiag_44[1] , \wNDiag_59[56] , 
        \wPDiag_38[18] , \wNDiag_39[52] , \wColumn_15[3] , \wPDiag_30[57] , 
        \wPDiag_47[2] , \wNDiag_24[30] , \wNDiag_44[34] , \wNDiag_24[29] , 
        \wPDiag_50[53] , \wNDiag_51[19] , \wPDiag_25[63] , \wColumn_39[27] , 
        \wReturn_2[0] , \wColumn_3[54] , \wPDiag_3[36] , \wColumn_7[56] , 
        \wPDiag_7[34] , \wColumn_59[23] , \wPDiag_20[5] , \wScan_27[2] , 
        \wPDiag_38[32] , \wNDiag_39[61] , \wPDiag_58[36] , \wNDiag_9[38] , 
        \wNDiag_9[21] , \wColumn_31[42] , \wPDiag_13[55] , \wPDiag_23[6] , 
        \wPDiag_25[50] , \wPDiag_25[49] , \wColumn_39[14] , \wScan_40[5] , 
        \wColumn_51[46] , \wScan_43[6] , \wColumn_59[10] , \wCall_45[0] , 
        \wNDiag_51[33] , \wPDiag_50[60] , \wNDiag_31[37] , \wPDiag_45[54] , 
        \wColumn_28[11] , \wNDiag_5[46] , \wPDiag_9[1] , \wNDiag_16[37] , 
        \wNDiag_20[32] , \wColumn_48[15] , \wPDiag_54[48] , \wPDiag_21[61] , 
        \wPDiag_54[51] , \wPDiag_34[55] , \wColumn_55[1] , \wNDiag_40[36] , 
        \wPDiag_62[54] , \wColumn_16[42] , \wPDiag_29[37] , \wNDiag_48[60] , 
        \wPDiag_49[33] , \wColumn_56[2] , \wScan_64[3] , \wPDiag_17[57] , 
        \wColumn_20[47] , \wColumn_40[43] , \wNDiag_35[35] , \wPDiag_41[56] , 
        \wNDiag_63[34] , \wReturn_47[0] , \wNDiag_20[18] , \wPDiag_21[52] , 
        \wNDiag_55[31] , \wColumn_28[22] , \wColumn_31[5] , \wNDiag_55[28] , 
        \wNDiag_36[9] , \wPDiag_54[62] , \wPDiag_63[4] , \wColumn_48[26] , 
        \wNDiag_28[57] , \wColumn_35[59] , \wColumn_55[44] , \wColumn_35[40] , 
        \wColumn_63[41] , \wColumn_63[58] , \wNDiag_28[5] , \wPDiag_8[10] , 
        \wColumn_15[32] , \wColumn_32[6] , \wColumn_43[33] , \wNDiag_48[53] , 
        \wPDiag_49[19] , \wPDiag_60[7] , \wNDiag_54[3] , \wColumn_23[37] , 
        \wColumn_2[47] , \wNDiag_6[36] , \wColumn_8[58] , \wColumn_8[41] , 
        \wPDiag_57[21] , \wPDiag_22[11] , \wPDiag_57[38] , \wPDiag_8[23] , 
        \wPDiag_14[14] , \wNDiag_23[42] , \wNDiag_57[0] , \wNDiag_43[46] , 
        \wPDiag_61[24] , \wNDiag_15[47] , \wPDiag_37[25] , \wPDiag_42[15] , 
        \wPDiag_14[27] , \wColumn_15[18] , \wScan_18[5] , \wColumn_56[34] , 
        \wColumn_36[30] , \wNDiag_30[7] , \wColumn_36[29] , \wColumn_60[28] , 
        \wColumn_43[19] , \wColumn_60[31] , \wNDiag_33[4] , \wPDiag_22[22] , 
        \wNDiag_36[45] , \wPDiag_37[16] , \wPDiag_61[17] , \wPDiag_42[26] , 
        \wNDiag_60[44] , \wColumn_29[7] , \wNDiag_56[58] , \wNDiag_56[41] , 
        \wPDiag_57[12] , \wNDiag_29[44] , \wColumn_34[8] , \wPDiag_2[16] , 
        \wColumn_17[62] , \wNDiag_25[0] , \wPDiag_28[17] , \wPDiag_48[13] , 
        \wNDiag_49[59] , \wNDiag_49[40] , \wColumn_54[57] , \wNDiag_26[3] , 
        \wColumn_34[53] , \wColumn_62[52] , \wColumn_41[63] , \wColumn_29[31] , 
        \wColumn_49[35] , \wPDiag_4[4] , \wPDiag_16[44] , \wNDiag_17[17] , 
        \wColumn_29[28] , \wPDiag_40[45] , \wNDiag_62[27] , \wColumn_17[51] , 
        \wPDiag_20[58] , \wNDiag_21[12] , \wNDiag_34[26] , \wNDiag_41[16] , 
        \wPDiag_20[41] , \wNDiag_54[22] , \wColumn_41[49] , \wColumn_62[61] , 
        \wColumn_17[48] , \wColumn_41[50] , \wNDiag_41[4] , \wColumn_21[54] , 
        \wColumn_34[60] , \wColumn_1[37] , \wScan_2[0] , \wPDiag_14[9] , 
        \wColumn_46[8] , \wPDiag_48[39] , \wPDiag_48[20] , \wNDiag_21[38] , 
        \wNDiag_21[21] , \wPDiag_28[24] , \wNDiag_54[11] , \wPDiag_55[42] , 
        \wPDiag_2[25] , \wPDiag_7[7] , \wNDiag_17[24] , \wPDiag_35[46] , 
        \wNDiag_62[14] , \wNDiag_34[15] , \wNDiag_41[25] , \wPDiag_63[47] , 
        \wNDiag_42[7] , \wNDiag_4[55] , \wNDiag_7[16] , \wColumn_58[4] , 
        \wColumn_9[61] , \wPDiag_15[34] , \wColumn_24[2] , \wNDiag_37[56] , 
        \wScan_16[3] , \wNDiag_61[57] , \wPDiag_23[31] , \wPDiag_43[35] , 
        \wNDiag_22[62] , \wPDiag_23[28] , \wPDiag_56[18] , \wNDiag_57[52] , 
        \wPDiag_1[55] , \wColumn_9[52] , \wPDiag_9[30] , \wScan_15[0] , 
        \wPDiag_9[29] , \wColumn_22[17] , \wColumn_14[12] , \wColumn_37[23] , 
        \wColumn_57[27] , \wColumn_42[13] , \wColumn_27[1] , \wPDiag_56[32] , 
        \wColumn_61[22] , \wNDiag_14[54] , \wNDiag_22[51] , \wNDiag_22[48] , 
        \wNDiag_57[61] , \wNDiag_42[55] , \wPDiag_60[37] , \wPDiag_36[36] , 
        \wPDiag_1[9] , \wNDiag_7[25] , \wPDiag_11[4] , \wPDiag_12[7] , 
        \wColumn_14[38] , \wReturn_35[0] , \wColumn_40[6] , \wColumn_37[10] , 
        \wColumn_42[20] , \wColumn_14[21] , \wColumn_42[39] , \wNDiag_59[6] , 
        \wColumn_61[11] , \wColumn_22[24] , \wColumn_43[5] , \wColumn_57[14] , 
        \wNDiag_44[9] , \wNDiag_3[14] , \wColumn_5[35] , \wColumn_10[10] , 
        \wColumn_33[21] , \wColumn_46[11] , \wNDiag_18[33] , \wPDiag_19[60] , 
        \wColumn_26[15] , \wColumn_33[38] , \wPDiag_35[2] , \wColumn_53[25] , 
        \wPDiag_11[36] , \wNDiag_26[60] , \wPDiag_27[33] , \wScan_55[2] , 
        \wNDiag_53[49] , \wNDiag_33[54] , \wNDiag_53[50] , \wPDiag_36[1] , 
        \wPDiag_47[37] , \wScan_56[1] , \wColumn_18[46] , \wNDiag_18[19] , 
        \wPDiag_19[53] , \wScan_31[6] , \wCall_37[0] , \wPDiag_51[6] , 
        \wColumn_53[16] , \wNDiag_3[27] , \wColumn_10[23] , \wNDiag_19[4] , 
        \wColumn_26[26] , \wColumn_33[12] , \wColumn_46[22] , \wPDiag_5[57] , 
        \wPDiag_52[5] , \wNDiag_46[57] , \wColumn_1[27] , \wColumn_1[14] , 
        \wPDiag_1[45] , \wPDiag_2[3] , \wNDiag_5[4] , \wColumn_6[45] , 
        \wPDiag_6[14] , \wNDiag_10[56] , \wPDiag_12[46] , \wNDiag_13[15] , 
        \wPDiag_24[43] , \wNDiag_25[10] , \wNDiag_26[53] , \wPDiag_27[19] , 
        \wScan_32[5] , \wPDiag_32[34] , \wPDiag_52[30] , \wPDiag_52[29] , 
        \wNDiag_53[63] , \wNDiag_50[20] , \wNDiag_50[39] , \wPDiag_44[47] , 
        \wNDiag_30[24] , \wNDiag_45[14] , \wNDiag_8[32] , \wColumn_13[60] , 
        \wColumn_30[48] , \wColumn_30[51] , \wPDiag_39[38] , \wPDiag_39[21] , 
        \wColumn_45[61] , \wColumn_50[55] , \wPDiag_59[25] , \wPDiag_6[27] , 
        \wColumn_18[6] , \wColumn_38[34] , \wColumn_58[30] , \wNDiag_6[7] , 
        \wColumn_58[29] , \wNDiag_13[26] , \wPDiag_31[44] , \wNDiag_25[23] , 
        \wNDiag_30[17] , \wNDiag_45[27] , \wNDiag_50[13] , \wPDiag_57[8] , 
        \wPDiag_51[59] , \wPDiag_51[40] , \wNDiag_58[45] , \wNDiag_8[18] , 
        \wColumn_25[56] , \wScan_29[4] , \wNDiag_38[58] , \wPDiag_59[16] , 
        \wNDiag_38[41] , \wPDiag_39[12] , \wPDiag_49[4] , \wColumn_13[53] , 
        \wNDiag_14[44] , \wColumn_30[62] , \wColumn_45[52] , \wPDiag_36[26] , 
        \wPDiag_43[16] , \wPDiag_15[17] , \wNDiag_42[45] , \wPDiag_60[27] , 
        \wNDiag_7[35] , \wColumn_9[42] , \wNDiag_22[41] , \wNDiag_47[3] , 
        \wPDiag_56[22] , \wNDiag_22[58] , \wPDiag_23[12] , \wScan_7[4] , 
        \wPDiag_9[13] , \wColumn_22[34] , \wColumn_14[31] , \wColumn_42[29] , 
        \wColumn_14[28] , \wColumn_37[19] , \wColumn_42[30] , \wColumn_61[18] , 
        \wPDiag_1[0] , \wNDiag_44[0] , \wPDiag_15[24] , \wPDiag_23[38] , 
        \wPDiag_23[21] , \wColumn_39[4] , \wNDiag_57[42] , \wNDiag_23[7] , 
        \wPDiag_36[15] , \wPDiag_56[11] , \wPDiag_43[25] , \wNDiag_61[47] , 
        \wNDiag_20[4] , \wNDiag_37[46] , \wPDiag_60[14] , \wColumn_2[57] , 
        \wPDiag_2[35] , \wNDiag_4[45] , \wPDiag_9[39] , \wColumn_27[8] , 
        \wColumn_37[33] , \wColumn_61[32] , \wPDiag_9[20] , \wColumn_57[37] , 
        \wPDiag_14[0] , \wColumn_17[58] , \wColumn_21[44] , \wColumn_41[40] , 
        \wColumn_17[41] , \wColumn_41[59] , \wPDiag_28[34] , \wPDiag_17[3] , 
        \wNDiag_41[35] , \wColumn_46[1] , \wPDiag_48[30] , \wPDiag_48[29] , 
        \wNDiag_49[63] , \wPDiag_63[57] , \wNDiag_17[34] , \wPDiag_20[62] , 
        \wPDiag_35[56] , \wColumn_45[2] , \wNDiag_54[18] , \wPDiag_55[52] , 
        \wNDiag_21[31] , \wNDiag_21[28] , \wColumn_49[16] , \wColumn_22[5] , 
        \wColumn_29[12] , \wNDiag_49[50] , \wNDiag_49[49] , \wNDiag_38[6] , 
        \wColumn_5[16] , \wColumn_6[55] , \wPDiag_6[37] , \wScan_10[4] , 
        \wNDiag_25[9] , \wNDiag_29[54] , \wReturn_54[0] , \wColumn_34[43] , 
        \wColumn_62[42] , \wPDiag_16[54] , \wPDiag_20[51] , \wColumn_29[38] , 
        \wColumn_54[47] , \wColumn_29[21] , \wColumn_49[25] , \wPDiag_20[48] , 
        \wColumn_21[6] , \wPDiag_55[61] , \wNDiag_34[36] , \wNDiag_54[32] , 
        \wPDiag_40[55] , \wNDiag_62[37] , \wNDiag_8[22] , \wNDiag_8[11] , 
        \wColumn_9[3] , \wNDiag_13[36] , \wPDiag_24[60] , \wScan_37[1] , 
        \wColumn_58[39] , \wColumn_38[24] , \wColumn_58[20] , \wPDiag_51[50] , 
        \wNDiag_25[33] , \wPDiag_51[49] , \wNDiag_45[37] , \wPDiag_31[54] , 
        \wPDiag_57[1] , \wNDiag_38[51] , \wNDiag_38[48] , \wPDiag_54[2] , 
        \wNDiag_58[55] , \wPDiag_12[56] , \wColumn_13[43] , \wScan_34[2] , 
        \wColumn_45[42] , \wColumn_25[46] , \wNDiag_30[34] , \wPDiag_24[53] , 
        \wNDiag_25[19] , \wPDiag_44[57] , \wColumn_30[41] , \wPDiag_33[5] , 
        \wNDiag_50[29] , \wPDiag_51[63] , \wColumn_61[4] , \wColumn_38[17] , 
        \wNDiag_50[30] , \wScan_50[6] , \wScan_53[5] , \wColumn_58[13] , 
        \wColumn_50[45] , \wColumn_30[58] , \wPDiag_59[35] , \wNDiag_18[10] , 
        \wPDiag_30[6] , \wNDiag_38[62] , \wPDiag_39[28] , \wPDiag_39[31] , 
        \wCall_56[0] , \wColumn_62[7] , \wPDiag_19[43] , \wColumn_10[33] , 
        \wColumn_46[32] , \wNDiag_3[37] , \wNDiag_3[3] , \wPDiag_5[47] , 
        \wColumn_26[36] , \wNDiag_26[43] , \wPDiag_52[39] , \wPDiag_27[10] , 
        \wPDiag_52[20] , \wPDiag_32[24] , \wPDiag_47[14] , \wNDiag_10[46] , 
        \wPDiag_11[15] , \wNDiag_46[47] , \wColumn_53[35] , \wNDiag_1[54] , 
        \wColumn_4[6] , \wColumn_5[25] , \wColumn_10[19] , \wColumn_33[31] , 
        \wColumn_33[28] , \wScan_48[4] , \wColumn_46[18] , \wNDiag_60[6] , 
        \wColumn_7[46] , \wPDiag_11[26] , \wNDiag_18[23] , \wPDiag_28[4] , 
        \wPDiag_32[17] , \wPDiag_47[27] , \wNDiag_63[5] , \wColumn_18[56] , 
        \wPDiag_27[23] , \wNDiag_33[44] , \wNDiag_53[40] , \wPDiag_52[13] , 
        \wNDiag_53[59] , \wPDiag_36[8] , \wPDiag_58[26] , \wPDiag_7[17] , 
        \wNDiag_9[31] , \wColumn_31[52] , \wPDiag_38[22] , \wColumn_51[56] , 
        \wNDiag_9[28] , \wColumn_12[63] , \wColumn_44[62] , \wColumn_59[19] , 
        \wNDiag_11[5] , \wNDiag_12[16] , \wPDiag_13[45] , \wNDiag_31[27] , 
        \wNDiag_44[17] , \wNDiag_24[13] , \wPDiag_25[59] , \wPDiag_25[40] , 
        \wPDiag_45[44] , \wColumn_44[51] , \wNDiag_51[23] , \wColumn_12[50] , 
        \wColumn_12[49] , \wColumn_31[61] , \wColumn_44[48] , \wPDiag_7[24] , 
        \wNDiag_8[8] , \wNDiag_12[25] , \wColumn_16[9] , \wColumn_24[55] , 
        \wPDiag_38[11] , \wNDiag_39[42] , \wPDiag_59[7] , \wPDiag_58[15] , 
        \wNDiag_24[39] , \wPDiag_44[8] , \wNDiag_59[46] , \wPDiag_50[43] , 
        \wNDiag_24[20] , \wNDiag_51[10] , \wPDiag_30[47] , \wNDiag_31[14] , 
        \wNDiag_44[24] , \wNDiag_12[6] , \wColumn_39[37] , \wColumn_59[33] , 
        \wColumn_2[8] , \wNDiag_2[17] , \wColumn_7[5] , \wColumn_19[45] , 
        \wColumn_4[36] , \wPDiag_10[35] , \wPDiag_26[2] , \wNDiag_32[57] , 
        \wScan_46[2] , \wPDiag_46[34] , \wPDiag_26[30] , \wPDiag_26[29] , 
        \wNDiag_27[63] , \wNDiag_52[53] , \wPDiag_53[19] , \wColumn_11[13] , 
        \wPDiag_18[63] , \wNDiag_19[30] , \wScan_45[1] , \wNDiag_19[29] , 
        \wColumn_27[16] , \wColumn_52[26] , \wNDiag_11[55] , \wScan_22[6] , 
        \wPDiag_25[1] , \wNDiag_27[50] , \wColumn_32[22] , \wColumn_47[12] , 
        \wNDiag_52[60] , \wNDiag_27[49] , \wPDiag_53[33] , \wPDiag_33[37] , 
        \wNDiag_47[54] , \wNDiag_2[24] , \wPDiag_4[54] , \wColumn_10[7] , 
        \wCall_24[0] , \wPDiag_42[6] , \wNDiag_6[15] , \wColumn_8[62] , 
        \wPDiag_8[33] , \wColumn_11[39] , \wColumn_11[20] , \wColumn_47[38] , 
        \wColumn_32[11] , \wColumn_47[21] , \wColumn_13[4] , \wColumn_27[25] , 
        \wColumn_52[15] , \wPDiag_41[5] , \wNDiag_14[8] , \wColumn_15[11] , 
        \wPDiag_18[50] , \wPDiag_18[49] , \wScan_21[5] , \wColumn_23[14] , 
        \wColumn_36[39] , \wColumn_36[20] , \wColumn_37[2] , \wColumn_60[21] , 
        \wColumn_43[10] , \wColumn_60[38] , \wColumn_56[24] , \wPDiag_22[32] , 
        \wNDiag_23[61] , \wNDiag_56[51] , \wNDiag_56[48] , \wPDiag_14[37] , 
        \wNDiag_36[55] , \wPDiag_42[36] , \wNDiag_60[54] , \wColumn_34[1] , 
        \wColumn_3[44] , \wPDiag_3[15] , \wNDiag_6[26] , \wPDiag_8[19] , 
        \wScan_9[2] , \wColumn_56[17] , \wColumn_15[22] , \wColumn_23[27] , 
        \wNDiag_49[5] , \wColumn_53[6] , \wColumn_60[12] , \wColumn_36[13] , 
        \wColumn_43[23] , \wColumn_50[5] , \wColumn_8[51] , \wColumn_8[48] , 
        \wNDiag_15[57] , \wReturn_26[0] , \wPDiag_37[35] , \wNDiag_43[56] , 
        \wNDiag_56[62] , \wPDiag_57[28] , \wPDiag_61[34] , \wPDiag_22[18] , 
        \wNDiag_23[52] , \wPDiag_57[31] , \wNDiag_16[14] , \wPDiag_17[47] , 
        \wNDiag_20[11] , \wPDiag_21[42] , \wNDiag_57[9] , \wScan_62[4] , 
        \wNDiag_55[38] , \wNDiag_55[21] , \wNDiag_35[25] , \wNDiag_40[15] , 
        \wPDiag_41[46] , \wNDiag_63[24] , \wColumn_16[61] , \wColumn_28[32] , 
        \wColumn_35[50] , \wNDiag_36[0] , \wColumn_48[36] , \wColumn_35[49] , 
        \wColumn_40[60] , \wColumn_63[48] , \wNDiag_35[3] , \wColumn_63[51] , 
        \wNDiag_48[43] , \wColumn_55[54] , \wPDiag_49[10] , \wPDiag_3[26] , 
        \wNDiag_5[56] , \wNDiag_28[47] , \wPDiag_29[14] , \wColumn_28[18] , 
        \wColumn_48[7] , \wNDiag_3[10] , \wNDiag_5[0] , \wColumn_6[58] , 
        \wColumn_6[41] , \wPDiag_9[8] , \wNDiag_16[27] , \wPDiag_34[45] , 
        \wNDiag_35[16] , \wNDiag_40[26] , \wNDiag_52[4] , \wPDiag_62[44] , 
        \wColumn_55[8] , \wNDiag_63[17] , \wNDiag_20[22] , \wPDiag_54[58] , 
        \wPDiag_54[41] , \wNDiag_55[12] , \wPDiag_29[27] , \wColumn_16[52] , 
        \wPDiag_19[5] , \wPDiag_49[23] , \wColumn_20[57] , \wColumn_35[63] , 
        \wColumn_40[53] , \wNDiag_51[7] , \wColumn_63[62] , \wPDiag_59[21] , 
        \wPDiag_59[38] , \wPDiag_6[10] , \wNDiag_8[36] , \wColumn_25[61] , 
        \wPDiag_39[25] , \wColumn_50[48] , \wColumn_30[55] , \wColumn_50[51] , 
        \wPDiag_12[42] , \wColumn_13[57] , \wNDiag_13[11] , \wNDiag_30[20] , 
        \wNDiag_45[10] , \wPDiag_24[47] , \wNDiag_30[39] , \wPDiag_44[43] , 
        \wNDiag_25[14] , \wPDiag_33[8] , \wColumn_45[56] , \wNDiag_50[24] , 
        \wColumn_61[9] , \wColumn_25[52] , \wColumn_50[62] , \wScan_29[0] , 
        \wNDiag_38[45] , \wPDiag_49[0] , \wPDiag_39[16] , \wPDiag_6[23] , 
        \wNDiag_6[3] , \wNDiag_25[27] , \wNDiag_50[17] , \wPDiag_51[44] , 
        \wNDiag_58[58] , \wNDiag_58[41] , \wPDiag_59[12] , \wNDiag_30[13] , 
        \wNDiag_45[23] , \wPDiag_31[59] , \wNDiag_13[22] , \wPDiag_31[40] , 
        \wColumn_18[42] , \wColumn_18[2] , \wColumn_38[30] , \wColumn_58[34] , 
        \wColumn_38[29] , \wColumn_5[31] , \wColumn_5[28] , \wPDiag_5[60] , 
        \wNDiag_10[61] , \wNDiag_33[49] , \wPDiag_36[5] , \wNDiag_63[8] , 
        \wPDiag_11[32] , \wNDiag_33[50] , \wPDiag_47[33] , \wScan_56[5] , 
        \wPDiag_27[37] , \wNDiag_46[60] , \wNDiag_53[54] , \wColumn_10[14] , 
        \wNDiag_18[37] , \wPDiag_28[9] , \wScan_55[6] , \wColumn_26[11] , 
        \wCall_53[0] , \wColumn_53[38] , \wColumn_53[21] , \wNDiag_10[52] , 
        \wPDiag_11[18] , \wNDiag_26[57] , \wColumn_33[25] , \wPDiag_35[6] , 
        \wColumn_46[15] , \wScan_32[1] , \wPDiag_52[34] , \wPDiag_32[30] , 
        \wPDiag_32[29] , \wNDiag_33[63] , \wNDiag_46[53] , \wPDiag_47[19] , 
        \wColumn_1[33] , \wNDiag_3[23] , \wPDiag_5[53] , \wPDiag_52[1] , 
        \wPDiag_9[34] , \wColumn_10[27] , \wNDiag_19[0] , \wColumn_14[16] , 
        \wPDiag_19[57] , \wColumn_26[22] , \wColumn_33[16] , \wColumn_46[26] , 
        \wColumn_53[12] , \wScan_31[2] , \wPDiag_51[2] , \wColumn_22[13] , 
        \wColumn_27[5] , \wColumn_37[27] , \wColumn_61[26] , \wColumn_42[17] , 
        \wReturn_51[0] , \wColumn_57[23] , \wNDiag_20[9] , \wColumn_1[19] , 
        \wPDiag_1[62] , \wNDiag_14[63] , \wScan_15[4] , \wPDiag_23[35] , 
        \wNDiag_57[56] , \wColumn_39[9] , \wPDiag_15[30] , \wPDiag_15[29] , 
        \wPDiag_36[18] , \wPDiag_43[31] , \wPDiag_60[19] , \wNDiag_61[53] , 
        \wNDiag_37[52] , \wNDiag_42[62] , \wPDiag_43[28] , \wNDiag_7[12] , 
        \wColumn_24[6] , \wPDiag_1[51] , \wPDiag_1[48] , \wNDiag_7[38] , 
        \wPDiag_11[0] , \wColumn_22[39] , \wColumn_22[20] , \wColumn_57[10] , 
        \wPDiag_12[3] , \wColumn_14[25] , \wColumn_43[1] , \wNDiag_59[2] , 
        \wColumn_61[15] , \wColumn_37[14] , \wColumn_42[24] , \wColumn_40[2] , 
        \wNDiag_7[21] , \wScan_2[4] , \wColumn_2[43] , \wPDiag_2[12] , 
        \wColumn_9[56] , \wNDiag_14[50] , \wNDiag_42[48] , \wNDiag_61[60] , 
        \wNDiag_14[49] , \wPDiag_36[32] , \wNDiag_42[51] , \wPDiag_60[33] , 
        \wNDiag_22[55] , \wNDiag_37[61] , \wPDiag_56[36] , \wPDiag_16[59] , 
        \wPDiag_16[40] , \wPDiag_20[45] , \wNDiag_21[16] , \wNDiag_54[26] , 
        \wNDiag_17[13] , \wNDiag_34[22] , \wPDiag_40[58] , \wNDiag_41[12] , 
        \wPDiag_40[41] , \wNDiag_62[23] , \wNDiag_4[62] , \wColumn_29[35] , 
        \wColumn_21[63] , \wNDiag_25[4] , \wNDiag_26[7] , \wColumn_49[31] , 
        \wColumn_34[57] , \wColumn_49[28] , \wColumn_62[56] , \wColumn_22[8] , 
        \wNDiag_49[44] , \wColumn_54[53] , \wPDiag_48[17] , \wPDiag_2[38] , 
        \wPDiag_2[21] , \wNDiag_4[51] , \wPDiag_28[13] , \wNDiag_29[59] , 
        \wNDiag_29[40] , \wNDiag_4[48] , \wColumn_58[0] , \wNDiag_42[3] , 
        \wPDiag_7[3] , \wNDiag_17[39] , \wNDiag_34[11] , \wNDiag_41[21] , 
        \wPDiag_63[43] , \wNDiag_17[20] , \wPDiag_35[42] , \wNDiag_41[38] , 
        \wNDiag_62[10] , \wPDiag_55[46] , \wPDiag_4[0] , \wColumn_21[50] , 
        \wColumn_21[49] , \wNDiag_21[25] , \wNDiag_54[15] , \wPDiag_28[39] , 
        \wPDiag_28[20] , \wPDiag_48[24] , \wColumn_54[60] , \wNDiag_6[32] , 
        \wColumn_8[45] , \wPDiag_14[10] , \wNDiag_15[43] , \wColumn_17[55] , 
        \wColumn_41[54] , \wNDiag_41[0] , \wPDiag_37[21] , \wPDiag_42[11] , 
        \wPDiag_61[39] , \wPDiag_37[38] , \wNDiag_43[42] , \wPDiag_61[20] , 
        \wNDiag_23[46] , \wNDiag_57[4] , \wPDiag_57[25] , \wPDiag_22[15] , 
        \wPDiag_8[14] , \wColumn_23[33] , \wColumn_50[8] , \wColumn_15[36] , 
        \wColumn_43[37] , \wNDiag_49[8] , \wNDiag_54[7] , \wColumn_1[6] , 
        \wNDiag_1[59] , \wNDiag_1[40] , \wColumn_3[63] , \wNDiag_6[18] , 
        \wPDiag_8[27] , \wPDiag_14[23] , \wPDiag_22[26] , \wColumn_29[3] , 
        \wNDiag_56[45] , \wNDiag_33[0] , \wNDiag_36[58] , \wPDiag_57[16] , 
        \wPDiag_37[12] , \wPDiag_42[22] , \wNDiag_60[40] , \wScan_18[1] , 
        \wNDiag_30[3] , \wNDiag_36[41] , \wNDiag_60[59] , \wPDiag_61[13] , 
        \wColumn_36[34] , \wColumn_60[35] , \wColumn_56[30] , \wColumn_16[46] , 
        \wPDiag_19[8] , \wColumn_23[19] , \wColumn_56[29] , \wColumn_20[43] , 
        \wColumn_40[47] , \wPDiag_29[33] , \wColumn_56[6] , \wColumn_3[50] , 
        \wPDiag_3[32] , \wNDiag_5[42] , \wPDiag_9[5] , \wNDiag_28[60] , 
        \wNDiag_16[33] , \wPDiag_17[60] , \wNDiag_40[32] , \wPDiag_49[37] , 
        \wPDiag_62[50] , \wPDiag_34[48] , \wPDiag_41[61] , \wPDiag_62[49] , 
        \wNDiag_20[36] , \wReturn_23[0] , \wPDiag_34[51] , \wColumn_55[5] , 
        \wPDiag_54[55] , \wColumn_48[11] , \wColumn_28[15] , \wNDiag_52[9] , 
        \wNDiag_28[1] , \wColumn_32[2] , \wNDiag_48[57] , \wPDiag_60[3] , 
        \wColumn_3[49] , \wPDiag_3[18] , \wColumn_28[26] , \wNDiag_28[53] , 
        \wPDiag_29[19] , \wColumn_35[44] , \wColumn_55[59] , \wColumn_63[45] , 
        \wColumn_55[40] , \wColumn_7[8] , \wPDiag_7[30] , \wNDiag_16[19] , 
        \wPDiag_17[53] , \wPDiag_21[56] , \wColumn_48[22] , \wColumn_31[1] , 
        \wNDiag_35[31] , \wNDiag_55[35] , \wPDiag_63[0] , \wPDiag_34[62] , 
        \wNDiag_35[28] , \wPDiag_62[63] , \wNDiag_63[29] , \wNDiag_40[18] , 
        \wPDiag_41[52] , \wNDiag_63[30] , \wPDiag_7[29] , \wScan_27[6] , 
        \wColumn_59[27] , \wColumn_39[23] , \wColumn_7[61] , \wNDiag_12[31] , 
        \wNDiag_12[28] , \wNDiag_24[34] , \wPDiag_50[57] , \wNDiag_44[30] , 
        \wPDiag_13[62] , \wCall_21[0] , \wNDiag_44[29] , \wPDiag_45[63] , 
        \wColumn_15[7] , \wPDiag_30[53] , \wPDiag_47[6] , \wColumn_16[4] , 
        \wNDiag_31[19] , \wNDiag_39[56] , \wPDiag_44[5] , \wColumn_7[52] , 
        \wNDiag_8[5] , \wNDiag_9[16] , \wPDiag_58[18] , \wNDiag_59[52] , 
        \wNDiag_11[8] , \wColumn_44[45] , \wColumn_12[44] , \wScan_24[5] , 
        \wColumn_24[58] , \wNDiag_9[25] , \wPDiag_13[51] , \wColumn_24[41] , 
        \wNDiag_31[33] , \wPDiag_13[48] , \wPDiag_30[60] , \wPDiag_45[49] , 
        \wPDiag_23[2] , \wPDiag_25[54] , \wPDiag_45[50] , \wColumn_31[46] , 
        \wColumn_39[10] , \wNDiag_51[37] , \wScan_40[1] , \wScan_43[2] , 
        \wColumn_59[14] , \wColumn_51[42] , \wPDiag_58[32] , \wNDiag_14[5] , 
        \wNDiag_19[17] , \wPDiag_20[1] , \wPDiag_38[36] , \wNDiag_59[61] , 
        \wPDiag_18[44] , \wColumn_2[5] , \wNDiag_2[30] , \wNDiag_2[29] , 
        \wColumn_4[11] , \wPDiag_4[59] , \wColumn_11[34] , \wColumn_13[9] , 
        \wColumn_27[31] , \wColumn_47[35] , \wColumn_27[28] , \wPDiag_41[8] , 
        \wColumn_52[18] , \wPDiag_4[40] , \wColumn_19[62] , \wNDiag_17[6] , 
        \wPDiag_26[17] , \wNDiag_27[44] , \wPDiag_53[27] , \wColumn_3[59] , 
        \wColumn_4[22] , \wPDiag_10[12] , \wNDiag_11[58] , \wNDiag_11[41] , 
        \wPDiag_33[23] , \wPDiag_46[13] , \wNDiag_47[59] , \wNDiag_47[40] , 
        \wColumn_32[36] , \wColumn_52[32] , \wScan_58[3] , \wPDiag_10[38] , 
        \wNDiag_19[24] , \wPDiag_38[3] , \wPDiag_10[21] , \wPDiag_33[10] , 
        \wPDiag_46[20] , \wColumn_19[51] , \wPDiag_26[24] , \wNDiag_32[43] , 
        \wPDiag_46[39] , \wNDiag_52[47] , \wPDiag_53[14] , \wColumn_19[48] , 
        \wNDiag_28[8] , \wColumn_3[40] , \wNDiag_28[43] , \wPDiag_3[22] , 
        \wPDiag_3[11] , \wNDiag_5[61] , \wColumn_20[60] , \wPDiag_29[10] , 
        \wNDiag_48[47] , \wPDiag_49[14] , \wColumn_35[54] , \wNDiag_35[7] , 
        \wColumn_55[50] , \wColumn_55[49] , \wColumn_63[55] , \wCall_18[0] , 
        \wNDiag_36[4] , \wColumn_48[32] , \wColumn_28[36] , \wReturn_7[0] , 
        \wColumn_16[56] , \wNDiag_16[10] , \wPDiag_17[43] , \wNDiag_35[38] , 
        \wPDiag_41[42] , \wNDiag_63[20] , \wNDiag_20[15] , \wNDiag_35[21] , 
        \wNDiag_40[11] , \wNDiag_63[39] , \wPDiag_21[46] , \wColumn_31[8] , 
        \wPDiag_63[9] , \wNDiag_55[25] , \wPDiag_19[1] , \wColumn_40[57] , 
        \wNDiag_51[3] , \wColumn_55[63] , \wColumn_20[53] , \wNDiag_20[26] , 
        \wPDiag_29[23] , \wPDiag_49[27] , \wNDiag_55[16] , \wPDiag_54[45] , 
        \wNDiag_16[23] , \wPDiag_34[41] , \wPDiag_62[59] , \wNDiag_63[13] , 
        \wPDiag_34[58] , \wNDiag_40[22] , \wPDiag_62[40] , \wNDiag_35[12] , 
        \wNDiag_52[0] , \wNDiag_5[52] , \wColumn_48[18] , \wNDiag_6[22] , 
        \wNDiag_6[11] , \wReturn_42[0] , \wColumn_48[3] , \wColumn_8[55] , 
        \wPDiag_8[37] , \wPDiag_14[33] , \wColumn_34[5] , \wNDiag_36[51] , 
        \wNDiag_15[60] , \wNDiag_33[9] , \wNDiag_43[61] , \wNDiag_60[49] , 
        \wNDiag_36[48] , \wPDiag_22[36] , \wPDiag_42[32] , \wNDiag_60[50] , 
        \wNDiag_56[55] , \wColumn_15[15] , \wColumn_23[10] , \wColumn_56[39] , 
        \wColumn_36[24] , \wColumn_56[20] , \wColumn_43[14] , \wColumn_37[6] , 
        \wPDiag_57[35] , \wColumn_60[25] , \wPDiag_14[19] , \wNDiag_15[53] , 
        \wNDiag_23[56] , \wScan_62[0] , \wNDiag_36[62] , \wPDiag_37[28] , 
        \wPDiag_42[18] , \wNDiag_43[52] , \wPDiag_61[30] , \wNDiag_60[63] , 
        \wPDiag_61[29] , \wPDiag_37[31] , \wScan_9[6] , \wColumn_15[26] , 
        \wColumn_36[17] , \wColumn_43[27] , \wColumn_50[1] , \wNDiag_49[1] , 
        \wColumn_60[16] , \wColumn_23[23] , \wColumn_53[2] , \wColumn_56[13] , 
        \wNDiag_1[63] , \wNDiag_2[39] , \wNDiag_2[20] , \wNDiag_2[13] , 
        \wColumn_4[32] , \wColumn_11[17] , \wColumn_32[26] , \wScan_61[3] , 
        \wColumn_47[16] , \wNDiag_19[34] , \wPDiag_25[5] , \wColumn_27[12] , 
        \wColumn_52[22] , \wPDiag_4[63] , \wPDiag_10[31] , \wPDiag_26[34] , 
        \wScan_45[5] , \wNDiag_32[53] , \wNDiag_52[57] , \wPDiag_33[19] , 
        \wPDiag_10[28] , \wPDiag_46[29] , \wNDiag_47[63] , \wNDiag_11[62] , 
        \wCall_40[0] , \wScan_46[6] , \wPDiag_46[30] , \wPDiag_26[6] , 
        \wColumn_4[18] , \wColumn_19[58] , \wColumn_19[41] , \wColumn_11[24] , 
        \wColumn_13[0] , \wPDiag_18[54] , \wScan_21[1] , \wColumn_27[38] , 
        \wPDiag_41[1] , \wColumn_27[21] , \wColumn_52[11] , \wColumn_32[15] , 
        \wColumn_47[25] , \wPDiag_42[2] , \wPDiag_4[50] , \wColumn_10[3] , 
        \wPDiag_4[49] , \wPDiag_7[13] , \wNDiag_11[51] , \wNDiag_11[48] , 
        \wNDiag_47[50] , \wNDiag_32[60] , \wNDiag_47[49] , \wNDiag_12[12] , 
        \wPDiag_13[58] , \wScan_22[2] , \wPDiag_33[33] , \wPDiag_53[37] , 
        \wNDiag_24[17] , \wNDiag_27[54] , \wPDiag_25[44] , \wNDiag_51[27] , 
        \wPDiag_13[41] , \wPDiag_45[40] , \wNDiag_31[23] , \wNDiag_44[13] , 
        \wPDiag_45[59] , \wColumn_39[19] , \wNDiag_1[50] , \wNDiag_1[49] , 
        \wColumn_7[42] , \wNDiag_9[35] , \wColumn_31[56] , \wPDiag_20[8] , 
        \wColumn_24[62] , \wPDiag_38[26] , \wColumn_51[52] , \wPDiag_58[22] , 
        \wColumn_7[1] , \wColumn_39[33] , \wNDiag_3[33] , \wColumn_4[2] , 
        \wPDiag_7[39] , \wNDiag_12[2] , \wPDiag_7[20] , \wColumn_59[37] , 
        \wNDiag_12[38] , \wNDiag_12[21] , \wPDiag_30[43] , \wNDiag_44[39] , 
        \wNDiag_31[10] , \wNDiag_44[20] , \wColumn_24[51] , \wNDiag_24[24] , 
        \wNDiag_51[14] , \wPDiag_38[15] , \wPDiag_50[47] , \wPDiag_58[11] , 
        \wNDiag_59[42] , \wScan_39[3] , \wNDiag_39[46] , \wColumn_51[61] , 
        \wPDiag_59[3] , \wNDiag_10[42] , \wPDiag_11[11] , \wNDiag_11[1] , 
        \wColumn_12[54] , \wColumn_24[48] , \wColumn_44[55] , \wPDiag_32[39] , 
        \wNDiag_46[43] , \wPDiag_32[20] , \wPDiag_47[10] , \wNDiag_26[47] , 
        \wPDiag_27[14] , \wPDiag_52[24] , \wNDiag_3[7] , \wPDiag_52[8] , 
        \wPDiag_5[43] , \wColumn_18[61] , \wNDiag_3[19] , \wColumn_5[12] , 
        \wColumn_10[37] , \wNDiag_19[9] , \wColumn_26[32] , \wColumn_46[36] , 
        \wNDiag_18[14] , \wPDiag_19[47] , \wColumn_5[38] , \wColumn_5[21] , 
        \wPDiag_11[22] , \wColumn_18[52] , \wPDiag_27[27] , \wPDiag_52[17] , 
        \wNDiag_53[44] , \wNDiag_63[1] , \wNDiag_18[27] , \wPDiag_28[0] , 
        \wPDiag_32[13] , \wNDiag_33[40] , \wNDiag_33[59] , \wPDiag_47[23] , 
        \wNDiag_60[2] , \wColumn_26[18] , \wColumn_33[35] , \wColumn_53[31] , 
        \wColumn_53[28] , \wColumn_1[23] , \wColumn_1[10] , \wPDiag_1[4] , 
        \wColumn_2[60] , \wPDiag_2[31] , \wPDiag_2[28] , \wNDiag_5[9] , 
        \wNDiag_8[15] , \wColumn_13[47] , \wColumn_25[42] , \wScan_48[0] , 
        \wScan_34[6] , \wPDiag_49[9] , \wColumn_9[7] , \wColumn_45[46] , 
        \wColumn_6[62] , \wCall_32[0] , \wNDiag_58[51] , \wPDiag_54[6] , 
        \wNDiag_58[48] , \wColumn_6[51] , \wColumn_6[48] , \wPDiag_6[33] , 
        \wPDiag_12[61] , \wNDiag_13[32] , \wNDiag_38[55] , \wPDiag_44[60] , 
        \wPDiag_31[50] , \wPDiag_57[5] , \wNDiag_45[33] , \wNDiag_25[37] , 
        \wPDiag_31[49] , \wColumn_38[39] , \wPDiag_51[54] , \wColumn_38[20] , 
        \wColumn_58[24] , \wPDiag_30[2] , \wScan_37[5] , \wPDiag_39[35] , 
        \wColumn_62[3] , \wNDiag_58[62] , \wPDiag_59[28] , \wPDiag_59[31] , 
        \wPDiag_6[19] , \wNDiag_8[26] , \wColumn_30[45] , \wScan_50[2] , 
        \wColumn_50[58] , \wColumn_50[41] , \wColumn_58[17] , \wPDiag_12[52] , 
        \wNDiag_13[18] , \wPDiag_24[57] , \wColumn_38[13] , \wScan_53[1] , 
        \wNDiag_50[34] , \wNDiag_30[30] , \wNDiag_30[29] , \wPDiag_31[63] , 
        \wPDiag_33[1] , \wColumn_61[0] , \wPDiag_44[53] , \wNDiag_45[19] , 
        \wColumn_29[16] , \wNDiag_4[58] , \wNDiag_4[41] , \wColumn_58[9] , 
        \wPDiag_14[4] , \wPDiag_16[63] , \wPDiag_17[7] , \wNDiag_21[35] , 
        \wColumn_49[12] , \wPDiag_40[62] , \wPDiag_55[56] , \wNDiag_41[28] , 
        \wNDiag_17[30] , \wNDiag_34[18] , \wPDiag_35[52] , \wColumn_45[6] , 
        \wNDiag_41[31] , \wNDiag_62[19] , \wPDiag_63[53] , \wNDiag_17[29] , 
        \wPDiag_28[30] , \wPDiag_28[29] , \wReturn_30[0] , \wPDiag_48[34] , 
        \wNDiag_29[63] , \wColumn_46[5] , \wColumn_2[53] , \wPDiag_4[9] , 
        \wScan_10[0] , \wScan_13[3] , \wPDiag_16[50] , \wPDiag_16[49] , 
        \wColumn_17[45] , \wNDiag_41[9] , \wColumn_21[59] , \wColumn_21[40] , 
        \wColumn_41[44] , \wPDiag_35[61] , \wNDiag_34[32] , \wPDiag_40[51] , 
        \wNDiag_62[33] , \wPDiag_20[55] , \wPDiag_40[48] , \wPDiag_63[60] , 
        \wNDiag_54[36] , \wColumn_21[2] , \wColumn_49[38] , \wColumn_29[25] , 
        \wColumn_49[21] , \wColumn_54[43] , \wNDiag_29[50] , \wColumn_34[47] , 
        \wColumn_62[46] , \wNDiag_38[2] , \wColumn_22[1] , \wNDiag_29[49] , 
        \wNDiag_44[4] , \wNDiag_49[54] , \wPDiag_1[58] , \wPDiag_1[41] , 
        \wScan_4[3] , \wColumn_14[35] , \wColumn_42[34] , \wPDiag_9[17] , 
        \wColumn_22[29] , \wColumn_57[19] , \wPDiag_11[9] , \wColumn_22[30] , 
        \wColumn_43[8] , \wScan_7[0] , \wPDiag_2[7] , \wNDiag_7[31] , 
        \wNDiag_7[28] , \wColumn_9[46] , \wPDiag_56[26] , \wPDiag_23[16] , 
        \wPDiag_9[24] , \wNDiag_14[59] , \wPDiag_15[13] , \wNDiag_22[45] , 
        \wNDiag_47[7] , \wNDiag_42[41] , \wPDiag_60[23] , \wNDiag_14[40] , 
        \wPDiag_36[22] , \wNDiag_42[58] , \wPDiag_43[12] , \wColumn_37[37] , 
        \wColumn_57[33] , \wColumn_61[36] , \wColumn_5[10] , \wPDiag_15[39] , 
        \wPDiag_15[20] , \wNDiag_20[0] , \wNDiag_23[3] , \wNDiag_37[42] , 
        \wPDiag_43[38] , \wPDiag_60[10] , \wNDiag_18[16] , \wPDiag_19[45] , 
        \wPDiag_23[25] , \wPDiag_36[11] , \wPDiag_43[21] , \wNDiag_61[43] , 
        \wColumn_39[0] , \wPDiag_56[15] , \wNDiag_57[46] , \wColumn_10[35] , 
        \wColumn_46[34] , \wColumn_26[30] , \wColumn_26[29] , \wColumn_53[19] , 
        \wPDiag_51[9] , \wNDiag_3[31] , \wPDiag_5[58] , \wPDiag_5[41] , 
        \wNDiag_3[28] , \wNDiag_3[5] , \wColumn_18[63] , \wNDiag_10[59] , 
        \wPDiag_11[13] , \wNDiag_26[45] , \wPDiag_27[16] , \wPDiag_52[26] , 
        \wNDiag_10[40] , \wNDiag_46[41] , \wPDiag_32[22] , \wNDiag_46[58] , 
        \wPDiag_47[12] , \wColumn_1[38] , \wColumn_1[21] , \wColumn_1[12] , 
        \wPDiag_1[43] , \wColumn_2[62] , \wColumn_5[23] , \wColumn_33[37] , 
        \wScan_48[2] , \wColumn_53[33] , \wColumn_6[60] , \wPDiag_6[31] , 
        \wPDiag_6[28] , \wPDiag_11[39] , \wPDiag_11[20] , \wNDiag_18[25] , 
        \wPDiag_28[2] , \wNDiag_60[0] , \wNDiag_33[42] , \wPDiag_47[38] , 
        \wNDiag_63[3] , \wPDiag_32[11] , \wPDiag_47[21] , \wColumn_18[50] , 
        \wColumn_18[49] , \wPDiag_27[25] , \wPDiag_52[15] , \wNDiag_53[46] , 
        \wColumn_58[26] , \wNDiag_6[8] , \wPDiag_12[63] , \wNDiag_13[30] , 
        \wColumn_18[9] , \wNDiag_25[35] , \wColumn_38[22] , \wNDiag_30[18] , 
        \wPDiag_51[56] , \wPDiag_31[52] , \wPDiag_57[7] , \wPDiag_44[62] , 
        \wNDiag_45[28] , \wNDiag_13[29] , \wColumn_9[5] , \wNDiag_38[57] , 
        \wNDiag_45[31] , \wNDiag_58[53] , \wPDiag_59[19] , \wPDiag_54[4] , 
        \wColumn_6[53] , \wNDiag_8[24] , \wNDiag_8[17] , \wColumn_13[45] , 
        \wScan_34[4] , \wPDiag_12[50] , \wPDiag_12[49] , \wColumn_25[59] , 
        \wColumn_25[40] , \wColumn_45[44] , \wPDiag_44[51] , \wPDiag_31[61] , 
        \wPDiag_44[48] , \wPDiag_24[55] , \wNDiag_30[32] , \wPDiag_33[3] , 
        \wNDiag_50[36] , \wColumn_61[2] , \wColumn_38[11] , \wScan_53[3] , 
        \wScan_50[0] , \wColumn_50[43] , \wColumn_58[15] , \wColumn_30[47] , 
        \wNDiag_58[60] , \wPDiag_59[33] , \wPDiag_14[6] , \wColumn_17[47] , 
        \wColumn_21[42] , \wPDiag_30[0] , \wPDiag_39[37] , \wColumn_62[1] , 
        \wNDiag_29[61] , \wColumn_41[46] , \wColumn_46[7] , \wColumn_2[51] , 
        \wColumn_2[48] , \wPDiag_2[33] , \wNDiag_4[43] , \wPDiag_16[61] , 
        \wPDiag_17[5] , \wNDiag_17[32] , \wPDiag_28[32] , \wPDiag_35[50] , 
        \wPDiag_48[36] , \wColumn_45[4] , \wPDiag_35[49] , \wPDiag_40[60] , 
        \wPDiag_63[48] , \wNDiag_21[37] , \wNDiag_41[33] , \wPDiag_63[51] , 
        \wPDiag_55[54] , \wColumn_29[14] , \wColumn_49[10] , \wNDiag_42[8] , 
        \wPDiag_7[8] , \wColumn_22[3] , \wPDiag_28[18] , \wNDiag_29[52] , 
        \wNDiag_49[56] , \wNDiag_38[0] , \wPDiag_2[19] , \wScan_10[2] , 
        \wColumn_34[45] , \wColumn_62[44] , \wColumn_54[58] , \wColumn_54[41] , 
        \wPDiag_2[5] , \wColumn_9[44] , \wScan_13[1] , \wColumn_29[27] , 
        \wNDiag_14[42] , \wPDiag_15[11] , \wPDiag_16[52] , \wNDiag_17[18] , 
        \wPDiag_20[57] , \wColumn_21[0] , \wColumn_49[23] , \wNDiag_54[34] , 
        \wNDiag_34[29] , \wPDiag_35[63] , \wPDiag_40[53] , \wNDiag_41[19] , 
        \wNDiag_62[31] , \wNDiag_62[28] , \wPDiag_63[62] , \wNDiag_34[30] , 
        \wPDiag_36[39] , \wNDiag_42[43] , \wPDiag_60[21] , \wPDiag_23[14] , 
        \wPDiag_36[20] , \wPDiag_43[10] , \wPDiag_60[38] , \wPDiag_56[24] , 
        \wNDiag_22[47] , \wScan_7[2] , \wNDiag_7[33] , \wPDiag_12[8] , 
        \wNDiag_47[5] , \wColumn_40[9] , \wScan_4[1] , \wPDiag_9[15] , 
        \wColumn_22[32] , \wColumn_42[36] , \wNDiag_59[9] , \wColumn_14[37] , 
        \wPDiag_1[6] , \wNDiag_44[6] , \wNDiag_7[19] , \wReturn_28[0] , 
        \wPDiag_15[22] , \wPDiag_23[27] , \wPDiag_56[17] , \wNDiag_23[1] , 
        \wColumn_39[2] , \wNDiag_57[44] , \wPDiag_60[12] , \wNDiag_61[58] , 
        \wNDiag_37[40] , \wPDiag_36[13] , \wPDiag_43[23] , \wNDiag_61[41] , 
        \wNDiag_37[59] , \wNDiag_20[2] , \wColumn_3[42] , \wPDiag_3[13] , 
        \wPDiag_9[26] , \wColumn_22[18] , \wColumn_37[35] , \wColumn_57[28] , 
        \wColumn_61[34] , \wNDiag_16[12] , \wPDiag_17[58] , \wNDiag_20[17] , 
        \wNDiag_55[27] , \wColumn_57[31] , \wPDiag_21[44] , \wPDiag_41[40] , 
        \wNDiag_63[22] , \wPDiag_17[41] , \wNDiag_35[23] , \wNDiag_40[13] , 
        \wPDiag_41[59] , \wColumn_28[34] , \wNDiag_5[63] , \wColumn_48[29] , 
        \wColumn_20[62] , \wColumn_35[56] , \wNDiag_36[6] , \wColumn_48[30] , 
        \wColumn_63[57] , \wNDiag_35[5] , \wColumn_55[52] , \wNDiag_28[58] , 
        \wNDiag_28[41] , \wColumn_32[9] , \wPDiag_49[16] , \wNDiag_48[45] , 
        \wPDiag_60[8] , \wPDiag_29[12] , \wPDiag_3[39] , \wNDiag_5[50] , 
        \wNDiag_5[49] , \wColumn_48[1] , \wPDiag_3[20] , \wNDiag_52[2] , 
        \wNDiag_6[13] , \wPDiag_8[35] , \wColumn_15[17] , \wColumn_16[54] , 
        \wNDiag_16[38] , \wNDiag_16[21] , \wPDiag_34[43] , \wNDiag_40[39] , 
        \wNDiag_63[11] , \wPDiag_19[3] , \wColumn_20[51] , \wNDiag_20[24] , 
        \wNDiag_35[10] , \wNDiag_40[20] , \wPDiag_62[42] , \wPDiag_29[38] , 
        \wPDiag_54[47] , \wNDiag_55[14] , \wPDiag_29[21] , \wPDiag_49[25] , 
        \wColumn_20[48] , \wColumn_55[61] , \wColumn_36[26] , \wColumn_40[55] , 
        \wColumn_43[16] , \wNDiag_51[1] , \wColumn_37[4] , \wColumn_60[27] , 
        \wPDiag_14[31] , \wPDiag_22[34] , \wColumn_23[12] , \wColumn_56[22] , 
        \wColumn_29[8] , \wNDiag_30[8] , \wPDiag_42[29] , \wNDiag_56[57] , 
        \wNDiag_43[63] , \wPDiag_14[28] , \wNDiag_36[53] , \wPDiag_37[19] , 
        \wPDiag_42[30] , \wNDiag_60[52] , \wPDiag_61[18] , \wNDiag_15[62] , 
        \wColumn_34[7] , \wScan_9[4] , \wScan_61[1] , \wColumn_1[4] , 
        \wNDiag_1[61] , \wNDiag_2[22] , \wNDiag_2[11] , \wNDiag_6[39] , 
        \wNDiag_6[20] , \wColumn_15[24] , \wColumn_23[38] , \wColumn_23[21] , 
        \wColumn_53[0] , \wColumn_36[15] , \wColumn_56[11] , \wColumn_43[25] , 
        \wNDiag_49[3] , \wColumn_60[14] , \wColumn_8[57] , \wNDiag_15[51] , 
        \wNDiag_15[48] , \wNDiag_36[60] , \wColumn_50[3] , \wPDiag_37[33] , 
        \wNDiag_43[50] , \wPDiag_61[32] , \wNDiag_43[49] , \wNDiag_60[61] , 
        \wPDiag_57[37] , \wScan_62[2] , \wNDiag_23[54] , \wColumn_4[30] , 
        \wPDiag_4[61] , \wColumn_19[43] , \wPDiag_10[33] , \wPDiag_26[4] , 
        \wNDiag_47[61] , \wNDiag_11[60] , \wNDiag_32[51] , \wScan_46[4] , 
        \wPDiag_46[32] , \wPDiag_26[36] , \wNDiag_32[48] , \wNDiag_52[55] , 
        \wColumn_4[29] , \wPDiag_4[52] , \wPDiag_10[19] , \wColumn_11[15] , 
        \wNDiag_19[36] , \wPDiag_38[8] , \wPDiag_25[7] , \wColumn_27[10] , 
        \wColumn_52[39] , \wColumn_52[20] , \wColumn_32[24] , \wColumn_47[14] , 
        \wNDiag_11[53] , \wScan_22[0] , \wNDiag_27[56] , \wPDiag_53[35] , 
        \wNDiag_32[62] , \wPDiag_33[28] , \wPDiag_33[31] , \wPDiag_46[18] , 
        \wNDiag_47[52] , \wColumn_7[59] , \wColumn_10[1] , \wColumn_11[26] , 
        \wColumn_32[17] , \wPDiag_42[0] , \wColumn_47[27] , \wColumn_13[2] , 
        \wPDiag_18[56] , \wColumn_27[23] , \wPDiag_41[3] , \wColumn_52[13] , 
        \wScan_21[3] , \wPDiag_58[39] , \wColumn_7[40] , \wPDiag_58[20] , 
        \wNDiag_9[37] , \wColumn_24[60] , \wPDiag_38[24] , \wColumn_51[50] , 
        \wColumn_51[49] , \wColumn_31[54] , \wNDiag_1[52] , \wCall_4[0] , 
        \wColumn_4[0] , \wPDiag_7[11] , \wCall_58[0] , \wNDiag_11[3] , 
        \wColumn_12[56] , \wNDiag_12[10] , \wNDiag_31[38] , \wPDiag_45[42] , 
        \wPDiag_13[43] , \wNDiag_31[21] , \wNDiag_44[11] , \wPDiag_23[9] , 
        \wNDiag_51[25] , \wNDiag_24[15] , \wPDiag_25[46] , \wColumn_24[53] , 
        \wColumn_44[57] , \wPDiag_59[1] , \wColumn_51[63] , \wColumn_7[3] , 
        \wPDiag_7[22] , \wNDiag_12[23] , \wNDiag_24[26] , \wPDiag_38[17] , 
        \wScan_39[1] , \wNDiag_39[44] , \wPDiag_58[13] , \wNDiag_59[40] , 
        \wNDiag_59[59] , \wPDiag_50[45] , \wNDiag_51[16] , \wNDiag_12[0] , 
        \wPDiag_30[58] , \wPDiag_30[41] , \wNDiag_31[12] , \wNDiag_44[22] , 
        \wColumn_59[35] , \wColumn_39[28] , \wNDiag_1[42] , \wColumn_3[61] , 
        \wPDiag_3[30] , \wNDiag_6[30] , \wNDiag_6[29] , \wPDiag_8[16] , 
        \wColumn_15[34] , \wColumn_39[31] , \wNDiag_54[5] , \wColumn_23[31] , 
        \wColumn_43[35] , \wColumn_53[9] , \wColumn_23[28] , \wColumn_56[18] , 
        \wColumn_8[47] , \wPDiag_22[17] , \wNDiag_23[44] , \wNDiag_57[6] , 
        \wPDiag_57[27] , \wPDiag_8[25] , \wPDiag_14[12] , \wNDiag_15[58] , 
        \wNDiag_15[41] , \wPDiag_37[23] , \wPDiag_42[13] , \wNDiag_43[59] , 
        \wScan_18[3] , \wNDiag_43[40] , \wPDiag_61[22] , \wColumn_56[32] , 
        \wPDiag_14[38] , \wNDiag_30[1] , \wColumn_36[36] , \wColumn_60[37] , 
        \wPDiag_37[10] , \wPDiag_42[20] , \wNDiag_60[42] , \wPDiag_14[21] , 
        \wNDiag_33[2] , \wPDiag_42[39] , \wPDiag_61[11] , \wNDiag_36[43] , 
        \wPDiag_22[24] , \wColumn_29[1] , \wNDiag_56[47] , \wPDiag_57[14] , 
        \wPDiag_3[29] , \wColumn_28[17] , \wNDiag_5[59] , \wNDiag_5[40] , 
        \wColumn_48[13] , \wPDiag_9[7] , \wNDiag_16[31] , \wNDiag_16[28] , 
        \wNDiag_20[34] , \wColumn_48[8] , \wPDiag_54[57] , \wPDiag_17[62] , 
        \wPDiag_34[53] , \wNDiag_40[30] , \wPDiag_62[52] , \wNDiag_63[18] , 
        \wNDiag_35[19] , \wColumn_55[7] , \wNDiag_40[29] , \wCall_61[0] , 
        \wPDiag_41[63] , \wPDiag_49[35] , \wColumn_56[4] , \wColumn_3[52] , 
        \wColumn_16[44] , \wNDiag_28[62] , \wPDiag_29[31] , \wPDiag_29[28] , 
        \wColumn_40[45] , \wScan_64[5] , \wPDiag_17[51] , \wColumn_20[58] , 
        \wNDiag_51[8] , \wColumn_20[41] , \wPDiag_41[49] , \wPDiag_62[61] , 
        \wPDiag_17[48] , \wNDiag_35[33] , \wPDiag_41[50] , \wNDiag_63[32] , 
        \wPDiag_21[54] , \wColumn_31[3] , \wPDiag_34[60] , \wPDiag_63[2] , 
        \wColumn_28[24] , \wColumn_48[39] , \wColumn_48[20] , \wNDiag_55[37] , 
        \wNDiag_28[48] , \wColumn_35[46] , \wColumn_55[42] , \wColumn_63[47] , 
        \wNDiag_28[3] , \wColumn_4[9] , \wColumn_24[43] , \wNDiag_28[51] , 
        \wColumn_32[0] , \wNDiag_48[55] , \wPDiag_60[1] , \wPDiag_59[8] , 
        \wColumn_7[63] , \wNDiag_8[7] , \wNDiag_9[14] , \wColumn_12[46] , 
        \wColumn_44[47] , \wColumn_16[6] , \wPDiag_44[7] , \wNDiag_59[49] , 
        \wNDiag_12[33] , \wPDiag_13[60] , \wPDiag_30[48] , \wNDiag_39[54] , 
        \wNDiag_59[50] , \wColumn_15[5] , \wNDiag_44[32] , \wPDiag_30[51] , 
        \wPDiag_47[4] , \wNDiag_24[36] , \wPDiag_45[61] , \wPDiag_50[55] , 
        \wReturn_63[0] , \wColumn_2[7] , \wColumn_7[50] , \wPDiag_7[32] , 
        \wNDiag_12[9] , \wScan_27[4] , \wColumn_39[38] , \wColumn_39[21] , 
        \wPDiag_20[3] , \wColumn_59[25] , \wPDiag_38[34] , \wPDiag_58[30] , 
        \wColumn_7[49] , \wPDiag_58[29] , \wNDiag_59[63] , \wPDiag_7[18] , 
        \wNDiag_9[27] , \wColumn_31[44] , \wScan_40[3] , \wColumn_51[59] , 
        \wColumn_51[40] , \wNDiag_11[43] , \wNDiag_12[19] , \wPDiag_13[53] , 
        \wPDiag_23[0] , \wColumn_39[12] , \wColumn_59[16] , \wScan_43[0] , 
        \wPDiag_25[56] , \wNDiag_51[35] , \wPDiag_30[62] , \wNDiag_31[31] , 
        \wNDiag_31[28] , \wNDiag_44[18] , \wPDiag_45[52] , \wPDiag_33[21] , 
        \wPDiag_46[11] , \wNDiag_2[32] , \wPDiag_10[10] , \wNDiag_17[4] , 
        \wNDiag_27[46] , \wPDiag_33[38] , \wCall_39[0] , \wNDiag_47[42] , 
        \wColumn_19[60] , \wPDiag_26[15] , \wPDiag_53[25] , \wPDiag_42[9] , 
        \wColumn_4[13] , \wPDiag_4[42] , \wColumn_10[8] , \wColumn_11[36] , 
        \wColumn_27[33] , \wColumn_47[37] , \wNDiag_2[18] , \wNDiag_14[7] , 
        \wNDiag_19[15] , \wPDiag_18[46] , \wColumn_19[53] , \wColumn_4[39] , 
        \wPDiag_10[23] , \wPDiag_26[26] , \wNDiag_52[45] , \wPDiag_53[16] , 
        \wNDiag_32[58] , \wPDiag_46[22] , \wNDiag_32[41] , \wPDiag_33[12] , 
        \wNDiag_19[26] , \wPDiag_38[1] , \wColumn_4[20] , \wPDiag_6[12] , 
        \wPDiag_12[59] , \wPDiag_12[40] , \wPDiag_24[45] , \wColumn_27[19] , 
        \wColumn_32[34] , \wColumn_52[30] , \wScan_58[1] , \wColumn_52[29] , 
        \wNDiag_25[16] , \wNDiag_50[26] , \wNDiag_30[22] , \wPDiag_44[58] , 
        \wNDiag_45[12] , \wNDiag_13[13] , \wPDiag_44[41] , \wNDiag_8[34] , 
        \wColumn_38[18] , \wColumn_25[63] , \wColumn_30[57] , \wColumn_50[53] , 
        \wPDiag_30[9] , \wColumn_62[8] , \wNDiag_3[38] , \wNDiag_3[12] , 
        \wColumn_5[33] , \wNDiag_5[2] , \wColumn_6[43] , \wPDiag_39[27] , 
        \wPDiag_59[23] , \wPDiag_6[38] , \wPDiag_6[21] , \wColumn_18[0] , 
        \wColumn_38[32] , \wColumn_58[36] , \wNDiag_6[1] , \wNDiag_13[39] , 
        \wNDiag_13[20] , \wNDiag_30[11] , \wNDiag_45[21] , \wPDiag_31[42] , 
        \wNDiag_25[25] , \wNDiag_45[38] , \wPDiag_51[46] , \wNDiag_50[15] , 
        \wPDiag_59[10] , \wColumn_10[16] , \wColumn_13[55] , \wColumn_25[50] , 
        \wColumn_25[49] , \wScan_29[2] , \wNDiag_58[43] , \wNDiag_38[47] , 
        \wPDiag_39[14] , \wPDiag_49[2] , \wColumn_45[54] , \wColumn_50[60] , 
        \wPDiag_35[4] , \wReturn_11[0] , \wColumn_26[13] , \wColumn_33[27] , 
        \wColumn_46[17] , \wColumn_53[23] , \wNDiag_18[35] , \wScan_55[4] , 
        \wNDiag_60[9] , \wPDiag_5[62] , \wNDiag_10[63] , \wPDiag_27[35] , 
        \wNDiag_53[56] , \wPDiag_47[31] , \wPDiag_11[30] , \wPDiag_11[29] , 
        \wNDiag_46[62] , \wPDiag_47[28] , \wPDiag_32[18] , \wNDiag_33[52] , 
        \wColumn_18[59] , \wColumn_18[40] , \wPDiag_36[7] , \wColumn_5[19] , 
        \wColumn_10[25] , \wPDiag_19[55] , \wScan_31[0] , \wColumn_26[39] , 
        \wColumn_26[20] , \wColumn_53[10] , \wPDiag_51[0] , \wNDiag_19[2] , 
        \wColumn_33[14] , \wColumn_46[24] , \wNDiag_3[21] , \wPDiag_52[3] , 
        \wPDiag_5[51] , \wPDiag_5[48] , \wNDiag_10[50] , \wPDiag_32[32] , 
        \wNDiag_46[48] , \wScan_1[5] , \wColumn_1[31] , \wColumn_1[28] , 
        \wPDiag_1[60] , \wNDiag_7[10] , \wNDiag_10[49] , \wNDiag_33[61] , 
        \wNDiag_26[55] , \wNDiag_46[51] , \wScan_32[3] , \wPDiag_52[36] , 
        \wNDiag_14[61] , \wScan_16[5] , \wColumn_24[4] , \wPDiag_43[33] , 
        \wNDiag_23[8] , \wNDiag_61[51] , \wPDiag_15[32] , \wNDiag_37[49] , 
        \wNDiag_42[60] , \wNDiag_61[48] , \wPDiag_23[37] , \wNDiag_37[50] , 
        \wNDiag_57[54] , \wScan_15[6] , \wPDiag_1[53] , \wColumn_9[54] , 
        \wPDiag_9[36] , \wColumn_22[11] , \wColumn_57[21] , \wColumn_57[38] , 
        \wCall_13[0] , \wColumn_27[7] , \wColumn_61[24] , \wColumn_14[14] , 
        \wNDiag_22[57] , \wColumn_37[25] , \wColumn_42[15] , \wPDiag_56[34] , 
        \wNDiag_14[52] , \wPDiag_15[18] , \wPDiag_36[30] , \wPDiag_36[29] , 
        \wNDiag_37[63] , \wPDiag_60[28] , \wNDiag_61[62] , \wNDiag_42[53] , 
        \wPDiag_43[19] , \wPDiag_60[31] , \wColumn_2[58] , \wColumn_2[41] , 
        \wNDiag_7[23] , \wPDiag_12[1] , \wColumn_40[0] , \wPDiag_11[2] , 
        \wColumn_14[27] , \wColumn_22[22] , \wColumn_37[16] , \wNDiag_59[0] , 
        \wColumn_61[17] , \wColumn_42[26] , \wColumn_43[3] , \wColumn_57[12] , 
        \wPDiag_28[11] , \wNDiag_29[42] , \wNDiag_38[9] , \wPDiag_2[10] , 
        \wNDiag_4[60] , \wColumn_21[61] , \wPDiag_48[15] , \wNDiag_49[46] , 
        \wReturn_49[0] , \wColumn_54[48] , \wColumn_54[51] , \wNDiag_25[6] , 
        \wColumn_34[55] , \wColumn_62[54] , \wNDiag_26[5] , \wColumn_49[33] , 
        \wPDiag_4[2] , \wPDiag_16[42] , \wColumn_29[37] , \wNDiag_34[20] , 
        \wNDiag_41[10] , \wNDiag_62[38] , \wNDiag_17[11] , \wNDiag_34[39] , 
        \wPDiag_40[43] , \wNDiag_62[21] , \wPDiag_20[47] , \wColumn_21[9] , 
        \wNDiag_54[24] , \wNDiag_21[14] , \wColumn_17[57] , \wColumn_41[56] , 
        \wNDiag_41[2] , \wColumn_21[52] , \wColumn_54[62] , \wColumn_1[9] , 
        \wNDiag_1[56] , \wScan_2[6] , \wPDiag_28[22] , \wPDiag_48[26] , 
        \wPDiag_2[23] , \wNDiag_17[22] , \wNDiag_21[27] , \wPDiag_55[44] , 
        \wNDiag_34[13] , \wNDiag_54[17] , \wPDiag_35[59] , \wNDiag_41[23] , 
        \wPDiag_63[41] , \wPDiag_35[40] , \wNDiag_62[12] , \wPDiag_63[58] , 
        \wNDiag_4[53] , \wPDiag_7[1] , \wNDiag_42[1] , \wColumn_7[44] , 
        \wPDiag_7[15] , \wNDiag_12[14] , \wPDiag_13[47] , \wNDiag_24[11] , 
        \wPDiag_25[42] , \wColumn_49[19] , \wColumn_58[2] , \wNDiag_51[38] , 
        \wNDiag_51[21] , \wNDiag_31[25] , \wNDiag_44[15] , \wPDiag_45[46] , 
        \wNDiag_9[33] , \wColumn_12[61] , \wColumn_31[50] , \wColumn_44[60] , 
        \wColumn_31[49] , \wPDiag_38[39] , \wColumn_51[54] , \wPDiag_38[20] , 
        \wPDiag_58[24] , \wNDiag_2[15] , \wColumn_4[34] , \wColumn_4[4] , 
        \wColumn_7[7] , \wColumn_39[35] , \wPDiag_7[26] , \wColumn_59[28] , 
        \wNDiag_12[27] , \wNDiag_12[4] , \wColumn_59[31] , \wColumn_15[8] , 
        \wPDiag_47[9] , \wNDiag_31[16] , \wNDiag_44[26] , \wNDiag_24[22] , 
        \wPDiag_30[45] , \wPDiag_50[41] , \wPDiag_38[13] , \wScan_39[5] , 
        \wPDiag_50[58] , \wNDiag_51[12] , \wPDiag_58[17] , \wNDiag_59[44] , 
        \wNDiag_39[40] , \wNDiag_39[59] , \wNDiag_9[19] , \wNDiag_11[7] , 
        \wColumn_24[57] , \wPDiag_59[5] , \wColumn_31[63] , \wColumn_12[52] , 
        \wColumn_44[53] , \wColumn_11[11] , \wPDiag_25[3] , \wColumn_32[39] , 
        \wPDiag_18[61] , \wNDiag_19[32] , \wColumn_27[14] , \wColumn_32[20] , 
        \wColumn_47[10] , \wColumn_52[24] , \wScan_45[3] , \wPDiag_10[37] , 
        \wPDiag_26[32] , \wNDiag_27[61] , \wNDiag_52[51] , \wNDiag_52[48] , 
        \wScan_46[0] , \wPDiag_46[36] , \wColumn_19[47] , \wPDiag_26[0] , 
        \wNDiag_32[55] , \wNDiag_2[26] , \wColumn_10[5] , \wColumn_11[22] , 
        \wColumn_13[6] , \wPDiag_18[52] , \wNDiag_19[18] , \wColumn_27[27] , 
        \wColumn_52[17] , \wPDiag_41[7] , \wColumn_32[13] , \wColumn_47[23] , 
        \wPDiag_42[4] , \wPDiag_4[56] , \wNDiag_6[24] , \wNDiag_6[17] , 
        \wNDiag_11[57] , \wPDiag_33[35] , \wNDiag_17[9] , \wScan_22[4] , 
        \wPDiag_26[18] , \wNDiag_27[52] , \wNDiag_47[56] , \wNDiag_52[62] , 
        \wPDiag_53[28] , \wPDiag_53[31] , \wColumn_8[60] , \wPDiag_14[35] , 
        \wColumn_34[3] , \wPDiag_42[34] , \wNDiag_60[56] , \wPDiag_22[29] , 
        \wNDiag_36[57] , \wNDiag_56[53] , \wPDiag_57[19] , \wNDiag_23[63] , 
        \wColumn_8[53] , \wPDiag_8[31] , \wPDiag_8[28] , \wPDiag_22[30] , 
        \wColumn_56[26] , \wColumn_23[16] , \wColumn_15[13] , \wColumn_37[0] , 
        \wColumn_60[23] , \wNDiag_23[50] , \wColumn_36[22] , \wColumn_43[12] , 
        \wNDiag_23[49] , \wNDiag_56[60] , \wScan_62[6] , \wPDiag_57[33] , 
        \wNDiag_15[55] , \wPDiag_37[37] , \wNDiag_43[54] , \wPDiag_61[36] , 
        \wColumn_50[7] , \wCall_64[0] , \wColumn_15[39] , \wColumn_15[20] , 
        \wColumn_43[38] , \wNDiag_49[7] , \wColumn_60[10] , \wColumn_23[25] , 
        \wColumn_36[11] , \wColumn_43[21] , \wColumn_53[4] , \wColumn_56[15] , 
        \wNDiag_54[8] , \wScan_61[5] , \wColumn_1[25] , \wColumn_1[16] , 
        \wPDiag_1[2] , \wColumn_3[46] , \wScan_9[0] , \wPDiag_29[16] , 
        \wPDiag_3[24] , \wPDiag_3[17] , \wColumn_16[63] , \wNDiag_28[45] , 
        \wColumn_35[52] , \wNDiag_35[1] , \wNDiag_48[58] , \wNDiag_48[41] , 
        \wPDiag_49[12] , \wColumn_55[56] , \wColumn_40[62] , \wColumn_63[53] , 
        \wColumn_28[29] , \wNDiag_36[2] , \wColumn_48[34] , \wColumn_16[50] , 
        \wColumn_16[49] , \wNDiag_16[16] , \wPDiag_17[45] , \wColumn_28[30] , 
        \wNDiag_35[27] , \wNDiag_40[17] , \wPDiag_41[44] , \wNDiag_63[26] , 
        \wNDiag_20[13] , \wPDiag_21[59] , \wPDiag_21[40] , \wNDiag_55[23] , 
        \wColumn_35[61] , \wColumn_40[51] , \wNDiag_51[5] , \wNDiag_16[25] , 
        \wPDiag_19[7] , \wColumn_20[55] , \wColumn_40[48] , \wColumn_63[60] , 
        \wNDiag_20[39] , \wPDiag_29[25] , \wPDiag_49[38] , \wPDiag_49[21] , 
        \wColumn_56[9] , \wNDiag_20[20] , \wPDiag_54[43] , \wNDiag_35[14] , 
        \wNDiag_55[10] , \wNDiag_40[24] , \wPDiag_62[46] , \wPDiag_34[47] , 
        \wNDiag_63[15] , \wNDiag_5[54] , \wNDiag_52[6] , \wNDiag_44[2] , 
        \wColumn_48[5] , \wPDiag_1[47] , \wScan_4[5] , \wScan_7[6] , 
        \wPDiag_9[11] , \wColumn_14[33] , \wColumn_22[36] , \wColumn_42[32] , 
        \wPDiag_2[1] , \wNDiag_7[37] , \wNDiag_22[43] , \wColumn_9[59] , 
        \wPDiag_56[39] , \wColumn_9[40] , \wPDiag_23[10] , \wNDiag_47[1] , 
        \wPDiag_56[20] , \wPDiag_9[22] , \wNDiag_14[46] , \wPDiag_15[15] , 
        \wPDiag_36[24] , \wPDiag_43[14] , \wNDiag_42[47] , \wColumn_57[35] , 
        \wPDiag_60[25] , \wColumn_14[19] , \wColumn_37[28] , \wColumn_42[18] , 
        \wColumn_61[30] , \wColumn_61[29] , \wNDiag_20[6] , \wColumn_37[31] , 
        \wColumn_2[55] , \wPDiag_2[37] , \wPDiag_15[26] , \wNDiag_23[5] , 
        \wPDiag_36[17] , \wPDiag_43[27] , \wNDiag_61[45] , \wPDiag_60[16] , 
        \wNDiag_37[44] , \wPDiag_23[23] , \wColumn_39[6] , \wNDiag_57[40] , 
        \wPDiag_56[13] , \wNDiag_57[59] , \wColumn_24[9] , \wNDiag_4[47] , 
        \wColumn_29[10] , \wReturn_9[0] , \wPDiag_14[2] , \wPDiag_17[1] , 
        \wNDiag_17[36] , \wPDiag_20[60] , \wColumn_49[14] , \wNDiag_21[33] , 
        \wPDiag_55[50] , \wPDiag_35[54] , \wNDiag_41[37] , \wPDiag_55[49] , 
        \wPDiag_63[55] , \wColumn_45[0] , \wColumn_46[3] , \wPDiag_48[32] , 
        \wNDiag_49[61] , \wPDiag_28[36] , \wScan_10[6] , \wScan_13[5] , 
        \wPDiag_16[56] , \wColumn_17[43] , \wColumn_41[42] , \wColumn_21[46] , 
        \wPDiag_20[53] , \wColumn_21[4] , \wNDiag_34[34] , \wPDiag_40[57] , 
        \wNDiag_62[35] , \wNDiag_21[19] , \wNDiag_54[29] , \wPDiag_55[63] , 
        \wColumn_49[27] , \wNDiag_54[30] , \wNDiag_26[8] , \wColumn_29[23] , 
        \wColumn_34[58] , \wColumn_34[41] , \wColumn_54[45] , \wColumn_62[59] , 
        \wColumn_62[40] , \wNDiag_38[4] , \wNDiag_3[35] , \wNDiag_3[1] , 
        \wColumn_6[57] , \wPDiag_6[35] , \wNDiag_8[13] , \wColumn_13[58] , 
        \wCall_16[0] , \wColumn_22[7] , \wNDiag_29[56] , \wPDiag_48[18] , 
        \wNDiag_49[52] , \wColumn_25[44] , \wColumn_9[1] , \wColumn_13[41] , 
        \wScan_34[0] , \wColumn_45[40] , \wColumn_45[59] , \wPDiag_54[0] , 
        \wNDiag_58[57] , \wNDiag_13[34] , \wPDiag_31[56] , \wNDiag_38[53] , 
        \wPDiag_39[19] , \wNDiag_45[35] , \wPDiag_57[3] , \wPDiag_24[62] , 
        \wNDiag_25[31] , \wNDiag_25[28] , \wNDiag_50[18] , \wPDiag_51[52] , 
        \wScan_37[3] , \wColumn_38[26] , \wPDiag_30[4] , \wNDiag_38[60] , 
        \wColumn_58[22] , \wPDiag_39[33] , \wPDiag_59[37] , \wColumn_62[5] , 
        \wNDiag_8[39] , \wNDiag_8[20] , \wReturn_14[0] , \wColumn_30[43] , 
        \wNDiag_10[44] , \wPDiag_12[54] , \wPDiag_24[51] , \wPDiag_33[7] , 
        \wColumn_38[15] , \wScan_50[4] , \wColumn_50[47] , \wColumn_58[11] , 
        \wPDiag_51[61] , \wColumn_61[6] , \wPDiag_24[48] , \wNDiag_50[32] , 
        \wNDiag_30[36] , \wPDiag_44[55] , \wPDiag_11[17] , \wPDiag_32[26] , 
        \wPDiag_47[16] , \wNDiag_26[58] , \wNDiag_26[41] , \wNDiag_46[45] , 
        \wPDiag_27[12] , \wPDiag_52[22] , \wPDiag_5[45] , \wColumn_26[34] , 
        \wColumn_5[27] , \wColumn_5[14] , \wColumn_10[31] , \wColumn_33[19] , 
        \wColumn_10[28] , \wColumn_46[29] , \wColumn_46[30] , \wPDiag_11[24] , 
        \wColumn_18[54] , \wNDiag_18[12] , \wPDiag_19[58] , \wPDiag_19[41] , 
        \wPDiag_27[38] , \wNDiag_53[42] , \wPDiag_27[21] , \wPDiag_52[11] , 
        \wPDiag_32[15] , \wPDiag_47[25] , \wNDiag_33[46] , \wNDiag_63[7] , 
        \wNDiag_18[38] , \wNDiag_18[21] , \wPDiag_28[6] , \wNDiag_60[4] , 
        \wColumn_33[33] , \wPDiag_35[9] , \wScan_1[1] , \wScan_2[2] , 
        \wColumn_2[45] , \wPDiag_2[14] , \wPDiag_16[46] , \wNDiag_17[15] , 
        \wPDiag_20[43] , \wNDiag_21[10] , \wScan_48[6] , \wColumn_53[37] , 
        \wNDiag_54[20] , \wNDiag_54[39] , \wPDiag_40[47] , \wNDiag_62[25] , 
        \wNDiag_34[24] , \wNDiag_41[14] , \wColumn_29[33] , \wColumn_17[60] , 
        \wNDiag_26[1] , \wColumn_49[37] , \wColumn_62[50] , \wNDiag_25[2] , 
        \wColumn_34[51] , \wColumn_34[48] , \wColumn_41[61] , \wColumn_62[49] , 
        \wColumn_54[55] , \wPDiag_28[15] , \wNDiag_29[46] , \wPDiag_48[11] , 
        \wNDiag_49[42] , \wPDiag_2[27] , \wNDiag_4[57] , \wPDiag_7[5] , 
        \wNDiag_42[5] , \wColumn_58[6] , \wPDiag_17[8] , \wNDiag_17[26] , 
        \wColumn_29[19] , \wPDiag_35[44] , \wNDiag_62[16] , \wNDiag_21[23] , 
        \wNDiag_34[17] , \wNDiag_41[27] , \wColumn_45[9] , \wPDiag_63[45] , 
        \wNDiag_54[13] , \wPDiag_55[59] , \wPDiag_28[26] , \wPDiag_55[40] , 
        \wColumn_1[35] , \wPDiag_4[6] , \wColumn_17[53] , \wColumn_21[56] , 
        \wPDiag_48[22] , \wColumn_34[62] , \wColumn_62[63] , \wPDiag_9[32] , 
        \wColumn_14[10] , \wColumn_27[3] , \wColumn_37[21] , \wColumn_41[52] , 
        \wNDiag_41[6] , \wColumn_42[11] , \wColumn_61[39] , \wColumn_37[38] , 
        \wColumn_61[20] , \wScan_15[2] , \wColumn_22[15] , \wColumn_57[25] , 
        \wPDiag_1[57] , \wNDiag_7[27] , \wNDiag_7[14] , \wColumn_9[63] , 
        \wNDiag_57[49] , \wPDiag_15[36] , \wNDiag_22[60] , \wPDiag_23[33] , 
        \wNDiag_57[50] , \wScan_16[1] , \wNDiag_37[54] , \wPDiag_43[37] , 
        \wColumn_24[0] , \wNDiag_61[55] , \wPDiag_9[18] , \wPDiag_11[6] , 
        \wColumn_43[7] , \wColumn_22[26] , \wColumn_14[23] , \wColumn_37[12] , 
        \wColumn_57[16] , \wColumn_42[22] , \wNDiag_59[4] , \wColumn_61[13] , 
        \wPDiag_12[5] , \wColumn_40[4] , \wPDiag_2[8] , \wNDiag_14[56] , 
        \wPDiag_36[34] , \wNDiag_42[57] , \wPDiag_60[35] , \wPDiag_56[30] , 
        \wNDiag_3[16] , \wColumn_9[50] , \wColumn_9[49] , \wNDiag_22[53] , 
        \wPDiag_23[19] , \wNDiag_47[8] , \wPDiag_56[29] , \wNDiag_57[63] , 
        \wColumn_5[37] , \wPDiag_11[34] , \wColumn_18[44] , \wPDiag_36[3] , 
        \wNDiag_26[62] , \wPDiag_27[31] , \wNDiag_33[56] , \wPDiag_47[35] , 
        \wScan_56[3] , \wPDiag_52[18] , \wNDiag_53[52] , \wPDiag_27[28] , 
        \wScan_55[0] , \wNDiag_18[31] , \wNDiag_18[28] , \wPDiag_19[62] , 
        \wColumn_10[12] , \wColumn_26[17] , \wColumn_53[27] , \wColumn_33[23] , 
        \wColumn_46[13] , \wPDiag_35[0] , \wNDiag_26[51] , \wNDiag_26[48] , 
        \wPDiag_52[32] , \wNDiag_53[61] , \wCall_1[0] , \wColumn_1[0] , 
        \wNDiag_3[25] , \wPDiag_5[55] , \wNDiag_10[54] , \wPDiag_32[36] , 
        \wNDiag_46[55] , \wNDiag_3[8] , \wColumn_4[17] , \wNDiag_5[6] , 
        \wColumn_6[47] , \wColumn_10[38] , \wPDiag_52[7] , \wColumn_10[21] , 
        \wColumn_33[10] , \wColumn_46[20] , \wPDiag_19[51] , \wNDiag_19[6] , 
        \wColumn_26[24] , \wColumn_46[39] , \wPDiag_51[4] , \wColumn_53[14] , 
        \wPDiag_19[48] , \wScan_31[4] , \wPDiag_59[27] , \wPDiag_6[16] , 
        \wNDiag_8[30] , \wNDiag_8[29] , \wPDiag_39[23] , \wColumn_50[57] , 
        \wColumn_13[62] , \wColumn_30[53] , \wColumn_45[63] , \wColumn_9[8] , 
        \wPDiag_12[44] , \wNDiag_13[17] , \wPDiag_44[45] , \wColumn_58[18] , 
        \wNDiag_30[26] , \wNDiag_45[16] , \wColumn_13[51] , \wPDiag_24[58] , 
        \wNDiag_25[12] , \wNDiag_50[22] , \wPDiag_24[41] , \wColumn_13[48] , 
        \wColumn_30[60] , \wColumn_45[49] , \wColumn_25[54] , \wColumn_45[50] , 
        \wPDiag_49[6] , \wScan_29[6] , \wPDiag_39[10] , \wNDiag_38[43] , 
        \wPDiag_54[9] , \wNDiag_58[47] , \wPDiag_59[14] , \wPDiag_6[25] , 
        \wNDiag_6[5] , \wNDiag_13[24] , \wNDiag_25[38] , \wNDiag_25[21] , 
        \wNDiag_50[11] , \wPDiag_51[42] , \wPDiag_31[46] , \wNDiag_30[15] , 
        \wNDiag_45[25] , \wColumn_58[32] , \wNDiag_14[3] , \wColumn_18[4] , 
        \wColumn_38[36] , \wPDiag_18[42] , \wNDiag_19[11] , \wNDiag_2[36] , 
        \wPDiag_4[46] , \wColumn_11[32] , \wColumn_47[33] , \wColumn_27[37] , 
        \wPDiag_10[14] , \wNDiag_17[0] , \wPDiag_26[11] , \wNDiag_27[42] , 
        \wPDiag_53[21] , \wPDiag_53[38] , \wNDiag_11[47] , \wNDiag_47[46] , 
        \wPDiag_33[25] , \wColumn_1[63] , \wColumn_1[50] , \wColumn_1[49] , 
        \wNDiag_1[46] , \wColumn_2[3] , \wPDiag_46[15] , \wColumn_4[24] , 
        \wColumn_11[18] , \wColumn_52[34] , \wScan_58[5] , \wColumn_32[30] , 
        \wColumn_32[29] , \wColumn_47[19] , \wPDiag_7[36] , \wPDiag_10[27] , 
        \wNDiag_19[22] , \wPDiag_38[5] , \wNDiag_32[45] , \wColumn_19[57] , 
        \wPDiag_26[22] , \wPDiag_33[16] , \wPDiag_46[26] , \wNDiag_52[58] , 
        \wPDiag_53[12] , \wNDiag_52[41] , \wPDiag_26[9] , \wScan_27[0] , 
        \wColumn_59[38] , \wColumn_59[21] , \wColumn_3[56] , \wPDiag_3[34] , 
        \wNDiag_5[44] , \wColumn_7[54] , \wNDiag_8[3] , \wNDiag_9[10] , 
        \wColumn_12[42] , \wNDiag_12[37] , \wColumn_15[1] , \wNDiag_24[32] , 
        \wColumn_39[25] , \wPDiag_25[61] , \wPDiag_50[48] , \wPDiag_50[51] , 
        \wPDiag_30[55] , \wPDiag_47[0] , \wColumn_16[2] , \wNDiag_39[50] , 
        \wNDiag_39[49] , \wNDiag_44[36] , \wNDiag_59[54] , \wScan_24[3] , 
        \wPDiag_44[3] , \wColumn_24[47] , \wColumn_44[43] , \wNDiag_9[23] , 
        \wPDiag_13[57] , \wPDiag_45[56] , \wPDiag_23[4] , \wNDiag_31[35] , 
        \wNDiag_51[31] , \wNDiag_24[18] , \wPDiag_25[52] , \wPDiag_50[62] , 
        \wNDiag_51[28] , \wColumn_31[59] , \wColumn_39[16] , \wScan_43[4] , 
        \wColumn_51[44] , \wColumn_59[12] , \wColumn_31[40] , \wPDiag_58[34] , 
        \wPDiag_9[3] , \wColumn_16[59] , \wColumn_16[40] , \wColumn_20[45] , 
        \wPDiag_20[7] , \wPDiag_38[30] , \wPDiag_38[29] , \wNDiag_39[63] , 
        \wScan_64[1] , \wColumn_40[58] , \wPDiag_29[35] , \wColumn_40[41] , 
        \wColumn_56[0] , \wPDiag_49[31] , \wNDiag_16[35] , \wPDiag_34[57] , 
        \wNDiag_48[62] , \wPDiag_49[28] , \wColumn_55[3] , \wNDiag_20[30] , 
        \wNDiag_40[34] , \wPDiag_62[56] , \wNDiag_20[29] , \wPDiag_21[63] , 
        \wPDiag_54[53] , \wNDiag_55[19] , \wColumn_28[13] , \wColumn_48[17] , 
        \wNDiag_28[55] , \wColumn_32[4] , \wPDiag_60[5] , \wNDiag_48[51] , 
        \wNDiag_48[48] , \wNDiag_28[7] , \wNDiag_3[59] , \wColumn_5[52] , 
        \wColumn_6[22] , \wNDiag_6[34] , \wColumn_8[43] , \wPDiag_14[16] , 
        \wPDiag_17[55] , \wPDiag_21[50] , \wPDiag_21[49] , \wColumn_28[39] , 
        \wColumn_28[20] , \wColumn_35[42] , \wColumn_63[43] , \wNDiag_35[8] , 
        \wColumn_55[46] , \wColumn_48[24] , \wNDiag_55[33] , \wColumn_31[7] , 
        \wPDiag_54[60] , \wPDiag_63[6] , \wPDiag_41[54] , \wNDiag_63[36] , 
        \wNDiag_35[37] , \wNDiag_15[45] , \wNDiag_43[44] , \wPDiag_61[26] , 
        \wPDiag_22[13] , \wNDiag_23[59] , \wPDiag_37[27] , \wPDiag_42[17] , 
        \wPDiag_57[23] , \wNDiag_23[40] , \wNDiag_57[2] , \wPDiag_8[38] , 
        \wPDiag_8[21] , \wPDiag_8[12] , \wPDiag_14[25] , \wColumn_15[30] , 
        \wColumn_15[29] , \wColumn_23[35] , \wColumn_36[18] , \wColumn_43[31] , 
        \wColumn_60[19] , \wPDiag_22[39] , \wPDiag_22[20] , \wColumn_43[28] , 
        \wNDiag_54[1] , \wPDiag_57[10] , \wColumn_29[5] , \wNDiag_56[43] , 
        \wNDiag_33[6] , \wPDiag_61[15] , \wNDiag_36[47] , \wNDiag_30[5] , 
        \wPDiag_37[14] , \wPDiag_42[24] , \wNDiag_60[46] , \wColumn_36[32] , 
        \wColumn_37[9] , \wColumn_60[33] , \wColumn_56[36] , \wNDiag_8[55] , 
        \wPDiag_18[3] , \wColumn_30[36] , \wNDiag_38[15] , \wColumn_50[32] , 
        \wPDiag_39[46] , \wColumn_6[11] , \wPDiag_12[38] , \wPDiag_12[21] , 
        \wPDiag_24[24] , \wNDiag_50[1] , \wPDiag_59[42] , \wPDiag_51[14] , 
        \wNDiag_58[11] , \wPDiag_44[39] , \wColumn_49[1] , \wNDiag_50[47] , 
        \wNDiag_30[43] , \wPDiag_44[20] , \wNDiag_53[2] , \wPDiag_31[10] , 
        \wColumn_38[60] , \wPDiag_6[59] , \wPDiag_6[40] , \wColumn_13[34] , 
        \wColumn_25[31] , \wColumn_25[28] , \wNDiag_34[5] , \wNDiag_38[26] , 
        \wNDiag_58[22] , \wColumn_33[9] , \wColumn_50[18] , \wPDiag_61[8] , 
        \wColumn_45[35] , \wColumn_38[53] , \wColumn_58[57] , \wScan_8[4] , 
        \wPDiag_11[51] , \wPDiag_11[48] , \wPDiag_12[12] , \wNDiag_13[58] , 
        \wNDiag_13[41] , \wPDiag_31[23] , \wNDiag_45[40] , \wPDiag_24[17] , 
        \wPDiag_44[13] , \wNDiag_45[59] , \wNDiag_25[44] , \wPDiag_51[27] , 
        \wPDiag_27[54] , \wNDiag_37[6] , \wColumn_51[3] , \wNDiag_53[37] , 
        \wPDiag_32[60] , \wPDiag_47[50] , \wNDiag_33[33] , \wPDiag_47[49] , 
        \wColumn_18[38] , \wColumn_18[21] , \wScan_63[2] , \wColumn_33[46] , 
        \wNDiag_18[54] , \wColumn_52[0] , \wColumn_53[42] , \wScan_60[1] , 
        \wColumn_28[8] , \wNDiag_48[3] , \wNDiag_3[40] , \wColumn_18[12] , 
        \wColumn_5[61] , \wPDiag_5[30] , \wPDiag_5[29] , \wNDiag_10[31] , 
        \wNDiag_10[28] , \wPDiag_32[53] , \wNDiag_33[19] , \wColumn_35[7] , 
        \wNDiag_46[29] , \wPDiag_47[63] , \wPDiag_11[62] , \wNDiag_26[34] , 
        \wNDiag_46[30] , \wPDiag_52[57] , \wColumn_10[44] , \wPDiag_19[34] , 
        \wColumn_36[4] , \wColumn_26[58] , \wColumn_26[41] , \wNDiag_31[8] , 
        \wColumn_46[45] , \wPDiag_1[18] , \wPDiag_9[57] , \wColumn_12[2] , 
        \wScan_20[3] , \wPDiag_40[3] , \wColumn_57[40] , \wColumn_57[59] , 
        \wScan_23[0] , \wColumn_37[44] , \wColumn_61[45] , \wColumn_11[1] , 
        \wNDiag_14[19] , \wPDiag_15[53] , \wPDiag_36[62] , \wNDiag_37[28] , 
        \wNDiag_42[18] , \wPDiag_43[52] , \wNDiag_61[30] , \wNDiag_37[31] , 
        \wPDiag_60[63] , \wNDiag_61[29] , \wNDiag_57[35] , \wColumn_14[46] , 
        \wPDiag_23[56] , \wPDiag_43[0] , \wColumn_22[43] , \wColumn_42[47] , 
        \wPDiag_39[8] , \wPDiag_1[32] , \wColumn_9[35] , \wNDiag_22[36] , 
        \wPDiag_24[7] , \wNDiag_14[33] , \wPDiag_27[4] , \wPDiag_56[55] , 
        \wPDiag_15[60] , \wPDiag_36[51] , \wPDiag_43[61] , \wPDiag_60[49] , 
        \wPDiag_36[48] , \wNDiag_42[32] , \wScan_47[4] , \wPDiag_60[50] , 
        \wColumn_2[39] , \wColumn_2[20] , \wNDiag_4[18] , \wNDiag_7[42] , 
        \wColumn_49[52] , \wCall_5[0] , \wNDiag_13[0] , \wPDiag_16[23] , 
        \wColumn_29[56] , \wNDiag_62[59] , \wPDiag_63[13] , \wNDiag_34[41] , 
        \wNDiag_34[58] , \wPDiag_40[22] , \wNDiag_62[40] , \wPDiag_35[12] , 
        \wPDiag_55[16] , \wColumn_6[3] , \wPDiag_20[26] , \wNDiag_54[45] , 
        \wNDiag_29[23] , \wColumn_5[0] , \wNDiag_10[3] , \wNDiag_49[27] , 
        \wPDiag_58[1] , \wPDiag_20[15] , \wColumn_21[19] , \wColumn_54[29] , 
        \wColumn_34[34] , \wScan_38[1] , \wColumn_54[30] , \wColumn_62[35] , 
        \wPDiag_55[25] , \wNDiag_1[23] , \wNDiag_1[6] , \wColumn_2[13] , 
        \wPDiag_2[42] , \wPDiag_16[10] , \wNDiag_21[46] , \wPDiag_35[38] , 
        \wNDiag_17[43] , \wPDiag_35[21] , \wNDiag_41[42] , \wPDiag_63[20] , 
        \wCall_59[0] , \wPDiag_40[11] , \wPDiag_63[39] , \wNDiag_4[32] , 
        \wColumn_49[61] , \wColumn_17[36] , \wPDiag_22[9] , \wColumn_41[37] , 
        \wColumn_21[33] , \wPDiag_48[47] , \wNDiag_49[14] , \wNDiag_2[5] , 
        \wNDiag_6[51] , \wNDiag_6[48] , \wPDiag_28[43] , \wNDiag_29[10] , 
        \wNDiag_62[3] , \wColumn_8[26] , \wNDiag_23[25] , \wNDiag_56[15] , 
        \wColumn_8[15] , \wPDiag_14[59] , \wColumn_15[55] , \wNDiag_15[39] , 
        \wNDiag_15[20] , \wPDiag_37[42] , \wPDiag_57[46] , \wNDiag_36[11] , 
        \wNDiag_43[38] , \wNDiag_60[10] , \wNDiag_43[21] , \wPDiag_61[43] , 
        \wScan_49[2] , \wNDiag_15[13] , \wColumn_23[50] , \wPDiag_29[2] , 
        \wColumn_43[54] , \wNDiag_61[0] , \wColumn_23[49] , \wColumn_56[60] , 
        \wPDiag_42[41] , \wNDiag_60[23] , \wPDiag_14[40] , \wPDiag_42[58] , 
        \wNDiag_43[12] , \wNDiag_23[16] , \wNDiag_36[22] , \wNDiag_56[26] , 
        \wNDiag_6[62] , \wPDiag_22[45] , \wPDiag_8[44] , \wColumn_23[63] , 
        \wColumn_56[53] , \wColumn_36[57] , \wColumn_60[56] , \wColumn_3[33] , 
        \wColumn_3[19] , \wPDiag_29[50] , \wPDiag_49[54] , \wPDiag_50[9] , 
        \wScan_51[0] , \wPDiag_3[51] , \wColumn_16[25] , \wPDiag_29[49] , 
        \wColumn_35[14] , \wColumn_40[24] , \wColumn_20[39] , \wPDiag_31[0] , 
        \wColumn_63[15] , \wColumn_63[1] , \wColumn_20[20] , \wColumn_55[10] , 
        \wPDiag_3[48] , \wNDiag_5[38] , \wNDiag_5[21] , \wPDiag_32[3] , 
        \wColumn_60[2] , \wColumn_8[5] , \wNDiag_16[50] , \wNDiag_16[49] , 
        \wNDiag_20[55] , \wScan_52[3] , \wPDiag_54[36] , \wNDiag_35[61] , 
        \wNDiag_40[51] , \wPDiag_62[33] , \wColumn_20[13] , \wPDiag_34[32] , 
        \wNDiag_40[48] , \wColumn_55[23] , \wNDiag_63[60] , \wColumn_40[17] , 
        \wColumn_16[16] , \wColumn_35[27] , \wPDiag_55[4] , \wColumn_63[26] , 
        \wNDiag_28[29] , \wPDiag_29[63] , \wScan_35[4] , \wPDiag_3[62] , 
        \wNDiag_5[12] , \wNDiag_16[63] , \wPDiag_17[30] , \wNDiag_28[30] , 
        \wPDiag_34[18] , \wNDiag_40[62] , \wNDiag_48[34] , \wPDiag_41[28] , 
        \wNDiag_35[52] , \wPDiag_41[31] , \wPDiag_62[19] , \wNDiag_63[53] , 
        \wPDiag_17[29] , \wColumn_19[9] , \wPDiag_21[35] , \wColumn_48[41] , 
        \wNDiag_55[56] , \wColumn_48[58] , \wPDiag_56[7] , \wNDiag_7[8] , 
        \wColumn_28[45] , \wScan_12[1] , \wNDiag_12[52] , \wPDiag_13[18] , 
        \wPDiag_30[29] , \wNDiag_31[63] , \wNDiag_44[53] , \wPDiag_45[19] , 
        \wPDiag_30[30] , \wNDiag_24[57] , \wPDiag_50[34] , \wNDiag_1[10] , 
        \wPDiag_7[60] , \wPDiag_7[53] , \wColumn_20[0] , \wColumn_39[40] , 
        \wColumn_39[59] , \wScan_11[2] , \wColumn_12[27] , \wColumn_23[3] , 
        \wColumn_59[44] , \wColumn_24[22] , \wColumn_31[16] , \wColumn_51[12] , 
        \wColumn_44[26] , \wNDiag_39[35] , \wNDiag_39[0] , \wPDiag_58[62] , 
        \wNDiag_59[28] , \wNDiag_59[31] , \wPDiag_16[5] , \wColumn_44[4] , 
        \wNDiag_2[60] , \wNDiag_2[53] , \wPDiag_6[8] , \wNDiag_12[61] , 
        \wPDiag_13[32] , \wPDiag_25[37] , \wNDiag_31[50] , \wNDiag_44[60] , 
        \wNDiag_51[54] , \wNDiag_31[49] , \wPDiag_45[33] , \wColumn_7[31] , 
        \wPDiag_38[55] , \wNDiag_43[8] , \wColumn_7[28] , \wPDiag_58[51] , 
        \wNDiag_9[46] , \wColumn_44[15] , \wPDiag_58[48] , \wColumn_11[57] , 
        \wColumn_12[14] , \wPDiag_15[6] , \wColumn_31[25] , \wColumn_47[7] , 
        \wColumn_24[11] , \wColumn_51[38] , \wColumn_51[21] , \wColumn_27[52] , 
        \wColumn_52[62] , \wNDiag_11[22] , \wPDiag_18[27] , \wNDiag_21[2] , 
        \wColumn_47[56] , \wPDiag_33[40] , \wNDiag_27[27] , \wNDiag_32[13] , 
        \wPDiag_33[59] , \wNDiag_47[23] , \wColumn_38[2] , \wNDiag_52[17] , 
        \wPDiag_53[44] , \wPDiag_3[5] , \wColumn_4[58] , \wPDiag_4[23] , 
        \wColumn_19[18] , \wNDiag_22[1] , \wPDiag_18[14] , \wNDiag_19[47] , 
        \wColumn_4[41] , \wScan_5[1] , \wNDiag_58[9] , \wPDiag_4[10] , 
        \wColumn_27[61] , \wColumn_32[55] , \wColumn_52[51] , \wReturn_29[0] , 
        \wNDiag_45[6] , \wColumn_52[48] , \wColumn_19[32] , \wNDiag_46[5] , 
        \wColumn_3[23] , \wNDiag_4[2] , \wScan_6[2] , \wPDiag_13[8] , 
        \wPDiag_26[47] , \wNDiag_27[14] , \wColumn_41[9] , \wNDiag_52[24] , 
        \wPDiag_46[43] , \wPDiag_10[42] , \wNDiag_11[11] , \wNDiag_32[39] , 
        \wNDiag_47[10] , \wNDiag_32[20] , \wColumn_63[36] , \wScan_28[2] , 
        \wColumn_35[37] , \wColumn_55[33] , \wNDiag_28[39] , \wNDiag_28[20] , 
        \wPDiag_48[2] , \wNDiag_48[24] , \wColumn_3[10] , \wNDiag_7[1] , 
        \wPDiag_17[39] , \wColumn_19[0] , \wPDiag_21[25] , \wPDiag_54[15] , 
        \wNDiag_55[46] , \wPDiag_41[21] , \wNDiag_63[43] , \wPDiag_17[20] , 
        \wPDiag_34[11] , \wPDiag_41[38] , \wPDiag_62[10] , \wColumn_28[55] , 
        \wNDiag_35[42] , \wNDiag_28[13] , \wPDiag_29[59] , \wColumn_48[51] , 
        \wColumn_48[48] , \wPDiag_3[58] , \wNDiag_5[31] , \wNDiag_5[28] , 
        \wColumn_16[35] , \wColumn_20[30] , \wPDiag_29[40] , \wPDiag_31[9] , 
        \wNDiag_48[17] , \wPDiag_49[44] , \wColumn_63[8] , \wColumn_20[29] , 
        \wColumn_55[19] , \wColumn_40[34] , \wColumn_48[62] , \wPDiag_3[41] , 
        \wColumn_4[51] , \wNDiag_6[58] , \wNDiag_6[41] , \wPDiag_8[54] , 
        \wPDiag_14[50] , \wNDiag_16[59] , \wNDiag_16[40] , \wPDiag_34[22] , 
        \wPDiag_17[13] , \wNDiag_40[58] , \wPDiag_41[12] , \wNDiag_20[45] , 
        \wNDiag_40[41] , \wPDiag_62[23] , \wPDiag_21[16] , \wPDiag_22[55] , 
        \wPDiag_53[3] , \wPDiag_54[26] , \wNDiag_36[32] , \wPDiag_42[48] , 
        \wNDiag_56[36] , \wPDiag_61[60] , \wPDiag_14[49] , \wPDiag_37[61] , 
        \wPDiag_42[51] , \wNDiag_60[33] , \wScan_30[0] , \wScan_33[3] , 
        \wColumn_36[47] , \wColumn_60[46] , \wNDiag_18[2] , \wPDiag_50[0] , 
        \wColumn_56[43] , \wColumn_8[36] , \wPDiag_14[63] , \wNDiag_15[30] , 
        \wNDiag_15[29] , \wPDiag_37[7] , \wNDiag_43[31] , \wNDiag_60[19] , 
        \wPDiag_61[53] , \wNDiag_36[18] , \wPDiag_37[52] , \wPDiag_42[62] , 
        \wNDiag_43[28] , \wReturn_10[0] , \wNDiag_23[35] , \wPDiag_57[56] , 
        \wPDiag_34[4] , \wColumn_15[45] , \wColumn_23[59] , \wColumn_23[40] , 
        \wColumn_43[44] , \wScan_54[4] , \wNDiag_61[9] , \wColumn_4[48] , 
        \wNDiag_58[0] , \wPDiag_4[19] , \wPDiag_10[2] , \wColumn_42[3] , 
        \wColumn_19[22] , \wNDiag_19[57] , \wColumn_32[45] , \wColumn_52[58] , 
        \wColumn_52[41] , \wPDiag_10[52] , \wNDiag_11[18] , \wNDiag_32[30] , 
        \wPDiag_13[1] , \wNDiag_32[29] , \wPDiag_33[63] , \wPDiag_46[53] , 
        \wNDiag_47[19] , \wColumn_41[0] , \wPDiag_26[57] , \wColumn_47[46] , 
        \wNDiag_52[34] , \wScan_0[5] , \wNDiag_1[19] , \wNDiag_2[43] , 
        \wColumn_4[62] , \wColumn_11[47] , \wScan_14[6] , \wPDiag_18[37] , 
        \wColumn_27[42] , \wPDiag_4[33] , \wPDiag_10[61] , \wCall_12[0] , 
        \wColumn_26[7] , \wNDiag_27[37] , \wPDiag_53[54] , \wNDiag_11[32] , 
        \wPDiag_33[49] , \wNDiag_47[33] , \wScan_17[5] , \wColumn_25[4] , 
        \wPDiag_33[50] , \wPDiag_46[60] , \wNDiag_22[8] , \wScan_3[6] , 
        \wColumn_19[11] , \wPDiag_5[2] , \wPDiag_6[1] , \wPDiag_30[13] , 
        \wColumn_39[63] , \wPDiag_45[23] , \wNDiag_31[59] , \wColumn_7[38] , 
        \wPDiag_13[22] , \wPDiag_25[27] , \wNDiag_31[40] , \wNDiag_43[1] , 
        \wPDiag_50[17] , \wNDiag_51[44] , \wColumn_59[2] , \wNDiag_40[2] , 
        \wColumn_7[21] , \wPDiag_58[58] , \wNDiag_59[12] , \wPDiag_38[45] , 
        \wPDiag_58[41] , \wNDiag_39[16] , \wColumn_51[31] , \wColumn_51[28] , 
        \wNDiag_1[33] , \wPDiag_7[43] , \wNDiag_9[56] , \wColumn_24[18] , 
        \wNDiag_12[42] , \wNDiag_24[47] , \wColumn_31[35] , \wPDiag_25[14] , 
        \wNDiag_27[5] , \wPDiag_30[20] , \wPDiag_50[24] , \wPDiag_13[11] , 
        \wPDiag_30[39] , \wPDiag_45[10] , \wNDiag_44[43] , \wColumn_59[54] , 
        \wColumn_20[9] , \wColumn_39[49] , \wNDiag_3[63] , \wNDiag_3[50] , 
        \wPDiag_5[39] , \wPDiag_5[20] , \wColumn_7[12] , \wColumn_12[37] , 
        \wColumn_39[50] , \wColumn_24[32] , \wNDiag_39[9] , \wColumn_44[36] , 
        \wNDiag_24[6] , \wNDiag_39[25] , \wReturn_48[0] , \wNDiag_59[21] , 
        \wNDiag_59[38] , \wNDiag_32[2] , \wColumn_28[1] , \wNDiag_3[49] , 
        \wColumn_10[54] , \wNDiag_10[38] , \wNDiag_26[24] , \wPDiag_52[47] , 
        \wNDiag_33[10] , \wNDiag_53[14] , \wNDiag_10[21] , \wPDiag_32[43] , 
        \wNDiag_46[20] , \wScan_19[3] , \wNDiag_46[39] , \wPDiag_19[24] , 
        \wNDiag_31[1] , \wColumn_46[55] , \wNDiag_10[12] , \wPDiag_11[58] , 
        \wPDiag_11[41] , \wColumn_26[51] , \wColumn_26[48] , \wNDiag_46[13] , 
        \wPDiag_47[59] , \wColumn_53[61] , \wNDiag_33[23] , \wPDiag_47[40] , 
        \wColumn_18[28] , \wNDiag_26[17] , \wPDiag_27[44] , \wNDiag_53[27] , 
        \wNDiag_56[6] , \wColumn_5[42] , \wPDiag_5[13] , \wColumn_18[31] , 
        \wColumn_26[62] , \wColumn_53[52] , \wNDiag_55[5] , \wColumn_33[56] , 
        \wColumn_6[18] , \wNDiag_18[44] , \wPDiag_19[17] , \wColumn_52[9] , 
        \wNDiag_38[36] , \wColumn_13[24] , \wNDiag_58[32] , \wPDiag_59[61] , 
        \wColumn_25[21] , \wNDiag_29[3] , \wColumn_30[15] , \wColumn_45[25] , 
        \wPDiag_6[50] , \wPDiag_6[49] , \wColumn_25[38] , \wColumn_33[0] , 
        \wColumn_50[11] , \wPDiag_61[1] , \wColumn_58[47] , \wNDiag_13[51] , 
        \wNDiag_25[54] , \wColumn_30[3] , \wPDiag_62[2] , \wColumn_38[43] , 
        \wPDiag_51[37] , \wNDiag_13[48] , \wPDiag_31[33] , \wNDiag_45[49] , 
        \wNDiag_30[60] , \wNDiag_45[50] , \wColumn_1[59] , \wColumn_1[40] , 
        \wPDiag_1[22] , \wColumn_2[30] , \wColumn_2[29] , \wPDiag_2[61] , 
        \wPDiag_2[52] , \wNDiag_4[22] , \wColumn_6[32] , \wPDiag_8[7] , 
        \wColumn_25[12] , \wColumn_50[22] , \wNDiag_8[45] , \wColumn_13[17] , 
        \wColumn_57[4] , \wColumn_45[16] , \wColumn_30[26] , \wPDiag_6[63] , 
        \wPDiag_12[31] , \wPDiag_12[28] , \wPDiag_39[56] , \wNDiag_50[8] , 
        \wNDiag_58[18] , \wPDiag_59[52] , \wPDiag_44[30] , \wNDiag_13[62] , 
        \wNDiag_30[53] , \wPDiag_44[29] , \wNDiag_45[63] , \wPDiag_31[19] , 
        \wPDiag_24[34] , \wColumn_49[8] , \wNDiag_50[57] , \wColumn_54[7] , 
        \wPDiag_16[19] , \wNDiag_17[53] , \wCall_60[0] , \wNDiag_21[56] , 
        \wNDiag_34[62] , \wPDiag_35[31] , \wPDiag_35[28] , \wNDiag_62[63] , 
        \wPDiag_63[29] , \wPDiag_40[18] , \wNDiag_41[52] , \wPDiag_63[30] , 
        \wPDiag_22[0] , \wScan_42[0] , \wPDiag_55[35] , \wColumn_14[5] , 
        \wColumn_17[26] , \wColumn_21[23] , \wPDiag_21[3] , \wColumn_54[13] , 
        \wPDiag_28[53] , \wNDiag_29[19] , \wColumn_34[17] , \wColumn_62[16] , 
        \wColumn_41[27] , \wColumn_29[46] , \wScan_41[3] , \wPDiag_48[57] , 
        \wPDiag_46[4] , \wNDiag_4[11] , \wColumn_49[42] , \wReturn_62[0] , 
        \wColumn_5[9] , \wNDiag_13[9] , \wNDiag_17[60] , \wPDiag_20[36] , 
        \wNDiag_54[55] , \wScan_26[4] , \wNDiag_62[50] , \wNDiag_34[48] , 
        \wPDiag_40[32] , \wPDiag_16[33] , \wNDiag_34[51] , \wNDiag_41[61] , 
        \wNDiag_62[49] , \wPDiag_58[8] , \wNDiag_9[7] , \wNDiag_49[37] , 
        \wNDiag_29[33] , \wPDiag_28[60] , \wNDiag_7[52] , \wColumn_9[25] , 
        \wColumn_14[56] , \wColumn_17[15] , \wColumn_17[6] , \wColumn_62[25] , 
        \wPDiag_45[7] , \wColumn_21[10] , \wColumn_34[24] , \wColumn_41[14] , 
        \wColumn_54[20] , \wColumn_22[53] , \wPDiag_39[1] , \wColumn_54[39] , 
        \wColumn_42[57] , \wColumn_57[63] , \wNDiag_14[23] , \wPDiag_36[58] , 
        \wScan_59[1] , \wPDiag_36[41] , \wNDiag_37[12] , \wNDiag_42[22] , 
        \wPDiag_60[40] , \wPDiag_60[59] , \wNDiag_61[13] , \wNDiag_22[26] , 
        \wPDiag_56[45] , \wNDiag_57[16] , \wPDiag_1[11] , \wPDiag_9[47] , 
        \wColumn_37[54] , \wColumn_57[49] , \wColumn_61[55] , \wNDiag_15[7] , 
        \wColumn_57[50] , \wColumn_22[60] , \wNDiag_1[27] , \wNDiag_2[57] , 
        \wColumn_3[7] , \wPDiag_4[27] , \wNDiag_7[61] , \wNDiag_16[4] , 
        \wCall_38[0] , \wColumn_9[16] , \wColumn_11[8] , \wPDiag_23[46] , 
        \wPDiag_43[9] , \wNDiag_14[10] , \wPDiag_15[43] , \wNDiag_22[15] , 
        \wNDiag_57[25] , \wNDiag_42[11] , \wNDiag_61[39] , \wNDiag_37[21] , 
        \wPDiag_43[42] , \wNDiag_61[20] , \wNDiag_37[38] , \wNDiag_22[5] , 
        \wColumn_38[6] , \wPDiag_3[1] , \wScan_6[6] , \wPDiag_10[46] , 
        \wColumn_11[53] , \wNDiag_11[26] , \wColumn_25[9] , \wNDiag_27[23] , 
        \wPDiag_53[40] , \wNDiag_32[17] , \wNDiag_52[13] , \wPDiag_53[59] , 
        \wPDiag_33[44] , \wNDiag_47[27] , \wPDiag_18[23] , \wNDiag_21[6] , 
        \wColumn_32[62] , \wColumn_47[52] , \wColumn_27[56] , \wNDiag_47[14] , 
        \wNDiag_32[24] , \wPDiag_46[47] , \wNDiag_11[15] , \wPDiag_26[43] , 
        \wNDiag_52[39] , \wNDiag_27[10] , \wNDiag_52[20] , \wNDiag_46[1] , 
        \wColumn_4[45] , \wPDiag_4[14] , \wColumn_19[36] , \wScan_5[5] , 
        \wColumn_11[60] , \wColumn_32[51] , \wNDiag_45[2] , \wColumn_52[55] , 
        \wColumn_47[61] , \wColumn_32[48] , \wPDiag_7[57] , \wScan_11[6] , 
        \wPDiag_18[10] , \wNDiag_19[43] , \wColumn_12[23] , \wPDiag_38[62] , 
        \wNDiag_39[28] , \wNDiag_39[31] , \wNDiag_59[35] , \wCall_17[0] , 
        \wColumn_23[7] , \wColumn_24[26] , \wColumn_31[12] , \wNDiag_39[4] , 
        \wColumn_44[22] , \wColumn_51[16] , \wColumn_59[59] , \wColumn_59[40] , 
        \wColumn_20[4] , \wNDiag_1[14] , \wColumn_7[35] , \wReturn_8[0] , 
        \wNDiag_9[42] , \wScan_12[5] , \wNDiag_24[53] , \wPDiag_25[19] , 
        \wColumn_39[44] , \wPDiag_50[29] , \wNDiag_51[63] , \wColumn_12[10] , 
        \wNDiag_12[56] , \wNDiag_27[8] , \wPDiag_50[30] , \wPDiag_15[2] , 
        \wColumn_24[15] , \wPDiag_30[34] , \wNDiag_44[57] , \wColumn_51[25] , 
        \wColumn_47[3] , \wColumn_31[38] , \wColumn_44[11] , \wColumn_31[21] , 
        \wPDiag_13[36] , \wNDiag_31[54] , \wPDiag_38[51] , \wPDiag_58[55] , 
        \wPDiag_38[48] , \wPDiag_45[37] , \wNDiag_24[60] , \wNDiag_51[50] , 
        \wPDiag_25[33] , \wNDiag_51[49] , \wNDiag_1[2] , \wColumn_3[37] , 
        \wPDiag_3[55] , \wNDiag_5[25] , \wPDiag_16[1] , \wColumn_44[0] , 
        \wNDiag_16[54] , \wNDiag_20[51] , \wPDiag_34[36] , \wNDiag_40[55] , 
        \wPDiag_62[37] , \wNDiag_20[48] , \wNDiag_55[61] , \wPDiag_32[7] , 
        \wPDiag_54[32] , \wColumn_60[6] , \wNDiag_5[16] , \wReturn_15[0] , 
        \wColumn_16[38] , \wColumn_16[21] , \wColumn_20[24] , \wPDiag_31[4] , 
        \wColumn_55[14] , \wColumn_63[5] , \wColumn_35[10] , \wColumn_40[39] , 
        \wColumn_63[11] , \wColumn_40[20] , \wColumn_28[58] , \wColumn_28[41] , 
        \wPDiag_29[54] , \wPDiag_49[50] , \wScan_51[4] , \wPDiag_49[49] , 
        \wPDiag_56[3] , \wColumn_48[45] , \wPDiag_17[34] , \wNDiag_20[62] , 
        \wPDiag_54[18] , \wNDiag_55[52] , \wPDiag_21[31] , \wPDiag_21[28] , 
        \wNDiag_35[56] , \wScan_36[3] , \wPDiag_41[35] , \wNDiag_63[57] , 
        \wNDiag_28[34] , \wNDiag_48[30] , \wNDiag_48[29] , \wPDiag_49[63] , 
        \wScan_35[0] , \wNDiag_6[55] , \wColumn_8[22] , \wColumn_8[1] , 
        \wColumn_16[12] , \wPDiag_55[0] , \wColumn_63[22] , \wColumn_35[23] , 
        \wColumn_40[13] , \wColumn_15[51] , \wColumn_15[48] , \wColumn_20[17] , 
        \wColumn_55[27] , \wColumn_23[54] , \wPDiag_29[6] , \wColumn_36[60] , 
        \wColumn_43[50] , \wNDiag_61[4] , \wNDiag_15[24] , \wPDiag_34[9] , 
        \wColumn_43[49] , \wColumn_60[61] , \wNDiag_36[15] , \wScan_49[6] , 
        \wPDiag_37[46] , \wNDiag_43[25] , \wPDiag_61[47] , \wNDiag_23[38] , 
        \wNDiag_60[14] , \wNDiag_23[21] , \wPDiag_57[42] , \wNDiag_56[11] , 
        \wNDiag_62[7] , \wColumn_2[24] , \wNDiag_2[1] , \wColumn_8[11] , 
        \wPDiag_8[59] , \wPDiag_8[40] , \wColumn_15[62] , \wColumn_36[53] , 
        \wColumn_43[63] , \wColumn_60[52] , \wColumn_56[57] , \wColumn_5[4] , 
        \wPDiag_14[44] , \wPDiag_22[58] , \wPDiag_22[41] , \wNDiag_23[12] , 
        \wNDiag_56[22] , \wNDiag_43[16] , \wNDiag_15[17] , \wNDiag_36[26] , 
        \wPDiag_42[45] , \wNDiag_60[27] , \wColumn_17[18] , \wColumn_34[30] , 
        \wColumn_34[29] , \wColumn_41[19] , \wColumn_62[31] , \wColumn_62[28] , 
        \wScan_38[5] , \wColumn_54[34] , \wNDiag_10[7] , \wNDiag_29[27] , 
        \wNDiag_49[23] , \wPDiag_58[5] , \wColumn_2[17] , \wColumn_6[7] , 
        \wPDiag_20[22] , \wNDiag_54[58] , \wNDiag_54[41] , \wPDiag_55[12] , 
        \wNDiag_13[4] , \wPDiag_16[27] , \wPDiag_35[16] , \wPDiag_40[26] , 
        \wNDiag_62[44] , \wPDiag_63[17] , \wNDiag_34[45] , \wColumn_14[8] , 
        \wPDiag_46[9] , \wColumn_29[52] , \wNDiag_29[14] , \wColumn_49[56] , 
        \wPDiag_2[46] , \wNDiag_4[36] , \wColumn_17[32] , \wColumn_21[37] , 
        \wPDiag_28[47] , \wPDiag_48[43] , \wNDiag_49[10] , \wColumn_41[33] , 
        \wColumn_29[61] , \wPDiag_16[14] , \wNDiag_17[47] , \wPDiag_35[25] , 
        \wPDiag_40[15] , \wNDiag_41[46] , \wPDiag_63[24] , \wColumn_1[54] , 
        \wPDiag_9[53] , \wColumn_11[5] , \wPDiag_20[11] , \wNDiag_21[42] , 
        \wPDiag_55[38] , \wPDiag_55[21] , \wPDiag_56[62] , \wNDiag_57[28] , 
        \wPDiag_15[57] , \wNDiag_22[18] , \wPDiag_23[52] , \wPDiag_43[4] , 
        \wNDiag_37[35] , \wNDiag_57[31] , \wNDiag_16[9] , \wScan_23[4] , 
        \wPDiag_43[56] , \wNDiag_61[34] , \wColumn_37[59] , \wColumn_37[40] , 
        \wColumn_61[58] , \wColumn_61[41] , \wColumn_12[6] , \wColumn_57[44] , 
        \wPDiag_40[7] , \wPDiag_1[36] , \wNDiag_7[46] , \wScan_47[0] , 
        \wNDiag_3[44] , \wColumn_5[56] , \wColumn_9[31] , \wNDiag_14[37] , 
        \wPDiag_27[0] , \wNDiag_42[36] , \wPDiag_60[54] , \wPDiag_23[61] , 
        \wPDiag_36[55] , \wColumn_9[28] , \wNDiag_22[32] , \wPDiag_56[51] , 
        \wPDiag_9[60] , \wPDiag_24[3] , \wPDiag_56[48] , \wColumn_14[42] , 
        \wColumn_22[47] , \wColumn_42[43] , \wScan_44[3] , \wPDiag_5[34] , 
        \wScan_8[0] , \wNDiag_18[50] , \wNDiag_18[49] , \wNDiag_48[7] , 
        \wColumn_52[4] , \wNDiag_55[8] , \wScan_60[5] , \wColumn_10[59] , 
        \wPDiag_11[55] , \wColumn_18[25] , \wColumn_33[42] , \wColumn_53[46] , 
        \wNDiag_33[37] , \wScan_63[6] , \wPDiag_27[50] , \wPDiag_47[54] , 
        \wColumn_51[7] , \wPDiag_52[60] , \wPDiag_27[49] , \wNDiag_53[33] , 
        \wColumn_10[40] , \wColumn_46[41] , \wNDiag_10[35] , \wNDiag_18[63] , 
        \wPDiag_19[30] , \wColumn_26[45] , \wColumn_46[58] , \wPDiag_19[29] , 
        \wNDiag_26[30] , \wNDiag_26[29] , \wColumn_36[0] , \wPDiag_27[63] , 
        \wPDiag_52[53] , \wNDiag_53[19] , \wNDiag_46[34] , \wPDiag_32[57] , 
        \wColumn_35[3] , \wColumn_6[26] , \wPDiag_12[25] , \wColumn_18[16] , 
        \wPDiag_31[14] , \wPDiag_44[24] , \wColumn_58[60] , \wPDiag_24[39] , 
        \wNDiag_30[47] , \wColumn_49[5] , \wNDiag_53[6] , \wNDiag_50[43] , 
        \wPDiag_24[20] , \wPDiag_51[10] , \wNDiag_50[5] , \wNDiag_58[15] , 
        \wPDiag_6[44] , \wNDiag_8[51] , \wNDiag_8[48] , \wPDiag_18[7] , 
        \wNDiag_38[11] , \wPDiag_39[42] , \wPDiag_59[46] , \wColumn_50[36] , 
        \wPDiag_12[16] , \wNDiag_13[45] , \wPDiag_24[13] , \wNDiag_25[59] , 
        \wNDiag_25[40] , \wColumn_30[32] , \wColumn_57[9] , \wNDiag_37[2] , 
        \wPDiag_31[27] , \wPDiag_51[23] , \wPDiag_44[17] , \wNDiag_45[44] , 
        \wColumn_58[53] , \wNDiag_8[62] , \wColumn_13[30] , \wColumn_38[57] , 
        \wColumn_13[29] , \wColumn_30[18] , \wColumn_45[28] , \wColumn_45[31] , 
        \wColumn_25[35] , \wCall_0[0] , \wPDiag_1[26] , \wColumn_6[15] , 
        \wNDiag_34[1] , \wNDiag_38[22] , \wNDiag_58[26] , \wPDiag_1[15] , 
        \wNDiag_7[56] , \wColumn_9[38] , \wNDiag_22[22] , \wColumn_9[21] , 
        \wPDiag_56[58] , \wNDiag_57[12] , \wColumn_9[12] , \wColumn_14[52] , 
        \wNDiag_14[27] , \wPDiag_36[45] , \wPDiag_56[41] , \wPDiag_27[9] , 
        \wNDiag_37[16] , \wNDiag_61[17] , \wNDiag_42[26] , \wPDiag_60[44] , 
        \wScan_59[5] , \wNDiag_14[14] , \wColumn_22[57] , \wColumn_37[63] , 
        \wColumn_61[62] , \wPDiag_39[5] , \wColumn_42[53] , \wPDiag_43[46] , 
        \wNDiag_61[24] , \wPDiag_15[47] , \wNDiag_42[15] , \wNDiag_22[11] , 
        \wNDiag_37[25] , \wNDiag_57[21] , \wNDiag_16[0] , \wPDiag_23[42] , 
        \wNDiag_57[38] , \wColumn_3[3] , \wColumn_1[44] , \wPDiag_9[43] , 
        \wNDiag_15[3] , \wColumn_57[54] , \wColumn_14[61] , \wColumn_37[49] , 
        \wColumn_61[51] , \wColumn_37[50] , \wColumn_42[60] , \wColumn_61[48] , 
        \wColumn_2[34] , \wPDiag_2[56] , \wColumn_17[22] , \wPDiag_28[57] , 
        \wPDiag_48[53] , \wNDiag_49[19] , \wColumn_34[13] , \wColumn_41[23] , 
        \wColumn_21[27] , \wPDiag_21[7] , \wColumn_62[12] , \wColumn_54[17] , 
        \wNDiag_4[26] , \wColumn_17[11] , \wColumn_17[2] , \wNDiag_17[57] , 
        \wPDiag_20[18] , \wNDiag_21[52] , \wPDiag_22[4] , \wScan_42[4] , 
        \wPDiag_55[31] , \wNDiag_41[56] , \wNDiag_54[62] , \wPDiag_55[28] , 
        \wPDiag_63[34] , \wColumn_21[14] , \wPDiag_35[35] , \wColumn_54[24] , 
        \wColumn_34[20] , \wColumn_41[10] , \wColumn_62[38] , \wColumn_62[21] , 
        \wPDiag_45[3] , \wScan_25[3] , \wColumn_34[39] , \wNDiag_4[15] , 
        \wNDiag_9[3] , \wNDiag_29[37] , \wPDiag_16[37] , \wNDiag_34[55] , 
        \wPDiag_48[60] , \wNDiag_49[33] , \wPDiag_20[32] , \wScan_26[0] , 
        \wNDiag_62[54] , \wPDiag_40[36] , \wNDiag_54[48] , \wNDiag_21[61] , 
        \wNDiag_54[51] , \wColumn_49[46] , \wPDiag_6[54] , \wNDiag_13[55] , 
        \wColumn_14[1] , \wColumn_29[42] , \wPDiag_46[0] , \wNDiag_45[54] , 
        \wNDiag_25[50] , \wNDiag_25[49] , \wPDiag_31[37] , \wPDiag_51[33] , 
        \wColumn_30[7] , \wColumn_38[47] , \wNDiag_50[60] , \wPDiag_62[6] , 
        \wColumn_25[25] , \wColumn_33[4] , \wColumn_58[43] , \wPDiag_61[5] , 
        \wColumn_6[36] , \wPDiag_12[35] , \wColumn_13[39] , \wColumn_30[11] , 
        \wColumn_50[15] , \wColumn_13[20] , \wColumn_45[21] , \wPDiag_24[30] , 
        \wNDiag_29[7] , \wColumn_45[38] , \wNDiag_34[8] , \wNDiag_38[32] , 
        \wNDiag_58[36] , \wPDiag_39[61] , \wColumn_54[3] , \wPDiag_24[29] , 
        \wNDiag_50[53] , \wPDiag_51[19] , \wNDiag_25[63] , \wNDiag_30[57] , 
        \wNDiag_38[18] , \wPDiag_44[34] , \wPDiag_39[52] , \wPDiag_8[3] , 
        \wNDiag_8[58] , \wNDiag_8[41] , \wColumn_45[12] , \wPDiag_59[56] , 
        \wColumn_30[22] , \wColumn_13[13] , \wColumn_57[0] , \wScan_0[1] , 
        \wNDiag_3[54] , \wColumn_10[50] , \wColumn_25[16] , \wColumn_50[26] , 
        \wColumn_26[55] , \wColumn_10[49] , \wColumn_46[48] , \wNDiag_10[25] , 
        \wPDiag_19[39] , \wNDiag_31[5] , \wColumn_33[61] , \wColumn_46[51] , 
        \wColumn_36[9] , \wPDiag_19[20] , \wPDiag_32[47] , \wNDiag_26[39] , 
        \wNDiag_26[20] , \wNDiag_33[14] , \wNDiag_46[24] , \wNDiag_53[10] , 
        \wColumn_28[5] , \wPDiag_52[43] , \wColumn_5[46] , \wPDiag_5[24] , 
        \wNDiag_32[6] , \wNDiag_18[59] , \wNDiag_18[40] , \wPDiag_19[13] , 
        \wPDiag_5[17] , \wColumn_10[63] , \wColumn_33[52] , \wColumn_46[62] , 
        \wColumn_53[56] , \wNDiag_55[1] , \wNDiag_9[52] , \wNDiag_10[16] , 
        \wColumn_18[35] , \wNDiag_26[13] , \wPDiag_27[59] , \wNDiag_53[23] , 
        \wNDiag_56[2] , \wPDiag_27[40] , \wPDiag_47[44] , \wPDiag_11[45] , 
        \wNDiag_46[17] , \wNDiag_33[27] , \wColumn_12[19] , \wColumn_31[31] , 
        \wColumn_31[28] , \wColumn_44[18] , \wNDiag_1[37] , \wScan_3[2] , 
        \wPDiag_5[6] , \wColumn_7[25] , \wPDiag_38[58] , \wColumn_51[35] , 
        \wPDiag_38[41] , \wNDiag_39[12] , \wNDiag_40[6] , \wPDiag_58[45] , 
        \wPDiag_6[5] , \wPDiag_25[23] , \wPDiag_50[13] , \wNDiag_59[16] , 
        \wNDiag_51[59] , \wNDiag_51[40] , \wColumn_59[6] , \wPDiag_13[26] , 
        \wPDiag_16[8] , \wPDiag_30[17] , \wNDiag_31[44] , \wNDiag_43[5] , 
        \wPDiag_45[27] , \wColumn_44[9] , \wColumn_59[63] , \wColumn_7[16] , 
        \wNDiag_9[61] , \wColumn_24[36] , \wNDiag_24[2] , \wNDiag_39[21] , 
        \wNDiag_59[25] , \wNDiag_39[38] , \wColumn_44[32] , \wColumn_12[33] , 
        \wNDiag_2[47] , \wPDiag_3[8] , \wPDiag_7[47] , \wColumn_39[54] , 
        \wColumn_59[49] , \wPDiag_10[56] , \wNDiag_12[46] , \wPDiag_13[15] , 
        \wColumn_59[50] , \wPDiag_30[24] , \wNDiag_44[47] , \wPDiag_13[5] , 
        \wNDiag_24[43] , \wPDiag_25[10] , \wPDiag_45[14] , \wPDiag_50[20] , 
        \wNDiag_27[1] , \wColumn_41[4] , \wPDiag_50[39] , \wNDiag_52[30] , 
        \wNDiag_52[29] , \wPDiag_53[63] , \wPDiag_26[53] , \wNDiag_27[19] , 
        \wNDiag_32[34] , \wPDiag_46[57] , \wColumn_19[26] , \wNDiag_46[8] , 
        \wColumn_4[55] , \wPDiag_10[6] , \wNDiag_19[53] , \wColumn_32[58] , 
        \wColumn_32[41] , \wColumn_42[7] , \wColumn_52[45] , \wPDiag_18[19] , 
        \wColumn_19[15] , \wNDiag_58[4] , \wPDiag_4[37] , \wScan_17[1] , 
        \wColumn_11[43] , \wNDiag_11[36] , \wPDiag_18[33] , \wNDiag_19[60] , 
        \wColumn_25[0] , \wPDiag_33[54] , \wColumn_26[3] , \wPDiag_26[60] , 
        \wNDiag_27[33] , \wNDiag_47[37] , \wPDiag_53[49] , \wPDiag_53[50] , 
        \wColumn_27[46] , \wScan_14[2] , \wColumn_47[42] , \wScan_0[3] , 
        \wNDiag_2[8] , \wColumn_8[18] , \wPDiag_8[50] , \wPDiag_8[49] , 
        \wNDiag_18[6] , \wPDiag_50[4] , \wColumn_56[47] , \wScan_30[4] , 
        \wPDiag_14[54] , \wColumn_36[43] , \wColumn_60[42] , \wNDiag_36[36] , 
        \wPDiag_42[55] , \wNDiag_60[37] , \wNDiag_56[32] , \wScan_3[0] , 
        \wColumn_3[27] , \wNDiag_6[45] , \wColumn_8[32] , \wPDiag_8[63] , 
        \wColumn_15[58] , \wColumn_15[41] , \wPDiag_22[51] , \wPDiag_22[48] , 
        \wPDiag_53[7] , \wPDiag_57[61] , \wColumn_43[59] , \wScan_54[0] , 
        \wColumn_23[44] , \wColumn_43[40] , \wPDiag_22[62] , \wNDiag_23[31] , 
        \wPDiag_34[0] , \wNDiag_23[28] , \wNDiag_15[34] , \wPDiag_37[3] , 
        \wNDiag_56[18] , \wPDiag_57[52] , \wPDiag_37[56] , \wNDiag_43[35] , 
        \wScan_57[3] , \wPDiag_61[57] , \wNDiag_7[5] , \wColumn_28[48] , 
        \wColumn_48[55] , \wPDiag_17[24] , \wColumn_28[51] , \wPDiag_62[14] , 
        \wColumn_19[4] , \wPDiag_21[21] , \wPDiag_34[15] , \wNDiag_35[46] , 
        \wPDiag_41[25] , \wNDiag_63[47] , \wPDiag_54[11] , \wPDiag_21[38] , 
        \wNDiag_55[42] , \wColumn_3[14] , \wPDiag_3[45] , \wNDiag_4[6] , 
        \wColumn_8[8] , \wScan_28[6] , \wNDiag_28[24] , \wPDiag_48[6] , 
        \wNDiag_48[39] , \wNDiag_48[20] , \wColumn_55[37] , \wColumn_35[33] , 
        \wPDiag_55[9] , \wColumn_63[32] , \wNDiag_16[44] , \wPDiag_17[17] , 
        \wNDiag_20[58] , \wPDiag_21[12] , \wNDiag_20[41] , \wPDiag_54[22] , 
        \wPDiag_34[26] , \wNDiag_40[45] , \wPDiag_62[27] , \wPDiag_41[16] , 
        \wNDiag_5[35] , \wColumn_28[62] , \wColumn_16[31] , \wColumn_16[28] , 
        \wColumn_40[30] , \wColumn_63[18] , \wColumn_20[34] , \wColumn_35[19] , 
        \wColumn_40[29] , \wNDiag_48[13] , \wPDiag_49[59] , \wPDiag_49[40] , 
        \wNDiag_28[17] , \wPDiag_29[44] , \wPDiag_5[4] , \wPDiag_6[7] , 
        \wPDiag_13[24] , \wNDiag_31[46] , \wColumn_59[61] , \wColumn_7[27] , 
        \wPDiag_25[38] , \wPDiag_25[21] , \wPDiag_30[15] , \wNDiag_43[7] , 
        \wPDiag_45[25] , \wPDiag_50[11] , \wNDiag_51[42] , \wColumn_59[4] , 
        \wNDiag_40[4] , \wPDiag_58[47] , \wNDiag_59[14] , \wPDiag_38[43] , 
        \wNDiag_39[10] , \wNDiag_1[35] , \wPDiag_7[45] , \wNDiag_9[50] , 
        \wColumn_31[33] , \wColumn_51[37] , \wNDiag_9[49] , \wPDiag_15[9] , 
        \wColumn_47[8] , \wNDiag_12[44] , \wPDiag_13[17] , \wNDiag_24[58] , 
        \wPDiag_25[12] , \wPDiag_50[22] , \wNDiag_24[41] , \wNDiag_27[3] , 
        \wNDiag_44[45] , \wPDiag_45[16] , \wPDiag_30[26] , \wColumn_39[56] , 
        \wColumn_59[52] , \wColumn_4[57] , \wColumn_7[14] , \wNDiag_9[63] , 
        \wColumn_44[30] , \wColumn_12[31] , \wColumn_12[28] , \wColumn_31[19] , 
        \wColumn_44[29] , \wColumn_24[34] , \wNDiag_24[0] , \wNDiag_39[23] , 
        \wReturn_34[0] , \wNDiag_59[27] , \wPDiag_10[54] , \wPDiag_10[4] , 
        \wNDiag_58[6] , \wColumn_19[24] , \wNDiag_19[51] , \wNDiag_19[48] , 
        \wColumn_42[5] , \wColumn_32[43] , \wNDiag_45[9] , \wColumn_52[47] , 
        \wPDiag_46[55] , \wColumn_11[41] , \wPDiag_13[7] , \wPDiag_26[51] , 
        \wPDiag_26[48] , \wNDiag_32[36] , \wNDiag_52[32] , \wColumn_41[6] , 
        \wPDiag_53[61] , \wColumn_47[59] , \wScan_14[0] , \wColumn_47[40] , 
        \wColumn_1[46] , \wPDiag_1[24] , \wNDiag_1[9] , \wNDiag_2[45] , 
        \wPDiag_4[35] , \wColumn_11[58] , \wNDiag_11[34] , \wPDiag_18[31] , 
        \wPDiag_18[28] , \wColumn_27[44] , \wNDiag_19[62] , \wColumn_25[2] , 
        \wColumn_26[1] , \wPDiag_26[62] , \wNDiag_27[31] , \wNDiag_52[18] , 
        \wPDiag_53[52] , \wNDiag_27[28] , \wPDiag_33[56] , \wNDiag_47[35] , 
        \wScan_17[3] , \wColumn_19[17] , \wPDiag_8[52] , \wPDiag_14[56] , 
        \wPDiag_22[53] , \wNDiag_23[19] , \wNDiag_56[30] , \wPDiag_42[57] , 
        \wPDiag_53[5] , \wNDiag_56[29] , \wPDiag_57[63] , \wNDiag_60[35] , 
        \wScan_33[5] , \wNDiag_36[34] , \wColumn_36[58] , \wColumn_36[41] , 
        \wColumn_60[40] , \wColumn_56[45] , \wColumn_60[59] , \wScan_30[6] , 
        \wCall_36[0] , \wPDiag_50[6] , \wColumn_3[25] , \wNDiag_4[4] , 
        \wNDiag_6[47] , \wNDiag_18[4] , \wColumn_8[30] , \wColumn_8[29] , 
        \wNDiag_15[36] , \wPDiag_37[54] , \wScan_57[1] , \wPDiag_37[1] , 
        \wNDiag_43[37] , \wPDiag_61[55] , \wNDiag_23[33] , \wPDiag_57[49] , 
        \wPDiag_8[61] , \wPDiag_22[60] , \wPDiag_57[50] , \wColumn_23[46] , 
        \wPDiag_34[2] , \wColumn_15[43] , \wColumn_16[19] , \wColumn_43[42] , 
        \wScan_54[2] , \wColumn_35[31] , \wColumn_63[29] , \wScan_28[4] , 
        \wColumn_35[28] , \wColumn_40[18] , \wColumn_63[30] , \wPDiag_48[4] , 
        \wNDiag_48[22] , \wColumn_55[35] , \wColumn_3[16] , \wNDiag_7[7] , 
        \wPDiag_17[26] , \wColumn_19[6] , \wPDiag_21[23] , \wNDiag_28[26] , 
        \wPDiag_54[13] , \wNDiag_55[59] , \wNDiag_35[44] , \wNDiag_55[40] , 
        \wPDiag_34[17] , \wPDiag_62[16] , \wPDiag_41[27] , \wNDiag_63[45] , 
        \wColumn_28[53] , \wPDiag_56[8] , \wPDiag_29[46] , \wColumn_48[57] , 
        \wPDiag_3[47] , \wNDiag_5[37] , \wColumn_16[33] , \wColumn_20[36] , 
        \wNDiag_28[15] , \wNDiag_48[11] , \wPDiag_49[42] , \wColumn_40[32] , 
        \wNDiag_7[54] , \wColumn_9[23] , \wColumn_14[50] , \wNDiag_16[46] , 
        \wPDiag_17[15] , \wColumn_28[60] , \wNDiag_40[47] , \wPDiag_62[25] , 
        \wPDiag_41[14] , \wNDiag_20[43] , \wPDiag_21[10] , \wPDiag_34[24] , 
        \wPDiag_54[20] , \wPDiag_54[39] , \wColumn_22[55] , \wPDiag_39[7] , 
        \wColumn_42[48] , \wColumn_61[60] , \wColumn_14[49] , \wColumn_37[61] , 
        \wColumn_42[51] , \wNDiag_14[25] , \wPDiag_24[8] , \wNDiag_61[15] , 
        \wNDiag_22[20] , \wPDiag_36[47] , \wNDiag_37[14] , \wNDiag_42[24] , 
        \wPDiag_60[46] , \wNDiag_57[10] , \wNDiag_22[39] , \wPDiag_56[43] , 
        \wPDiag_1[17] , \wColumn_3[1] , \wPDiag_9[58] , \wColumn_14[63] , 
        \wNDiag_15[1] , \wColumn_37[52] , \wColumn_61[53] , \wColumn_42[62] , 
        \wPDiag_9[41] , \wColumn_57[56] , \wColumn_2[36] , \wPDiag_2[54] , 
        \wNDiag_4[24] , \wColumn_9[10] , \wNDiag_16[2] , \wNDiag_22[13] , 
        \wPDiag_23[59] , \wPDiag_23[40] , \wNDiag_57[23] , \wNDiag_14[16] , 
        \wPDiag_15[45] , \wNDiag_37[27] , \wPDiag_43[44] , \wNDiag_61[26] , 
        \wNDiag_17[55] , \wPDiag_35[37] , \wNDiag_41[54] , \wNDiag_42[17] , 
        \wPDiag_63[36] , \wNDiag_21[50] , \wNDiag_21[49] , \wScan_42[6] , 
        \wPDiag_55[33] , \wNDiag_54[60] , \wPDiag_22[6] , \wCall_44[0] , 
        \wNDiag_4[17] , \wColumn_14[3] , \wColumn_17[39] , \wColumn_21[25] , 
        \wPDiag_21[5] , \wColumn_54[15] , \wColumn_41[21] , \wColumn_17[20] , 
        \wColumn_34[11] , \wColumn_41[38] , \wColumn_62[10] , \wPDiag_28[55] , 
        \wScan_41[5] , \wPDiag_48[51] , \wPDiag_48[48] , \wPDiag_46[2] , 
        \wColumn_29[59] , \wColumn_29[40] , \wColumn_49[44] , \wNDiag_9[1] , 
        \wPDiag_16[35] , \wPDiag_20[30] , \wPDiag_20[29] , \wNDiag_21[63] , 
        \wNDiag_54[53] , \wPDiag_55[19] , \wScan_26[2] , \wNDiag_34[57] , 
        \wPDiag_40[34] , \wNDiag_49[31] , \wNDiag_62[56] , \wPDiag_48[62] , 
        \wNDiag_49[28] , \wColumn_13[22] , \wColumn_17[13] , \wScan_25[1] , 
        \wNDiag_29[35] , \wColumn_34[22] , \wColumn_41[12] , \wColumn_17[0] , 
        \wPDiag_45[1] , \wColumn_62[23] , \wColumn_21[16] , \wNDiag_29[5] , 
        \wColumn_30[13] , \wNDiag_38[30] , \wColumn_54[26] , \wNDiag_38[29] , 
        \wPDiag_39[63] , \wColumn_45[23] , \wNDiag_58[34] , \wColumn_33[6] , 
        \wPDiag_61[7] , \wPDiag_6[56] , \wColumn_25[27] , \wColumn_50[17] , 
        \wPDiag_8[1] , \wNDiag_13[57] , \wPDiag_24[18] , \wNDiag_25[52] , 
        \wColumn_30[5] , \wColumn_38[45] , \wReturn_46[0] , \wColumn_58[58] , 
        \wColumn_58[41] , \wNDiag_37[9] , \wPDiag_62[4] , \wNDiag_50[62] , 
        \wPDiag_51[31] , \wPDiag_51[28] , \wPDiag_31[35] , \wNDiag_45[56] , 
        \wColumn_25[14] , \wColumn_1[56] , \wColumn_2[26] , \wReturn_3[0] , 
        \wNDiag_3[56] , \wPDiag_5[26] , \wColumn_6[34] , \wNDiag_8[43] , 
        \wColumn_30[20] , \wColumn_50[24] , \wColumn_45[10] , \wColumn_13[11] , 
        \wColumn_30[39] , \wColumn_57[2] , \wPDiag_12[37] , \wPDiag_39[50] , 
        \wPDiag_39[49] , \wPDiag_59[54] , \wPDiag_24[32] , \wNDiag_30[55] , 
        \wPDiag_44[36] , \wNDiag_25[61] , \wNDiag_50[48] , \wNDiag_32[4] , 
        \wNDiag_50[51] , \wColumn_54[1] , \wColumn_28[7] , \wColumn_10[52] , 
        \wNDiag_10[27] , \wNDiag_26[22] , \wPDiag_52[58] , \wNDiag_53[12] , 
        \wPDiag_52[41] , \wScan_19[5] , \wPDiag_19[22] , \wPDiag_32[45] , 
        \wNDiag_33[16] , \wNDiag_46[26] , \wColumn_35[8] , \wNDiag_10[14] , 
        \wColumn_26[57] , \wNDiag_31[7] , \wColumn_33[63] , \wColumn_46[53] , 
        \wColumn_5[44] , \wPDiag_5[15] , \wPDiag_11[47] , \wNDiag_33[25] , 
        \wPDiag_47[46] , \wColumn_18[37] , \wNDiag_26[11] , \wNDiag_46[15] , 
        \wPDiag_27[42] , \wNDiag_53[21] , \wNDiag_53[38] , \wNDiag_56[0] , 
        \wColumn_10[61] , \wColumn_53[54] , \wNDiag_55[3] , \wColumn_33[50] , 
        \wColumn_33[49] , \wColumn_46[60] , \wColumn_6[5] , \wNDiag_13[6] , 
        \wPDiag_16[25] , \wNDiag_18[42] , \wPDiag_19[11] , \wColumn_29[50] , 
        \wColumn_49[54] , \wColumn_29[49] , \wNDiag_34[47] , \wPDiag_35[14] , 
        \wPDiag_40[24] , \wNDiag_62[46] , \wPDiag_20[39] , \wPDiag_63[15] , 
        \wNDiag_54[43] , \wNDiag_10[5] , \wPDiag_20[20] , \wPDiag_55[10] , 
        \wNDiag_29[25] , \wColumn_2[15] , \wPDiag_2[44] , \wColumn_5[6] , 
        \wNDiag_9[8] , \wNDiag_49[38] , \wPDiag_16[16] , \wColumn_17[9] , 
        \wColumn_34[32] , \wNDiag_49[21] , \wColumn_54[36] , \wPDiag_58[7] , 
        \wColumn_62[33] , \wNDiag_17[45] , \wPDiag_20[13] , \wNDiag_21[59] , 
        \wNDiag_21[40] , \wPDiag_45[8] , \wPDiag_55[23] , \wPDiag_40[17] , 
        \wPDiag_35[27] , \wNDiag_41[44] , \wPDiag_63[26] , \wColumn_29[63] , 
        \wNDiag_4[34] , \wColumn_17[30] , \wColumn_34[18] , \wColumn_41[28] , 
        \wColumn_17[29] , \wColumn_41[31] , \wColumn_62[19] , \wColumn_21[35] , 
        \wPDiag_28[45] , \wNDiag_29[16] , \wPDiag_48[58] , \wPDiag_48[41] , 
        \wNDiag_49[12] , \wPDiag_1[34] , \wColumn_3[8] , \wPDiag_9[51] , 
        \wColumn_12[4] , \wPDiag_40[5] , \wPDiag_9[48] , \wNDiag_15[8] , 
        \wScan_20[5] , \wScan_23[6] , \wColumn_37[42] , \wColumn_57[46] , 
        \wColumn_61[43] , \wColumn_9[33] , \wColumn_9[19] , \wColumn_11[7] , 
        \wPDiag_15[55] , \wPDiag_23[50] , \wNDiag_37[37] , \wPDiag_43[54] , 
        \wNDiag_61[36] , \wCall_25[0] , \wPDiag_43[6] , \wPDiag_23[49] , 
        \wPDiag_56[60] , \wPDiag_9[62] , \wColumn_14[59] , \wColumn_42[41] , 
        \wNDiag_57[33] , \wColumn_14[40] , \wColumn_42[58] , \wScan_44[1] , 
        \wColumn_22[45] , \wPDiag_24[1] , \wNDiag_14[35] , \wNDiag_22[30] , 
        \wNDiag_22[29] , \wPDiag_56[53] , \wNDiag_57[19] , \wPDiag_23[63] , 
        \wPDiag_36[57] , \wNDiag_42[34] , \wPDiag_60[56] , \wPDiag_27[2] , 
        \wNDiag_3[46] , \wColumn_5[54] , \wNDiag_7[44] , \wScan_47[2] , 
        \wScan_8[2] , \wPDiag_11[57] , \wNDiag_26[18] , \wPDiag_27[52] , 
        \wColumn_51[5] , \wNDiag_53[28] , \wPDiag_52[62] , \wNDiag_53[31] , 
        \wColumn_18[27] , \wReturn_27[0] , \wNDiag_33[35] , \wPDiag_47[56] , 
        \wNDiag_56[9] , \wColumn_33[59] , \wColumn_33[40] , \wScan_63[4] , 
        \wNDiag_18[52] , \wPDiag_19[18] , \wColumn_53[44] , \wColumn_52[6] , 
        \wNDiag_48[5] , \wPDiag_5[36] , \wColumn_18[14] , \wPDiag_8[8] , 
        \wNDiag_8[53] , \wColumn_10[42] , \wNDiag_10[37] , \wPDiag_32[55] , 
        \wColumn_35[1] , \wNDiag_46[36] , \wNDiag_18[61] , \wPDiag_19[32] , 
        \wNDiag_26[32] , \wPDiag_27[61] , \wPDiag_52[51] , \wPDiag_52[48] , 
        \wColumn_36[2] , \wColumn_26[47] , \wColumn_46[43] , \wColumn_13[18] , 
        \wColumn_30[29] , \wColumn_45[19] , \wColumn_30[30] , \wColumn_50[34] , 
        \wColumn_6[24] , \wPDiag_18[5] , \wNDiag_38[13] , \wPDiag_39[40] , 
        \wPDiag_39[59] , \wNDiag_50[7] , \wNDiag_58[17] , \wColumn_6[17] , 
        \wPDiag_12[27] , \wPDiag_24[22] , \wColumn_49[7] , \wPDiag_59[44] , 
        \wNDiag_50[41] , \wNDiag_30[45] , \wPDiag_31[16] , \wNDiag_50[58] , 
        \wPDiag_51[12] , \wPDiag_44[26] , \wNDiag_53[4] , \wColumn_54[8] , 
        \wColumn_58[62] , \wNDiag_58[24] , \wPDiag_6[46] , \wNDiag_8[60] , 
        \wColumn_13[32] , \wColumn_25[37] , \wNDiag_34[3] , \wNDiag_38[39] , 
        \wNDiag_38[20] , \wColumn_45[33] , \wColumn_38[55] , \wColumn_58[51] , 
        \wColumn_11[48] , \wPDiag_12[14] , \wNDiag_13[47] , \wPDiag_44[15] , 
        \wColumn_58[48] , \wPDiag_31[25] , \wNDiag_45[46] , \wNDiag_21[4] , 
        \wPDiag_24[11] , \wNDiag_25[42] , \wNDiag_37[0] , \wPDiag_51[38] , 
        \wPDiag_51[21] , \wColumn_27[54] , \wColumn_32[60] , \wColumn_47[50] , 
        \wColumn_47[49] , \wNDiag_1[25] , \wNDiag_2[55] , \wColumn_11[51] , 
        \wNDiag_11[24] , \wPDiag_18[38] , \wPDiag_18[21] , \wColumn_26[8] , 
        \wNDiag_32[15] , \wNDiag_47[25] , \wNDiag_27[38] , \wPDiag_33[46] , 
        \wPDiag_53[42] , \wNDiag_27[21] , \wNDiag_52[11] , \wColumn_38[4] , 
        \wPDiag_3[3] , \wColumn_4[47] , \wPDiag_4[25] , \wPDiag_18[12] , 
        \wNDiag_19[58] , \wNDiag_22[7] , \wNDiag_19[41] , \wPDiag_4[16] , 
        \wColumn_11[62] , \wColumn_32[53] , \wColumn_47[63] , \wNDiag_45[0] , 
        \wColumn_52[57] , \wNDiag_46[3] , \wScan_6[4] , \wPDiag_10[44] , 
        \wColumn_19[34] , \wPDiag_26[58] , \wPDiag_26[41] , \wNDiag_27[12] , 
        \wNDiag_32[26] , \wNDiag_52[22] , \wNDiag_11[17] , \wNDiag_47[16] , 
        \wPDiag_46[45] , \wNDiag_12[54] , \wPDiag_30[36] , \wColumn_20[6] , 
        \wNDiag_24[51] , \wNDiag_44[55] , \wNDiag_51[61] , \wNDiag_24[48] , 
        \wPDiag_50[32] , \wColumn_39[46] , \wNDiag_1[16] , \wPDiag_7[55] , 
        \wColumn_59[42] , \wScan_11[4] , \wColumn_12[38] , \wColumn_12[21] , 
        \wColumn_23[5] , \wColumn_24[24] , \wColumn_51[14] , \wNDiag_39[6] , 
        \wColumn_44[39] , \wColumn_44[20] , \wReturn_55[0] , \wNDiag_24[9] , 
        \wColumn_31[10] , \wPDiag_38[60] , \wNDiag_59[37] , \wPDiag_16[3] , 
        \wNDiag_39[33] , \wColumn_44[2] , \wNDiag_1[0] , \wNDiag_2[3] , 
        \wColumn_3[35] , \wPDiag_3[57] , \wColumn_7[37] , \wPDiag_13[34] , 
        \wNDiag_24[62] , \wPDiag_25[31] , \wPDiag_25[28] , \wPDiag_50[18] , 
        \wNDiag_51[52] , \wPDiag_45[35] , \wNDiag_31[56] , \wPDiag_38[53] , 
        \wNDiag_39[19] , \wNDiag_9[59] , \wColumn_12[12] , \wPDiag_58[57] , 
        \wPDiag_15[0] , \wNDiag_9[40] , \wColumn_31[23] , \wColumn_47[1] , 
        \wColumn_44[13] , \wColumn_16[23] , \wColumn_24[17] , \wPDiag_29[56] , 
        \wNDiag_48[18] , \wPDiag_49[52] , \wColumn_51[27] , \wScan_51[6] , 
        \wColumn_63[13] , \wColumn_20[26] , \wColumn_35[12] , \wColumn_40[22] , 
        \wColumn_55[16] , \wPDiag_31[6] , \wCall_57[0] , \wColumn_63[7] , 
        \wNDiag_5[27] , \wPDiag_32[5] , \wColumn_60[4] , \wColumn_8[3] , 
        \wColumn_16[10] , \wNDiag_16[56] , \wNDiag_20[53] , \wPDiag_21[19] , 
        \wPDiag_54[29] , \wNDiag_55[63] , \wPDiag_34[34] , \wScan_52[5] , 
        \wPDiag_54[30] , \wColumn_20[15] , \wNDiag_40[57] , \wPDiag_62[35] , 
        \wColumn_35[38] , \wColumn_55[25] , \wPDiag_55[2] , \wColumn_63[20] , 
        \wNDiag_28[36] , \wColumn_35[21] , \wColumn_40[11] , \wColumn_63[39] , 
        \wNDiag_5[14] , \wPDiag_17[36] , \wScan_35[2] , \wScan_36[1] , 
        \wNDiag_48[32] , \wPDiag_49[61] , \wPDiag_41[37] , \wNDiag_63[55] , 
        \wNDiag_20[60] , \wNDiag_35[54] , \wPDiag_21[33] , \wNDiag_55[50] , 
        \wColumn_48[47] , \wNDiag_55[49] , \wNDiag_6[57] , \wColumn_28[43] , 
        \wPDiag_56[1] , \wNDiag_62[5] , \wColumn_8[39] , \wColumn_8[20] , 
        \wPDiag_57[40] , \wPDiag_14[46] , \wColumn_15[53] , \wNDiag_15[26] , 
        \wNDiag_23[23] , \wNDiag_56[13] , \wPDiag_57[59] , \wNDiag_36[17] , 
        \wPDiag_37[8] , \wNDiag_43[27] , \wPDiag_61[45] , \wNDiag_60[16] , 
        \wColumn_36[62] , \wPDiag_37[44] , \wColumn_43[52] , \wScan_49[4] , 
        \wNDiag_61[6] , \wColumn_60[63] , \wColumn_23[56] , \wPDiag_29[4] , 
        \wNDiag_36[24] , \wNDiag_15[15] , \wNDiag_43[14] , \wPDiag_42[47] , 
        \wNDiag_60[25] , \wColumn_8[13] , \wPDiag_22[43] , \wPDiag_8[42] , 
        \wNDiag_23[10] , \wNDiag_56[39] , \wNDiag_56[20] , \wColumn_15[60] , 
        \wColumn_36[51] , \wColumn_56[55] , \wColumn_43[61] , \wColumn_60[49] , 
        \wColumn_36[48] , \wColumn_60[50] , \wNDiag_3[61] , \wNDiag_3[52] , 
        \wColumn_10[56] , \wColumn_26[53] , \wColumn_53[63] , \wNDiag_31[3] , 
        \wColumn_46[57] , \wNDiag_10[23] , \wScan_19[1] , \wPDiag_19[26] , 
        \wPDiag_32[58] , \wNDiag_46[22] , \wNDiag_33[12] , \wColumn_18[19] , 
        \wNDiag_26[26] , \wPDiag_32[41] , \wPDiag_52[45] , \wNDiag_53[16] , 
        \wColumn_28[3] , \wColumn_5[59] , \wColumn_5[40] , \wPDiag_5[22] , 
        \wNDiag_18[46] , \wPDiag_19[15] , \wNDiag_32[0] , \wPDiag_5[11] , 
        \wColumn_26[60] , \wColumn_33[54] , \wNDiag_48[8] , \wColumn_53[49] , 
        \wColumn_53[50] , \wNDiag_55[7] , \wNDiag_56[4] , \wPDiag_6[52] , 
        \wNDiag_10[10] , \wPDiag_11[43] , \wColumn_18[33] , \wNDiag_26[15] , 
        \wPDiag_27[46] , \wNDiag_33[21] , \wColumn_51[8] , \wNDiag_53[25] , 
        \wNDiag_33[38] , \wNDiag_46[11] , \wPDiag_12[19] , \wNDiag_13[53] , 
        \wPDiag_31[31] , \wPDiag_47[42] , \wNDiag_25[56] , \wNDiag_30[62] , 
        \wPDiag_31[28] , \wPDiag_44[18] , \wNDiag_45[52] , \wColumn_30[1] , 
        \wColumn_38[58] , \wPDiag_51[35] , \wColumn_38[41] , \wPDiag_62[0] , 
        \wColumn_58[45] , \wColumn_6[30] , \wColumn_6[29] , \wPDiag_6[61] , 
        \wColumn_13[26] , \wColumn_25[23] , \wColumn_50[13] , \wNDiag_29[1] , 
        \wColumn_33[2] , \wPDiag_61[3] , \wColumn_30[17] , \wColumn_45[27] , 
        \wNDiag_38[34] , \wNDiag_58[30] , \wNDiag_58[29] , \wPDiag_59[63] , 
        \wColumn_54[5] , \wPDiag_12[33] , \wNDiag_13[60] , \wReturn_22[0] , 
        \wPDiag_24[36] , \wNDiag_50[55] , \wNDiag_30[48] , \wPDiag_44[32] , 
        \wNDiag_53[9] , \wPDiag_18[8] , \wNDiag_30[51] , \wPDiag_39[54] , 
        \wNDiag_45[61] , \wPDiag_59[49] , \wNDiag_8[47] , \wColumn_13[15] , 
        \wPDiag_59[50] , \wColumn_30[24] , \wColumn_57[6] , \wColumn_45[14] , 
        \wColumn_25[10] , \wColumn_1[42] , \wPDiag_1[39] , \wPDiag_1[20] , 
        \wColumn_2[32] , \wColumn_2[18] , \wPDiag_8[5] , \wColumn_50[20] , 
        \wPDiag_28[48] , \wScan_41[1] , \wPDiag_48[55] , \wColumn_50[39] , 
        \wPDiag_2[50] , \wPDiag_2[49] , \wColumn_17[24] , \wPDiag_28[51] , 
        \wColumn_62[14] , \wColumn_21[38] , \wColumn_21[21] , \wColumn_34[15] , 
        \wColumn_41[25] , \wColumn_54[11] , \wPDiag_21[1] , \wNDiag_4[39] , 
        \wNDiag_4[20] , \wPDiag_22[2] , \wColumn_17[17] , \wNDiag_17[51] , 
        \wNDiag_21[54] , \wPDiag_35[33] , \wNDiag_41[49] , \wScan_42[2] , 
        \wPDiag_55[37] , \wNDiag_62[61] , \wNDiag_17[48] , \wNDiag_34[60] , 
        \wNDiag_41[50] , \wPDiag_63[32] , \wColumn_21[12] , \wColumn_54[22] , 
        \wColumn_17[4] , \wPDiag_45[5] , \wColumn_62[27] , \wNDiag_29[31] , 
        \wColumn_34[26] , \wColumn_41[16] , \wPDiag_2[63] , \wNDiag_4[13] , 
        \wColumn_6[8] , \wNDiag_9[5] , \wNDiag_10[8] , \wScan_25[5] , 
        \wPDiag_28[62] , \wNDiag_29[28] , \wPDiag_16[31] , \wPDiag_16[28] , 
        \wNDiag_49[35] , \wNDiag_17[62] , \wScan_26[6] , \wPDiag_40[30] , 
        \wNDiag_62[52] , \wPDiag_63[18] , \wNDiag_34[53] , \wPDiag_35[19] , 
        \wPDiag_40[29] , \wNDiag_41[63] , \wPDiag_20[34] , \wNDiag_54[57] , 
        \wColumn_49[59] , \wColumn_49[40] , \wColumn_14[7] , \wCall_20[0] , 
        \wColumn_29[44] , \wPDiag_46[6] , \wPDiag_1[13] , \wColumn_3[5] , 
        \wNDiag_7[63] , \wNDiag_7[50] , \wNDiag_7[49] , \wColumn_9[27] , 
        \wColumn_9[14] , \wColumn_14[54] , \wNDiag_14[38] , \wNDiag_22[24] , 
        \wPDiag_56[47] , \wNDiag_57[14] , \wNDiag_42[20] , \wPDiag_60[42] , 
        \wNDiag_14[21] , \wNDiag_37[10] , \wNDiag_42[39] , \wNDiag_61[11] , 
        \wPDiag_36[43] , \wColumn_42[55] , \wScan_59[3] , \wNDiag_14[12] , 
        \wPDiag_15[58] , \wPDiag_15[41] , \wColumn_22[51] , \wColumn_22[48] , 
        \wColumn_57[61] , \wNDiag_37[23] , \wPDiag_39[3] , \wNDiag_42[13] , 
        \wPDiag_43[59] , \wPDiag_23[44] , \wPDiag_43[40] , \wNDiag_61[22] , 
        \wNDiag_16[6] , \wNDiag_22[17] , \wNDiag_57[27] , \wPDiag_9[45] , 
        \wNDiag_15[5] , \wColumn_22[62] , \wColumn_37[56] , \wColumn_57[52] , 
        \wColumn_61[57] , \wNDiag_2[58] , \wNDiag_2[41] , \wColumn_3[38] , 
        \wNDiag_5[19] , \wColumn_12[9] , \wPDiag_40[8] , \wNDiag_7[3] , 
        \wColumn_28[57] , \wColumn_48[53] , \wPDiag_17[22] , \wPDiag_34[13] , 
        \wNDiag_35[59] , \wNDiag_35[40] , \wPDiag_41[23] , \wNDiag_63[41] , 
        \wColumn_19[2] , \wPDiag_62[12] , \wNDiag_63[58] , \wPDiag_21[27] , 
        \wNDiag_55[44] , \wPDiag_54[17] , \wColumn_3[21] , \wNDiag_28[22] , 
        \wColumn_3[12] , \wPDiag_3[43] , \wNDiag_4[0] , \wColumn_20[18] , 
        \wScan_28[0] , \wPDiag_48[0] , \wNDiag_48[26] , \wColumn_55[31] , 
        \wColumn_55[28] , \wNDiag_16[42] , \wNDiag_20[47] , \wColumn_35[35] , 
        \wColumn_63[34] , \wPDiag_21[14] , \wPDiag_54[24] , \wPDiag_41[10] , 
        \wPDiag_62[38] , \wPDiag_17[11] , \wPDiag_34[20] , \wNDiag_40[43] , 
        \wPDiag_62[21] , \wPDiag_34[39] , \wNDiag_5[33] , \wPDiag_32[8] , 
        \wColumn_48[60] , \wColumn_60[9] , \wColumn_16[37] , \wColumn_20[32] , 
        \wColumn_40[36] , \wNDiag_28[11] , \wNDiag_48[15] , \wPDiag_49[46] , 
        \wPDiag_29[42] , \wColumn_4[53] , \wNDiag_6[43] , \wColumn_8[34] , 
        \wPDiag_8[56] , \wNDiag_18[0] , \wPDiag_50[2] , \wPDiag_14[52] , 
        \wNDiag_15[18] , \wScan_30[2] , \wScan_33[1] , \wColumn_36[45] , 
        \wColumn_56[58] , \wColumn_56[41] , \wColumn_60[44] , \wColumn_15[47] , 
        \wPDiag_22[57] , \wNDiag_36[30] , \wNDiag_36[29] , \wPDiag_37[63] , 
        \wNDiag_60[28] , \wPDiag_61[62] , \wPDiag_42[53] , \wNDiag_43[19] , 
        \wNDiag_60[31] , \wColumn_43[46] , \wPDiag_53[1] , \wNDiag_56[34] , 
        \wColumn_23[42] , \wPDiag_29[9] , \wScan_54[6] , \wPDiag_34[6] , 
        \wCall_52[0] , \wPDiag_14[61] , \wNDiag_23[37] , \wPDiag_57[54] , 
        \wPDiag_37[49] , \wNDiag_43[33] , \wPDiag_61[51] , \wNDiag_15[32] , 
        \wPDiag_37[50] , \wPDiag_42[60] , \wPDiag_61[48] , \wPDiag_37[5] , 
        \wScan_57[5] , \wNDiag_62[8] , \wPDiag_10[50] , \wPDiag_13[3] , 
        \wPDiag_26[55] , \wColumn_41[2] , \wNDiag_52[36] , \wPDiag_10[49] , 
        \wNDiag_32[32] , \wPDiag_46[48] , \wPDiag_10[0] , \wColumn_19[39] , 
        \wPDiag_33[61] , \wPDiag_46[51] , \wColumn_19[20] , \wNDiag_19[55] , 
        \wColumn_32[47] , \wColumn_52[43] , \wColumn_42[1] , \wNDiag_58[2] , 
        \wColumn_19[13] , \wColumn_38[9] , \wColumn_4[60] , \wPDiag_4[31] , 
        \wPDiag_4[28] , \wPDiag_10[63] , \wNDiag_47[31] , \wNDiag_11[30] , 
        \wNDiag_11[29] , \wColumn_25[6] , \wNDiag_32[18] , \wPDiag_46[62] , 
        \wNDiag_47[28] , \wPDiag_33[52] , \wNDiag_27[35] , \wPDiag_53[56] , 
        \wPDiag_18[35] , \wColumn_26[5] , \wReturn_50[0] , \wColumn_27[59] , 
        \wColumn_27[40] , \wColumn_47[44] , \wColumn_1[61] , \wColumn_1[52] , 
        \wNDiag_1[38] , \wNDiag_1[31] , \wNDiag_1[28] , \wScan_3[4] , 
        \wPDiag_5[0] , \wNDiag_9[54] , \wColumn_11[45] , \wNDiag_21[9] , 
        \wScan_14[4] , \wColumn_31[37] , \wPDiag_38[47] , \wColumn_51[33] , 
        \wNDiag_39[14] , \wNDiag_40[0] , \wNDiag_59[10] , \wPDiag_6[3] , 
        \wColumn_7[23] , \wPDiag_13[39] , \wPDiag_25[25] , \wNDiag_51[46] , 
        \wPDiag_58[43] , \wColumn_59[0] , \wPDiag_30[11] , \wPDiag_50[15] , 
        \wPDiag_13[20] , \wNDiag_31[42] , \wPDiag_45[21] , \wNDiag_43[3] , 
        \wPDiag_45[38] , \wColumn_7[10] , \wColumn_39[61] , \wNDiag_59[23] , 
        \wColumn_12[35] , \wColumn_23[8] , \wNDiag_24[4] , \wNDiag_39[27] , 
        \wColumn_24[30] , \wColumn_24[29] , \wColumn_51[19] , \wColumn_44[34] , 
        \wColumn_39[52] , \wNDiag_1[21] , \wNDiag_1[4] , \wNDiag_6[53] , 
        \wPDiag_7[58] , \wPDiag_7[41] , \wColumn_59[56] , \wColumn_8[24] , 
        \wNDiag_12[59] , \wNDiag_12[40] , \wNDiag_44[58] , \wPDiag_45[12] , 
        \wPDiag_13[13] , \wPDiag_30[22] , \wNDiag_44[41] , \wColumn_15[57] , 
        \wColumn_23[52] , \wNDiag_24[45] , \wNDiag_27[7] , \wPDiag_25[16] , 
        \wPDiag_50[26] , \wColumn_56[62] , \wPDiag_29[0] , \wNDiag_15[22] , 
        \wColumn_43[56] , \wScan_49[0] , \wNDiag_61[2] , \wNDiag_60[12] , 
        \wPDiag_61[58] , \wNDiag_23[27] , \wNDiag_36[13] , \wPDiag_37[40] , 
        \wNDiag_43[23] , \wPDiag_61[41] , \wPDiag_37[59] , \wNDiag_56[17] , 
        \wPDiag_57[44] , \wNDiag_62[1] , \wNDiag_2[7] , \wNDiag_6[60] , 
        \wPDiag_8[46] , \wNDiag_18[9] , \wColumn_23[61] , \wColumn_36[55] , 
        \wColumn_60[54] , \wColumn_56[51] , \wColumn_56[48] , \wNDiag_23[14] , 
        \wPDiag_53[8] , \wNDiag_56[24] , \wColumn_3[31] , \wPDiag_3[60] , 
        \wPDiag_3[53] , \wNDiag_5[23] , \wColumn_8[17] , \wPDiag_22[47] , 
        \wPDiag_14[42] , \wNDiag_15[11] , \wNDiag_36[39] , \wNDiag_36[20] , 
        \wPDiag_42[43] , \wNDiag_60[21] , \wNDiag_16[52] , \wPDiag_17[18] , 
        \wPDiag_34[30] , \wPDiag_34[29] , \wNDiag_35[63] , \wNDiag_40[53] , 
        \wPDiag_41[19] , \wNDiag_43[10] , \wNDiag_60[38] , \wPDiag_62[31] , 
        \wPDiag_62[28] , \wNDiag_63[62] , \wNDiag_20[57] , \wScan_52[1] , 
        \wPDiag_54[34] , \wPDiag_32[1] , \wColumn_60[0] , \wColumn_16[27] , 
        \wColumn_20[22] , \wPDiag_31[2] , \wColumn_63[3] , \wColumn_55[12] , 
        \wColumn_35[16] , \wColumn_40[26] , \wColumn_63[17] , \wNDiag_28[18] , 
        \wPDiag_29[52] , \wPDiag_49[56] , \wScan_51[2] , \wPDiag_56[5] , 
        \wNDiag_5[10] , \wColumn_28[47] , \wColumn_48[43] , \wNDiag_16[61] , 
        \wPDiag_17[32] , \wPDiag_21[37] , \wNDiag_55[54] , \wNDiag_35[50] , 
        \wNDiag_40[60] , \wNDiag_63[48] , \wNDiag_35[49] , \wScan_36[5] , 
        \wPDiag_41[33] , \wPDiag_48[9] , \wNDiag_48[36] , \wNDiag_63[51] , 
        \wColumn_3[28] , \wPDiag_29[61] , \wScan_35[6] , \wNDiag_4[9] , 
        \wColumn_8[7] , \wNDiag_28[32] , \wColumn_35[25] , \wColumn_7[19] , 
        \wScan_11[0] , \wColumn_16[14] , \wColumn_40[15] , \wColumn_20[11] , 
        \wCall_33[0] , \wColumn_55[38] , \wPDiag_55[6] , \wColumn_63[24] , 
        \wNDiag_39[37] , \wColumn_55[21] , \wPDiag_58[60] , \wPDiag_7[51] , 
        \wColumn_12[25] , \wColumn_31[14] , \wColumn_44[24] , \wNDiag_59[33] , 
        \wNDiag_39[2] , \wColumn_23[1] , \wColumn_24[39] , \wColumn_24[20] , 
        \wColumn_51[10] , \wPDiag_7[48] , \wColumn_39[42] , \wColumn_59[46] , 
        \wColumn_20[2] , \wNDiag_1[12] , \wPDiag_5[9] , \wColumn_7[33] , 
        \wNDiag_9[44] , \wScan_12[3] , \wPDiag_50[36] , \wNDiag_12[50] , 
        \wNDiag_12[49] , \wNDiag_24[55] , \wNDiag_31[61] , \wNDiag_44[51] , 
        \wPDiag_30[32] , \wNDiag_44[48] , \wColumn_24[13] , \wReturn_31[0] , 
        \wColumn_31[27] , \wColumn_51[23] , \wColumn_44[17] , \wColumn_12[16] , 
        \wPDiag_15[4] , \wNDiag_40[9] , \wColumn_47[5] , \wNDiag_12[63] , 
        \wPDiag_13[30] , \wPDiag_38[57] , \wPDiag_58[53] , \wNDiag_59[19] , 
        \wPDiag_30[18] , \wNDiag_31[52] , \wNDiag_44[62] , \wPDiag_45[28] , 
        \wPDiag_13[29] , \wPDiag_25[35] , \wPDiag_45[31] , \wNDiag_51[56] , 
        \wColumn_59[9] , \wNDiag_2[62] , \wNDiag_2[51] , \wNDiag_2[48] , 
        \wPDiag_4[38] , \wPDiag_7[62] , \wPDiag_16[7] , \wColumn_44[6] , 
        \wPDiag_4[21] , \wNDiag_22[3] , \wColumn_38[0] , \wScan_6[0] , 
        \wPDiag_10[59] , \wColumn_11[55] , \wNDiag_11[39] , \wNDiag_11[20] , 
        \wNDiag_27[25] , \wNDiag_52[15] , \wNDiag_47[38] , \wPDiag_53[46] , 
        \wPDiag_33[42] , \wNDiag_47[21] , \wPDiag_18[25] , \wNDiag_32[11] , 
        \wNDiag_11[13] , \wNDiag_21[0] , \wColumn_27[50] , \wColumn_47[54] , 
        \wColumn_52[60] , \wColumn_27[49] , \wPDiag_46[41] , \wPDiag_10[40] , 
        \wNDiag_32[22] , \wColumn_19[30] , \wPDiag_26[45] , \wNDiag_27[16] , 
        \wPDiag_46[58] , \wNDiag_47[12] , \wNDiag_52[26] , \wNDiag_46[7] , 
        \wPDiag_3[7] , \wNDiag_3[42] , \wColumn_4[43] , \wPDiag_4[12] , 
        \wColumn_19[29] , \wColumn_27[63] , \wNDiag_45[4] , \wColumn_32[57] , 
        \wColumn_52[53] , \wScan_5[3] , \wColumn_5[63] , \wColumn_5[50] , 
        \wColumn_5[49] , \wReturn_6[0] , \wPDiag_10[9] , \wNDiag_19[45] , 
        \wColumn_42[8] , \wPDiag_18[16] , \wColumn_38[62] , \wColumn_6[39] , 
        \wColumn_6[20] , \wPDiag_12[23] , \wNDiag_30[41] , \wPDiag_24[26] , 
        \wNDiag_30[58] , \wNDiag_53[0] , \wPDiag_31[12] , \wPDiag_44[22] , 
        \wColumn_49[3] , \wPDiag_51[16] , \wNDiag_50[45] , \wPDiag_59[40] , 
        \wColumn_6[13] , \wPDiag_6[42] , \wNDiag_8[57] , \wPDiag_18[1] , 
        \wNDiag_38[17] , \wNDiag_50[3] , \wNDiag_58[13] , \wPDiag_59[59] , 
        \wColumn_25[19] , \wPDiag_39[44] , \wColumn_30[34] , \wColumn_50[30] , 
        \wColumn_50[29] , \wPDiag_12[10] , \wCall_19[0] , \wPDiag_24[15] , 
        \wPDiag_51[25] , \wNDiag_25[46] , \wNDiag_37[4] , \wNDiag_45[42] , 
        \wNDiag_13[43] , \wPDiag_31[38] , \wPDiag_44[11] , \wPDiag_31[21] , 
        \wColumn_13[36] , \wNDiag_29[8] , \wColumn_30[8] , \wColumn_38[51] , 
        \wColumn_58[55] , \wPDiag_62[9] , \wColumn_38[48] , \wColumn_45[37] , 
        \wColumn_25[33] , \wNDiag_34[7] , \wNDiag_38[24] , \wNDiag_58[39] , 
        \wNDiag_58[20] , \wPDiag_5[18] , \wScan_8[6] , \wNDiag_18[56] , 
        \wNDiag_48[1] , \wColumn_52[2] , \wColumn_18[23] , \wColumn_33[44] , 
        \wColumn_53[59] , \wColumn_53[40] , \wScan_60[3] , \wScan_63[0] , 
        \wColumn_10[46] , \wNDiag_10[19] , \wPDiag_11[53] , \wPDiag_32[62] , 
        \wNDiag_33[28] , \wNDiag_46[18] , \wPDiag_47[52] , \wPDiag_27[56] , 
        \wNDiag_33[31] , \wNDiag_53[35] , \wColumn_51[1] , \wPDiag_19[36] , 
        \wColumn_26[43] , \wColumn_46[47] , \wPDiag_5[32] , \wNDiag_10[33] , 
        \wNDiag_26[36] , \wColumn_36[6] , \wReturn_43[0] , \wPDiag_32[51] , 
        \wColumn_35[5] , \wPDiag_47[61] , \wPDiag_52[55] , \wPDiag_11[60] , 
        \wPDiag_32[48] , \wNDiag_46[32] , \wNDiag_32[9] , \wColumn_18[10] , 
        \wPDiag_9[55] , \wColumn_11[3] , \wPDiag_23[54] , \wNDiag_57[37] , 
        \wPDiag_43[2] , \wPDiag_15[51] , \wPDiag_15[48] , \wPDiag_36[60] , 
        \wPDiag_43[50] , \wNDiag_61[32] , \wScan_23[2] , \wNDiag_37[33] , 
        \wPDiag_43[49] , \wPDiag_60[61] , \wColumn_37[46] , \wColumn_61[47] , 
        \wColumn_57[42] , \wColumn_12[0] , \wScan_20[1] , \wPDiag_40[1] , 
        \wPDiag_1[30] , \wPDiag_1[29] , \wNDiag_7[59] , \wNDiag_7[40] , 
        \wColumn_9[37] , \wNDiag_14[31] , \wPDiag_36[53] , \wCall_41[0] , 
        \wScan_47[6] , \wNDiag_42[29] , \wPDiag_43[63] , \wNDiag_37[19] , 
        \wNDiag_14[28] , \wPDiag_27[6] , \wNDiag_42[30] , \wPDiag_60[52] , 
        \wNDiag_61[18] , \wPDiag_15[62] , \wNDiag_22[34] , \wPDiag_56[57] , 
        \wColumn_2[22] , \wColumn_5[2] , \wColumn_14[44] , \wColumn_22[58] , 
        \wColumn_22[41] , \wPDiag_24[5] , \wColumn_34[36] , \wColumn_42[45] , 
        \wScan_44[5] , \wScan_38[3] , \wColumn_62[37] , \wNDiag_49[25] , 
        \wColumn_54[32] , \wPDiag_58[3] , \wColumn_2[11] , \wColumn_6[1] , 
        \wNDiag_10[1] , \wNDiag_29[38] , \wNDiag_29[21] , \wNDiag_13[2] , 
        \wPDiag_16[21] , \wPDiag_20[24] , \wNDiag_34[43] , \wNDiag_54[47] , 
        \wPDiag_55[14] , \wPDiag_16[38] , \wPDiag_35[10] , \wPDiag_40[39] , 
        \wPDiag_63[11] , \wPDiag_28[41] , \wColumn_29[54] , \wPDiag_40[20] , 
        \wNDiag_62[42] , \wColumn_49[50] , \wColumn_49[49] , \wPDiag_2[59] , 
        \wPDiag_2[40] , \wNDiag_4[30] , \wColumn_17[34] , \wColumn_21[31] , 
        \wColumn_21[28] , \wPDiag_28[58] , \wNDiag_29[12] , \wPDiag_48[45] , 
        \wNDiag_49[16] , \wColumn_54[18] , \wPDiag_21[8] , \wColumn_41[35] , 
        \wColumn_49[63] , \wNDiag_4[29] , \wPDiag_16[12] , \wNDiag_17[58] , 
        \wNDiag_41[40] , \wPDiag_63[22] , \wNDiag_17[41] , \wPDiag_40[13] , 
        \wNDiag_41[59] , \wPDiag_20[17] , \wPDiag_35[23] , \wPDiag_55[27] , 
        \wNDiag_21[44] ;
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_12 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_13[6] , \wScan_13[5] , \wScan_13[4] , 
        \wScan_13[3] , \wScan_13[2] , \wScan_13[1] , \wScan_13[0] }), 
        .ScanOut({\wScan_12[6] , \wScan_12[5] , \wScan_12[4] , \wScan_12[3] , 
        \wScan_12[2] , \wScan_12[1] , \wScan_12[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_12[0] ), .ReturnIn(\wReturn_13[0] ), .ColIn({
        \wColumn_12[63] , \wColumn_12[62] , \wColumn_12[61] , \wColumn_12[60] , 
        \wColumn_12[59] , \wColumn_12[58] , \wColumn_12[57] , \wColumn_12[56] , 
        \wColumn_12[55] , \wColumn_12[54] , \wColumn_12[53] , \wColumn_12[52] , 
        \wColumn_12[51] , \wColumn_12[50] , \wColumn_12[49] , \wColumn_12[48] , 
        \wColumn_12[47] , \wColumn_12[46] , \wColumn_12[45] , \wColumn_12[44] , 
        \wColumn_12[43] , \wColumn_12[42] , \wColumn_12[41] , \wColumn_12[40] , 
        \wColumn_12[39] , \wColumn_12[38] , \wColumn_12[37] , \wColumn_12[36] , 
        \wColumn_12[35] , \wColumn_12[34] , \wColumn_12[33] , \wColumn_12[32] , 
        \wColumn_12[31] , \wColumn_12[30] , \wColumn_12[29] , \wColumn_12[28] , 
        \wColumn_12[27] , \wColumn_12[26] , \wColumn_12[25] , \wColumn_12[24] , 
        \wColumn_12[23] , \wColumn_12[22] , \wColumn_12[21] , \wColumn_12[20] , 
        \wColumn_12[19] , \wColumn_12[18] , \wColumn_12[17] , \wColumn_12[16] , 
        \wColumn_12[15] , \wColumn_12[14] , \wColumn_12[13] , \wColumn_12[12] , 
        \wColumn_12[11] , \wColumn_12[10] , \wColumn_12[9] , \wColumn_12[8] , 
        \wColumn_12[7] , \wColumn_12[6] , \wColumn_12[5] , \wColumn_12[4] , 
        \wColumn_12[3] , \wColumn_12[2] , \wColumn_12[1] , \wColumn_12[0] }), 
        .PDiagIn({\wPDiag_12[63] , \wPDiag_12[62] , \wPDiag_12[61] , 
        \wPDiag_12[60] , \wPDiag_12[59] , \wPDiag_12[58] , \wPDiag_12[57] , 
        \wPDiag_12[56] , \wPDiag_12[55] , \wPDiag_12[54] , \wPDiag_12[53] , 
        \wPDiag_12[52] , \wPDiag_12[51] , \wPDiag_12[50] , \wPDiag_12[49] , 
        \wPDiag_12[48] , \wPDiag_12[47] , \wPDiag_12[46] , \wPDiag_12[45] , 
        \wPDiag_12[44] , \wPDiag_12[43] , \wPDiag_12[42] , \wPDiag_12[41] , 
        \wPDiag_12[40] , \wPDiag_12[39] , \wPDiag_12[38] , \wPDiag_12[37] , 
        \wPDiag_12[36] , \wPDiag_12[35] , \wPDiag_12[34] , \wPDiag_12[33] , 
        \wPDiag_12[32] , \wPDiag_12[31] , \wPDiag_12[30] , \wPDiag_12[29] , 
        \wPDiag_12[28] , \wPDiag_12[27] , \wPDiag_12[26] , \wPDiag_12[25] , 
        \wPDiag_12[24] , \wPDiag_12[23] , \wPDiag_12[22] , \wPDiag_12[21] , 
        \wPDiag_12[20] , \wPDiag_12[19] , \wPDiag_12[18] , \wPDiag_12[17] , 
        \wPDiag_12[16] , \wPDiag_12[15] , \wPDiag_12[14] , \wPDiag_12[13] , 
        \wPDiag_12[12] , \wPDiag_12[11] , \wPDiag_12[10] , \wPDiag_12[9] , 
        \wPDiag_12[8] , \wPDiag_12[7] , \wPDiag_12[6] , \wPDiag_12[5] , 
        \wPDiag_12[4] , \wPDiag_12[3] , \wPDiag_12[2] , \wPDiag_12[1] , 
        \wPDiag_12[0] }), .NDiagIn({\wNDiag_12[63] , \wNDiag_12[62] , 
        \wNDiag_12[61] , \wNDiag_12[60] , \wNDiag_12[59] , \wNDiag_12[58] , 
        \wNDiag_12[57] , \wNDiag_12[56] , \wNDiag_12[55] , \wNDiag_12[54] , 
        \wNDiag_12[53] , \wNDiag_12[52] , \wNDiag_12[51] , \wNDiag_12[50] , 
        \wNDiag_12[49] , \wNDiag_12[48] , \wNDiag_12[47] , \wNDiag_12[46] , 
        \wNDiag_12[45] , \wNDiag_12[44] , \wNDiag_12[43] , \wNDiag_12[42] , 
        \wNDiag_12[41] , \wNDiag_12[40] , \wNDiag_12[39] , \wNDiag_12[38] , 
        \wNDiag_12[37] , \wNDiag_12[36] , \wNDiag_12[35] , \wNDiag_12[34] , 
        \wNDiag_12[33] , \wNDiag_12[32] , \wNDiag_12[31] , \wNDiag_12[30] , 
        \wNDiag_12[29] , \wNDiag_12[28] , \wNDiag_12[27] , \wNDiag_12[26] , 
        \wNDiag_12[25] , \wNDiag_12[24] , \wNDiag_12[23] , \wNDiag_12[22] , 
        \wNDiag_12[21] , \wNDiag_12[20] , \wNDiag_12[19] , \wNDiag_12[18] , 
        \wNDiag_12[17] , \wNDiag_12[16] , \wNDiag_12[15] , \wNDiag_12[14] , 
        \wNDiag_12[13] , \wNDiag_12[12] , \wNDiag_12[11] , \wNDiag_12[10] , 
        \wNDiag_12[9] , \wNDiag_12[8] , \wNDiag_12[7] , \wNDiag_12[6] , 
        \wNDiag_12[5] , \wNDiag_12[4] , \wNDiag_12[3] , \wNDiag_12[2] , 
        \wNDiag_12[1] , \wNDiag_12[0] }), .CallOut(\wCall_13[0] ), .ReturnOut(
        \wReturn_12[0] ), .ColOut({\wColumn_13[63] , \wColumn_13[62] , 
        \wColumn_13[61] , \wColumn_13[60] , \wColumn_13[59] , \wColumn_13[58] , 
        \wColumn_13[57] , \wColumn_13[56] , \wColumn_13[55] , \wColumn_13[54] , 
        \wColumn_13[53] , \wColumn_13[52] , \wColumn_13[51] , \wColumn_13[50] , 
        \wColumn_13[49] , \wColumn_13[48] , \wColumn_13[47] , \wColumn_13[46] , 
        \wColumn_13[45] , \wColumn_13[44] , \wColumn_13[43] , \wColumn_13[42] , 
        \wColumn_13[41] , \wColumn_13[40] , \wColumn_13[39] , \wColumn_13[38] , 
        \wColumn_13[37] , \wColumn_13[36] , \wColumn_13[35] , \wColumn_13[34] , 
        \wColumn_13[33] , \wColumn_13[32] , \wColumn_13[31] , \wColumn_13[30] , 
        \wColumn_13[29] , \wColumn_13[28] , \wColumn_13[27] , \wColumn_13[26] , 
        \wColumn_13[25] , \wColumn_13[24] , \wColumn_13[23] , \wColumn_13[22] , 
        \wColumn_13[21] , \wColumn_13[20] , \wColumn_13[19] , \wColumn_13[18] , 
        \wColumn_13[17] , \wColumn_13[16] , \wColumn_13[15] , \wColumn_13[14] , 
        \wColumn_13[13] , \wColumn_13[12] , \wColumn_13[11] , \wColumn_13[10] , 
        \wColumn_13[9] , \wColumn_13[8] , \wColumn_13[7] , \wColumn_13[6] , 
        \wColumn_13[5] , \wColumn_13[4] , \wColumn_13[3] , \wColumn_13[2] , 
        \wColumn_13[1] , \wColumn_13[0] }), .PDiagOut({\wPDiag_13[63] , 
        \wPDiag_13[62] , \wPDiag_13[61] , \wPDiag_13[60] , \wPDiag_13[59] , 
        \wPDiag_13[58] , \wPDiag_13[57] , \wPDiag_13[56] , \wPDiag_13[55] , 
        \wPDiag_13[54] , \wPDiag_13[53] , \wPDiag_13[52] , \wPDiag_13[51] , 
        \wPDiag_13[50] , \wPDiag_13[49] , \wPDiag_13[48] , \wPDiag_13[47] , 
        \wPDiag_13[46] , \wPDiag_13[45] , \wPDiag_13[44] , \wPDiag_13[43] , 
        \wPDiag_13[42] , \wPDiag_13[41] , \wPDiag_13[40] , \wPDiag_13[39] , 
        \wPDiag_13[38] , \wPDiag_13[37] , \wPDiag_13[36] , \wPDiag_13[35] , 
        \wPDiag_13[34] , \wPDiag_13[33] , \wPDiag_13[32] , \wPDiag_13[31] , 
        \wPDiag_13[30] , \wPDiag_13[29] , \wPDiag_13[28] , \wPDiag_13[27] , 
        \wPDiag_13[26] , \wPDiag_13[25] , \wPDiag_13[24] , \wPDiag_13[23] , 
        \wPDiag_13[22] , \wPDiag_13[21] , \wPDiag_13[20] , \wPDiag_13[19] , 
        \wPDiag_13[18] , \wPDiag_13[17] , \wPDiag_13[16] , \wPDiag_13[15] , 
        \wPDiag_13[14] , \wPDiag_13[13] , \wPDiag_13[12] , \wPDiag_13[11] , 
        \wPDiag_13[10] , \wPDiag_13[9] , \wPDiag_13[8] , \wPDiag_13[7] , 
        \wPDiag_13[6] , \wPDiag_13[5] , \wPDiag_13[4] , \wPDiag_13[3] , 
        \wPDiag_13[2] , \wPDiag_13[1] , \wPDiag_13[0] }), .NDiagOut({
        \wNDiag_13[63] , \wNDiag_13[62] , \wNDiag_13[61] , \wNDiag_13[60] , 
        \wNDiag_13[59] , \wNDiag_13[58] , \wNDiag_13[57] , \wNDiag_13[56] , 
        \wNDiag_13[55] , \wNDiag_13[54] , \wNDiag_13[53] , \wNDiag_13[52] , 
        \wNDiag_13[51] , \wNDiag_13[50] , \wNDiag_13[49] , \wNDiag_13[48] , 
        \wNDiag_13[47] , \wNDiag_13[46] , \wNDiag_13[45] , \wNDiag_13[44] , 
        \wNDiag_13[43] , \wNDiag_13[42] , \wNDiag_13[41] , \wNDiag_13[40] , 
        \wNDiag_13[39] , \wNDiag_13[38] , \wNDiag_13[37] , \wNDiag_13[36] , 
        \wNDiag_13[35] , \wNDiag_13[34] , \wNDiag_13[33] , \wNDiag_13[32] , 
        \wNDiag_13[31] , \wNDiag_13[30] , \wNDiag_13[29] , \wNDiag_13[28] , 
        \wNDiag_13[27] , \wNDiag_13[26] , \wNDiag_13[25] , \wNDiag_13[24] , 
        \wNDiag_13[23] , \wNDiag_13[22] , \wNDiag_13[21] , \wNDiag_13[20] , 
        \wNDiag_13[19] , \wNDiag_13[18] , \wNDiag_13[17] , \wNDiag_13[16] , 
        \wNDiag_13[15] , \wNDiag_13[14] , \wNDiag_13[13] , \wNDiag_13[12] , 
        \wNDiag_13[11] , \wNDiag_13[10] , \wNDiag_13[9] , \wNDiag_13[8] , 
        \wNDiag_13[7] , \wNDiag_13[6] , \wNDiag_13[5] , \wNDiag_13[4] , 
        \wNDiag_13[3] , \wNDiag_13[2] , \wNDiag_13[1] , \wNDiag_13[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_35 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_36[6] , \wScan_36[5] , \wScan_36[4] , 
        \wScan_36[3] , \wScan_36[2] , \wScan_36[1] , \wScan_36[0] }), 
        .ScanOut({\wScan_35[6] , \wScan_35[5] , \wScan_35[4] , \wScan_35[3] , 
        \wScan_35[2] , \wScan_35[1] , \wScan_35[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_35[0] ), .ReturnIn(\wReturn_36[0] ), .ColIn({
        \wColumn_35[63] , \wColumn_35[62] , \wColumn_35[61] , \wColumn_35[60] , 
        \wColumn_35[59] , \wColumn_35[58] , \wColumn_35[57] , \wColumn_35[56] , 
        \wColumn_35[55] , \wColumn_35[54] , \wColumn_35[53] , \wColumn_35[52] , 
        \wColumn_35[51] , \wColumn_35[50] , \wColumn_35[49] , \wColumn_35[48] , 
        \wColumn_35[47] , \wColumn_35[46] , \wColumn_35[45] , \wColumn_35[44] , 
        \wColumn_35[43] , \wColumn_35[42] , \wColumn_35[41] , \wColumn_35[40] , 
        \wColumn_35[39] , \wColumn_35[38] , \wColumn_35[37] , \wColumn_35[36] , 
        \wColumn_35[35] , \wColumn_35[34] , \wColumn_35[33] , \wColumn_35[32] , 
        \wColumn_35[31] , \wColumn_35[30] , \wColumn_35[29] , \wColumn_35[28] , 
        \wColumn_35[27] , \wColumn_35[26] , \wColumn_35[25] , \wColumn_35[24] , 
        \wColumn_35[23] , \wColumn_35[22] , \wColumn_35[21] , \wColumn_35[20] , 
        \wColumn_35[19] , \wColumn_35[18] , \wColumn_35[17] , \wColumn_35[16] , 
        \wColumn_35[15] , \wColumn_35[14] , \wColumn_35[13] , \wColumn_35[12] , 
        \wColumn_35[11] , \wColumn_35[10] , \wColumn_35[9] , \wColumn_35[8] , 
        \wColumn_35[7] , \wColumn_35[6] , \wColumn_35[5] , \wColumn_35[4] , 
        \wColumn_35[3] , \wColumn_35[2] , \wColumn_35[1] , \wColumn_35[0] }), 
        .PDiagIn({\wPDiag_35[63] , \wPDiag_35[62] , \wPDiag_35[61] , 
        \wPDiag_35[60] , \wPDiag_35[59] , \wPDiag_35[58] , \wPDiag_35[57] , 
        \wPDiag_35[56] , \wPDiag_35[55] , \wPDiag_35[54] , \wPDiag_35[53] , 
        \wPDiag_35[52] , \wPDiag_35[51] , \wPDiag_35[50] , \wPDiag_35[49] , 
        \wPDiag_35[48] , \wPDiag_35[47] , \wPDiag_35[46] , \wPDiag_35[45] , 
        \wPDiag_35[44] , \wPDiag_35[43] , \wPDiag_35[42] , \wPDiag_35[41] , 
        \wPDiag_35[40] , \wPDiag_35[39] , \wPDiag_35[38] , \wPDiag_35[37] , 
        \wPDiag_35[36] , \wPDiag_35[35] , \wPDiag_35[34] , \wPDiag_35[33] , 
        \wPDiag_35[32] , \wPDiag_35[31] , \wPDiag_35[30] , \wPDiag_35[29] , 
        \wPDiag_35[28] , \wPDiag_35[27] , \wPDiag_35[26] , \wPDiag_35[25] , 
        \wPDiag_35[24] , \wPDiag_35[23] , \wPDiag_35[22] , \wPDiag_35[21] , 
        \wPDiag_35[20] , \wPDiag_35[19] , \wPDiag_35[18] , \wPDiag_35[17] , 
        \wPDiag_35[16] , \wPDiag_35[15] , \wPDiag_35[14] , \wPDiag_35[13] , 
        \wPDiag_35[12] , \wPDiag_35[11] , \wPDiag_35[10] , \wPDiag_35[9] , 
        \wPDiag_35[8] , \wPDiag_35[7] , \wPDiag_35[6] , \wPDiag_35[5] , 
        \wPDiag_35[4] , \wPDiag_35[3] , \wPDiag_35[2] , \wPDiag_35[1] , 
        \wPDiag_35[0] }), .NDiagIn({\wNDiag_35[63] , \wNDiag_35[62] , 
        \wNDiag_35[61] , \wNDiag_35[60] , \wNDiag_35[59] , \wNDiag_35[58] , 
        \wNDiag_35[57] , \wNDiag_35[56] , \wNDiag_35[55] , \wNDiag_35[54] , 
        \wNDiag_35[53] , \wNDiag_35[52] , \wNDiag_35[51] , \wNDiag_35[50] , 
        \wNDiag_35[49] , \wNDiag_35[48] , \wNDiag_35[47] , \wNDiag_35[46] , 
        \wNDiag_35[45] , \wNDiag_35[44] , \wNDiag_35[43] , \wNDiag_35[42] , 
        \wNDiag_35[41] , \wNDiag_35[40] , \wNDiag_35[39] , \wNDiag_35[38] , 
        \wNDiag_35[37] , \wNDiag_35[36] , \wNDiag_35[35] , \wNDiag_35[34] , 
        \wNDiag_35[33] , \wNDiag_35[32] , \wNDiag_35[31] , \wNDiag_35[30] , 
        \wNDiag_35[29] , \wNDiag_35[28] , \wNDiag_35[27] , \wNDiag_35[26] , 
        \wNDiag_35[25] , \wNDiag_35[24] , \wNDiag_35[23] , \wNDiag_35[22] , 
        \wNDiag_35[21] , \wNDiag_35[20] , \wNDiag_35[19] , \wNDiag_35[18] , 
        \wNDiag_35[17] , \wNDiag_35[16] , \wNDiag_35[15] , \wNDiag_35[14] , 
        \wNDiag_35[13] , \wNDiag_35[12] , \wNDiag_35[11] , \wNDiag_35[10] , 
        \wNDiag_35[9] , \wNDiag_35[8] , \wNDiag_35[7] , \wNDiag_35[6] , 
        \wNDiag_35[5] , \wNDiag_35[4] , \wNDiag_35[3] , \wNDiag_35[2] , 
        \wNDiag_35[1] , \wNDiag_35[0] }), .CallOut(\wCall_36[0] ), .ReturnOut(
        \wReturn_35[0] ), .ColOut({\wColumn_36[63] , \wColumn_36[62] , 
        \wColumn_36[61] , \wColumn_36[60] , \wColumn_36[59] , \wColumn_36[58] , 
        \wColumn_36[57] , \wColumn_36[56] , \wColumn_36[55] , \wColumn_36[54] , 
        \wColumn_36[53] , \wColumn_36[52] , \wColumn_36[51] , \wColumn_36[50] , 
        \wColumn_36[49] , \wColumn_36[48] , \wColumn_36[47] , \wColumn_36[46] , 
        \wColumn_36[45] , \wColumn_36[44] , \wColumn_36[43] , \wColumn_36[42] , 
        \wColumn_36[41] , \wColumn_36[40] , \wColumn_36[39] , \wColumn_36[38] , 
        \wColumn_36[37] , \wColumn_36[36] , \wColumn_36[35] , \wColumn_36[34] , 
        \wColumn_36[33] , \wColumn_36[32] , \wColumn_36[31] , \wColumn_36[30] , 
        \wColumn_36[29] , \wColumn_36[28] , \wColumn_36[27] , \wColumn_36[26] , 
        \wColumn_36[25] , \wColumn_36[24] , \wColumn_36[23] , \wColumn_36[22] , 
        \wColumn_36[21] , \wColumn_36[20] , \wColumn_36[19] , \wColumn_36[18] , 
        \wColumn_36[17] , \wColumn_36[16] , \wColumn_36[15] , \wColumn_36[14] , 
        \wColumn_36[13] , \wColumn_36[12] , \wColumn_36[11] , \wColumn_36[10] , 
        \wColumn_36[9] , \wColumn_36[8] , \wColumn_36[7] , \wColumn_36[6] , 
        \wColumn_36[5] , \wColumn_36[4] , \wColumn_36[3] , \wColumn_36[2] , 
        \wColumn_36[1] , \wColumn_36[0] }), .PDiagOut({\wPDiag_36[63] , 
        \wPDiag_36[62] , \wPDiag_36[61] , \wPDiag_36[60] , \wPDiag_36[59] , 
        \wPDiag_36[58] , \wPDiag_36[57] , \wPDiag_36[56] , \wPDiag_36[55] , 
        \wPDiag_36[54] , \wPDiag_36[53] , \wPDiag_36[52] , \wPDiag_36[51] , 
        \wPDiag_36[50] , \wPDiag_36[49] , \wPDiag_36[48] , \wPDiag_36[47] , 
        \wPDiag_36[46] , \wPDiag_36[45] , \wPDiag_36[44] , \wPDiag_36[43] , 
        \wPDiag_36[42] , \wPDiag_36[41] , \wPDiag_36[40] , \wPDiag_36[39] , 
        \wPDiag_36[38] , \wPDiag_36[37] , \wPDiag_36[36] , \wPDiag_36[35] , 
        \wPDiag_36[34] , \wPDiag_36[33] , \wPDiag_36[32] , \wPDiag_36[31] , 
        \wPDiag_36[30] , \wPDiag_36[29] , \wPDiag_36[28] , \wPDiag_36[27] , 
        \wPDiag_36[26] , \wPDiag_36[25] , \wPDiag_36[24] , \wPDiag_36[23] , 
        \wPDiag_36[22] , \wPDiag_36[21] , \wPDiag_36[20] , \wPDiag_36[19] , 
        \wPDiag_36[18] , \wPDiag_36[17] , \wPDiag_36[16] , \wPDiag_36[15] , 
        \wPDiag_36[14] , \wPDiag_36[13] , \wPDiag_36[12] , \wPDiag_36[11] , 
        \wPDiag_36[10] , \wPDiag_36[9] , \wPDiag_36[8] , \wPDiag_36[7] , 
        \wPDiag_36[6] , \wPDiag_36[5] , \wPDiag_36[4] , \wPDiag_36[3] , 
        \wPDiag_36[2] , \wPDiag_36[1] , \wPDiag_36[0] }), .NDiagOut({
        \wNDiag_36[63] , \wNDiag_36[62] , \wNDiag_36[61] , \wNDiag_36[60] , 
        \wNDiag_36[59] , \wNDiag_36[58] , \wNDiag_36[57] , \wNDiag_36[56] , 
        \wNDiag_36[55] , \wNDiag_36[54] , \wNDiag_36[53] , \wNDiag_36[52] , 
        \wNDiag_36[51] , \wNDiag_36[50] , \wNDiag_36[49] , \wNDiag_36[48] , 
        \wNDiag_36[47] , \wNDiag_36[46] , \wNDiag_36[45] , \wNDiag_36[44] , 
        \wNDiag_36[43] , \wNDiag_36[42] , \wNDiag_36[41] , \wNDiag_36[40] , 
        \wNDiag_36[39] , \wNDiag_36[38] , \wNDiag_36[37] , \wNDiag_36[36] , 
        \wNDiag_36[35] , \wNDiag_36[34] , \wNDiag_36[33] , \wNDiag_36[32] , 
        \wNDiag_36[31] , \wNDiag_36[30] , \wNDiag_36[29] , \wNDiag_36[28] , 
        \wNDiag_36[27] , \wNDiag_36[26] , \wNDiag_36[25] , \wNDiag_36[24] , 
        \wNDiag_36[23] , \wNDiag_36[22] , \wNDiag_36[21] , \wNDiag_36[20] , 
        \wNDiag_36[19] , \wNDiag_36[18] , \wNDiag_36[17] , \wNDiag_36[16] , 
        \wNDiag_36[15] , \wNDiag_36[14] , \wNDiag_36[13] , \wNDiag_36[12] , 
        \wNDiag_36[11] , \wNDiag_36[10] , \wNDiag_36[9] , \wNDiag_36[8] , 
        \wNDiag_36[7] , \wNDiag_36[6] , \wNDiag_36[5] , \wNDiag_36[4] , 
        \wNDiag_36[3] , \wNDiag_36[2] , \wNDiag_36[1] , \wNDiag_36[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_40 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_41[6] , \wScan_41[5] , \wScan_41[4] , 
        \wScan_41[3] , \wScan_41[2] , \wScan_41[1] , \wScan_41[0] }), 
        .ScanOut({\wScan_40[6] , \wScan_40[5] , \wScan_40[4] , \wScan_40[3] , 
        \wScan_40[2] , \wScan_40[1] , \wScan_40[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_40[0] ), .ReturnIn(\wReturn_41[0] ), .ColIn({
        \wColumn_40[63] , \wColumn_40[62] , \wColumn_40[61] , \wColumn_40[60] , 
        \wColumn_40[59] , \wColumn_40[58] , \wColumn_40[57] , \wColumn_40[56] , 
        \wColumn_40[55] , \wColumn_40[54] , \wColumn_40[53] , \wColumn_40[52] , 
        \wColumn_40[51] , \wColumn_40[50] , \wColumn_40[49] , \wColumn_40[48] , 
        \wColumn_40[47] , \wColumn_40[46] , \wColumn_40[45] , \wColumn_40[44] , 
        \wColumn_40[43] , \wColumn_40[42] , \wColumn_40[41] , \wColumn_40[40] , 
        \wColumn_40[39] , \wColumn_40[38] , \wColumn_40[37] , \wColumn_40[36] , 
        \wColumn_40[35] , \wColumn_40[34] , \wColumn_40[33] , \wColumn_40[32] , 
        \wColumn_40[31] , \wColumn_40[30] , \wColumn_40[29] , \wColumn_40[28] , 
        \wColumn_40[27] , \wColumn_40[26] , \wColumn_40[25] , \wColumn_40[24] , 
        \wColumn_40[23] , \wColumn_40[22] , \wColumn_40[21] , \wColumn_40[20] , 
        \wColumn_40[19] , \wColumn_40[18] , \wColumn_40[17] , \wColumn_40[16] , 
        \wColumn_40[15] , \wColumn_40[14] , \wColumn_40[13] , \wColumn_40[12] , 
        \wColumn_40[11] , \wColumn_40[10] , \wColumn_40[9] , \wColumn_40[8] , 
        \wColumn_40[7] , \wColumn_40[6] , \wColumn_40[5] , \wColumn_40[4] , 
        \wColumn_40[3] , \wColumn_40[2] , \wColumn_40[1] , \wColumn_40[0] }), 
        .PDiagIn({\wPDiag_40[63] , \wPDiag_40[62] , \wPDiag_40[61] , 
        \wPDiag_40[60] , \wPDiag_40[59] , \wPDiag_40[58] , \wPDiag_40[57] , 
        \wPDiag_40[56] , \wPDiag_40[55] , \wPDiag_40[54] , \wPDiag_40[53] , 
        \wPDiag_40[52] , \wPDiag_40[51] , \wPDiag_40[50] , \wPDiag_40[49] , 
        \wPDiag_40[48] , \wPDiag_40[47] , \wPDiag_40[46] , \wPDiag_40[45] , 
        \wPDiag_40[44] , \wPDiag_40[43] , \wPDiag_40[42] , \wPDiag_40[41] , 
        \wPDiag_40[40] , \wPDiag_40[39] , \wPDiag_40[38] , \wPDiag_40[37] , 
        \wPDiag_40[36] , \wPDiag_40[35] , \wPDiag_40[34] , \wPDiag_40[33] , 
        \wPDiag_40[32] , \wPDiag_40[31] , \wPDiag_40[30] , \wPDiag_40[29] , 
        \wPDiag_40[28] , \wPDiag_40[27] , \wPDiag_40[26] , \wPDiag_40[25] , 
        \wPDiag_40[24] , \wPDiag_40[23] , \wPDiag_40[22] , \wPDiag_40[21] , 
        \wPDiag_40[20] , \wPDiag_40[19] , \wPDiag_40[18] , \wPDiag_40[17] , 
        \wPDiag_40[16] , \wPDiag_40[15] , \wPDiag_40[14] , \wPDiag_40[13] , 
        \wPDiag_40[12] , \wPDiag_40[11] , \wPDiag_40[10] , \wPDiag_40[9] , 
        \wPDiag_40[8] , \wPDiag_40[7] , \wPDiag_40[6] , \wPDiag_40[5] , 
        \wPDiag_40[4] , \wPDiag_40[3] , \wPDiag_40[2] , \wPDiag_40[1] , 
        \wPDiag_40[0] }), .NDiagIn({\wNDiag_40[63] , \wNDiag_40[62] , 
        \wNDiag_40[61] , \wNDiag_40[60] , \wNDiag_40[59] , \wNDiag_40[58] , 
        \wNDiag_40[57] , \wNDiag_40[56] , \wNDiag_40[55] , \wNDiag_40[54] , 
        \wNDiag_40[53] , \wNDiag_40[52] , \wNDiag_40[51] , \wNDiag_40[50] , 
        \wNDiag_40[49] , \wNDiag_40[48] , \wNDiag_40[47] , \wNDiag_40[46] , 
        \wNDiag_40[45] , \wNDiag_40[44] , \wNDiag_40[43] , \wNDiag_40[42] , 
        \wNDiag_40[41] , \wNDiag_40[40] , \wNDiag_40[39] , \wNDiag_40[38] , 
        \wNDiag_40[37] , \wNDiag_40[36] , \wNDiag_40[35] , \wNDiag_40[34] , 
        \wNDiag_40[33] , \wNDiag_40[32] , \wNDiag_40[31] , \wNDiag_40[30] , 
        \wNDiag_40[29] , \wNDiag_40[28] , \wNDiag_40[27] , \wNDiag_40[26] , 
        \wNDiag_40[25] , \wNDiag_40[24] , \wNDiag_40[23] , \wNDiag_40[22] , 
        \wNDiag_40[21] , \wNDiag_40[20] , \wNDiag_40[19] , \wNDiag_40[18] , 
        \wNDiag_40[17] , \wNDiag_40[16] , \wNDiag_40[15] , \wNDiag_40[14] , 
        \wNDiag_40[13] , \wNDiag_40[12] , \wNDiag_40[11] , \wNDiag_40[10] , 
        \wNDiag_40[9] , \wNDiag_40[8] , \wNDiag_40[7] , \wNDiag_40[6] , 
        \wNDiag_40[5] , \wNDiag_40[4] , \wNDiag_40[3] , \wNDiag_40[2] , 
        \wNDiag_40[1] , \wNDiag_40[0] }), .CallOut(\wCall_41[0] ), .ReturnOut(
        \wReturn_40[0] ), .ColOut({\wColumn_41[63] , \wColumn_41[62] , 
        \wColumn_41[61] , \wColumn_41[60] , \wColumn_41[59] , \wColumn_41[58] , 
        \wColumn_41[57] , \wColumn_41[56] , \wColumn_41[55] , \wColumn_41[54] , 
        \wColumn_41[53] , \wColumn_41[52] , \wColumn_41[51] , \wColumn_41[50] , 
        \wColumn_41[49] , \wColumn_41[48] , \wColumn_41[47] , \wColumn_41[46] , 
        \wColumn_41[45] , \wColumn_41[44] , \wColumn_41[43] , \wColumn_41[42] , 
        \wColumn_41[41] , \wColumn_41[40] , \wColumn_41[39] , \wColumn_41[38] , 
        \wColumn_41[37] , \wColumn_41[36] , \wColumn_41[35] , \wColumn_41[34] , 
        \wColumn_41[33] , \wColumn_41[32] , \wColumn_41[31] , \wColumn_41[30] , 
        \wColumn_41[29] , \wColumn_41[28] , \wColumn_41[27] , \wColumn_41[26] , 
        \wColumn_41[25] , \wColumn_41[24] , \wColumn_41[23] , \wColumn_41[22] , 
        \wColumn_41[21] , \wColumn_41[20] , \wColumn_41[19] , \wColumn_41[18] , 
        \wColumn_41[17] , \wColumn_41[16] , \wColumn_41[15] , \wColumn_41[14] , 
        \wColumn_41[13] , \wColumn_41[12] , \wColumn_41[11] , \wColumn_41[10] , 
        \wColumn_41[9] , \wColumn_41[8] , \wColumn_41[7] , \wColumn_41[6] , 
        \wColumn_41[5] , \wColumn_41[4] , \wColumn_41[3] , \wColumn_41[2] , 
        \wColumn_41[1] , \wColumn_41[0] }), .PDiagOut({\wPDiag_41[63] , 
        \wPDiag_41[62] , \wPDiag_41[61] , \wPDiag_41[60] , \wPDiag_41[59] , 
        \wPDiag_41[58] , \wPDiag_41[57] , \wPDiag_41[56] , \wPDiag_41[55] , 
        \wPDiag_41[54] , \wPDiag_41[53] , \wPDiag_41[52] , \wPDiag_41[51] , 
        \wPDiag_41[50] , \wPDiag_41[49] , \wPDiag_41[48] , \wPDiag_41[47] , 
        \wPDiag_41[46] , \wPDiag_41[45] , \wPDiag_41[44] , \wPDiag_41[43] , 
        \wPDiag_41[42] , \wPDiag_41[41] , \wPDiag_41[40] , \wPDiag_41[39] , 
        \wPDiag_41[38] , \wPDiag_41[37] , \wPDiag_41[36] , \wPDiag_41[35] , 
        \wPDiag_41[34] , \wPDiag_41[33] , \wPDiag_41[32] , \wPDiag_41[31] , 
        \wPDiag_41[30] , \wPDiag_41[29] , \wPDiag_41[28] , \wPDiag_41[27] , 
        \wPDiag_41[26] , \wPDiag_41[25] , \wPDiag_41[24] , \wPDiag_41[23] , 
        \wPDiag_41[22] , \wPDiag_41[21] , \wPDiag_41[20] , \wPDiag_41[19] , 
        \wPDiag_41[18] , \wPDiag_41[17] , \wPDiag_41[16] , \wPDiag_41[15] , 
        \wPDiag_41[14] , \wPDiag_41[13] , \wPDiag_41[12] , \wPDiag_41[11] , 
        \wPDiag_41[10] , \wPDiag_41[9] , \wPDiag_41[8] , \wPDiag_41[7] , 
        \wPDiag_41[6] , \wPDiag_41[5] , \wPDiag_41[4] , \wPDiag_41[3] , 
        \wPDiag_41[2] , \wPDiag_41[1] , \wPDiag_41[0] }), .NDiagOut({
        \wNDiag_41[63] , \wNDiag_41[62] , \wNDiag_41[61] , \wNDiag_41[60] , 
        \wNDiag_41[59] , \wNDiag_41[58] , \wNDiag_41[57] , \wNDiag_41[56] , 
        \wNDiag_41[55] , \wNDiag_41[54] , \wNDiag_41[53] , \wNDiag_41[52] , 
        \wNDiag_41[51] , \wNDiag_41[50] , \wNDiag_41[49] , \wNDiag_41[48] , 
        \wNDiag_41[47] , \wNDiag_41[46] , \wNDiag_41[45] , \wNDiag_41[44] , 
        \wNDiag_41[43] , \wNDiag_41[42] , \wNDiag_41[41] , \wNDiag_41[40] , 
        \wNDiag_41[39] , \wNDiag_41[38] , \wNDiag_41[37] , \wNDiag_41[36] , 
        \wNDiag_41[35] , \wNDiag_41[34] , \wNDiag_41[33] , \wNDiag_41[32] , 
        \wNDiag_41[31] , \wNDiag_41[30] , \wNDiag_41[29] , \wNDiag_41[28] , 
        \wNDiag_41[27] , \wNDiag_41[26] , \wNDiag_41[25] , \wNDiag_41[24] , 
        \wNDiag_41[23] , \wNDiag_41[22] , \wNDiag_41[21] , \wNDiag_41[20] , 
        \wNDiag_41[19] , \wNDiag_41[18] , \wNDiag_41[17] , \wNDiag_41[16] , 
        \wNDiag_41[15] , \wNDiag_41[14] , \wNDiag_41[13] , \wNDiag_41[12] , 
        \wNDiag_41[11] , \wNDiag_41[10] , \wNDiag_41[9] , \wNDiag_41[8] , 
        \wNDiag_41[7] , \wNDiag_41[6] , \wNDiag_41[5] , \wNDiag_41[4] , 
        \wNDiag_41[3] , \wNDiag_41[2] , \wNDiag_41[1] , \wNDiag_41[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_0 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_1[6] , \wScan_1[5] , \wScan_1[4] , 
        \wScan_1[3] , \wScan_1[2] , \wScan_1[1] , \wScan_1[0] }), .ScanOut({
        \wScan_0[6] , \wScan_0[5] , \wScan_0[4] , \wScan_0[3] , \wScan_0[2] , 
        \wScan_0[1] , \wScan_0[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_0[0] ), 
        .ReturnIn(\wReturn_1[0] ), .ColIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .PDiagIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .NDiagIn({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallOut(\wCall_1[0] ), .ReturnOut(\wReturn_0[0] ), .ColOut({
        \wColumn_1[63] , \wColumn_1[62] , \wColumn_1[61] , \wColumn_1[60] , 
        \wColumn_1[59] , \wColumn_1[58] , \wColumn_1[57] , \wColumn_1[56] , 
        \wColumn_1[55] , \wColumn_1[54] , \wColumn_1[53] , \wColumn_1[52] , 
        \wColumn_1[51] , \wColumn_1[50] , \wColumn_1[49] , \wColumn_1[48] , 
        \wColumn_1[47] , \wColumn_1[46] , \wColumn_1[45] , \wColumn_1[44] , 
        \wColumn_1[43] , \wColumn_1[42] , \wColumn_1[41] , \wColumn_1[40] , 
        \wColumn_1[39] , \wColumn_1[38] , \wColumn_1[37] , \wColumn_1[36] , 
        \wColumn_1[35] , \wColumn_1[34] , \wColumn_1[33] , \wColumn_1[32] , 
        \wColumn_1[31] , \wColumn_1[30] , \wColumn_1[29] , \wColumn_1[28] , 
        \wColumn_1[27] , \wColumn_1[26] , \wColumn_1[25] , \wColumn_1[24] , 
        \wColumn_1[23] , \wColumn_1[22] , \wColumn_1[21] , \wColumn_1[20] , 
        \wColumn_1[19] , \wColumn_1[18] , \wColumn_1[17] , \wColumn_1[16] , 
        \wColumn_1[15] , \wColumn_1[14] , \wColumn_1[13] , \wColumn_1[12] , 
        \wColumn_1[11] , \wColumn_1[10] , \wColumn_1[9] , \wColumn_1[8] , 
        \wColumn_1[7] , \wColumn_1[6] , \wColumn_1[5] , \wColumn_1[4] , 
        \wColumn_1[3] , \wColumn_1[2] , \wColumn_1[1] , \wColumn_1[0] }), 
        .PDiagOut({\wPDiag_1[63] , \wPDiag_1[62] , \wPDiag_1[61] , 
        \wPDiag_1[60] , \wPDiag_1[59] , \wPDiag_1[58] , \wPDiag_1[57] , 
        \wPDiag_1[56] , \wPDiag_1[55] , \wPDiag_1[54] , \wPDiag_1[53] , 
        \wPDiag_1[52] , \wPDiag_1[51] , \wPDiag_1[50] , \wPDiag_1[49] , 
        \wPDiag_1[48] , \wPDiag_1[47] , \wPDiag_1[46] , \wPDiag_1[45] , 
        \wPDiag_1[44] , \wPDiag_1[43] , \wPDiag_1[42] , \wPDiag_1[41] , 
        \wPDiag_1[40] , \wPDiag_1[39] , \wPDiag_1[38] , \wPDiag_1[37] , 
        \wPDiag_1[36] , \wPDiag_1[35] , \wPDiag_1[34] , \wPDiag_1[33] , 
        \wPDiag_1[32] , \wPDiag_1[31] , \wPDiag_1[30] , \wPDiag_1[29] , 
        \wPDiag_1[28] , \wPDiag_1[27] , \wPDiag_1[26] , \wPDiag_1[25] , 
        \wPDiag_1[24] , \wPDiag_1[23] , \wPDiag_1[22] , \wPDiag_1[21] , 
        \wPDiag_1[20] , \wPDiag_1[19] , \wPDiag_1[18] , \wPDiag_1[17] , 
        \wPDiag_1[16] , \wPDiag_1[15] , \wPDiag_1[14] , \wPDiag_1[13] , 
        \wPDiag_1[12] , \wPDiag_1[11] , \wPDiag_1[10] , \wPDiag_1[9] , 
        \wPDiag_1[8] , \wPDiag_1[7] , \wPDiag_1[6] , \wPDiag_1[5] , 
        \wPDiag_1[4] , \wPDiag_1[3] , \wPDiag_1[2] , \wPDiag_1[1] , 
        \wPDiag_1[0] }), .NDiagOut({\wNDiag_1[63] , \wNDiag_1[62] , 
        \wNDiag_1[61] , \wNDiag_1[60] , \wNDiag_1[59] , \wNDiag_1[58] , 
        \wNDiag_1[57] , \wNDiag_1[56] , \wNDiag_1[55] , \wNDiag_1[54] , 
        \wNDiag_1[53] , \wNDiag_1[52] , \wNDiag_1[51] , \wNDiag_1[50] , 
        \wNDiag_1[49] , \wNDiag_1[48] , \wNDiag_1[47] , \wNDiag_1[46] , 
        \wNDiag_1[45] , \wNDiag_1[44] , \wNDiag_1[43] , \wNDiag_1[42] , 
        \wNDiag_1[41] , \wNDiag_1[40] , \wNDiag_1[39] , \wNDiag_1[38] , 
        \wNDiag_1[37] , \wNDiag_1[36] , \wNDiag_1[35] , \wNDiag_1[34] , 
        \wNDiag_1[33] , \wNDiag_1[32] , \wNDiag_1[31] , \wNDiag_1[30] , 
        \wNDiag_1[29] , \wNDiag_1[28] , \wNDiag_1[27] , \wNDiag_1[26] , 
        \wNDiag_1[25] , \wNDiag_1[24] , \wNDiag_1[23] , \wNDiag_1[22] , 
        \wNDiag_1[21] , \wNDiag_1[20] , \wNDiag_1[19] , \wNDiag_1[18] , 
        \wNDiag_1[17] , \wNDiag_1[16] , \wNDiag_1[15] , \wNDiag_1[14] , 
        \wNDiag_1[13] , \wNDiag_1[12] , \wNDiag_1[11] , \wNDiag_1[10] , 
        \wNDiag_1[9] , \wNDiag_1[8] , \wNDiag_1[7] , \wNDiag_1[6] , 
        \wNDiag_1[5] , \wNDiag_1[4] , \wNDiag_1[3] , \wNDiag_1[2] , 
        \wNDiag_1[1] , \wNDiag_1[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_2 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_3[6] , \wScan_3[5] , \wScan_3[4] , 
        \wScan_3[3] , \wScan_3[2] , \wScan_3[1] , \wScan_3[0] }), .ScanOut({
        \wScan_2[6] , \wScan_2[5] , \wScan_2[4] , \wScan_2[3] , \wScan_2[2] , 
        \wScan_2[1] , \wScan_2[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_2[0] ), 
        .ReturnIn(\wReturn_3[0] ), .ColIn({\wColumn_2[63] , \wColumn_2[62] , 
        \wColumn_2[61] , \wColumn_2[60] , \wColumn_2[59] , \wColumn_2[58] , 
        \wColumn_2[57] , \wColumn_2[56] , \wColumn_2[55] , \wColumn_2[54] , 
        \wColumn_2[53] , \wColumn_2[52] , \wColumn_2[51] , \wColumn_2[50] , 
        \wColumn_2[49] , \wColumn_2[48] , \wColumn_2[47] , \wColumn_2[46] , 
        \wColumn_2[45] , \wColumn_2[44] , \wColumn_2[43] , \wColumn_2[42] , 
        \wColumn_2[41] , \wColumn_2[40] , \wColumn_2[39] , \wColumn_2[38] , 
        \wColumn_2[37] , \wColumn_2[36] , \wColumn_2[35] , \wColumn_2[34] , 
        \wColumn_2[33] , \wColumn_2[32] , \wColumn_2[31] , \wColumn_2[30] , 
        \wColumn_2[29] , \wColumn_2[28] , \wColumn_2[27] , \wColumn_2[26] , 
        \wColumn_2[25] , \wColumn_2[24] , \wColumn_2[23] , \wColumn_2[22] , 
        \wColumn_2[21] , \wColumn_2[20] , \wColumn_2[19] , \wColumn_2[18] , 
        \wColumn_2[17] , \wColumn_2[16] , \wColumn_2[15] , \wColumn_2[14] , 
        \wColumn_2[13] , \wColumn_2[12] , \wColumn_2[11] , \wColumn_2[10] , 
        \wColumn_2[9] , \wColumn_2[8] , \wColumn_2[7] , \wColumn_2[6] , 
        \wColumn_2[5] , \wColumn_2[4] , \wColumn_2[3] , \wColumn_2[2] , 
        \wColumn_2[1] , \wColumn_2[0] }), .PDiagIn({\wPDiag_2[63] , 
        \wPDiag_2[62] , \wPDiag_2[61] , \wPDiag_2[60] , \wPDiag_2[59] , 
        \wPDiag_2[58] , \wPDiag_2[57] , \wPDiag_2[56] , \wPDiag_2[55] , 
        \wPDiag_2[54] , \wPDiag_2[53] , \wPDiag_2[52] , \wPDiag_2[51] , 
        \wPDiag_2[50] , \wPDiag_2[49] , \wPDiag_2[48] , \wPDiag_2[47] , 
        \wPDiag_2[46] , \wPDiag_2[45] , \wPDiag_2[44] , \wPDiag_2[43] , 
        \wPDiag_2[42] , \wPDiag_2[41] , \wPDiag_2[40] , \wPDiag_2[39] , 
        \wPDiag_2[38] , \wPDiag_2[37] , \wPDiag_2[36] , \wPDiag_2[35] , 
        \wPDiag_2[34] , \wPDiag_2[33] , \wPDiag_2[32] , \wPDiag_2[31] , 
        \wPDiag_2[30] , \wPDiag_2[29] , \wPDiag_2[28] , \wPDiag_2[27] , 
        \wPDiag_2[26] , \wPDiag_2[25] , \wPDiag_2[24] , \wPDiag_2[23] , 
        \wPDiag_2[22] , \wPDiag_2[21] , \wPDiag_2[20] , \wPDiag_2[19] , 
        \wPDiag_2[18] , \wPDiag_2[17] , \wPDiag_2[16] , \wPDiag_2[15] , 
        \wPDiag_2[14] , \wPDiag_2[13] , \wPDiag_2[12] , \wPDiag_2[11] , 
        \wPDiag_2[10] , \wPDiag_2[9] , \wPDiag_2[8] , \wPDiag_2[7] , 
        \wPDiag_2[6] , \wPDiag_2[5] , \wPDiag_2[4] , \wPDiag_2[3] , 
        \wPDiag_2[2] , \wPDiag_2[1] , \wPDiag_2[0] }), .NDiagIn({
        \wNDiag_2[63] , \wNDiag_2[62] , \wNDiag_2[61] , \wNDiag_2[60] , 
        \wNDiag_2[59] , \wNDiag_2[58] , \wNDiag_2[57] , \wNDiag_2[56] , 
        \wNDiag_2[55] , \wNDiag_2[54] , \wNDiag_2[53] , \wNDiag_2[52] , 
        \wNDiag_2[51] , \wNDiag_2[50] , \wNDiag_2[49] , \wNDiag_2[48] , 
        \wNDiag_2[47] , \wNDiag_2[46] , \wNDiag_2[45] , \wNDiag_2[44] , 
        \wNDiag_2[43] , \wNDiag_2[42] , \wNDiag_2[41] , \wNDiag_2[40] , 
        \wNDiag_2[39] , \wNDiag_2[38] , \wNDiag_2[37] , \wNDiag_2[36] , 
        \wNDiag_2[35] , \wNDiag_2[34] , \wNDiag_2[33] , \wNDiag_2[32] , 
        \wNDiag_2[31] , \wNDiag_2[30] , \wNDiag_2[29] , \wNDiag_2[28] , 
        \wNDiag_2[27] , \wNDiag_2[26] , \wNDiag_2[25] , \wNDiag_2[24] , 
        \wNDiag_2[23] , \wNDiag_2[22] , \wNDiag_2[21] , \wNDiag_2[20] , 
        \wNDiag_2[19] , \wNDiag_2[18] , \wNDiag_2[17] , \wNDiag_2[16] , 
        \wNDiag_2[15] , \wNDiag_2[14] , \wNDiag_2[13] , \wNDiag_2[12] , 
        \wNDiag_2[11] , \wNDiag_2[10] , \wNDiag_2[9] , \wNDiag_2[8] , 
        \wNDiag_2[7] , \wNDiag_2[6] , \wNDiag_2[5] , \wNDiag_2[4] , 
        \wNDiag_2[3] , \wNDiag_2[2] , \wNDiag_2[1] , \wNDiag_2[0] }), 
        .CallOut(\wCall_3[0] ), .ReturnOut(\wReturn_2[0] ), .ColOut({
        \wColumn_3[63] , \wColumn_3[62] , \wColumn_3[61] , \wColumn_3[60] , 
        \wColumn_3[59] , \wColumn_3[58] , \wColumn_3[57] , \wColumn_3[56] , 
        \wColumn_3[55] , \wColumn_3[54] , \wColumn_3[53] , \wColumn_3[52] , 
        \wColumn_3[51] , \wColumn_3[50] , \wColumn_3[49] , \wColumn_3[48] , 
        \wColumn_3[47] , \wColumn_3[46] , \wColumn_3[45] , \wColumn_3[44] , 
        \wColumn_3[43] , \wColumn_3[42] , \wColumn_3[41] , \wColumn_3[40] , 
        \wColumn_3[39] , \wColumn_3[38] , \wColumn_3[37] , \wColumn_3[36] , 
        \wColumn_3[35] , \wColumn_3[34] , \wColumn_3[33] , \wColumn_3[32] , 
        \wColumn_3[31] , \wColumn_3[30] , \wColumn_3[29] , \wColumn_3[28] , 
        \wColumn_3[27] , \wColumn_3[26] , \wColumn_3[25] , \wColumn_3[24] , 
        \wColumn_3[23] , \wColumn_3[22] , \wColumn_3[21] , \wColumn_3[20] , 
        \wColumn_3[19] , \wColumn_3[18] , \wColumn_3[17] , \wColumn_3[16] , 
        \wColumn_3[15] , \wColumn_3[14] , \wColumn_3[13] , \wColumn_3[12] , 
        \wColumn_3[11] , \wColumn_3[10] , \wColumn_3[9] , \wColumn_3[8] , 
        \wColumn_3[7] , \wColumn_3[6] , \wColumn_3[5] , \wColumn_3[4] , 
        \wColumn_3[3] , \wColumn_3[2] , \wColumn_3[1] , \wColumn_3[0] }), 
        .PDiagOut({\wPDiag_3[63] , \wPDiag_3[62] , \wPDiag_3[61] , 
        \wPDiag_3[60] , \wPDiag_3[59] , \wPDiag_3[58] , \wPDiag_3[57] , 
        \wPDiag_3[56] , \wPDiag_3[55] , \wPDiag_3[54] , \wPDiag_3[53] , 
        \wPDiag_3[52] , \wPDiag_3[51] , \wPDiag_3[50] , \wPDiag_3[49] , 
        \wPDiag_3[48] , \wPDiag_3[47] , \wPDiag_3[46] , \wPDiag_3[45] , 
        \wPDiag_3[44] , \wPDiag_3[43] , \wPDiag_3[42] , \wPDiag_3[41] , 
        \wPDiag_3[40] , \wPDiag_3[39] , \wPDiag_3[38] , \wPDiag_3[37] , 
        \wPDiag_3[36] , \wPDiag_3[35] , \wPDiag_3[34] , \wPDiag_3[33] , 
        \wPDiag_3[32] , \wPDiag_3[31] , \wPDiag_3[30] , \wPDiag_3[29] , 
        \wPDiag_3[28] , \wPDiag_3[27] , \wPDiag_3[26] , \wPDiag_3[25] , 
        \wPDiag_3[24] , \wPDiag_3[23] , \wPDiag_3[22] , \wPDiag_3[21] , 
        \wPDiag_3[20] , \wPDiag_3[19] , \wPDiag_3[18] , \wPDiag_3[17] , 
        \wPDiag_3[16] , \wPDiag_3[15] , \wPDiag_3[14] , \wPDiag_3[13] , 
        \wPDiag_3[12] , \wPDiag_3[11] , \wPDiag_3[10] , \wPDiag_3[9] , 
        \wPDiag_3[8] , \wPDiag_3[7] , \wPDiag_3[6] , \wPDiag_3[5] , 
        \wPDiag_3[4] , \wPDiag_3[3] , \wPDiag_3[2] , \wPDiag_3[1] , 
        \wPDiag_3[0] }), .NDiagOut({\wNDiag_3[63] , \wNDiag_3[62] , 
        \wNDiag_3[61] , \wNDiag_3[60] , \wNDiag_3[59] , \wNDiag_3[58] , 
        \wNDiag_3[57] , \wNDiag_3[56] , \wNDiag_3[55] , \wNDiag_3[54] , 
        \wNDiag_3[53] , \wNDiag_3[52] , \wNDiag_3[51] , \wNDiag_3[50] , 
        \wNDiag_3[49] , \wNDiag_3[48] , \wNDiag_3[47] , \wNDiag_3[46] , 
        \wNDiag_3[45] , \wNDiag_3[44] , \wNDiag_3[43] , \wNDiag_3[42] , 
        \wNDiag_3[41] , \wNDiag_3[40] , \wNDiag_3[39] , \wNDiag_3[38] , 
        \wNDiag_3[37] , \wNDiag_3[36] , \wNDiag_3[35] , \wNDiag_3[34] , 
        \wNDiag_3[33] , \wNDiag_3[32] , \wNDiag_3[31] , \wNDiag_3[30] , 
        \wNDiag_3[29] , \wNDiag_3[28] , \wNDiag_3[27] , \wNDiag_3[26] , 
        \wNDiag_3[25] , \wNDiag_3[24] , \wNDiag_3[23] , \wNDiag_3[22] , 
        \wNDiag_3[21] , \wNDiag_3[20] , \wNDiag_3[19] , \wNDiag_3[18] , 
        \wNDiag_3[17] , \wNDiag_3[16] , \wNDiag_3[15] , \wNDiag_3[14] , 
        \wNDiag_3[13] , \wNDiag_3[12] , \wNDiag_3[11] , \wNDiag_3[10] , 
        \wNDiag_3[9] , \wNDiag_3[8] , \wNDiag_3[7] , \wNDiag_3[6] , 
        \wNDiag_3[5] , \wNDiag_3[4] , \wNDiag_3[3] , \wNDiag_3[2] , 
        \wNDiag_3[1] , \wNDiag_3[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_3 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_4[6] , \wScan_4[5] , \wScan_4[4] , 
        \wScan_4[3] , \wScan_4[2] , \wScan_4[1] , \wScan_4[0] }), .ScanOut({
        \wScan_3[6] , \wScan_3[5] , \wScan_3[4] , \wScan_3[3] , \wScan_3[2] , 
        \wScan_3[1] , \wScan_3[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_3[0] ), 
        .ReturnIn(\wReturn_4[0] ), .ColIn({\wColumn_3[63] , \wColumn_3[62] , 
        \wColumn_3[61] , \wColumn_3[60] , \wColumn_3[59] , \wColumn_3[58] , 
        \wColumn_3[57] , \wColumn_3[56] , \wColumn_3[55] , \wColumn_3[54] , 
        \wColumn_3[53] , \wColumn_3[52] , \wColumn_3[51] , \wColumn_3[50] , 
        \wColumn_3[49] , \wColumn_3[48] , \wColumn_3[47] , \wColumn_3[46] , 
        \wColumn_3[45] , \wColumn_3[44] , \wColumn_3[43] , \wColumn_3[42] , 
        \wColumn_3[41] , \wColumn_3[40] , \wColumn_3[39] , \wColumn_3[38] , 
        \wColumn_3[37] , \wColumn_3[36] , \wColumn_3[35] , \wColumn_3[34] , 
        \wColumn_3[33] , \wColumn_3[32] , \wColumn_3[31] , \wColumn_3[30] , 
        \wColumn_3[29] , \wColumn_3[28] , \wColumn_3[27] , \wColumn_3[26] , 
        \wColumn_3[25] , \wColumn_3[24] , \wColumn_3[23] , \wColumn_3[22] , 
        \wColumn_3[21] , \wColumn_3[20] , \wColumn_3[19] , \wColumn_3[18] , 
        \wColumn_3[17] , \wColumn_3[16] , \wColumn_3[15] , \wColumn_3[14] , 
        \wColumn_3[13] , \wColumn_3[12] , \wColumn_3[11] , \wColumn_3[10] , 
        \wColumn_3[9] , \wColumn_3[8] , \wColumn_3[7] , \wColumn_3[6] , 
        \wColumn_3[5] , \wColumn_3[4] , \wColumn_3[3] , \wColumn_3[2] , 
        \wColumn_3[1] , \wColumn_3[0] }), .PDiagIn({\wPDiag_3[63] , 
        \wPDiag_3[62] , \wPDiag_3[61] , \wPDiag_3[60] , \wPDiag_3[59] , 
        \wPDiag_3[58] , \wPDiag_3[57] , \wPDiag_3[56] , \wPDiag_3[55] , 
        \wPDiag_3[54] , \wPDiag_3[53] , \wPDiag_3[52] , \wPDiag_3[51] , 
        \wPDiag_3[50] , \wPDiag_3[49] , \wPDiag_3[48] , \wPDiag_3[47] , 
        \wPDiag_3[46] , \wPDiag_3[45] , \wPDiag_3[44] , \wPDiag_3[43] , 
        \wPDiag_3[42] , \wPDiag_3[41] , \wPDiag_3[40] , \wPDiag_3[39] , 
        \wPDiag_3[38] , \wPDiag_3[37] , \wPDiag_3[36] , \wPDiag_3[35] , 
        \wPDiag_3[34] , \wPDiag_3[33] , \wPDiag_3[32] , \wPDiag_3[31] , 
        \wPDiag_3[30] , \wPDiag_3[29] , \wPDiag_3[28] , \wPDiag_3[27] , 
        \wPDiag_3[26] , \wPDiag_3[25] , \wPDiag_3[24] , \wPDiag_3[23] , 
        \wPDiag_3[22] , \wPDiag_3[21] , \wPDiag_3[20] , \wPDiag_3[19] , 
        \wPDiag_3[18] , \wPDiag_3[17] , \wPDiag_3[16] , \wPDiag_3[15] , 
        \wPDiag_3[14] , \wPDiag_3[13] , \wPDiag_3[12] , \wPDiag_3[11] , 
        \wPDiag_3[10] , \wPDiag_3[9] , \wPDiag_3[8] , \wPDiag_3[7] , 
        \wPDiag_3[6] , \wPDiag_3[5] , \wPDiag_3[4] , \wPDiag_3[3] , 
        \wPDiag_3[2] , \wPDiag_3[1] , \wPDiag_3[0] }), .NDiagIn({
        \wNDiag_3[63] , \wNDiag_3[62] , \wNDiag_3[61] , \wNDiag_3[60] , 
        \wNDiag_3[59] , \wNDiag_3[58] , \wNDiag_3[57] , \wNDiag_3[56] , 
        \wNDiag_3[55] , \wNDiag_3[54] , \wNDiag_3[53] , \wNDiag_3[52] , 
        \wNDiag_3[51] , \wNDiag_3[50] , \wNDiag_3[49] , \wNDiag_3[48] , 
        \wNDiag_3[47] , \wNDiag_3[46] , \wNDiag_3[45] , \wNDiag_3[44] , 
        \wNDiag_3[43] , \wNDiag_3[42] , \wNDiag_3[41] , \wNDiag_3[40] , 
        \wNDiag_3[39] , \wNDiag_3[38] , \wNDiag_3[37] , \wNDiag_3[36] , 
        \wNDiag_3[35] , \wNDiag_3[34] , \wNDiag_3[33] , \wNDiag_3[32] , 
        \wNDiag_3[31] , \wNDiag_3[30] , \wNDiag_3[29] , \wNDiag_3[28] , 
        \wNDiag_3[27] , \wNDiag_3[26] , \wNDiag_3[25] , \wNDiag_3[24] , 
        \wNDiag_3[23] , \wNDiag_3[22] , \wNDiag_3[21] , \wNDiag_3[20] , 
        \wNDiag_3[19] , \wNDiag_3[18] , \wNDiag_3[17] , \wNDiag_3[16] , 
        \wNDiag_3[15] , \wNDiag_3[14] , \wNDiag_3[13] , \wNDiag_3[12] , 
        \wNDiag_3[11] , \wNDiag_3[10] , \wNDiag_3[9] , \wNDiag_3[8] , 
        \wNDiag_3[7] , \wNDiag_3[6] , \wNDiag_3[5] , \wNDiag_3[4] , 
        \wNDiag_3[3] , \wNDiag_3[2] , \wNDiag_3[1] , \wNDiag_3[0] }), 
        .CallOut(\wCall_4[0] ), .ReturnOut(\wReturn_3[0] ), .ColOut({
        \wColumn_4[63] , \wColumn_4[62] , \wColumn_4[61] , \wColumn_4[60] , 
        \wColumn_4[59] , \wColumn_4[58] , \wColumn_4[57] , \wColumn_4[56] , 
        \wColumn_4[55] , \wColumn_4[54] , \wColumn_4[53] , \wColumn_4[52] , 
        \wColumn_4[51] , \wColumn_4[50] , \wColumn_4[49] , \wColumn_4[48] , 
        \wColumn_4[47] , \wColumn_4[46] , \wColumn_4[45] , \wColumn_4[44] , 
        \wColumn_4[43] , \wColumn_4[42] , \wColumn_4[41] , \wColumn_4[40] , 
        \wColumn_4[39] , \wColumn_4[38] , \wColumn_4[37] , \wColumn_4[36] , 
        \wColumn_4[35] , \wColumn_4[34] , \wColumn_4[33] , \wColumn_4[32] , 
        \wColumn_4[31] , \wColumn_4[30] , \wColumn_4[29] , \wColumn_4[28] , 
        \wColumn_4[27] , \wColumn_4[26] , \wColumn_4[25] , \wColumn_4[24] , 
        \wColumn_4[23] , \wColumn_4[22] , \wColumn_4[21] , \wColumn_4[20] , 
        \wColumn_4[19] , \wColumn_4[18] , \wColumn_4[17] , \wColumn_4[16] , 
        \wColumn_4[15] , \wColumn_4[14] , \wColumn_4[13] , \wColumn_4[12] , 
        \wColumn_4[11] , \wColumn_4[10] , \wColumn_4[9] , \wColumn_4[8] , 
        \wColumn_4[7] , \wColumn_4[6] , \wColumn_4[5] , \wColumn_4[4] , 
        \wColumn_4[3] , \wColumn_4[2] , \wColumn_4[1] , \wColumn_4[0] }), 
        .PDiagOut({\wPDiag_4[63] , \wPDiag_4[62] , \wPDiag_4[61] , 
        \wPDiag_4[60] , \wPDiag_4[59] , \wPDiag_4[58] , \wPDiag_4[57] , 
        \wPDiag_4[56] , \wPDiag_4[55] , \wPDiag_4[54] , \wPDiag_4[53] , 
        \wPDiag_4[52] , \wPDiag_4[51] , \wPDiag_4[50] , \wPDiag_4[49] , 
        \wPDiag_4[48] , \wPDiag_4[47] , \wPDiag_4[46] , \wPDiag_4[45] , 
        \wPDiag_4[44] , \wPDiag_4[43] , \wPDiag_4[42] , \wPDiag_4[41] , 
        \wPDiag_4[40] , \wPDiag_4[39] , \wPDiag_4[38] , \wPDiag_4[37] , 
        \wPDiag_4[36] , \wPDiag_4[35] , \wPDiag_4[34] , \wPDiag_4[33] , 
        \wPDiag_4[32] , \wPDiag_4[31] , \wPDiag_4[30] , \wPDiag_4[29] , 
        \wPDiag_4[28] , \wPDiag_4[27] , \wPDiag_4[26] , \wPDiag_4[25] , 
        \wPDiag_4[24] , \wPDiag_4[23] , \wPDiag_4[22] , \wPDiag_4[21] , 
        \wPDiag_4[20] , \wPDiag_4[19] , \wPDiag_4[18] , \wPDiag_4[17] , 
        \wPDiag_4[16] , \wPDiag_4[15] , \wPDiag_4[14] , \wPDiag_4[13] , 
        \wPDiag_4[12] , \wPDiag_4[11] , \wPDiag_4[10] , \wPDiag_4[9] , 
        \wPDiag_4[8] , \wPDiag_4[7] , \wPDiag_4[6] , \wPDiag_4[5] , 
        \wPDiag_4[4] , \wPDiag_4[3] , \wPDiag_4[2] , \wPDiag_4[1] , 
        \wPDiag_4[0] }), .NDiagOut({\wNDiag_4[63] , \wNDiag_4[62] , 
        \wNDiag_4[61] , \wNDiag_4[60] , \wNDiag_4[59] , \wNDiag_4[58] , 
        \wNDiag_4[57] , \wNDiag_4[56] , \wNDiag_4[55] , \wNDiag_4[54] , 
        \wNDiag_4[53] , \wNDiag_4[52] , \wNDiag_4[51] , \wNDiag_4[50] , 
        \wNDiag_4[49] , \wNDiag_4[48] , \wNDiag_4[47] , \wNDiag_4[46] , 
        \wNDiag_4[45] , \wNDiag_4[44] , \wNDiag_4[43] , \wNDiag_4[42] , 
        \wNDiag_4[41] , \wNDiag_4[40] , \wNDiag_4[39] , \wNDiag_4[38] , 
        \wNDiag_4[37] , \wNDiag_4[36] , \wNDiag_4[35] , \wNDiag_4[34] , 
        \wNDiag_4[33] , \wNDiag_4[32] , \wNDiag_4[31] , \wNDiag_4[30] , 
        \wNDiag_4[29] , \wNDiag_4[28] , \wNDiag_4[27] , \wNDiag_4[26] , 
        \wNDiag_4[25] , \wNDiag_4[24] , \wNDiag_4[23] , \wNDiag_4[22] , 
        \wNDiag_4[21] , \wNDiag_4[20] , \wNDiag_4[19] , \wNDiag_4[18] , 
        \wNDiag_4[17] , \wNDiag_4[16] , \wNDiag_4[15] , \wNDiag_4[14] , 
        \wNDiag_4[13] , \wNDiag_4[12] , \wNDiag_4[11] , \wNDiag_4[10] , 
        \wNDiag_4[9] , \wNDiag_4[8] , \wNDiag_4[7] , \wNDiag_4[6] , 
        \wNDiag_4[5] , \wNDiag_4[4] , \wNDiag_4[3] , \wNDiag_4[2] , 
        \wNDiag_4[1] , \wNDiag_4[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_27 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_28[6] , \wScan_28[5] , \wScan_28[4] , 
        \wScan_28[3] , \wScan_28[2] , \wScan_28[1] , \wScan_28[0] }), 
        .ScanOut({\wScan_27[6] , \wScan_27[5] , \wScan_27[4] , \wScan_27[3] , 
        \wScan_27[2] , \wScan_27[1] , \wScan_27[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_27[0] ), .ReturnIn(\wReturn_28[0] ), .ColIn({
        \wColumn_27[63] , \wColumn_27[62] , \wColumn_27[61] , \wColumn_27[60] , 
        \wColumn_27[59] , \wColumn_27[58] , \wColumn_27[57] , \wColumn_27[56] , 
        \wColumn_27[55] , \wColumn_27[54] , \wColumn_27[53] , \wColumn_27[52] , 
        \wColumn_27[51] , \wColumn_27[50] , \wColumn_27[49] , \wColumn_27[48] , 
        \wColumn_27[47] , \wColumn_27[46] , \wColumn_27[45] , \wColumn_27[44] , 
        \wColumn_27[43] , \wColumn_27[42] , \wColumn_27[41] , \wColumn_27[40] , 
        \wColumn_27[39] , \wColumn_27[38] , \wColumn_27[37] , \wColumn_27[36] , 
        \wColumn_27[35] , \wColumn_27[34] , \wColumn_27[33] , \wColumn_27[32] , 
        \wColumn_27[31] , \wColumn_27[30] , \wColumn_27[29] , \wColumn_27[28] , 
        \wColumn_27[27] , \wColumn_27[26] , \wColumn_27[25] , \wColumn_27[24] , 
        \wColumn_27[23] , \wColumn_27[22] , \wColumn_27[21] , \wColumn_27[20] , 
        \wColumn_27[19] , \wColumn_27[18] , \wColumn_27[17] , \wColumn_27[16] , 
        \wColumn_27[15] , \wColumn_27[14] , \wColumn_27[13] , \wColumn_27[12] , 
        \wColumn_27[11] , \wColumn_27[10] , \wColumn_27[9] , \wColumn_27[8] , 
        \wColumn_27[7] , \wColumn_27[6] , \wColumn_27[5] , \wColumn_27[4] , 
        \wColumn_27[3] , \wColumn_27[2] , \wColumn_27[1] , \wColumn_27[0] }), 
        .PDiagIn({\wPDiag_27[63] , \wPDiag_27[62] , \wPDiag_27[61] , 
        \wPDiag_27[60] , \wPDiag_27[59] , \wPDiag_27[58] , \wPDiag_27[57] , 
        \wPDiag_27[56] , \wPDiag_27[55] , \wPDiag_27[54] , \wPDiag_27[53] , 
        \wPDiag_27[52] , \wPDiag_27[51] , \wPDiag_27[50] , \wPDiag_27[49] , 
        \wPDiag_27[48] , \wPDiag_27[47] , \wPDiag_27[46] , \wPDiag_27[45] , 
        \wPDiag_27[44] , \wPDiag_27[43] , \wPDiag_27[42] , \wPDiag_27[41] , 
        \wPDiag_27[40] , \wPDiag_27[39] , \wPDiag_27[38] , \wPDiag_27[37] , 
        \wPDiag_27[36] , \wPDiag_27[35] , \wPDiag_27[34] , \wPDiag_27[33] , 
        \wPDiag_27[32] , \wPDiag_27[31] , \wPDiag_27[30] , \wPDiag_27[29] , 
        \wPDiag_27[28] , \wPDiag_27[27] , \wPDiag_27[26] , \wPDiag_27[25] , 
        \wPDiag_27[24] , \wPDiag_27[23] , \wPDiag_27[22] , \wPDiag_27[21] , 
        \wPDiag_27[20] , \wPDiag_27[19] , \wPDiag_27[18] , \wPDiag_27[17] , 
        \wPDiag_27[16] , \wPDiag_27[15] , \wPDiag_27[14] , \wPDiag_27[13] , 
        \wPDiag_27[12] , \wPDiag_27[11] , \wPDiag_27[10] , \wPDiag_27[9] , 
        \wPDiag_27[8] , \wPDiag_27[7] , \wPDiag_27[6] , \wPDiag_27[5] , 
        \wPDiag_27[4] , \wPDiag_27[3] , \wPDiag_27[2] , \wPDiag_27[1] , 
        \wPDiag_27[0] }), .NDiagIn({\wNDiag_27[63] , \wNDiag_27[62] , 
        \wNDiag_27[61] , \wNDiag_27[60] , \wNDiag_27[59] , \wNDiag_27[58] , 
        \wNDiag_27[57] , \wNDiag_27[56] , \wNDiag_27[55] , \wNDiag_27[54] , 
        \wNDiag_27[53] , \wNDiag_27[52] , \wNDiag_27[51] , \wNDiag_27[50] , 
        \wNDiag_27[49] , \wNDiag_27[48] , \wNDiag_27[47] , \wNDiag_27[46] , 
        \wNDiag_27[45] , \wNDiag_27[44] , \wNDiag_27[43] , \wNDiag_27[42] , 
        \wNDiag_27[41] , \wNDiag_27[40] , \wNDiag_27[39] , \wNDiag_27[38] , 
        \wNDiag_27[37] , \wNDiag_27[36] , \wNDiag_27[35] , \wNDiag_27[34] , 
        \wNDiag_27[33] , \wNDiag_27[32] , \wNDiag_27[31] , \wNDiag_27[30] , 
        \wNDiag_27[29] , \wNDiag_27[28] , \wNDiag_27[27] , \wNDiag_27[26] , 
        \wNDiag_27[25] , \wNDiag_27[24] , \wNDiag_27[23] , \wNDiag_27[22] , 
        \wNDiag_27[21] , \wNDiag_27[20] , \wNDiag_27[19] , \wNDiag_27[18] , 
        \wNDiag_27[17] , \wNDiag_27[16] , \wNDiag_27[15] , \wNDiag_27[14] , 
        \wNDiag_27[13] , \wNDiag_27[12] , \wNDiag_27[11] , \wNDiag_27[10] , 
        \wNDiag_27[9] , \wNDiag_27[8] , \wNDiag_27[7] , \wNDiag_27[6] , 
        \wNDiag_27[5] , \wNDiag_27[4] , \wNDiag_27[3] , \wNDiag_27[2] , 
        \wNDiag_27[1] , \wNDiag_27[0] }), .CallOut(\wCall_28[0] ), .ReturnOut(
        \wReturn_27[0] ), .ColOut({\wColumn_28[63] , \wColumn_28[62] , 
        \wColumn_28[61] , \wColumn_28[60] , \wColumn_28[59] , \wColumn_28[58] , 
        \wColumn_28[57] , \wColumn_28[56] , \wColumn_28[55] , \wColumn_28[54] , 
        \wColumn_28[53] , \wColumn_28[52] , \wColumn_28[51] , \wColumn_28[50] , 
        \wColumn_28[49] , \wColumn_28[48] , \wColumn_28[47] , \wColumn_28[46] , 
        \wColumn_28[45] , \wColumn_28[44] , \wColumn_28[43] , \wColumn_28[42] , 
        \wColumn_28[41] , \wColumn_28[40] , \wColumn_28[39] , \wColumn_28[38] , 
        \wColumn_28[37] , \wColumn_28[36] , \wColumn_28[35] , \wColumn_28[34] , 
        \wColumn_28[33] , \wColumn_28[32] , \wColumn_28[31] , \wColumn_28[30] , 
        \wColumn_28[29] , \wColumn_28[28] , \wColumn_28[27] , \wColumn_28[26] , 
        \wColumn_28[25] , \wColumn_28[24] , \wColumn_28[23] , \wColumn_28[22] , 
        \wColumn_28[21] , \wColumn_28[20] , \wColumn_28[19] , \wColumn_28[18] , 
        \wColumn_28[17] , \wColumn_28[16] , \wColumn_28[15] , \wColumn_28[14] , 
        \wColumn_28[13] , \wColumn_28[12] , \wColumn_28[11] , \wColumn_28[10] , 
        \wColumn_28[9] , \wColumn_28[8] , \wColumn_28[7] , \wColumn_28[6] , 
        \wColumn_28[5] , \wColumn_28[4] , \wColumn_28[3] , \wColumn_28[2] , 
        \wColumn_28[1] , \wColumn_28[0] }), .PDiagOut({\wPDiag_28[63] , 
        \wPDiag_28[62] , \wPDiag_28[61] , \wPDiag_28[60] , \wPDiag_28[59] , 
        \wPDiag_28[58] , \wPDiag_28[57] , \wPDiag_28[56] , \wPDiag_28[55] , 
        \wPDiag_28[54] , \wPDiag_28[53] , \wPDiag_28[52] , \wPDiag_28[51] , 
        \wPDiag_28[50] , \wPDiag_28[49] , \wPDiag_28[48] , \wPDiag_28[47] , 
        \wPDiag_28[46] , \wPDiag_28[45] , \wPDiag_28[44] , \wPDiag_28[43] , 
        \wPDiag_28[42] , \wPDiag_28[41] , \wPDiag_28[40] , \wPDiag_28[39] , 
        \wPDiag_28[38] , \wPDiag_28[37] , \wPDiag_28[36] , \wPDiag_28[35] , 
        \wPDiag_28[34] , \wPDiag_28[33] , \wPDiag_28[32] , \wPDiag_28[31] , 
        \wPDiag_28[30] , \wPDiag_28[29] , \wPDiag_28[28] , \wPDiag_28[27] , 
        \wPDiag_28[26] , \wPDiag_28[25] , \wPDiag_28[24] , \wPDiag_28[23] , 
        \wPDiag_28[22] , \wPDiag_28[21] , \wPDiag_28[20] , \wPDiag_28[19] , 
        \wPDiag_28[18] , \wPDiag_28[17] , \wPDiag_28[16] , \wPDiag_28[15] , 
        \wPDiag_28[14] , \wPDiag_28[13] , \wPDiag_28[12] , \wPDiag_28[11] , 
        \wPDiag_28[10] , \wPDiag_28[9] , \wPDiag_28[8] , \wPDiag_28[7] , 
        \wPDiag_28[6] , \wPDiag_28[5] , \wPDiag_28[4] , \wPDiag_28[3] , 
        \wPDiag_28[2] , \wPDiag_28[1] , \wPDiag_28[0] }), .NDiagOut({
        \wNDiag_28[63] , \wNDiag_28[62] , \wNDiag_28[61] , \wNDiag_28[60] , 
        \wNDiag_28[59] , \wNDiag_28[58] , \wNDiag_28[57] , \wNDiag_28[56] , 
        \wNDiag_28[55] , \wNDiag_28[54] , \wNDiag_28[53] , \wNDiag_28[52] , 
        \wNDiag_28[51] , \wNDiag_28[50] , \wNDiag_28[49] , \wNDiag_28[48] , 
        \wNDiag_28[47] , \wNDiag_28[46] , \wNDiag_28[45] , \wNDiag_28[44] , 
        \wNDiag_28[43] , \wNDiag_28[42] , \wNDiag_28[41] , \wNDiag_28[40] , 
        \wNDiag_28[39] , \wNDiag_28[38] , \wNDiag_28[37] , \wNDiag_28[36] , 
        \wNDiag_28[35] , \wNDiag_28[34] , \wNDiag_28[33] , \wNDiag_28[32] , 
        \wNDiag_28[31] , \wNDiag_28[30] , \wNDiag_28[29] , \wNDiag_28[28] , 
        \wNDiag_28[27] , \wNDiag_28[26] , \wNDiag_28[25] , \wNDiag_28[24] , 
        \wNDiag_28[23] , \wNDiag_28[22] , \wNDiag_28[21] , \wNDiag_28[20] , 
        \wNDiag_28[19] , \wNDiag_28[18] , \wNDiag_28[17] , \wNDiag_28[16] , 
        \wNDiag_28[15] , \wNDiag_28[14] , \wNDiag_28[13] , \wNDiag_28[12] , 
        \wNDiag_28[11] , \wNDiag_28[10] , \wNDiag_28[9] , \wNDiag_28[8] , 
        \wNDiag_28[7] , \wNDiag_28[6] , \wNDiag_28[5] , \wNDiag_28[4] , 
        \wNDiag_28[3] , \wNDiag_28[2] , \wNDiag_28[1] , \wNDiag_28[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_49 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_50[6] , \wScan_50[5] , \wScan_50[4] , 
        \wScan_50[3] , \wScan_50[2] , \wScan_50[1] , \wScan_50[0] }), 
        .ScanOut({\wScan_49[6] , \wScan_49[5] , \wScan_49[4] , \wScan_49[3] , 
        \wScan_49[2] , \wScan_49[1] , \wScan_49[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_49[0] ), .ReturnIn(\wReturn_50[0] ), .ColIn({
        \wColumn_49[63] , \wColumn_49[62] , \wColumn_49[61] , \wColumn_49[60] , 
        \wColumn_49[59] , \wColumn_49[58] , \wColumn_49[57] , \wColumn_49[56] , 
        \wColumn_49[55] , \wColumn_49[54] , \wColumn_49[53] , \wColumn_49[52] , 
        \wColumn_49[51] , \wColumn_49[50] , \wColumn_49[49] , \wColumn_49[48] , 
        \wColumn_49[47] , \wColumn_49[46] , \wColumn_49[45] , \wColumn_49[44] , 
        \wColumn_49[43] , \wColumn_49[42] , \wColumn_49[41] , \wColumn_49[40] , 
        \wColumn_49[39] , \wColumn_49[38] , \wColumn_49[37] , \wColumn_49[36] , 
        \wColumn_49[35] , \wColumn_49[34] , \wColumn_49[33] , \wColumn_49[32] , 
        \wColumn_49[31] , \wColumn_49[30] , \wColumn_49[29] , \wColumn_49[28] , 
        \wColumn_49[27] , \wColumn_49[26] , \wColumn_49[25] , \wColumn_49[24] , 
        \wColumn_49[23] , \wColumn_49[22] , \wColumn_49[21] , \wColumn_49[20] , 
        \wColumn_49[19] , \wColumn_49[18] , \wColumn_49[17] , \wColumn_49[16] , 
        \wColumn_49[15] , \wColumn_49[14] , \wColumn_49[13] , \wColumn_49[12] , 
        \wColumn_49[11] , \wColumn_49[10] , \wColumn_49[9] , \wColumn_49[8] , 
        \wColumn_49[7] , \wColumn_49[6] , \wColumn_49[5] , \wColumn_49[4] , 
        \wColumn_49[3] , \wColumn_49[2] , \wColumn_49[1] , \wColumn_49[0] }), 
        .PDiagIn({\wPDiag_49[63] , \wPDiag_49[62] , \wPDiag_49[61] , 
        \wPDiag_49[60] , \wPDiag_49[59] , \wPDiag_49[58] , \wPDiag_49[57] , 
        \wPDiag_49[56] , \wPDiag_49[55] , \wPDiag_49[54] , \wPDiag_49[53] , 
        \wPDiag_49[52] , \wPDiag_49[51] , \wPDiag_49[50] , \wPDiag_49[49] , 
        \wPDiag_49[48] , \wPDiag_49[47] , \wPDiag_49[46] , \wPDiag_49[45] , 
        \wPDiag_49[44] , \wPDiag_49[43] , \wPDiag_49[42] , \wPDiag_49[41] , 
        \wPDiag_49[40] , \wPDiag_49[39] , \wPDiag_49[38] , \wPDiag_49[37] , 
        \wPDiag_49[36] , \wPDiag_49[35] , \wPDiag_49[34] , \wPDiag_49[33] , 
        \wPDiag_49[32] , \wPDiag_49[31] , \wPDiag_49[30] , \wPDiag_49[29] , 
        \wPDiag_49[28] , \wPDiag_49[27] , \wPDiag_49[26] , \wPDiag_49[25] , 
        \wPDiag_49[24] , \wPDiag_49[23] , \wPDiag_49[22] , \wPDiag_49[21] , 
        \wPDiag_49[20] , \wPDiag_49[19] , \wPDiag_49[18] , \wPDiag_49[17] , 
        \wPDiag_49[16] , \wPDiag_49[15] , \wPDiag_49[14] , \wPDiag_49[13] , 
        \wPDiag_49[12] , \wPDiag_49[11] , \wPDiag_49[10] , \wPDiag_49[9] , 
        \wPDiag_49[8] , \wPDiag_49[7] , \wPDiag_49[6] , \wPDiag_49[5] , 
        \wPDiag_49[4] , \wPDiag_49[3] , \wPDiag_49[2] , \wPDiag_49[1] , 
        \wPDiag_49[0] }), .NDiagIn({\wNDiag_49[63] , \wNDiag_49[62] , 
        \wNDiag_49[61] , \wNDiag_49[60] , \wNDiag_49[59] , \wNDiag_49[58] , 
        \wNDiag_49[57] , \wNDiag_49[56] , \wNDiag_49[55] , \wNDiag_49[54] , 
        \wNDiag_49[53] , \wNDiag_49[52] , \wNDiag_49[51] , \wNDiag_49[50] , 
        \wNDiag_49[49] , \wNDiag_49[48] , \wNDiag_49[47] , \wNDiag_49[46] , 
        \wNDiag_49[45] , \wNDiag_49[44] , \wNDiag_49[43] , \wNDiag_49[42] , 
        \wNDiag_49[41] , \wNDiag_49[40] , \wNDiag_49[39] , \wNDiag_49[38] , 
        \wNDiag_49[37] , \wNDiag_49[36] , \wNDiag_49[35] , \wNDiag_49[34] , 
        \wNDiag_49[33] , \wNDiag_49[32] , \wNDiag_49[31] , \wNDiag_49[30] , 
        \wNDiag_49[29] , \wNDiag_49[28] , \wNDiag_49[27] , \wNDiag_49[26] , 
        \wNDiag_49[25] , \wNDiag_49[24] , \wNDiag_49[23] , \wNDiag_49[22] , 
        \wNDiag_49[21] , \wNDiag_49[20] , \wNDiag_49[19] , \wNDiag_49[18] , 
        \wNDiag_49[17] , \wNDiag_49[16] , \wNDiag_49[15] , \wNDiag_49[14] , 
        \wNDiag_49[13] , \wNDiag_49[12] , \wNDiag_49[11] , \wNDiag_49[10] , 
        \wNDiag_49[9] , \wNDiag_49[8] , \wNDiag_49[7] , \wNDiag_49[6] , 
        \wNDiag_49[5] , \wNDiag_49[4] , \wNDiag_49[3] , \wNDiag_49[2] , 
        \wNDiag_49[1] , \wNDiag_49[0] }), .CallOut(\wCall_50[0] ), .ReturnOut(
        \wReturn_49[0] ), .ColOut({\wColumn_50[63] , \wColumn_50[62] , 
        \wColumn_50[61] , \wColumn_50[60] , \wColumn_50[59] , \wColumn_50[58] , 
        \wColumn_50[57] , \wColumn_50[56] , \wColumn_50[55] , \wColumn_50[54] , 
        \wColumn_50[53] , \wColumn_50[52] , \wColumn_50[51] , \wColumn_50[50] , 
        \wColumn_50[49] , \wColumn_50[48] , \wColumn_50[47] , \wColumn_50[46] , 
        \wColumn_50[45] , \wColumn_50[44] , \wColumn_50[43] , \wColumn_50[42] , 
        \wColumn_50[41] , \wColumn_50[40] , \wColumn_50[39] , \wColumn_50[38] , 
        \wColumn_50[37] , \wColumn_50[36] , \wColumn_50[35] , \wColumn_50[34] , 
        \wColumn_50[33] , \wColumn_50[32] , \wColumn_50[31] , \wColumn_50[30] , 
        \wColumn_50[29] , \wColumn_50[28] , \wColumn_50[27] , \wColumn_50[26] , 
        \wColumn_50[25] , \wColumn_50[24] , \wColumn_50[23] , \wColumn_50[22] , 
        \wColumn_50[21] , \wColumn_50[20] , \wColumn_50[19] , \wColumn_50[18] , 
        \wColumn_50[17] , \wColumn_50[16] , \wColumn_50[15] , \wColumn_50[14] , 
        \wColumn_50[13] , \wColumn_50[12] , \wColumn_50[11] , \wColumn_50[10] , 
        \wColumn_50[9] , \wColumn_50[8] , \wColumn_50[7] , \wColumn_50[6] , 
        \wColumn_50[5] , \wColumn_50[4] , \wColumn_50[3] , \wColumn_50[2] , 
        \wColumn_50[1] , \wColumn_50[0] }), .PDiagOut({\wPDiag_50[63] , 
        \wPDiag_50[62] , \wPDiag_50[61] , \wPDiag_50[60] , \wPDiag_50[59] , 
        \wPDiag_50[58] , \wPDiag_50[57] , \wPDiag_50[56] , \wPDiag_50[55] , 
        \wPDiag_50[54] , \wPDiag_50[53] , \wPDiag_50[52] , \wPDiag_50[51] , 
        \wPDiag_50[50] , \wPDiag_50[49] , \wPDiag_50[48] , \wPDiag_50[47] , 
        \wPDiag_50[46] , \wPDiag_50[45] , \wPDiag_50[44] , \wPDiag_50[43] , 
        \wPDiag_50[42] , \wPDiag_50[41] , \wPDiag_50[40] , \wPDiag_50[39] , 
        \wPDiag_50[38] , \wPDiag_50[37] , \wPDiag_50[36] , \wPDiag_50[35] , 
        \wPDiag_50[34] , \wPDiag_50[33] , \wPDiag_50[32] , \wPDiag_50[31] , 
        \wPDiag_50[30] , \wPDiag_50[29] , \wPDiag_50[28] , \wPDiag_50[27] , 
        \wPDiag_50[26] , \wPDiag_50[25] , \wPDiag_50[24] , \wPDiag_50[23] , 
        \wPDiag_50[22] , \wPDiag_50[21] , \wPDiag_50[20] , \wPDiag_50[19] , 
        \wPDiag_50[18] , \wPDiag_50[17] , \wPDiag_50[16] , \wPDiag_50[15] , 
        \wPDiag_50[14] , \wPDiag_50[13] , \wPDiag_50[12] , \wPDiag_50[11] , 
        \wPDiag_50[10] , \wPDiag_50[9] , \wPDiag_50[8] , \wPDiag_50[7] , 
        \wPDiag_50[6] , \wPDiag_50[5] , \wPDiag_50[4] , \wPDiag_50[3] , 
        \wPDiag_50[2] , \wPDiag_50[1] , \wPDiag_50[0] }), .NDiagOut({
        \wNDiag_50[63] , \wNDiag_50[62] , \wNDiag_50[61] , \wNDiag_50[60] , 
        \wNDiag_50[59] , \wNDiag_50[58] , \wNDiag_50[57] , \wNDiag_50[56] , 
        \wNDiag_50[55] , \wNDiag_50[54] , \wNDiag_50[53] , \wNDiag_50[52] , 
        \wNDiag_50[51] , \wNDiag_50[50] , \wNDiag_50[49] , \wNDiag_50[48] , 
        \wNDiag_50[47] , \wNDiag_50[46] , \wNDiag_50[45] , \wNDiag_50[44] , 
        \wNDiag_50[43] , \wNDiag_50[42] , \wNDiag_50[41] , \wNDiag_50[40] , 
        \wNDiag_50[39] , \wNDiag_50[38] , \wNDiag_50[37] , \wNDiag_50[36] , 
        \wNDiag_50[35] , \wNDiag_50[34] , \wNDiag_50[33] , \wNDiag_50[32] , 
        \wNDiag_50[31] , \wNDiag_50[30] , \wNDiag_50[29] , \wNDiag_50[28] , 
        \wNDiag_50[27] , \wNDiag_50[26] , \wNDiag_50[25] , \wNDiag_50[24] , 
        \wNDiag_50[23] , \wNDiag_50[22] , \wNDiag_50[21] , \wNDiag_50[20] , 
        \wNDiag_50[19] , \wNDiag_50[18] , \wNDiag_50[17] , \wNDiag_50[16] , 
        \wNDiag_50[15] , \wNDiag_50[14] , \wNDiag_50[13] , \wNDiag_50[12] , 
        \wNDiag_50[11] , \wNDiag_50[10] , \wNDiag_50[9] , \wNDiag_50[8] , 
        \wNDiag_50[7] , \wNDiag_50[6] , \wNDiag_50[5] , \wNDiag_50[4] , 
        \wNDiag_50[3] , \wNDiag_50[2] , \wNDiag_50[1] , \wNDiag_50[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_52 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_53[6] , \wScan_53[5] , \wScan_53[4] , 
        \wScan_53[3] , \wScan_53[2] , \wScan_53[1] , \wScan_53[0] }), 
        .ScanOut({\wScan_52[6] , \wScan_52[5] , \wScan_52[4] , \wScan_52[3] , 
        \wScan_52[2] , \wScan_52[1] , \wScan_52[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_52[0] ), .ReturnIn(\wReturn_53[0] ), .ColIn({
        \wColumn_52[63] , \wColumn_52[62] , \wColumn_52[61] , \wColumn_52[60] , 
        \wColumn_52[59] , \wColumn_52[58] , \wColumn_52[57] , \wColumn_52[56] , 
        \wColumn_52[55] , \wColumn_52[54] , \wColumn_52[53] , \wColumn_52[52] , 
        \wColumn_52[51] , \wColumn_52[50] , \wColumn_52[49] , \wColumn_52[48] , 
        \wColumn_52[47] , \wColumn_52[46] , \wColumn_52[45] , \wColumn_52[44] , 
        \wColumn_52[43] , \wColumn_52[42] , \wColumn_52[41] , \wColumn_52[40] , 
        \wColumn_52[39] , \wColumn_52[38] , \wColumn_52[37] , \wColumn_52[36] , 
        \wColumn_52[35] , \wColumn_52[34] , \wColumn_52[33] , \wColumn_52[32] , 
        \wColumn_52[31] , \wColumn_52[30] , \wColumn_52[29] , \wColumn_52[28] , 
        \wColumn_52[27] , \wColumn_52[26] , \wColumn_52[25] , \wColumn_52[24] , 
        \wColumn_52[23] , \wColumn_52[22] , \wColumn_52[21] , \wColumn_52[20] , 
        \wColumn_52[19] , \wColumn_52[18] , \wColumn_52[17] , \wColumn_52[16] , 
        \wColumn_52[15] , \wColumn_52[14] , \wColumn_52[13] , \wColumn_52[12] , 
        \wColumn_52[11] , \wColumn_52[10] , \wColumn_52[9] , \wColumn_52[8] , 
        \wColumn_52[7] , \wColumn_52[6] , \wColumn_52[5] , \wColumn_52[4] , 
        \wColumn_52[3] , \wColumn_52[2] , \wColumn_52[1] , \wColumn_52[0] }), 
        .PDiagIn({\wPDiag_52[63] , \wPDiag_52[62] , \wPDiag_52[61] , 
        \wPDiag_52[60] , \wPDiag_52[59] , \wPDiag_52[58] , \wPDiag_52[57] , 
        \wPDiag_52[56] , \wPDiag_52[55] , \wPDiag_52[54] , \wPDiag_52[53] , 
        \wPDiag_52[52] , \wPDiag_52[51] , \wPDiag_52[50] , \wPDiag_52[49] , 
        \wPDiag_52[48] , \wPDiag_52[47] , \wPDiag_52[46] , \wPDiag_52[45] , 
        \wPDiag_52[44] , \wPDiag_52[43] , \wPDiag_52[42] , \wPDiag_52[41] , 
        \wPDiag_52[40] , \wPDiag_52[39] , \wPDiag_52[38] , \wPDiag_52[37] , 
        \wPDiag_52[36] , \wPDiag_52[35] , \wPDiag_52[34] , \wPDiag_52[33] , 
        \wPDiag_52[32] , \wPDiag_52[31] , \wPDiag_52[30] , \wPDiag_52[29] , 
        \wPDiag_52[28] , \wPDiag_52[27] , \wPDiag_52[26] , \wPDiag_52[25] , 
        \wPDiag_52[24] , \wPDiag_52[23] , \wPDiag_52[22] , \wPDiag_52[21] , 
        \wPDiag_52[20] , \wPDiag_52[19] , \wPDiag_52[18] , \wPDiag_52[17] , 
        \wPDiag_52[16] , \wPDiag_52[15] , \wPDiag_52[14] , \wPDiag_52[13] , 
        \wPDiag_52[12] , \wPDiag_52[11] , \wPDiag_52[10] , \wPDiag_52[9] , 
        \wPDiag_52[8] , \wPDiag_52[7] , \wPDiag_52[6] , \wPDiag_52[5] , 
        \wPDiag_52[4] , \wPDiag_52[3] , \wPDiag_52[2] , \wPDiag_52[1] , 
        \wPDiag_52[0] }), .NDiagIn({\wNDiag_52[63] , \wNDiag_52[62] , 
        \wNDiag_52[61] , \wNDiag_52[60] , \wNDiag_52[59] , \wNDiag_52[58] , 
        \wNDiag_52[57] , \wNDiag_52[56] , \wNDiag_52[55] , \wNDiag_52[54] , 
        \wNDiag_52[53] , \wNDiag_52[52] , \wNDiag_52[51] , \wNDiag_52[50] , 
        \wNDiag_52[49] , \wNDiag_52[48] , \wNDiag_52[47] , \wNDiag_52[46] , 
        \wNDiag_52[45] , \wNDiag_52[44] , \wNDiag_52[43] , \wNDiag_52[42] , 
        \wNDiag_52[41] , \wNDiag_52[40] , \wNDiag_52[39] , \wNDiag_52[38] , 
        \wNDiag_52[37] , \wNDiag_52[36] , \wNDiag_52[35] , \wNDiag_52[34] , 
        \wNDiag_52[33] , \wNDiag_52[32] , \wNDiag_52[31] , \wNDiag_52[30] , 
        \wNDiag_52[29] , \wNDiag_52[28] , \wNDiag_52[27] , \wNDiag_52[26] , 
        \wNDiag_52[25] , \wNDiag_52[24] , \wNDiag_52[23] , \wNDiag_52[22] , 
        \wNDiag_52[21] , \wNDiag_52[20] , \wNDiag_52[19] , \wNDiag_52[18] , 
        \wNDiag_52[17] , \wNDiag_52[16] , \wNDiag_52[15] , \wNDiag_52[14] , 
        \wNDiag_52[13] , \wNDiag_52[12] , \wNDiag_52[11] , \wNDiag_52[10] , 
        \wNDiag_52[9] , \wNDiag_52[8] , \wNDiag_52[7] , \wNDiag_52[6] , 
        \wNDiag_52[5] , \wNDiag_52[4] , \wNDiag_52[3] , \wNDiag_52[2] , 
        \wNDiag_52[1] , \wNDiag_52[0] }), .CallOut(\wCall_53[0] ), .ReturnOut(
        \wReturn_52[0] ), .ColOut({\wColumn_53[63] , \wColumn_53[62] , 
        \wColumn_53[61] , \wColumn_53[60] , \wColumn_53[59] , \wColumn_53[58] , 
        \wColumn_53[57] , \wColumn_53[56] , \wColumn_53[55] , \wColumn_53[54] , 
        \wColumn_53[53] , \wColumn_53[52] , \wColumn_53[51] , \wColumn_53[50] , 
        \wColumn_53[49] , \wColumn_53[48] , \wColumn_53[47] , \wColumn_53[46] , 
        \wColumn_53[45] , \wColumn_53[44] , \wColumn_53[43] , \wColumn_53[42] , 
        \wColumn_53[41] , \wColumn_53[40] , \wColumn_53[39] , \wColumn_53[38] , 
        \wColumn_53[37] , \wColumn_53[36] , \wColumn_53[35] , \wColumn_53[34] , 
        \wColumn_53[33] , \wColumn_53[32] , \wColumn_53[31] , \wColumn_53[30] , 
        \wColumn_53[29] , \wColumn_53[28] , \wColumn_53[27] , \wColumn_53[26] , 
        \wColumn_53[25] , \wColumn_53[24] , \wColumn_53[23] , \wColumn_53[22] , 
        \wColumn_53[21] , \wColumn_53[20] , \wColumn_53[19] , \wColumn_53[18] , 
        \wColumn_53[17] , \wColumn_53[16] , \wColumn_53[15] , \wColumn_53[14] , 
        \wColumn_53[13] , \wColumn_53[12] , \wColumn_53[11] , \wColumn_53[10] , 
        \wColumn_53[9] , \wColumn_53[8] , \wColumn_53[7] , \wColumn_53[6] , 
        \wColumn_53[5] , \wColumn_53[4] , \wColumn_53[3] , \wColumn_53[2] , 
        \wColumn_53[1] , \wColumn_53[0] }), .PDiagOut({\wPDiag_53[63] , 
        \wPDiag_53[62] , \wPDiag_53[61] , \wPDiag_53[60] , \wPDiag_53[59] , 
        \wPDiag_53[58] , \wPDiag_53[57] , \wPDiag_53[56] , \wPDiag_53[55] , 
        \wPDiag_53[54] , \wPDiag_53[53] , \wPDiag_53[52] , \wPDiag_53[51] , 
        \wPDiag_53[50] , \wPDiag_53[49] , \wPDiag_53[48] , \wPDiag_53[47] , 
        \wPDiag_53[46] , \wPDiag_53[45] , \wPDiag_53[44] , \wPDiag_53[43] , 
        \wPDiag_53[42] , \wPDiag_53[41] , \wPDiag_53[40] , \wPDiag_53[39] , 
        \wPDiag_53[38] , \wPDiag_53[37] , \wPDiag_53[36] , \wPDiag_53[35] , 
        \wPDiag_53[34] , \wPDiag_53[33] , \wPDiag_53[32] , \wPDiag_53[31] , 
        \wPDiag_53[30] , \wPDiag_53[29] , \wPDiag_53[28] , \wPDiag_53[27] , 
        \wPDiag_53[26] , \wPDiag_53[25] , \wPDiag_53[24] , \wPDiag_53[23] , 
        \wPDiag_53[22] , \wPDiag_53[21] , \wPDiag_53[20] , \wPDiag_53[19] , 
        \wPDiag_53[18] , \wPDiag_53[17] , \wPDiag_53[16] , \wPDiag_53[15] , 
        \wPDiag_53[14] , \wPDiag_53[13] , \wPDiag_53[12] , \wPDiag_53[11] , 
        \wPDiag_53[10] , \wPDiag_53[9] , \wPDiag_53[8] , \wPDiag_53[7] , 
        \wPDiag_53[6] , \wPDiag_53[5] , \wPDiag_53[4] , \wPDiag_53[3] , 
        \wPDiag_53[2] , \wPDiag_53[1] , \wPDiag_53[0] }), .NDiagOut({
        \wNDiag_53[63] , \wNDiag_53[62] , \wNDiag_53[61] , \wNDiag_53[60] , 
        \wNDiag_53[59] , \wNDiag_53[58] , \wNDiag_53[57] , \wNDiag_53[56] , 
        \wNDiag_53[55] , \wNDiag_53[54] , \wNDiag_53[53] , \wNDiag_53[52] , 
        \wNDiag_53[51] , \wNDiag_53[50] , \wNDiag_53[49] , \wNDiag_53[48] , 
        \wNDiag_53[47] , \wNDiag_53[46] , \wNDiag_53[45] , \wNDiag_53[44] , 
        \wNDiag_53[43] , \wNDiag_53[42] , \wNDiag_53[41] , \wNDiag_53[40] , 
        \wNDiag_53[39] , \wNDiag_53[38] , \wNDiag_53[37] , \wNDiag_53[36] , 
        \wNDiag_53[35] , \wNDiag_53[34] , \wNDiag_53[33] , \wNDiag_53[32] , 
        \wNDiag_53[31] , \wNDiag_53[30] , \wNDiag_53[29] , \wNDiag_53[28] , 
        \wNDiag_53[27] , \wNDiag_53[26] , \wNDiag_53[25] , \wNDiag_53[24] , 
        \wNDiag_53[23] , \wNDiag_53[22] , \wNDiag_53[21] , \wNDiag_53[20] , 
        \wNDiag_53[19] , \wNDiag_53[18] , \wNDiag_53[17] , \wNDiag_53[16] , 
        \wNDiag_53[15] , \wNDiag_53[14] , \wNDiag_53[13] , \wNDiag_53[12] , 
        \wNDiag_53[11] , \wNDiag_53[10] , \wNDiag_53[9] , \wNDiag_53[8] , 
        \wNDiag_53[7] , \wNDiag_53[6] , \wNDiag_53[5] , \wNDiag_53[4] , 
        \wNDiag_53[3] , \wNDiag_53[2] , \wNDiag_53[1] , \wNDiag_53[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_4 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_5[6] , \wScan_5[5] , \wScan_5[4] , 
        \wScan_5[3] , \wScan_5[2] , \wScan_5[1] , \wScan_5[0] }), .ScanOut({
        \wScan_4[6] , \wScan_4[5] , \wScan_4[4] , \wScan_4[3] , \wScan_4[2] , 
        \wScan_4[1] , \wScan_4[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_4[0] ), 
        .ReturnIn(\wReturn_5[0] ), .ColIn({\wColumn_4[63] , \wColumn_4[62] , 
        \wColumn_4[61] , \wColumn_4[60] , \wColumn_4[59] , \wColumn_4[58] , 
        \wColumn_4[57] , \wColumn_4[56] , \wColumn_4[55] , \wColumn_4[54] , 
        \wColumn_4[53] , \wColumn_4[52] , \wColumn_4[51] , \wColumn_4[50] , 
        \wColumn_4[49] , \wColumn_4[48] , \wColumn_4[47] , \wColumn_4[46] , 
        \wColumn_4[45] , \wColumn_4[44] , \wColumn_4[43] , \wColumn_4[42] , 
        \wColumn_4[41] , \wColumn_4[40] , \wColumn_4[39] , \wColumn_4[38] , 
        \wColumn_4[37] , \wColumn_4[36] , \wColumn_4[35] , \wColumn_4[34] , 
        \wColumn_4[33] , \wColumn_4[32] , \wColumn_4[31] , \wColumn_4[30] , 
        \wColumn_4[29] , \wColumn_4[28] , \wColumn_4[27] , \wColumn_4[26] , 
        \wColumn_4[25] , \wColumn_4[24] , \wColumn_4[23] , \wColumn_4[22] , 
        \wColumn_4[21] , \wColumn_4[20] , \wColumn_4[19] , \wColumn_4[18] , 
        \wColumn_4[17] , \wColumn_4[16] , \wColumn_4[15] , \wColumn_4[14] , 
        \wColumn_4[13] , \wColumn_4[12] , \wColumn_4[11] , \wColumn_4[10] , 
        \wColumn_4[9] , \wColumn_4[8] , \wColumn_4[7] , \wColumn_4[6] , 
        \wColumn_4[5] , \wColumn_4[4] , \wColumn_4[3] , \wColumn_4[2] , 
        \wColumn_4[1] , \wColumn_4[0] }), .PDiagIn({\wPDiag_4[63] , 
        \wPDiag_4[62] , \wPDiag_4[61] , \wPDiag_4[60] , \wPDiag_4[59] , 
        \wPDiag_4[58] , \wPDiag_4[57] , \wPDiag_4[56] , \wPDiag_4[55] , 
        \wPDiag_4[54] , \wPDiag_4[53] , \wPDiag_4[52] , \wPDiag_4[51] , 
        \wPDiag_4[50] , \wPDiag_4[49] , \wPDiag_4[48] , \wPDiag_4[47] , 
        \wPDiag_4[46] , \wPDiag_4[45] , \wPDiag_4[44] , \wPDiag_4[43] , 
        \wPDiag_4[42] , \wPDiag_4[41] , \wPDiag_4[40] , \wPDiag_4[39] , 
        \wPDiag_4[38] , \wPDiag_4[37] , \wPDiag_4[36] , \wPDiag_4[35] , 
        \wPDiag_4[34] , \wPDiag_4[33] , \wPDiag_4[32] , \wPDiag_4[31] , 
        \wPDiag_4[30] , \wPDiag_4[29] , \wPDiag_4[28] , \wPDiag_4[27] , 
        \wPDiag_4[26] , \wPDiag_4[25] , \wPDiag_4[24] , \wPDiag_4[23] , 
        \wPDiag_4[22] , \wPDiag_4[21] , \wPDiag_4[20] , \wPDiag_4[19] , 
        \wPDiag_4[18] , \wPDiag_4[17] , \wPDiag_4[16] , \wPDiag_4[15] , 
        \wPDiag_4[14] , \wPDiag_4[13] , \wPDiag_4[12] , \wPDiag_4[11] , 
        \wPDiag_4[10] , \wPDiag_4[9] , \wPDiag_4[8] , \wPDiag_4[7] , 
        \wPDiag_4[6] , \wPDiag_4[5] , \wPDiag_4[4] , \wPDiag_4[3] , 
        \wPDiag_4[2] , \wPDiag_4[1] , \wPDiag_4[0] }), .NDiagIn({
        \wNDiag_4[63] , \wNDiag_4[62] , \wNDiag_4[61] , \wNDiag_4[60] , 
        \wNDiag_4[59] , \wNDiag_4[58] , \wNDiag_4[57] , \wNDiag_4[56] , 
        \wNDiag_4[55] , \wNDiag_4[54] , \wNDiag_4[53] , \wNDiag_4[52] , 
        \wNDiag_4[51] , \wNDiag_4[50] , \wNDiag_4[49] , \wNDiag_4[48] , 
        \wNDiag_4[47] , \wNDiag_4[46] , \wNDiag_4[45] , \wNDiag_4[44] , 
        \wNDiag_4[43] , \wNDiag_4[42] , \wNDiag_4[41] , \wNDiag_4[40] , 
        \wNDiag_4[39] , \wNDiag_4[38] , \wNDiag_4[37] , \wNDiag_4[36] , 
        \wNDiag_4[35] , \wNDiag_4[34] , \wNDiag_4[33] , \wNDiag_4[32] , 
        \wNDiag_4[31] , \wNDiag_4[30] , \wNDiag_4[29] , \wNDiag_4[28] , 
        \wNDiag_4[27] , \wNDiag_4[26] , \wNDiag_4[25] , \wNDiag_4[24] , 
        \wNDiag_4[23] , \wNDiag_4[22] , \wNDiag_4[21] , \wNDiag_4[20] , 
        \wNDiag_4[19] , \wNDiag_4[18] , \wNDiag_4[17] , \wNDiag_4[16] , 
        \wNDiag_4[15] , \wNDiag_4[14] , \wNDiag_4[13] , \wNDiag_4[12] , 
        \wNDiag_4[11] , \wNDiag_4[10] , \wNDiag_4[9] , \wNDiag_4[8] , 
        \wNDiag_4[7] , \wNDiag_4[6] , \wNDiag_4[5] , \wNDiag_4[4] , 
        \wNDiag_4[3] , \wNDiag_4[2] , \wNDiag_4[1] , \wNDiag_4[0] }), 
        .CallOut(\wCall_5[0] ), .ReturnOut(\wReturn_4[0] ), .ColOut({
        \wColumn_5[63] , \wColumn_5[62] , \wColumn_5[61] , \wColumn_5[60] , 
        \wColumn_5[59] , \wColumn_5[58] , \wColumn_5[57] , \wColumn_5[56] , 
        \wColumn_5[55] , \wColumn_5[54] , \wColumn_5[53] , \wColumn_5[52] , 
        \wColumn_5[51] , \wColumn_5[50] , \wColumn_5[49] , \wColumn_5[48] , 
        \wColumn_5[47] , \wColumn_5[46] , \wColumn_5[45] , \wColumn_5[44] , 
        \wColumn_5[43] , \wColumn_5[42] , \wColumn_5[41] , \wColumn_5[40] , 
        \wColumn_5[39] , \wColumn_5[38] , \wColumn_5[37] , \wColumn_5[36] , 
        \wColumn_5[35] , \wColumn_5[34] , \wColumn_5[33] , \wColumn_5[32] , 
        \wColumn_5[31] , \wColumn_5[30] , \wColumn_5[29] , \wColumn_5[28] , 
        \wColumn_5[27] , \wColumn_5[26] , \wColumn_5[25] , \wColumn_5[24] , 
        \wColumn_5[23] , \wColumn_5[22] , \wColumn_5[21] , \wColumn_5[20] , 
        \wColumn_5[19] , \wColumn_5[18] , \wColumn_5[17] , \wColumn_5[16] , 
        \wColumn_5[15] , \wColumn_5[14] , \wColumn_5[13] , \wColumn_5[12] , 
        \wColumn_5[11] , \wColumn_5[10] , \wColumn_5[9] , \wColumn_5[8] , 
        \wColumn_5[7] , \wColumn_5[6] , \wColumn_5[5] , \wColumn_5[4] , 
        \wColumn_5[3] , \wColumn_5[2] , \wColumn_5[1] , \wColumn_5[0] }), 
        .PDiagOut({\wPDiag_5[63] , \wPDiag_5[62] , \wPDiag_5[61] , 
        \wPDiag_5[60] , \wPDiag_5[59] , \wPDiag_5[58] , \wPDiag_5[57] , 
        \wPDiag_5[56] , \wPDiag_5[55] , \wPDiag_5[54] , \wPDiag_5[53] , 
        \wPDiag_5[52] , \wPDiag_5[51] , \wPDiag_5[50] , \wPDiag_5[49] , 
        \wPDiag_5[48] , \wPDiag_5[47] , \wPDiag_5[46] , \wPDiag_5[45] , 
        \wPDiag_5[44] , \wPDiag_5[43] , \wPDiag_5[42] , \wPDiag_5[41] , 
        \wPDiag_5[40] , \wPDiag_5[39] , \wPDiag_5[38] , \wPDiag_5[37] , 
        \wPDiag_5[36] , \wPDiag_5[35] , \wPDiag_5[34] , \wPDiag_5[33] , 
        \wPDiag_5[32] , \wPDiag_5[31] , \wPDiag_5[30] , \wPDiag_5[29] , 
        \wPDiag_5[28] , \wPDiag_5[27] , \wPDiag_5[26] , \wPDiag_5[25] , 
        \wPDiag_5[24] , \wPDiag_5[23] , \wPDiag_5[22] , \wPDiag_5[21] , 
        \wPDiag_5[20] , \wPDiag_5[19] , \wPDiag_5[18] , \wPDiag_5[17] , 
        \wPDiag_5[16] , \wPDiag_5[15] , \wPDiag_5[14] , \wPDiag_5[13] , 
        \wPDiag_5[12] , \wPDiag_5[11] , \wPDiag_5[10] , \wPDiag_5[9] , 
        \wPDiag_5[8] , \wPDiag_5[7] , \wPDiag_5[6] , \wPDiag_5[5] , 
        \wPDiag_5[4] , \wPDiag_5[3] , \wPDiag_5[2] , \wPDiag_5[1] , 
        \wPDiag_5[0] }), .NDiagOut({\wNDiag_5[63] , \wNDiag_5[62] , 
        \wNDiag_5[61] , \wNDiag_5[60] , \wNDiag_5[59] , \wNDiag_5[58] , 
        \wNDiag_5[57] , \wNDiag_5[56] , \wNDiag_5[55] , \wNDiag_5[54] , 
        \wNDiag_5[53] , \wNDiag_5[52] , \wNDiag_5[51] , \wNDiag_5[50] , 
        \wNDiag_5[49] , \wNDiag_5[48] , \wNDiag_5[47] , \wNDiag_5[46] , 
        \wNDiag_5[45] , \wNDiag_5[44] , \wNDiag_5[43] , \wNDiag_5[42] , 
        \wNDiag_5[41] , \wNDiag_5[40] , \wNDiag_5[39] , \wNDiag_5[38] , 
        \wNDiag_5[37] , \wNDiag_5[36] , \wNDiag_5[35] , \wNDiag_5[34] , 
        \wNDiag_5[33] , \wNDiag_5[32] , \wNDiag_5[31] , \wNDiag_5[30] , 
        \wNDiag_5[29] , \wNDiag_5[28] , \wNDiag_5[27] , \wNDiag_5[26] , 
        \wNDiag_5[25] , \wNDiag_5[24] , \wNDiag_5[23] , \wNDiag_5[22] , 
        \wNDiag_5[21] , \wNDiag_5[20] , \wNDiag_5[19] , \wNDiag_5[18] , 
        \wNDiag_5[17] , \wNDiag_5[16] , \wNDiag_5[15] , \wNDiag_5[14] , 
        \wNDiag_5[13] , \wNDiag_5[12] , \wNDiag_5[11] , \wNDiag_5[10] , 
        \wNDiag_5[9] , \wNDiag_5[8] , \wNDiag_5[7] , \wNDiag_5[6] , 
        \wNDiag_5[5] , \wNDiag_5[4] , \wNDiag_5[3] , \wNDiag_5[2] , 
        \wNDiag_5[1] , \wNDiag_5[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_5 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_6[6] , \wScan_6[5] , \wScan_6[4] , 
        \wScan_6[3] , \wScan_6[2] , \wScan_6[1] , \wScan_6[0] }), .ScanOut({
        \wScan_5[6] , \wScan_5[5] , \wScan_5[4] , \wScan_5[3] , \wScan_5[2] , 
        \wScan_5[1] , \wScan_5[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_5[0] ), 
        .ReturnIn(\wReturn_6[0] ), .ColIn({\wColumn_5[63] , \wColumn_5[62] , 
        \wColumn_5[61] , \wColumn_5[60] , \wColumn_5[59] , \wColumn_5[58] , 
        \wColumn_5[57] , \wColumn_5[56] , \wColumn_5[55] , \wColumn_5[54] , 
        \wColumn_5[53] , \wColumn_5[52] , \wColumn_5[51] , \wColumn_5[50] , 
        \wColumn_5[49] , \wColumn_5[48] , \wColumn_5[47] , \wColumn_5[46] , 
        \wColumn_5[45] , \wColumn_5[44] , \wColumn_5[43] , \wColumn_5[42] , 
        \wColumn_5[41] , \wColumn_5[40] , \wColumn_5[39] , \wColumn_5[38] , 
        \wColumn_5[37] , \wColumn_5[36] , \wColumn_5[35] , \wColumn_5[34] , 
        \wColumn_5[33] , \wColumn_5[32] , \wColumn_5[31] , \wColumn_5[30] , 
        \wColumn_5[29] , \wColumn_5[28] , \wColumn_5[27] , \wColumn_5[26] , 
        \wColumn_5[25] , \wColumn_5[24] , \wColumn_5[23] , \wColumn_5[22] , 
        \wColumn_5[21] , \wColumn_5[20] , \wColumn_5[19] , \wColumn_5[18] , 
        \wColumn_5[17] , \wColumn_5[16] , \wColumn_5[15] , \wColumn_5[14] , 
        \wColumn_5[13] , \wColumn_5[12] , \wColumn_5[11] , \wColumn_5[10] , 
        \wColumn_5[9] , \wColumn_5[8] , \wColumn_5[7] , \wColumn_5[6] , 
        \wColumn_5[5] , \wColumn_5[4] , \wColumn_5[3] , \wColumn_5[2] , 
        \wColumn_5[1] , \wColumn_5[0] }), .PDiagIn({\wPDiag_5[63] , 
        \wPDiag_5[62] , \wPDiag_5[61] , \wPDiag_5[60] , \wPDiag_5[59] , 
        \wPDiag_5[58] , \wPDiag_5[57] , \wPDiag_5[56] , \wPDiag_5[55] , 
        \wPDiag_5[54] , \wPDiag_5[53] , \wPDiag_5[52] , \wPDiag_5[51] , 
        \wPDiag_5[50] , \wPDiag_5[49] , \wPDiag_5[48] , \wPDiag_5[47] , 
        \wPDiag_5[46] , \wPDiag_5[45] , \wPDiag_5[44] , \wPDiag_5[43] , 
        \wPDiag_5[42] , \wPDiag_5[41] , \wPDiag_5[40] , \wPDiag_5[39] , 
        \wPDiag_5[38] , \wPDiag_5[37] , \wPDiag_5[36] , \wPDiag_5[35] , 
        \wPDiag_5[34] , \wPDiag_5[33] , \wPDiag_5[32] , \wPDiag_5[31] , 
        \wPDiag_5[30] , \wPDiag_5[29] , \wPDiag_5[28] , \wPDiag_5[27] , 
        \wPDiag_5[26] , \wPDiag_5[25] , \wPDiag_5[24] , \wPDiag_5[23] , 
        \wPDiag_5[22] , \wPDiag_5[21] , \wPDiag_5[20] , \wPDiag_5[19] , 
        \wPDiag_5[18] , \wPDiag_5[17] , \wPDiag_5[16] , \wPDiag_5[15] , 
        \wPDiag_5[14] , \wPDiag_5[13] , \wPDiag_5[12] , \wPDiag_5[11] , 
        \wPDiag_5[10] , \wPDiag_5[9] , \wPDiag_5[8] , \wPDiag_5[7] , 
        \wPDiag_5[6] , \wPDiag_5[5] , \wPDiag_5[4] , \wPDiag_5[3] , 
        \wPDiag_5[2] , \wPDiag_5[1] , \wPDiag_5[0] }), .NDiagIn({
        \wNDiag_5[63] , \wNDiag_5[62] , \wNDiag_5[61] , \wNDiag_5[60] , 
        \wNDiag_5[59] , \wNDiag_5[58] , \wNDiag_5[57] , \wNDiag_5[56] , 
        \wNDiag_5[55] , \wNDiag_5[54] , \wNDiag_5[53] , \wNDiag_5[52] , 
        \wNDiag_5[51] , \wNDiag_5[50] , \wNDiag_5[49] , \wNDiag_5[48] , 
        \wNDiag_5[47] , \wNDiag_5[46] , \wNDiag_5[45] , \wNDiag_5[44] , 
        \wNDiag_5[43] , \wNDiag_5[42] , \wNDiag_5[41] , \wNDiag_5[40] , 
        \wNDiag_5[39] , \wNDiag_5[38] , \wNDiag_5[37] , \wNDiag_5[36] , 
        \wNDiag_5[35] , \wNDiag_5[34] , \wNDiag_5[33] , \wNDiag_5[32] , 
        \wNDiag_5[31] , \wNDiag_5[30] , \wNDiag_5[29] , \wNDiag_5[28] , 
        \wNDiag_5[27] , \wNDiag_5[26] , \wNDiag_5[25] , \wNDiag_5[24] , 
        \wNDiag_5[23] , \wNDiag_5[22] , \wNDiag_5[21] , \wNDiag_5[20] , 
        \wNDiag_5[19] , \wNDiag_5[18] , \wNDiag_5[17] , \wNDiag_5[16] , 
        \wNDiag_5[15] , \wNDiag_5[14] , \wNDiag_5[13] , \wNDiag_5[12] , 
        \wNDiag_5[11] , \wNDiag_5[10] , \wNDiag_5[9] , \wNDiag_5[8] , 
        \wNDiag_5[7] , \wNDiag_5[6] , \wNDiag_5[5] , \wNDiag_5[4] , 
        \wNDiag_5[3] , \wNDiag_5[2] , \wNDiag_5[1] , \wNDiag_5[0] }), 
        .CallOut(\wCall_6[0] ), .ReturnOut(\wReturn_5[0] ), .ColOut({
        \wColumn_6[63] , \wColumn_6[62] , \wColumn_6[61] , \wColumn_6[60] , 
        \wColumn_6[59] , \wColumn_6[58] , \wColumn_6[57] , \wColumn_6[56] , 
        \wColumn_6[55] , \wColumn_6[54] , \wColumn_6[53] , \wColumn_6[52] , 
        \wColumn_6[51] , \wColumn_6[50] , \wColumn_6[49] , \wColumn_6[48] , 
        \wColumn_6[47] , \wColumn_6[46] , \wColumn_6[45] , \wColumn_6[44] , 
        \wColumn_6[43] , \wColumn_6[42] , \wColumn_6[41] , \wColumn_6[40] , 
        \wColumn_6[39] , \wColumn_6[38] , \wColumn_6[37] , \wColumn_6[36] , 
        \wColumn_6[35] , \wColumn_6[34] , \wColumn_6[33] , \wColumn_6[32] , 
        \wColumn_6[31] , \wColumn_6[30] , \wColumn_6[29] , \wColumn_6[28] , 
        \wColumn_6[27] , \wColumn_6[26] , \wColumn_6[25] , \wColumn_6[24] , 
        \wColumn_6[23] , \wColumn_6[22] , \wColumn_6[21] , \wColumn_6[20] , 
        \wColumn_6[19] , \wColumn_6[18] , \wColumn_6[17] , \wColumn_6[16] , 
        \wColumn_6[15] , \wColumn_6[14] , \wColumn_6[13] , \wColumn_6[12] , 
        \wColumn_6[11] , \wColumn_6[10] , \wColumn_6[9] , \wColumn_6[8] , 
        \wColumn_6[7] , \wColumn_6[6] , \wColumn_6[5] , \wColumn_6[4] , 
        \wColumn_6[3] , \wColumn_6[2] , \wColumn_6[1] , \wColumn_6[0] }), 
        .PDiagOut({\wPDiag_6[63] , \wPDiag_6[62] , \wPDiag_6[61] , 
        \wPDiag_6[60] , \wPDiag_6[59] , \wPDiag_6[58] , \wPDiag_6[57] , 
        \wPDiag_6[56] , \wPDiag_6[55] , \wPDiag_6[54] , \wPDiag_6[53] , 
        \wPDiag_6[52] , \wPDiag_6[51] , \wPDiag_6[50] , \wPDiag_6[49] , 
        \wPDiag_6[48] , \wPDiag_6[47] , \wPDiag_6[46] , \wPDiag_6[45] , 
        \wPDiag_6[44] , \wPDiag_6[43] , \wPDiag_6[42] , \wPDiag_6[41] , 
        \wPDiag_6[40] , \wPDiag_6[39] , \wPDiag_6[38] , \wPDiag_6[37] , 
        \wPDiag_6[36] , \wPDiag_6[35] , \wPDiag_6[34] , \wPDiag_6[33] , 
        \wPDiag_6[32] , \wPDiag_6[31] , \wPDiag_6[30] , \wPDiag_6[29] , 
        \wPDiag_6[28] , \wPDiag_6[27] , \wPDiag_6[26] , \wPDiag_6[25] , 
        \wPDiag_6[24] , \wPDiag_6[23] , \wPDiag_6[22] , \wPDiag_6[21] , 
        \wPDiag_6[20] , \wPDiag_6[19] , \wPDiag_6[18] , \wPDiag_6[17] , 
        \wPDiag_6[16] , \wPDiag_6[15] , \wPDiag_6[14] , \wPDiag_6[13] , 
        \wPDiag_6[12] , \wPDiag_6[11] , \wPDiag_6[10] , \wPDiag_6[9] , 
        \wPDiag_6[8] , \wPDiag_6[7] , \wPDiag_6[6] , \wPDiag_6[5] , 
        \wPDiag_6[4] , \wPDiag_6[3] , \wPDiag_6[2] , \wPDiag_6[1] , 
        \wPDiag_6[0] }), .NDiagOut({\wNDiag_6[63] , \wNDiag_6[62] , 
        \wNDiag_6[61] , \wNDiag_6[60] , \wNDiag_6[59] , \wNDiag_6[58] , 
        \wNDiag_6[57] , \wNDiag_6[56] , \wNDiag_6[55] , \wNDiag_6[54] , 
        \wNDiag_6[53] , \wNDiag_6[52] , \wNDiag_6[51] , \wNDiag_6[50] , 
        \wNDiag_6[49] , \wNDiag_6[48] , \wNDiag_6[47] , \wNDiag_6[46] , 
        \wNDiag_6[45] , \wNDiag_6[44] , \wNDiag_6[43] , \wNDiag_6[42] , 
        \wNDiag_6[41] , \wNDiag_6[40] , \wNDiag_6[39] , \wNDiag_6[38] , 
        \wNDiag_6[37] , \wNDiag_6[36] , \wNDiag_6[35] , \wNDiag_6[34] , 
        \wNDiag_6[33] , \wNDiag_6[32] , \wNDiag_6[31] , \wNDiag_6[30] , 
        \wNDiag_6[29] , \wNDiag_6[28] , \wNDiag_6[27] , \wNDiag_6[26] , 
        \wNDiag_6[25] , \wNDiag_6[24] , \wNDiag_6[23] , \wNDiag_6[22] , 
        \wNDiag_6[21] , \wNDiag_6[20] , \wNDiag_6[19] , \wNDiag_6[18] , 
        \wNDiag_6[17] , \wNDiag_6[16] , \wNDiag_6[15] , \wNDiag_6[14] , 
        \wNDiag_6[13] , \wNDiag_6[12] , \wNDiag_6[11] , \wNDiag_6[10] , 
        \wNDiag_6[9] , \wNDiag_6[8] , \wNDiag_6[7] , \wNDiag_6[6] , 
        \wNDiag_6[5] , \wNDiag_6[4] , \wNDiag_6[3] , \wNDiag_6[2] , 
        \wNDiag_6[1] , \wNDiag_6[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_15 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_16[6] , \wScan_16[5] , \wScan_16[4] , 
        \wScan_16[3] , \wScan_16[2] , \wScan_16[1] , \wScan_16[0] }), 
        .ScanOut({\wScan_15[6] , \wScan_15[5] , \wScan_15[4] , \wScan_15[3] , 
        \wScan_15[2] , \wScan_15[1] , \wScan_15[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_15[0] ), .ReturnIn(\wReturn_16[0] ), .ColIn({
        \wColumn_15[63] , \wColumn_15[62] , \wColumn_15[61] , \wColumn_15[60] , 
        \wColumn_15[59] , \wColumn_15[58] , \wColumn_15[57] , \wColumn_15[56] , 
        \wColumn_15[55] , \wColumn_15[54] , \wColumn_15[53] , \wColumn_15[52] , 
        \wColumn_15[51] , \wColumn_15[50] , \wColumn_15[49] , \wColumn_15[48] , 
        \wColumn_15[47] , \wColumn_15[46] , \wColumn_15[45] , \wColumn_15[44] , 
        \wColumn_15[43] , \wColumn_15[42] , \wColumn_15[41] , \wColumn_15[40] , 
        \wColumn_15[39] , \wColumn_15[38] , \wColumn_15[37] , \wColumn_15[36] , 
        \wColumn_15[35] , \wColumn_15[34] , \wColumn_15[33] , \wColumn_15[32] , 
        \wColumn_15[31] , \wColumn_15[30] , \wColumn_15[29] , \wColumn_15[28] , 
        \wColumn_15[27] , \wColumn_15[26] , \wColumn_15[25] , \wColumn_15[24] , 
        \wColumn_15[23] , \wColumn_15[22] , \wColumn_15[21] , \wColumn_15[20] , 
        \wColumn_15[19] , \wColumn_15[18] , \wColumn_15[17] , \wColumn_15[16] , 
        \wColumn_15[15] , \wColumn_15[14] , \wColumn_15[13] , \wColumn_15[12] , 
        \wColumn_15[11] , \wColumn_15[10] , \wColumn_15[9] , \wColumn_15[8] , 
        \wColumn_15[7] , \wColumn_15[6] , \wColumn_15[5] , \wColumn_15[4] , 
        \wColumn_15[3] , \wColumn_15[2] , \wColumn_15[1] , \wColumn_15[0] }), 
        .PDiagIn({\wPDiag_15[63] , \wPDiag_15[62] , \wPDiag_15[61] , 
        \wPDiag_15[60] , \wPDiag_15[59] , \wPDiag_15[58] , \wPDiag_15[57] , 
        \wPDiag_15[56] , \wPDiag_15[55] , \wPDiag_15[54] , \wPDiag_15[53] , 
        \wPDiag_15[52] , \wPDiag_15[51] , \wPDiag_15[50] , \wPDiag_15[49] , 
        \wPDiag_15[48] , \wPDiag_15[47] , \wPDiag_15[46] , \wPDiag_15[45] , 
        \wPDiag_15[44] , \wPDiag_15[43] , \wPDiag_15[42] , \wPDiag_15[41] , 
        \wPDiag_15[40] , \wPDiag_15[39] , \wPDiag_15[38] , \wPDiag_15[37] , 
        \wPDiag_15[36] , \wPDiag_15[35] , \wPDiag_15[34] , \wPDiag_15[33] , 
        \wPDiag_15[32] , \wPDiag_15[31] , \wPDiag_15[30] , \wPDiag_15[29] , 
        \wPDiag_15[28] , \wPDiag_15[27] , \wPDiag_15[26] , \wPDiag_15[25] , 
        \wPDiag_15[24] , \wPDiag_15[23] , \wPDiag_15[22] , \wPDiag_15[21] , 
        \wPDiag_15[20] , \wPDiag_15[19] , \wPDiag_15[18] , \wPDiag_15[17] , 
        \wPDiag_15[16] , \wPDiag_15[15] , \wPDiag_15[14] , \wPDiag_15[13] , 
        \wPDiag_15[12] , \wPDiag_15[11] , \wPDiag_15[10] , \wPDiag_15[9] , 
        \wPDiag_15[8] , \wPDiag_15[7] , \wPDiag_15[6] , \wPDiag_15[5] , 
        \wPDiag_15[4] , \wPDiag_15[3] , \wPDiag_15[2] , \wPDiag_15[1] , 
        \wPDiag_15[0] }), .NDiagIn({\wNDiag_15[63] , \wNDiag_15[62] , 
        \wNDiag_15[61] , \wNDiag_15[60] , \wNDiag_15[59] , \wNDiag_15[58] , 
        \wNDiag_15[57] , \wNDiag_15[56] , \wNDiag_15[55] , \wNDiag_15[54] , 
        \wNDiag_15[53] , \wNDiag_15[52] , \wNDiag_15[51] , \wNDiag_15[50] , 
        \wNDiag_15[49] , \wNDiag_15[48] , \wNDiag_15[47] , \wNDiag_15[46] , 
        \wNDiag_15[45] , \wNDiag_15[44] , \wNDiag_15[43] , \wNDiag_15[42] , 
        \wNDiag_15[41] , \wNDiag_15[40] , \wNDiag_15[39] , \wNDiag_15[38] , 
        \wNDiag_15[37] , \wNDiag_15[36] , \wNDiag_15[35] , \wNDiag_15[34] , 
        \wNDiag_15[33] , \wNDiag_15[32] , \wNDiag_15[31] , \wNDiag_15[30] , 
        \wNDiag_15[29] , \wNDiag_15[28] , \wNDiag_15[27] , \wNDiag_15[26] , 
        \wNDiag_15[25] , \wNDiag_15[24] , \wNDiag_15[23] , \wNDiag_15[22] , 
        \wNDiag_15[21] , \wNDiag_15[20] , \wNDiag_15[19] , \wNDiag_15[18] , 
        \wNDiag_15[17] , \wNDiag_15[16] , \wNDiag_15[15] , \wNDiag_15[14] , 
        \wNDiag_15[13] , \wNDiag_15[12] , \wNDiag_15[11] , \wNDiag_15[10] , 
        \wNDiag_15[9] , \wNDiag_15[8] , \wNDiag_15[7] , \wNDiag_15[6] , 
        \wNDiag_15[5] , \wNDiag_15[4] , \wNDiag_15[3] , \wNDiag_15[2] , 
        \wNDiag_15[1] , \wNDiag_15[0] }), .CallOut(\wCall_16[0] ), .ReturnOut(
        \wReturn_15[0] ), .ColOut({\wColumn_16[63] , \wColumn_16[62] , 
        \wColumn_16[61] , \wColumn_16[60] , \wColumn_16[59] , \wColumn_16[58] , 
        \wColumn_16[57] , \wColumn_16[56] , \wColumn_16[55] , \wColumn_16[54] , 
        \wColumn_16[53] , \wColumn_16[52] , \wColumn_16[51] , \wColumn_16[50] , 
        \wColumn_16[49] , \wColumn_16[48] , \wColumn_16[47] , \wColumn_16[46] , 
        \wColumn_16[45] , \wColumn_16[44] , \wColumn_16[43] , \wColumn_16[42] , 
        \wColumn_16[41] , \wColumn_16[40] , \wColumn_16[39] , \wColumn_16[38] , 
        \wColumn_16[37] , \wColumn_16[36] , \wColumn_16[35] , \wColumn_16[34] , 
        \wColumn_16[33] , \wColumn_16[32] , \wColumn_16[31] , \wColumn_16[30] , 
        \wColumn_16[29] , \wColumn_16[28] , \wColumn_16[27] , \wColumn_16[26] , 
        \wColumn_16[25] , \wColumn_16[24] , \wColumn_16[23] , \wColumn_16[22] , 
        \wColumn_16[21] , \wColumn_16[20] , \wColumn_16[19] , \wColumn_16[18] , 
        \wColumn_16[17] , \wColumn_16[16] , \wColumn_16[15] , \wColumn_16[14] , 
        \wColumn_16[13] , \wColumn_16[12] , \wColumn_16[11] , \wColumn_16[10] , 
        \wColumn_16[9] , \wColumn_16[8] , \wColumn_16[7] , \wColumn_16[6] , 
        \wColumn_16[5] , \wColumn_16[4] , \wColumn_16[3] , \wColumn_16[2] , 
        \wColumn_16[1] , \wColumn_16[0] }), .PDiagOut({\wPDiag_16[63] , 
        \wPDiag_16[62] , \wPDiag_16[61] , \wPDiag_16[60] , \wPDiag_16[59] , 
        \wPDiag_16[58] , \wPDiag_16[57] , \wPDiag_16[56] , \wPDiag_16[55] , 
        \wPDiag_16[54] , \wPDiag_16[53] , \wPDiag_16[52] , \wPDiag_16[51] , 
        \wPDiag_16[50] , \wPDiag_16[49] , \wPDiag_16[48] , \wPDiag_16[47] , 
        \wPDiag_16[46] , \wPDiag_16[45] , \wPDiag_16[44] , \wPDiag_16[43] , 
        \wPDiag_16[42] , \wPDiag_16[41] , \wPDiag_16[40] , \wPDiag_16[39] , 
        \wPDiag_16[38] , \wPDiag_16[37] , \wPDiag_16[36] , \wPDiag_16[35] , 
        \wPDiag_16[34] , \wPDiag_16[33] , \wPDiag_16[32] , \wPDiag_16[31] , 
        \wPDiag_16[30] , \wPDiag_16[29] , \wPDiag_16[28] , \wPDiag_16[27] , 
        \wPDiag_16[26] , \wPDiag_16[25] , \wPDiag_16[24] , \wPDiag_16[23] , 
        \wPDiag_16[22] , \wPDiag_16[21] , \wPDiag_16[20] , \wPDiag_16[19] , 
        \wPDiag_16[18] , \wPDiag_16[17] , \wPDiag_16[16] , \wPDiag_16[15] , 
        \wPDiag_16[14] , \wPDiag_16[13] , \wPDiag_16[12] , \wPDiag_16[11] , 
        \wPDiag_16[10] , \wPDiag_16[9] , \wPDiag_16[8] , \wPDiag_16[7] , 
        \wPDiag_16[6] , \wPDiag_16[5] , \wPDiag_16[4] , \wPDiag_16[3] , 
        \wPDiag_16[2] , \wPDiag_16[1] , \wPDiag_16[0] }), .NDiagOut({
        \wNDiag_16[63] , \wNDiag_16[62] , \wNDiag_16[61] , \wNDiag_16[60] , 
        \wNDiag_16[59] , \wNDiag_16[58] , \wNDiag_16[57] , \wNDiag_16[56] , 
        \wNDiag_16[55] , \wNDiag_16[54] , \wNDiag_16[53] , \wNDiag_16[52] , 
        \wNDiag_16[51] , \wNDiag_16[50] , \wNDiag_16[49] , \wNDiag_16[48] , 
        \wNDiag_16[47] , \wNDiag_16[46] , \wNDiag_16[45] , \wNDiag_16[44] , 
        \wNDiag_16[43] , \wNDiag_16[42] , \wNDiag_16[41] , \wNDiag_16[40] , 
        \wNDiag_16[39] , \wNDiag_16[38] , \wNDiag_16[37] , \wNDiag_16[36] , 
        \wNDiag_16[35] , \wNDiag_16[34] , \wNDiag_16[33] , \wNDiag_16[32] , 
        \wNDiag_16[31] , \wNDiag_16[30] , \wNDiag_16[29] , \wNDiag_16[28] , 
        \wNDiag_16[27] , \wNDiag_16[26] , \wNDiag_16[25] , \wNDiag_16[24] , 
        \wNDiag_16[23] , \wNDiag_16[22] , \wNDiag_16[21] , \wNDiag_16[20] , 
        \wNDiag_16[19] , \wNDiag_16[18] , \wNDiag_16[17] , \wNDiag_16[16] , 
        \wNDiag_16[15] , \wNDiag_16[14] , \wNDiag_16[13] , \wNDiag_16[12] , 
        \wNDiag_16[11] , \wNDiag_16[10] , \wNDiag_16[9] , \wNDiag_16[8] , 
        \wNDiag_16[7] , \wNDiag_16[6] , \wNDiag_16[5] , \wNDiag_16[4] , 
        \wNDiag_16[3] , \wNDiag_16[2] , \wNDiag_16[1] , \wNDiag_16[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_20 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_21[6] , \wScan_21[5] , \wScan_21[4] , 
        \wScan_21[3] , \wScan_21[2] , \wScan_21[1] , \wScan_21[0] }), 
        .ScanOut({\wScan_20[6] , \wScan_20[5] , \wScan_20[4] , \wScan_20[3] , 
        \wScan_20[2] , \wScan_20[1] , \wScan_20[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_20[0] ), .ReturnIn(\wReturn_21[0] ), .ColIn({
        \wColumn_20[63] , \wColumn_20[62] , \wColumn_20[61] , \wColumn_20[60] , 
        \wColumn_20[59] , \wColumn_20[58] , \wColumn_20[57] , \wColumn_20[56] , 
        \wColumn_20[55] , \wColumn_20[54] , \wColumn_20[53] , \wColumn_20[52] , 
        \wColumn_20[51] , \wColumn_20[50] , \wColumn_20[49] , \wColumn_20[48] , 
        \wColumn_20[47] , \wColumn_20[46] , \wColumn_20[45] , \wColumn_20[44] , 
        \wColumn_20[43] , \wColumn_20[42] , \wColumn_20[41] , \wColumn_20[40] , 
        \wColumn_20[39] , \wColumn_20[38] , \wColumn_20[37] , \wColumn_20[36] , 
        \wColumn_20[35] , \wColumn_20[34] , \wColumn_20[33] , \wColumn_20[32] , 
        \wColumn_20[31] , \wColumn_20[30] , \wColumn_20[29] , \wColumn_20[28] , 
        \wColumn_20[27] , \wColumn_20[26] , \wColumn_20[25] , \wColumn_20[24] , 
        \wColumn_20[23] , \wColumn_20[22] , \wColumn_20[21] , \wColumn_20[20] , 
        \wColumn_20[19] , \wColumn_20[18] , \wColumn_20[17] , \wColumn_20[16] , 
        \wColumn_20[15] , \wColumn_20[14] , \wColumn_20[13] , \wColumn_20[12] , 
        \wColumn_20[11] , \wColumn_20[10] , \wColumn_20[9] , \wColumn_20[8] , 
        \wColumn_20[7] , \wColumn_20[6] , \wColumn_20[5] , \wColumn_20[4] , 
        \wColumn_20[3] , \wColumn_20[2] , \wColumn_20[1] , \wColumn_20[0] }), 
        .PDiagIn({\wPDiag_20[63] , \wPDiag_20[62] , \wPDiag_20[61] , 
        \wPDiag_20[60] , \wPDiag_20[59] , \wPDiag_20[58] , \wPDiag_20[57] , 
        \wPDiag_20[56] , \wPDiag_20[55] , \wPDiag_20[54] , \wPDiag_20[53] , 
        \wPDiag_20[52] , \wPDiag_20[51] , \wPDiag_20[50] , \wPDiag_20[49] , 
        \wPDiag_20[48] , \wPDiag_20[47] , \wPDiag_20[46] , \wPDiag_20[45] , 
        \wPDiag_20[44] , \wPDiag_20[43] , \wPDiag_20[42] , \wPDiag_20[41] , 
        \wPDiag_20[40] , \wPDiag_20[39] , \wPDiag_20[38] , \wPDiag_20[37] , 
        \wPDiag_20[36] , \wPDiag_20[35] , \wPDiag_20[34] , \wPDiag_20[33] , 
        \wPDiag_20[32] , \wPDiag_20[31] , \wPDiag_20[30] , \wPDiag_20[29] , 
        \wPDiag_20[28] , \wPDiag_20[27] , \wPDiag_20[26] , \wPDiag_20[25] , 
        \wPDiag_20[24] , \wPDiag_20[23] , \wPDiag_20[22] , \wPDiag_20[21] , 
        \wPDiag_20[20] , \wPDiag_20[19] , \wPDiag_20[18] , \wPDiag_20[17] , 
        \wPDiag_20[16] , \wPDiag_20[15] , \wPDiag_20[14] , \wPDiag_20[13] , 
        \wPDiag_20[12] , \wPDiag_20[11] , \wPDiag_20[10] , \wPDiag_20[9] , 
        \wPDiag_20[8] , \wPDiag_20[7] , \wPDiag_20[6] , \wPDiag_20[5] , 
        \wPDiag_20[4] , \wPDiag_20[3] , \wPDiag_20[2] , \wPDiag_20[1] , 
        \wPDiag_20[0] }), .NDiagIn({\wNDiag_20[63] , \wNDiag_20[62] , 
        \wNDiag_20[61] , \wNDiag_20[60] , \wNDiag_20[59] , \wNDiag_20[58] , 
        \wNDiag_20[57] , \wNDiag_20[56] , \wNDiag_20[55] , \wNDiag_20[54] , 
        \wNDiag_20[53] , \wNDiag_20[52] , \wNDiag_20[51] , \wNDiag_20[50] , 
        \wNDiag_20[49] , \wNDiag_20[48] , \wNDiag_20[47] , \wNDiag_20[46] , 
        \wNDiag_20[45] , \wNDiag_20[44] , \wNDiag_20[43] , \wNDiag_20[42] , 
        \wNDiag_20[41] , \wNDiag_20[40] , \wNDiag_20[39] , \wNDiag_20[38] , 
        \wNDiag_20[37] , \wNDiag_20[36] , \wNDiag_20[35] , \wNDiag_20[34] , 
        \wNDiag_20[33] , \wNDiag_20[32] , \wNDiag_20[31] , \wNDiag_20[30] , 
        \wNDiag_20[29] , \wNDiag_20[28] , \wNDiag_20[27] , \wNDiag_20[26] , 
        \wNDiag_20[25] , \wNDiag_20[24] , \wNDiag_20[23] , \wNDiag_20[22] , 
        \wNDiag_20[21] , \wNDiag_20[20] , \wNDiag_20[19] , \wNDiag_20[18] , 
        \wNDiag_20[17] , \wNDiag_20[16] , \wNDiag_20[15] , \wNDiag_20[14] , 
        \wNDiag_20[13] , \wNDiag_20[12] , \wNDiag_20[11] , \wNDiag_20[10] , 
        \wNDiag_20[9] , \wNDiag_20[8] , \wNDiag_20[7] , \wNDiag_20[6] , 
        \wNDiag_20[5] , \wNDiag_20[4] , \wNDiag_20[3] , \wNDiag_20[2] , 
        \wNDiag_20[1] , \wNDiag_20[0] }), .CallOut(\wCall_21[0] ), .ReturnOut(
        \wReturn_20[0] ), .ColOut({\wColumn_21[63] , \wColumn_21[62] , 
        \wColumn_21[61] , \wColumn_21[60] , \wColumn_21[59] , \wColumn_21[58] , 
        \wColumn_21[57] , \wColumn_21[56] , \wColumn_21[55] , \wColumn_21[54] , 
        \wColumn_21[53] , \wColumn_21[52] , \wColumn_21[51] , \wColumn_21[50] , 
        \wColumn_21[49] , \wColumn_21[48] , \wColumn_21[47] , \wColumn_21[46] , 
        \wColumn_21[45] , \wColumn_21[44] , \wColumn_21[43] , \wColumn_21[42] , 
        \wColumn_21[41] , \wColumn_21[40] , \wColumn_21[39] , \wColumn_21[38] , 
        \wColumn_21[37] , \wColumn_21[36] , \wColumn_21[35] , \wColumn_21[34] , 
        \wColumn_21[33] , \wColumn_21[32] , \wColumn_21[31] , \wColumn_21[30] , 
        \wColumn_21[29] , \wColumn_21[28] , \wColumn_21[27] , \wColumn_21[26] , 
        \wColumn_21[25] , \wColumn_21[24] , \wColumn_21[23] , \wColumn_21[22] , 
        \wColumn_21[21] , \wColumn_21[20] , \wColumn_21[19] , \wColumn_21[18] , 
        \wColumn_21[17] , \wColumn_21[16] , \wColumn_21[15] , \wColumn_21[14] , 
        \wColumn_21[13] , \wColumn_21[12] , \wColumn_21[11] , \wColumn_21[10] , 
        \wColumn_21[9] , \wColumn_21[8] , \wColumn_21[7] , \wColumn_21[6] , 
        \wColumn_21[5] , \wColumn_21[4] , \wColumn_21[3] , \wColumn_21[2] , 
        \wColumn_21[1] , \wColumn_21[0] }), .PDiagOut({\wPDiag_21[63] , 
        \wPDiag_21[62] , \wPDiag_21[61] , \wPDiag_21[60] , \wPDiag_21[59] , 
        \wPDiag_21[58] , \wPDiag_21[57] , \wPDiag_21[56] , \wPDiag_21[55] , 
        \wPDiag_21[54] , \wPDiag_21[53] , \wPDiag_21[52] , \wPDiag_21[51] , 
        \wPDiag_21[50] , \wPDiag_21[49] , \wPDiag_21[48] , \wPDiag_21[47] , 
        \wPDiag_21[46] , \wPDiag_21[45] , \wPDiag_21[44] , \wPDiag_21[43] , 
        \wPDiag_21[42] , \wPDiag_21[41] , \wPDiag_21[40] , \wPDiag_21[39] , 
        \wPDiag_21[38] , \wPDiag_21[37] , \wPDiag_21[36] , \wPDiag_21[35] , 
        \wPDiag_21[34] , \wPDiag_21[33] , \wPDiag_21[32] , \wPDiag_21[31] , 
        \wPDiag_21[30] , \wPDiag_21[29] , \wPDiag_21[28] , \wPDiag_21[27] , 
        \wPDiag_21[26] , \wPDiag_21[25] , \wPDiag_21[24] , \wPDiag_21[23] , 
        \wPDiag_21[22] , \wPDiag_21[21] , \wPDiag_21[20] , \wPDiag_21[19] , 
        \wPDiag_21[18] , \wPDiag_21[17] , \wPDiag_21[16] , \wPDiag_21[15] , 
        \wPDiag_21[14] , \wPDiag_21[13] , \wPDiag_21[12] , \wPDiag_21[11] , 
        \wPDiag_21[10] , \wPDiag_21[9] , \wPDiag_21[8] , \wPDiag_21[7] , 
        \wPDiag_21[6] , \wPDiag_21[5] , \wPDiag_21[4] , \wPDiag_21[3] , 
        \wPDiag_21[2] , \wPDiag_21[1] , \wPDiag_21[0] }), .NDiagOut({
        \wNDiag_21[63] , \wNDiag_21[62] , \wNDiag_21[61] , \wNDiag_21[60] , 
        \wNDiag_21[59] , \wNDiag_21[58] , \wNDiag_21[57] , \wNDiag_21[56] , 
        \wNDiag_21[55] , \wNDiag_21[54] , \wNDiag_21[53] , \wNDiag_21[52] , 
        \wNDiag_21[51] , \wNDiag_21[50] , \wNDiag_21[49] , \wNDiag_21[48] , 
        \wNDiag_21[47] , \wNDiag_21[46] , \wNDiag_21[45] , \wNDiag_21[44] , 
        \wNDiag_21[43] , \wNDiag_21[42] , \wNDiag_21[41] , \wNDiag_21[40] , 
        \wNDiag_21[39] , \wNDiag_21[38] , \wNDiag_21[37] , \wNDiag_21[36] , 
        \wNDiag_21[35] , \wNDiag_21[34] , \wNDiag_21[33] , \wNDiag_21[32] , 
        \wNDiag_21[31] , \wNDiag_21[30] , \wNDiag_21[29] , \wNDiag_21[28] , 
        \wNDiag_21[27] , \wNDiag_21[26] , \wNDiag_21[25] , \wNDiag_21[24] , 
        \wNDiag_21[23] , \wNDiag_21[22] , \wNDiag_21[21] , \wNDiag_21[20] , 
        \wNDiag_21[19] , \wNDiag_21[18] , \wNDiag_21[17] , \wNDiag_21[16] , 
        \wNDiag_21[15] , \wNDiag_21[14] , \wNDiag_21[13] , \wNDiag_21[12] , 
        \wNDiag_21[11] , \wNDiag_21[10] , \wNDiag_21[9] , \wNDiag_21[8] , 
        \wNDiag_21[7] , \wNDiag_21[6] , \wNDiag_21[5] , \wNDiag_21[4] , 
        \wNDiag_21[3] , \wNDiag_21[2] , \wNDiag_21[1] , \wNDiag_21[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_55 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_56[6] , \wScan_56[5] , \wScan_56[4] , 
        \wScan_56[3] , \wScan_56[2] , \wScan_56[1] , \wScan_56[0] }), 
        .ScanOut({\wScan_55[6] , \wScan_55[5] , \wScan_55[4] , \wScan_55[3] , 
        \wScan_55[2] , \wScan_55[1] , \wScan_55[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_55[0] ), .ReturnIn(\wReturn_56[0] ), .ColIn({
        \wColumn_55[63] , \wColumn_55[62] , \wColumn_55[61] , \wColumn_55[60] , 
        \wColumn_55[59] , \wColumn_55[58] , \wColumn_55[57] , \wColumn_55[56] , 
        \wColumn_55[55] , \wColumn_55[54] , \wColumn_55[53] , \wColumn_55[52] , 
        \wColumn_55[51] , \wColumn_55[50] , \wColumn_55[49] , \wColumn_55[48] , 
        \wColumn_55[47] , \wColumn_55[46] , \wColumn_55[45] , \wColumn_55[44] , 
        \wColumn_55[43] , \wColumn_55[42] , \wColumn_55[41] , \wColumn_55[40] , 
        \wColumn_55[39] , \wColumn_55[38] , \wColumn_55[37] , \wColumn_55[36] , 
        \wColumn_55[35] , \wColumn_55[34] , \wColumn_55[33] , \wColumn_55[32] , 
        \wColumn_55[31] , \wColumn_55[30] , \wColumn_55[29] , \wColumn_55[28] , 
        \wColumn_55[27] , \wColumn_55[26] , \wColumn_55[25] , \wColumn_55[24] , 
        \wColumn_55[23] , \wColumn_55[22] , \wColumn_55[21] , \wColumn_55[20] , 
        \wColumn_55[19] , \wColumn_55[18] , \wColumn_55[17] , \wColumn_55[16] , 
        \wColumn_55[15] , \wColumn_55[14] , \wColumn_55[13] , \wColumn_55[12] , 
        \wColumn_55[11] , \wColumn_55[10] , \wColumn_55[9] , \wColumn_55[8] , 
        \wColumn_55[7] , \wColumn_55[6] , \wColumn_55[5] , \wColumn_55[4] , 
        \wColumn_55[3] , \wColumn_55[2] , \wColumn_55[1] , \wColumn_55[0] }), 
        .PDiagIn({\wPDiag_55[63] , \wPDiag_55[62] , \wPDiag_55[61] , 
        \wPDiag_55[60] , \wPDiag_55[59] , \wPDiag_55[58] , \wPDiag_55[57] , 
        \wPDiag_55[56] , \wPDiag_55[55] , \wPDiag_55[54] , \wPDiag_55[53] , 
        \wPDiag_55[52] , \wPDiag_55[51] , \wPDiag_55[50] , \wPDiag_55[49] , 
        \wPDiag_55[48] , \wPDiag_55[47] , \wPDiag_55[46] , \wPDiag_55[45] , 
        \wPDiag_55[44] , \wPDiag_55[43] , \wPDiag_55[42] , \wPDiag_55[41] , 
        \wPDiag_55[40] , \wPDiag_55[39] , \wPDiag_55[38] , \wPDiag_55[37] , 
        \wPDiag_55[36] , \wPDiag_55[35] , \wPDiag_55[34] , \wPDiag_55[33] , 
        \wPDiag_55[32] , \wPDiag_55[31] , \wPDiag_55[30] , \wPDiag_55[29] , 
        \wPDiag_55[28] , \wPDiag_55[27] , \wPDiag_55[26] , \wPDiag_55[25] , 
        \wPDiag_55[24] , \wPDiag_55[23] , \wPDiag_55[22] , \wPDiag_55[21] , 
        \wPDiag_55[20] , \wPDiag_55[19] , \wPDiag_55[18] , \wPDiag_55[17] , 
        \wPDiag_55[16] , \wPDiag_55[15] , \wPDiag_55[14] , \wPDiag_55[13] , 
        \wPDiag_55[12] , \wPDiag_55[11] , \wPDiag_55[10] , \wPDiag_55[9] , 
        \wPDiag_55[8] , \wPDiag_55[7] , \wPDiag_55[6] , \wPDiag_55[5] , 
        \wPDiag_55[4] , \wPDiag_55[3] , \wPDiag_55[2] , \wPDiag_55[1] , 
        \wPDiag_55[0] }), .NDiagIn({\wNDiag_55[63] , \wNDiag_55[62] , 
        \wNDiag_55[61] , \wNDiag_55[60] , \wNDiag_55[59] , \wNDiag_55[58] , 
        \wNDiag_55[57] , \wNDiag_55[56] , \wNDiag_55[55] , \wNDiag_55[54] , 
        \wNDiag_55[53] , \wNDiag_55[52] , \wNDiag_55[51] , \wNDiag_55[50] , 
        \wNDiag_55[49] , \wNDiag_55[48] , \wNDiag_55[47] , \wNDiag_55[46] , 
        \wNDiag_55[45] , \wNDiag_55[44] , \wNDiag_55[43] , \wNDiag_55[42] , 
        \wNDiag_55[41] , \wNDiag_55[40] , \wNDiag_55[39] , \wNDiag_55[38] , 
        \wNDiag_55[37] , \wNDiag_55[36] , \wNDiag_55[35] , \wNDiag_55[34] , 
        \wNDiag_55[33] , \wNDiag_55[32] , \wNDiag_55[31] , \wNDiag_55[30] , 
        \wNDiag_55[29] , \wNDiag_55[28] , \wNDiag_55[27] , \wNDiag_55[26] , 
        \wNDiag_55[25] , \wNDiag_55[24] , \wNDiag_55[23] , \wNDiag_55[22] , 
        \wNDiag_55[21] , \wNDiag_55[20] , \wNDiag_55[19] , \wNDiag_55[18] , 
        \wNDiag_55[17] , \wNDiag_55[16] , \wNDiag_55[15] , \wNDiag_55[14] , 
        \wNDiag_55[13] , \wNDiag_55[12] , \wNDiag_55[11] , \wNDiag_55[10] , 
        \wNDiag_55[9] , \wNDiag_55[8] , \wNDiag_55[7] , \wNDiag_55[6] , 
        \wNDiag_55[5] , \wNDiag_55[4] , \wNDiag_55[3] , \wNDiag_55[2] , 
        \wNDiag_55[1] , \wNDiag_55[0] }), .CallOut(\wCall_56[0] ), .ReturnOut(
        \wReturn_55[0] ), .ColOut({\wColumn_56[63] , \wColumn_56[62] , 
        \wColumn_56[61] , \wColumn_56[60] , \wColumn_56[59] , \wColumn_56[58] , 
        \wColumn_56[57] , \wColumn_56[56] , \wColumn_56[55] , \wColumn_56[54] , 
        \wColumn_56[53] , \wColumn_56[52] , \wColumn_56[51] , \wColumn_56[50] , 
        \wColumn_56[49] , \wColumn_56[48] , \wColumn_56[47] , \wColumn_56[46] , 
        \wColumn_56[45] , \wColumn_56[44] , \wColumn_56[43] , \wColumn_56[42] , 
        \wColumn_56[41] , \wColumn_56[40] , \wColumn_56[39] , \wColumn_56[38] , 
        \wColumn_56[37] , \wColumn_56[36] , \wColumn_56[35] , \wColumn_56[34] , 
        \wColumn_56[33] , \wColumn_56[32] , \wColumn_56[31] , \wColumn_56[30] , 
        \wColumn_56[29] , \wColumn_56[28] , \wColumn_56[27] , \wColumn_56[26] , 
        \wColumn_56[25] , \wColumn_56[24] , \wColumn_56[23] , \wColumn_56[22] , 
        \wColumn_56[21] , \wColumn_56[20] , \wColumn_56[19] , \wColumn_56[18] , 
        \wColumn_56[17] , \wColumn_56[16] , \wColumn_56[15] , \wColumn_56[14] , 
        \wColumn_56[13] , \wColumn_56[12] , \wColumn_56[11] , \wColumn_56[10] , 
        \wColumn_56[9] , \wColumn_56[8] , \wColumn_56[7] , \wColumn_56[6] , 
        \wColumn_56[5] , \wColumn_56[4] , \wColumn_56[3] , \wColumn_56[2] , 
        \wColumn_56[1] , \wColumn_56[0] }), .PDiagOut({\wPDiag_56[63] , 
        \wPDiag_56[62] , \wPDiag_56[61] , \wPDiag_56[60] , \wPDiag_56[59] , 
        \wPDiag_56[58] , \wPDiag_56[57] , \wPDiag_56[56] , \wPDiag_56[55] , 
        \wPDiag_56[54] , \wPDiag_56[53] , \wPDiag_56[52] , \wPDiag_56[51] , 
        \wPDiag_56[50] , \wPDiag_56[49] , \wPDiag_56[48] , \wPDiag_56[47] , 
        \wPDiag_56[46] , \wPDiag_56[45] , \wPDiag_56[44] , \wPDiag_56[43] , 
        \wPDiag_56[42] , \wPDiag_56[41] , \wPDiag_56[40] , \wPDiag_56[39] , 
        \wPDiag_56[38] , \wPDiag_56[37] , \wPDiag_56[36] , \wPDiag_56[35] , 
        \wPDiag_56[34] , \wPDiag_56[33] , \wPDiag_56[32] , \wPDiag_56[31] , 
        \wPDiag_56[30] , \wPDiag_56[29] , \wPDiag_56[28] , \wPDiag_56[27] , 
        \wPDiag_56[26] , \wPDiag_56[25] , \wPDiag_56[24] , \wPDiag_56[23] , 
        \wPDiag_56[22] , \wPDiag_56[21] , \wPDiag_56[20] , \wPDiag_56[19] , 
        \wPDiag_56[18] , \wPDiag_56[17] , \wPDiag_56[16] , \wPDiag_56[15] , 
        \wPDiag_56[14] , \wPDiag_56[13] , \wPDiag_56[12] , \wPDiag_56[11] , 
        \wPDiag_56[10] , \wPDiag_56[9] , \wPDiag_56[8] , \wPDiag_56[7] , 
        \wPDiag_56[6] , \wPDiag_56[5] , \wPDiag_56[4] , \wPDiag_56[3] , 
        \wPDiag_56[2] , \wPDiag_56[1] , \wPDiag_56[0] }), .NDiagOut({
        \wNDiag_56[63] , \wNDiag_56[62] , \wNDiag_56[61] , \wNDiag_56[60] , 
        \wNDiag_56[59] , \wNDiag_56[58] , \wNDiag_56[57] , \wNDiag_56[56] , 
        \wNDiag_56[55] , \wNDiag_56[54] , \wNDiag_56[53] , \wNDiag_56[52] , 
        \wNDiag_56[51] , \wNDiag_56[50] , \wNDiag_56[49] , \wNDiag_56[48] , 
        \wNDiag_56[47] , \wNDiag_56[46] , \wNDiag_56[45] , \wNDiag_56[44] , 
        \wNDiag_56[43] , \wNDiag_56[42] , \wNDiag_56[41] , \wNDiag_56[40] , 
        \wNDiag_56[39] , \wNDiag_56[38] , \wNDiag_56[37] , \wNDiag_56[36] , 
        \wNDiag_56[35] , \wNDiag_56[34] , \wNDiag_56[33] , \wNDiag_56[32] , 
        \wNDiag_56[31] , \wNDiag_56[30] , \wNDiag_56[29] , \wNDiag_56[28] , 
        \wNDiag_56[27] , \wNDiag_56[26] , \wNDiag_56[25] , \wNDiag_56[24] , 
        \wNDiag_56[23] , \wNDiag_56[22] , \wNDiag_56[21] , \wNDiag_56[20] , 
        \wNDiag_56[19] , \wNDiag_56[18] , \wNDiag_56[17] , \wNDiag_56[16] , 
        \wNDiag_56[15] , \wNDiag_56[14] , \wNDiag_56[13] , \wNDiag_56[12] , 
        \wNDiag_56[11] , \wNDiag_56[10] , \wNDiag_56[9] , \wNDiag_56[8] , 
        \wNDiag_56[7] , \wNDiag_56[6] , \wNDiag_56[5] , \wNDiag_56[4] , 
        \wNDiag_56[3] , \wNDiag_56[2] , \wNDiag_56[1] , \wNDiag_56[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_21 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_22[6] , \wScan_22[5] , \wScan_22[4] , 
        \wScan_22[3] , \wScan_22[2] , \wScan_22[1] , \wScan_22[0] }), 
        .ScanOut({\wScan_21[6] , \wScan_21[5] , \wScan_21[4] , \wScan_21[3] , 
        \wScan_21[2] , \wScan_21[1] , \wScan_21[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_21[0] ), .ReturnIn(\wReturn_22[0] ), .ColIn({
        \wColumn_21[63] , \wColumn_21[62] , \wColumn_21[61] , \wColumn_21[60] , 
        \wColumn_21[59] , \wColumn_21[58] , \wColumn_21[57] , \wColumn_21[56] , 
        \wColumn_21[55] , \wColumn_21[54] , \wColumn_21[53] , \wColumn_21[52] , 
        \wColumn_21[51] , \wColumn_21[50] , \wColumn_21[49] , \wColumn_21[48] , 
        \wColumn_21[47] , \wColumn_21[46] , \wColumn_21[45] , \wColumn_21[44] , 
        \wColumn_21[43] , \wColumn_21[42] , \wColumn_21[41] , \wColumn_21[40] , 
        \wColumn_21[39] , \wColumn_21[38] , \wColumn_21[37] , \wColumn_21[36] , 
        \wColumn_21[35] , \wColumn_21[34] , \wColumn_21[33] , \wColumn_21[32] , 
        \wColumn_21[31] , \wColumn_21[30] , \wColumn_21[29] , \wColumn_21[28] , 
        \wColumn_21[27] , \wColumn_21[26] , \wColumn_21[25] , \wColumn_21[24] , 
        \wColumn_21[23] , \wColumn_21[22] , \wColumn_21[21] , \wColumn_21[20] , 
        \wColumn_21[19] , \wColumn_21[18] , \wColumn_21[17] , \wColumn_21[16] , 
        \wColumn_21[15] , \wColumn_21[14] , \wColumn_21[13] , \wColumn_21[12] , 
        \wColumn_21[11] , \wColumn_21[10] , \wColumn_21[9] , \wColumn_21[8] , 
        \wColumn_21[7] , \wColumn_21[6] , \wColumn_21[5] , \wColumn_21[4] , 
        \wColumn_21[3] , \wColumn_21[2] , \wColumn_21[1] , \wColumn_21[0] }), 
        .PDiagIn({\wPDiag_21[63] , \wPDiag_21[62] , \wPDiag_21[61] , 
        \wPDiag_21[60] , \wPDiag_21[59] , \wPDiag_21[58] , \wPDiag_21[57] , 
        \wPDiag_21[56] , \wPDiag_21[55] , \wPDiag_21[54] , \wPDiag_21[53] , 
        \wPDiag_21[52] , \wPDiag_21[51] , \wPDiag_21[50] , \wPDiag_21[49] , 
        \wPDiag_21[48] , \wPDiag_21[47] , \wPDiag_21[46] , \wPDiag_21[45] , 
        \wPDiag_21[44] , \wPDiag_21[43] , \wPDiag_21[42] , \wPDiag_21[41] , 
        \wPDiag_21[40] , \wPDiag_21[39] , \wPDiag_21[38] , \wPDiag_21[37] , 
        \wPDiag_21[36] , \wPDiag_21[35] , \wPDiag_21[34] , \wPDiag_21[33] , 
        \wPDiag_21[32] , \wPDiag_21[31] , \wPDiag_21[30] , \wPDiag_21[29] , 
        \wPDiag_21[28] , \wPDiag_21[27] , \wPDiag_21[26] , \wPDiag_21[25] , 
        \wPDiag_21[24] , \wPDiag_21[23] , \wPDiag_21[22] , \wPDiag_21[21] , 
        \wPDiag_21[20] , \wPDiag_21[19] , \wPDiag_21[18] , \wPDiag_21[17] , 
        \wPDiag_21[16] , \wPDiag_21[15] , \wPDiag_21[14] , \wPDiag_21[13] , 
        \wPDiag_21[12] , \wPDiag_21[11] , \wPDiag_21[10] , \wPDiag_21[9] , 
        \wPDiag_21[8] , \wPDiag_21[7] , \wPDiag_21[6] , \wPDiag_21[5] , 
        \wPDiag_21[4] , \wPDiag_21[3] , \wPDiag_21[2] , \wPDiag_21[1] , 
        \wPDiag_21[0] }), .NDiagIn({\wNDiag_21[63] , \wNDiag_21[62] , 
        \wNDiag_21[61] , \wNDiag_21[60] , \wNDiag_21[59] , \wNDiag_21[58] , 
        \wNDiag_21[57] , \wNDiag_21[56] , \wNDiag_21[55] , \wNDiag_21[54] , 
        \wNDiag_21[53] , \wNDiag_21[52] , \wNDiag_21[51] , \wNDiag_21[50] , 
        \wNDiag_21[49] , \wNDiag_21[48] , \wNDiag_21[47] , \wNDiag_21[46] , 
        \wNDiag_21[45] , \wNDiag_21[44] , \wNDiag_21[43] , \wNDiag_21[42] , 
        \wNDiag_21[41] , \wNDiag_21[40] , \wNDiag_21[39] , \wNDiag_21[38] , 
        \wNDiag_21[37] , \wNDiag_21[36] , \wNDiag_21[35] , \wNDiag_21[34] , 
        \wNDiag_21[33] , \wNDiag_21[32] , \wNDiag_21[31] , \wNDiag_21[30] , 
        \wNDiag_21[29] , \wNDiag_21[28] , \wNDiag_21[27] , \wNDiag_21[26] , 
        \wNDiag_21[25] , \wNDiag_21[24] , \wNDiag_21[23] , \wNDiag_21[22] , 
        \wNDiag_21[21] , \wNDiag_21[20] , \wNDiag_21[19] , \wNDiag_21[18] , 
        \wNDiag_21[17] , \wNDiag_21[16] , \wNDiag_21[15] , \wNDiag_21[14] , 
        \wNDiag_21[13] , \wNDiag_21[12] , \wNDiag_21[11] , \wNDiag_21[10] , 
        \wNDiag_21[9] , \wNDiag_21[8] , \wNDiag_21[7] , \wNDiag_21[6] , 
        \wNDiag_21[5] , \wNDiag_21[4] , \wNDiag_21[3] , \wNDiag_21[2] , 
        \wNDiag_21[1] , \wNDiag_21[0] }), .CallOut(\wCall_22[0] ), .ReturnOut(
        \wReturn_21[0] ), .ColOut({\wColumn_22[63] , \wColumn_22[62] , 
        \wColumn_22[61] , \wColumn_22[60] , \wColumn_22[59] , \wColumn_22[58] , 
        \wColumn_22[57] , \wColumn_22[56] , \wColumn_22[55] , \wColumn_22[54] , 
        \wColumn_22[53] , \wColumn_22[52] , \wColumn_22[51] , \wColumn_22[50] , 
        \wColumn_22[49] , \wColumn_22[48] , \wColumn_22[47] , \wColumn_22[46] , 
        \wColumn_22[45] , \wColumn_22[44] , \wColumn_22[43] , \wColumn_22[42] , 
        \wColumn_22[41] , \wColumn_22[40] , \wColumn_22[39] , \wColumn_22[38] , 
        \wColumn_22[37] , \wColumn_22[36] , \wColumn_22[35] , \wColumn_22[34] , 
        \wColumn_22[33] , \wColumn_22[32] , \wColumn_22[31] , \wColumn_22[30] , 
        \wColumn_22[29] , \wColumn_22[28] , \wColumn_22[27] , \wColumn_22[26] , 
        \wColumn_22[25] , \wColumn_22[24] , \wColumn_22[23] , \wColumn_22[22] , 
        \wColumn_22[21] , \wColumn_22[20] , \wColumn_22[19] , \wColumn_22[18] , 
        \wColumn_22[17] , \wColumn_22[16] , \wColumn_22[15] , \wColumn_22[14] , 
        \wColumn_22[13] , \wColumn_22[12] , \wColumn_22[11] , \wColumn_22[10] , 
        \wColumn_22[9] , \wColumn_22[8] , \wColumn_22[7] , \wColumn_22[6] , 
        \wColumn_22[5] , \wColumn_22[4] , \wColumn_22[3] , \wColumn_22[2] , 
        \wColumn_22[1] , \wColumn_22[0] }), .PDiagOut({\wPDiag_22[63] , 
        \wPDiag_22[62] , \wPDiag_22[61] , \wPDiag_22[60] , \wPDiag_22[59] , 
        \wPDiag_22[58] , \wPDiag_22[57] , \wPDiag_22[56] , \wPDiag_22[55] , 
        \wPDiag_22[54] , \wPDiag_22[53] , \wPDiag_22[52] , \wPDiag_22[51] , 
        \wPDiag_22[50] , \wPDiag_22[49] , \wPDiag_22[48] , \wPDiag_22[47] , 
        \wPDiag_22[46] , \wPDiag_22[45] , \wPDiag_22[44] , \wPDiag_22[43] , 
        \wPDiag_22[42] , \wPDiag_22[41] , \wPDiag_22[40] , \wPDiag_22[39] , 
        \wPDiag_22[38] , \wPDiag_22[37] , \wPDiag_22[36] , \wPDiag_22[35] , 
        \wPDiag_22[34] , \wPDiag_22[33] , \wPDiag_22[32] , \wPDiag_22[31] , 
        \wPDiag_22[30] , \wPDiag_22[29] , \wPDiag_22[28] , \wPDiag_22[27] , 
        \wPDiag_22[26] , \wPDiag_22[25] , \wPDiag_22[24] , \wPDiag_22[23] , 
        \wPDiag_22[22] , \wPDiag_22[21] , \wPDiag_22[20] , \wPDiag_22[19] , 
        \wPDiag_22[18] , \wPDiag_22[17] , \wPDiag_22[16] , \wPDiag_22[15] , 
        \wPDiag_22[14] , \wPDiag_22[13] , \wPDiag_22[12] , \wPDiag_22[11] , 
        \wPDiag_22[10] , \wPDiag_22[9] , \wPDiag_22[8] , \wPDiag_22[7] , 
        \wPDiag_22[6] , \wPDiag_22[5] , \wPDiag_22[4] , \wPDiag_22[3] , 
        \wPDiag_22[2] , \wPDiag_22[1] , \wPDiag_22[0] }), .NDiagOut({
        \wNDiag_22[63] , \wNDiag_22[62] , \wNDiag_22[61] , \wNDiag_22[60] , 
        \wNDiag_22[59] , \wNDiag_22[58] , \wNDiag_22[57] , \wNDiag_22[56] , 
        \wNDiag_22[55] , \wNDiag_22[54] , \wNDiag_22[53] , \wNDiag_22[52] , 
        \wNDiag_22[51] , \wNDiag_22[50] , \wNDiag_22[49] , \wNDiag_22[48] , 
        \wNDiag_22[47] , \wNDiag_22[46] , \wNDiag_22[45] , \wNDiag_22[44] , 
        \wNDiag_22[43] , \wNDiag_22[42] , \wNDiag_22[41] , \wNDiag_22[40] , 
        \wNDiag_22[39] , \wNDiag_22[38] , \wNDiag_22[37] , \wNDiag_22[36] , 
        \wNDiag_22[35] , \wNDiag_22[34] , \wNDiag_22[33] , \wNDiag_22[32] , 
        \wNDiag_22[31] , \wNDiag_22[30] , \wNDiag_22[29] , \wNDiag_22[28] , 
        \wNDiag_22[27] , \wNDiag_22[26] , \wNDiag_22[25] , \wNDiag_22[24] , 
        \wNDiag_22[23] , \wNDiag_22[22] , \wNDiag_22[21] , \wNDiag_22[20] , 
        \wNDiag_22[19] , \wNDiag_22[18] , \wNDiag_22[17] , \wNDiag_22[16] , 
        \wNDiag_22[15] , \wNDiag_22[14] , \wNDiag_22[13] , \wNDiag_22[12] , 
        \wNDiag_22[11] , \wNDiag_22[10] , \wNDiag_22[9] , \wNDiag_22[8] , 
        \wNDiag_22[7] , \wNDiag_22[6] , \wNDiag_22[5] , \wNDiag_22[4] , 
        \wNDiag_22[3] , \wNDiag_22[2] , \wNDiag_22[1] , \wNDiag_22[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_29 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_30[6] , \wScan_30[5] , \wScan_30[4] , 
        \wScan_30[3] , \wScan_30[2] , \wScan_30[1] , \wScan_30[0] }), 
        .ScanOut({\wScan_29[6] , \wScan_29[5] , \wScan_29[4] , \wScan_29[3] , 
        \wScan_29[2] , \wScan_29[1] , \wScan_29[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_29[0] ), .ReturnIn(\wReturn_30[0] ), .ColIn({
        \wColumn_29[63] , \wColumn_29[62] , \wColumn_29[61] , \wColumn_29[60] , 
        \wColumn_29[59] , \wColumn_29[58] , \wColumn_29[57] , \wColumn_29[56] , 
        \wColumn_29[55] , \wColumn_29[54] , \wColumn_29[53] , \wColumn_29[52] , 
        \wColumn_29[51] , \wColumn_29[50] , \wColumn_29[49] , \wColumn_29[48] , 
        \wColumn_29[47] , \wColumn_29[46] , \wColumn_29[45] , \wColumn_29[44] , 
        \wColumn_29[43] , \wColumn_29[42] , \wColumn_29[41] , \wColumn_29[40] , 
        \wColumn_29[39] , \wColumn_29[38] , \wColumn_29[37] , \wColumn_29[36] , 
        \wColumn_29[35] , \wColumn_29[34] , \wColumn_29[33] , \wColumn_29[32] , 
        \wColumn_29[31] , \wColumn_29[30] , \wColumn_29[29] , \wColumn_29[28] , 
        \wColumn_29[27] , \wColumn_29[26] , \wColumn_29[25] , \wColumn_29[24] , 
        \wColumn_29[23] , \wColumn_29[22] , \wColumn_29[21] , \wColumn_29[20] , 
        \wColumn_29[19] , \wColumn_29[18] , \wColumn_29[17] , \wColumn_29[16] , 
        \wColumn_29[15] , \wColumn_29[14] , \wColumn_29[13] , \wColumn_29[12] , 
        \wColumn_29[11] , \wColumn_29[10] , \wColumn_29[9] , \wColumn_29[8] , 
        \wColumn_29[7] , \wColumn_29[6] , \wColumn_29[5] , \wColumn_29[4] , 
        \wColumn_29[3] , \wColumn_29[2] , \wColumn_29[1] , \wColumn_29[0] }), 
        .PDiagIn({\wPDiag_29[63] , \wPDiag_29[62] , \wPDiag_29[61] , 
        \wPDiag_29[60] , \wPDiag_29[59] , \wPDiag_29[58] , \wPDiag_29[57] , 
        \wPDiag_29[56] , \wPDiag_29[55] , \wPDiag_29[54] , \wPDiag_29[53] , 
        \wPDiag_29[52] , \wPDiag_29[51] , \wPDiag_29[50] , \wPDiag_29[49] , 
        \wPDiag_29[48] , \wPDiag_29[47] , \wPDiag_29[46] , \wPDiag_29[45] , 
        \wPDiag_29[44] , \wPDiag_29[43] , \wPDiag_29[42] , \wPDiag_29[41] , 
        \wPDiag_29[40] , \wPDiag_29[39] , \wPDiag_29[38] , \wPDiag_29[37] , 
        \wPDiag_29[36] , \wPDiag_29[35] , \wPDiag_29[34] , \wPDiag_29[33] , 
        \wPDiag_29[32] , \wPDiag_29[31] , \wPDiag_29[30] , \wPDiag_29[29] , 
        \wPDiag_29[28] , \wPDiag_29[27] , \wPDiag_29[26] , \wPDiag_29[25] , 
        \wPDiag_29[24] , \wPDiag_29[23] , \wPDiag_29[22] , \wPDiag_29[21] , 
        \wPDiag_29[20] , \wPDiag_29[19] , \wPDiag_29[18] , \wPDiag_29[17] , 
        \wPDiag_29[16] , \wPDiag_29[15] , \wPDiag_29[14] , \wPDiag_29[13] , 
        \wPDiag_29[12] , \wPDiag_29[11] , \wPDiag_29[10] , \wPDiag_29[9] , 
        \wPDiag_29[8] , \wPDiag_29[7] , \wPDiag_29[6] , \wPDiag_29[5] , 
        \wPDiag_29[4] , \wPDiag_29[3] , \wPDiag_29[2] , \wPDiag_29[1] , 
        \wPDiag_29[0] }), .NDiagIn({\wNDiag_29[63] , \wNDiag_29[62] , 
        \wNDiag_29[61] , \wNDiag_29[60] , \wNDiag_29[59] , \wNDiag_29[58] , 
        \wNDiag_29[57] , \wNDiag_29[56] , \wNDiag_29[55] , \wNDiag_29[54] , 
        \wNDiag_29[53] , \wNDiag_29[52] , \wNDiag_29[51] , \wNDiag_29[50] , 
        \wNDiag_29[49] , \wNDiag_29[48] , \wNDiag_29[47] , \wNDiag_29[46] , 
        \wNDiag_29[45] , \wNDiag_29[44] , \wNDiag_29[43] , \wNDiag_29[42] , 
        \wNDiag_29[41] , \wNDiag_29[40] , \wNDiag_29[39] , \wNDiag_29[38] , 
        \wNDiag_29[37] , \wNDiag_29[36] , \wNDiag_29[35] , \wNDiag_29[34] , 
        \wNDiag_29[33] , \wNDiag_29[32] , \wNDiag_29[31] , \wNDiag_29[30] , 
        \wNDiag_29[29] , \wNDiag_29[28] , \wNDiag_29[27] , \wNDiag_29[26] , 
        \wNDiag_29[25] , \wNDiag_29[24] , \wNDiag_29[23] , \wNDiag_29[22] , 
        \wNDiag_29[21] , \wNDiag_29[20] , \wNDiag_29[19] , \wNDiag_29[18] , 
        \wNDiag_29[17] , \wNDiag_29[16] , \wNDiag_29[15] , \wNDiag_29[14] , 
        \wNDiag_29[13] , \wNDiag_29[12] , \wNDiag_29[11] , \wNDiag_29[10] , 
        \wNDiag_29[9] , \wNDiag_29[8] , \wNDiag_29[7] , \wNDiag_29[6] , 
        \wNDiag_29[5] , \wNDiag_29[4] , \wNDiag_29[3] , \wNDiag_29[2] , 
        \wNDiag_29[1] , \wNDiag_29[0] }), .CallOut(\wCall_30[0] ), .ReturnOut(
        \wReturn_29[0] ), .ColOut({\wColumn_30[63] , \wColumn_30[62] , 
        \wColumn_30[61] , \wColumn_30[60] , \wColumn_30[59] , \wColumn_30[58] , 
        \wColumn_30[57] , \wColumn_30[56] , \wColumn_30[55] , \wColumn_30[54] , 
        \wColumn_30[53] , \wColumn_30[52] , \wColumn_30[51] , \wColumn_30[50] , 
        \wColumn_30[49] , \wColumn_30[48] , \wColumn_30[47] , \wColumn_30[46] , 
        \wColumn_30[45] , \wColumn_30[44] , \wColumn_30[43] , \wColumn_30[42] , 
        \wColumn_30[41] , \wColumn_30[40] , \wColumn_30[39] , \wColumn_30[38] , 
        \wColumn_30[37] , \wColumn_30[36] , \wColumn_30[35] , \wColumn_30[34] , 
        \wColumn_30[33] , \wColumn_30[32] , \wColumn_30[31] , \wColumn_30[30] , 
        \wColumn_30[29] , \wColumn_30[28] , \wColumn_30[27] , \wColumn_30[26] , 
        \wColumn_30[25] , \wColumn_30[24] , \wColumn_30[23] , \wColumn_30[22] , 
        \wColumn_30[21] , \wColumn_30[20] , \wColumn_30[19] , \wColumn_30[18] , 
        \wColumn_30[17] , \wColumn_30[16] , \wColumn_30[15] , \wColumn_30[14] , 
        \wColumn_30[13] , \wColumn_30[12] , \wColumn_30[11] , \wColumn_30[10] , 
        \wColumn_30[9] , \wColumn_30[8] , \wColumn_30[7] , \wColumn_30[6] , 
        \wColumn_30[5] , \wColumn_30[4] , \wColumn_30[3] , \wColumn_30[2] , 
        \wColumn_30[1] , \wColumn_30[0] }), .PDiagOut({\wPDiag_30[63] , 
        \wPDiag_30[62] , \wPDiag_30[61] , \wPDiag_30[60] , \wPDiag_30[59] , 
        \wPDiag_30[58] , \wPDiag_30[57] , \wPDiag_30[56] , \wPDiag_30[55] , 
        \wPDiag_30[54] , \wPDiag_30[53] , \wPDiag_30[52] , \wPDiag_30[51] , 
        \wPDiag_30[50] , \wPDiag_30[49] , \wPDiag_30[48] , \wPDiag_30[47] , 
        \wPDiag_30[46] , \wPDiag_30[45] , \wPDiag_30[44] , \wPDiag_30[43] , 
        \wPDiag_30[42] , \wPDiag_30[41] , \wPDiag_30[40] , \wPDiag_30[39] , 
        \wPDiag_30[38] , \wPDiag_30[37] , \wPDiag_30[36] , \wPDiag_30[35] , 
        \wPDiag_30[34] , \wPDiag_30[33] , \wPDiag_30[32] , \wPDiag_30[31] , 
        \wPDiag_30[30] , \wPDiag_30[29] , \wPDiag_30[28] , \wPDiag_30[27] , 
        \wPDiag_30[26] , \wPDiag_30[25] , \wPDiag_30[24] , \wPDiag_30[23] , 
        \wPDiag_30[22] , \wPDiag_30[21] , \wPDiag_30[20] , \wPDiag_30[19] , 
        \wPDiag_30[18] , \wPDiag_30[17] , \wPDiag_30[16] , \wPDiag_30[15] , 
        \wPDiag_30[14] , \wPDiag_30[13] , \wPDiag_30[12] , \wPDiag_30[11] , 
        \wPDiag_30[10] , \wPDiag_30[9] , \wPDiag_30[8] , \wPDiag_30[7] , 
        \wPDiag_30[6] , \wPDiag_30[5] , \wPDiag_30[4] , \wPDiag_30[3] , 
        \wPDiag_30[2] , \wPDiag_30[1] , \wPDiag_30[0] }), .NDiagOut({
        \wNDiag_30[63] , \wNDiag_30[62] , \wNDiag_30[61] , \wNDiag_30[60] , 
        \wNDiag_30[59] , \wNDiag_30[58] , \wNDiag_30[57] , \wNDiag_30[56] , 
        \wNDiag_30[55] , \wNDiag_30[54] , \wNDiag_30[53] , \wNDiag_30[52] , 
        \wNDiag_30[51] , \wNDiag_30[50] , \wNDiag_30[49] , \wNDiag_30[48] , 
        \wNDiag_30[47] , \wNDiag_30[46] , \wNDiag_30[45] , \wNDiag_30[44] , 
        \wNDiag_30[43] , \wNDiag_30[42] , \wNDiag_30[41] , \wNDiag_30[40] , 
        \wNDiag_30[39] , \wNDiag_30[38] , \wNDiag_30[37] , \wNDiag_30[36] , 
        \wNDiag_30[35] , \wNDiag_30[34] , \wNDiag_30[33] , \wNDiag_30[32] , 
        \wNDiag_30[31] , \wNDiag_30[30] , \wNDiag_30[29] , \wNDiag_30[28] , 
        \wNDiag_30[27] , \wNDiag_30[26] , \wNDiag_30[25] , \wNDiag_30[24] , 
        \wNDiag_30[23] , \wNDiag_30[22] , \wNDiag_30[21] , \wNDiag_30[20] , 
        \wNDiag_30[19] , \wNDiag_30[18] , \wNDiag_30[17] , \wNDiag_30[16] , 
        \wNDiag_30[15] , \wNDiag_30[14] , \wNDiag_30[13] , \wNDiag_30[12] , 
        \wNDiag_30[11] , \wNDiag_30[10] , \wNDiag_30[9] , \wNDiag_30[8] , 
        \wNDiag_30[7] , \wNDiag_30[6] , \wNDiag_30[5] , \wNDiag_30[4] , 
        \wNDiag_30[3] , \wNDiag_30[2] , \wNDiag_30[1] , \wNDiag_30[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_32 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_33[6] , \wScan_33[5] , \wScan_33[4] , 
        \wScan_33[3] , \wScan_33[2] , \wScan_33[1] , \wScan_33[0] }), 
        .ScanOut({\wScan_32[6] , \wScan_32[5] , \wScan_32[4] , \wScan_32[3] , 
        \wScan_32[2] , \wScan_32[1] , \wScan_32[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_32[0] ), .ReturnIn(\wReturn_33[0] ), .ColIn({
        \wColumn_32[63] , \wColumn_32[62] , \wColumn_32[61] , \wColumn_32[60] , 
        \wColumn_32[59] , \wColumn_32[58] , \wColumn_32[57] , \wColumn_32[56] , 
        \wColumn_32[55] , \wColumn_32[54] , \wColumn_32[53] , \wColumn_32[52] , 
        \wColumn_32[51] , \wColumn_32[50] , \wColumn_32[49] , \wColumn_32[48] , 
        \wColumn_32[47] , \wColumn_32[46] , \wColumn_32[45] , \wColumn_32[44] , 
        \wColumn_32[43] , \wColumn_32[42] , \wColumn_32[41] , \wColumn_32[40] , 
        \wColumn_32[39] , \wColumn_32[38] , \wColumn_32[37] , \wColumn_32[36] , 
        \wColumn_32[35] , \wColumn_32[34] , \wColumn_32[33] , \wColumn_32[32] , 
        \wColumn_32[31] , \wColumn_32[30] , \wColumn_32[29] , \wColumn_32[28] , 
        \wColumn_32[27] , \wColumn_32[26] , \wColumn_32[25] , \wColumn_32[24] , 
        \wColumn_32[23] , \wColumn_32[22] , \wColumn_32[21] , \wColumn_32[20] , 
        \wColumn_32[19] , \wColumn_32[18] , \wColumn_32[17] , \wColumn_32[16] , 
        \wColumn_32[15] , \wColumn_32[14] , \wColumn_32[13] , \wColumn_32[12] , 
        \wColumn_32[11] , \wColumn_32[10] , \wColumn_32[9] , \wColumn_32[8] , 
        \wColumn_32[7] , \wColumn_32[6] , \wColumn_32[5] , \wColumn_32[4] , 
        \wColumn_32[3] , \wColumn_32[2] , \wColumn_32[1] , \wColumn_32[0] }), 
        .PDiagIn({\wPDiag_32[63] , \wPDiag_32[62] , \wPDiag_32[61] , 
        \wPDiag_32[60] , \wPDiag_32[59] , \wPDiag_32[58] , \wPDiag_32[57] , 
        \wPDiag_32[56] , \wPDiag_32[55] , \wPDiag_32[54] , \wPDiag_32[53] , 
        \wPDiag_32[52] , \wPDiag_32[51] , \wPDiag_32[50] , \wPDiag_32[49] , 
        \wPDiag_32[48] , \wPDiag_32[47] , \wPDiag_32[46] , \wPDiag_32[45] , 
        \wPDiag_32[44] , \wPDiag_32[43] , \wPDiag_32[42] , \wPDiag_32[41] , 
        \wPDiag_32[40] , \wPDiag_32[39] , \wPDiag_32[38] , \wPDiag_32[37] , 
        \wPDiag_32[36] , \wPDiag_32[35] , \wPDiag_32[34] , \wPDiag_32[33] , 
        \wPDiag_32[32] , \wPDiag_32[31] , \wPDiag_32[30] , \wPDiag_32[29] , 
        \wPDiag_32[28] , \wPDiag_32[27] , \wPDiag_32[26] , \wPDiag_32[25] , 
        \wPDiag_32[24] , \wPDiag_32[23] , \wPDiag_32[22] , \wPDiag_32[21] , 
        \wPDiag_32[20] , \wPDiag_32[19] , \wPDiag_32[18] , \wPDiag_32[17] , 
        \wPDiag_32[16] , \wPDiag_32[15] , \wPDiag_32[14] , \wPDiag_32[13] , 
        \wPDiag_32[12] , \wPDiag_32[11] , \wPDiag_32[10] , \wPDiag_32[9] , 
        \wPDiag_32[8] , \wPDiag_32[7] , \wPDiag_32[6] , \wPDiag_32[5] , 
        \wPDiag_32[4] , \wPDiag_32[3] , \wPDiag_32[2] , \wPDiag_32[1] , 
        \wPDiag_32[0] }), .NDiagIn({\wNDiag_32[63] , \wNDiag_32[62] , 
        \wNDiag_32[61] , \wNDiag_32[60] , \wNDiag_32[59] , \wNDiag_32[58] , 
        \wNDiag_32[57] , \wNDiag_32[56] , \wNDiag_32[55] , \wNDiag_32[54] , 
        \wNDiag_32[53] , \wNDiag_32[52] , \wNDiag_32[51] , \wNDiag_32[50] , 
        \wNDiag_32[49] , \wNDiag_32[48] , \wNDiag_32[47] , \wNDiag_32[46] , 
        \wNDiag_32[45] , \wNDiag_32[44] , \wNDiag_32[43] , \wNDiag_32[42] , 
        \wNDiag_32[41] , \wNDiag_32[40] , \wNDiag_32[39] , \wNDiag_32[38] , 
        \wNDiag_32[37] , \wNDiag_32[36] , \wNDiag_32[35] , \wNDiag_32[34] , 
        \wNDiag_32[33] , \wNDiag_32[32] , \wNDiag_32[31] , \wNDiag_32[30] , 
        \wNDiag_32[29] , \wNDiag_32[28] , \wNDiag_32[27] , \wNDiag_32[26] , 
        \wNDiag_32[25] , \wNDiag_32[24] , \wNDiag_32[23] , \wNDiag_32[22] , 
        \wNDiag_32[21] , \wNDiag_32[20] , \wNDiag_32[19] , \wNDiag_32[18] , 
        \wNDiag_32[17] , \wNDiag_32[16] , \wNDiag_32[15] , \wNDiag_32[14] , 
        \wNDiag_32[13] , \wNDiag_32[12] , \wNDiag_32[11] , \wNDiag_32[10] , 
        \wNDiag_32[9] , \wNDiag_32[8] , \wNDiag_32[7] , \wNDiag_32[6] , 
        \wNDiag_32[5] , \wNDiag_32[4] , \wNDiag_32[3] , \wNDiag_32[2] , 
        \wNDiag_32[1] , \wNDiag_32[0] }), .CallOut(\wCall_33[0] ), .ReturnOut(
        \wReturn_32[0] ), .ColOut({\wColumn_33[63] , \wColumn_33[62] , 
        \wColumn_33[61] , \wColumn_33[60] , \wColumn_33[59] , \wColumn_33[58] , 
        \wColumn_33[57] , \wColumn_33[56] , \wColumn_33[55] , \wColumn_33[54] , 
        \wColumn_33[53] , \wColumn_33[52] , \wColumn_33[51] , \wColumn_33[50] , 
        \wColumn_33[49] , \wColumn_33[48] , \wColumn_33[47] , \wColumn_33[46] , 
        \wColumn_33[45] , \wColumn_33[44] , \wColumn_33[43] , \wColumn_33[42] , 
        \wColumn_33[41] , \wColumn_33[40] , \wColumn_33[39] , \wColumn_33[38] , 
        \wColumn_33[37] , \wColumn_33[36] , \wColumn_33[35] , \wColumn_33[34] , 
        \wColumn_33[33] , \wColumn_33[32] , \wColumn_33[31] , \wColumn_33[30] , 
        \wColumn_33[29] , \wColumn_33[28] , \wColumn_33[27] , \wColumn_33[26] , 
        \wColumn_33[25] , \wColumn_33[24] , \wColumn_33[23] , \wColumn_33[22] , 
        \wColumn_33[21] , \wColumn_33[20] , \wColumn_33[19] , \wColumn_33[18] , 
        \wColumn_33[17] , \wColumn_33[16] , \wColumn_33[15] , \wColumn_33[14] , 
        \wColumn_33[13] , \wColumn_33[12] , \wColumn_33[11] , \wColumn_33[10] , 
        \wColumn_33[9] , \wColumn_33[8] , \wColumn_33[7] , \wColumn_33[6] , 
        \wColumn_33[5] , \wColumn_33[4] , \wColumn_33[3] , \wColumn_33[2] , 
        \wColumn_33[1] , \wColumn_33[0] }), .PDiagOut({\wPDiag_33[63] , 
        \wPDiag_33[62] , \wPDiag_33[61] , \wPDiag_33[60] , \wPDiag_33[59] , 
        \wPDiag_33[58] , \wPDiag_33[57] , \wPDiag_33[56] , \wPDiag_33[55] , 
        \wPDiag_33[54] , \wPDiag_33[53] , \wPDiag_33[52] , \wPDiag_33[51] , 
        \wPDiag_33[50] , \wPDiag_33[49] , \wPDiag_33[48] , \wPDiag_33[47] , 
        \wPDiag_33[46] , \wPDiag_33[45] , \wPDiag_33[44] , \wPDiag_33[43] , 
        \wPDiag_33[42] , \wPDiag_33[41] , \wPDiag_33[40] , \wPDiag_33[39] , 
        \wPDiag_33[38] , \wPDiag_33[37] , \wPDiag_33[36] , \wPDiag_33[35] , 
        \wPDiag_33[34] , \wPDiag_33[33] , \wPDiag_33[32] , \wPDiag_33[31] , 
        \wPDiag_33[30] , \wPDiag_33[29] , \wPDiag_33[28] , \wPDiag_33[27] , 
        \wPDiag_33[26] , \wPDiag_33[25] , \wPDiag_33[24] , \wPDiag_33[23] , 
        \wPDiag_33[22] , \wPDiag_33[21] , \wPDiag_33[20] , \wPDiag_33[19] , 
        \wPDiag_33[18] , \wPDiag_33[17] , \wPDiag_33[16] , \wPDiag_33[15] , 
        \wPDiag_33[14] , \wPDiag_33[13] , \wPDiag_33[12] , \wPDiag_33[11] , 
        \wPDiag_33[10] , \wPDiag_33[9] , \wPDiag_33[8] , \wPDiag_33[7] , 
        \wPDiag_33[6] , \wPDiag_33[5] , \wPDiag_33[4] , \wPDiag_33[3] , 
        \wPDiag_33[2] , \wPDiag_33[1] , \wPDiag_33[0] }), .NDiagOut({
        \wNDiag_33[63] , \wNDiag_33[62] , \wNDiag_33[61] , \wNDiag_33[60] , 
        \wNDiag_33[59] , \wNDiag_33[58] , \wNDiag_33[57] , \wNDiag_33[56] , 
        \wNDiag_33[55] , \wNDiag_33[54] , \wNDiag_33[53] , \wNDiag_33[52] , 
        \wNDiag_33[51] , \wNDiag_33[50] , \wNDiag_33[49] , \wNDiag_33[48] , 
        \wNDiag_33[47] , \wNDiag_33[46] , \wNDiag_33[45] , \wNDiag_33[44] , 
        \wNDiag_33[43] , \wNDiag_33[42] , \wNDiag_33[41] , \wNDiag_33[40] , 
        \wNDiag_33[39] , \wNDiag_33[38] , \wNDiag_33[37] , \wNDiag_33[36] , 
        \wNDiag_33[35] , \wNDiag_33[34] , \wNDiag_33[33] , \wNDiag_33[32] , 
        \wNDiag_33[31] , \wNDiag_33[30] , \wNDiag_33[29] , \wNDiag_33[28] , 
        \wNDiag_33[27] , \wNDiag_33[26] , \wNDiag_33[25] , \wNDiag_33[24] , 
        \wNDiag_33[23] , \wNDiag_33[22] , \wNDiag_33[21] , \wNDiag_33[20] , 
        \wNDiag_33[19] , \wNDiag_33[18] , \wNDiag_33[17] , \wNDiag_33[16] , 
        \wNDiag_33[15] , \wNDiag_33[14] , \wNDiag_33[13] , \wNDiag_33[12] , 
        \wNDiag_33[11] , \wNDiag_33[10] , \wNDiag_33[9] , \wNDiag_33[8] , 
        \wNDiag_33[7] , \wNDiag_33[6] , \wNDiag_33[5] , \wNDiag_33[4] , 
        \wNDiag_33[3] , \wNDiag_33[2] , \wNDiag_33[1] , \wNDiag_33[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_47 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_48[6] , \wScan_48[5] , \wScan_48[4] , 
        \wScan_48[3] , \wScan_48[2] , \wScan_48[1] , \wScan_48[0] }), 
        .ScanOut({\wScan_47[6] , \wScan_47[5] , \wScan_47[4] , \wScan_47[3] , 
        \wScan_47[2] , \wScan_47[1] , \wScan_47[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_47[0] ), .ReturnIn(\wReturn_48[0] ), .ColIn({
        \wColumn_47[63] , \wColumn_47[62] , \wColumn_47[61] , \wColumn_47[60] , 
        \wColumn_47[59] , \wColumn_47[58] , \wColumn_47[57] , \wColumn_47[56] , 
        \wColumn_47[55] , \wColumn_47[54] , \wColumn_47[53] , \wColumn_47[52] , 
        \wColumn_47[51] , \wColumn_47[50] , \wColumn_47[49] , \wColumn_47[48] , 
        \wColumn_47[47] , \wColumn_47[46] , \wColumn_47[45] , \wColumn_47[44] , 
        \wColumn_47[43] , \wColumn_47[42] , \wColumn_47[41] , \wColumn_47[40] , 
        \wColumn_47[39] , \wColumn_47[38] , \wColumn_47[37] , \wColumn_47[36] , 
        \wColumn_47[35] , \wColumn_47[34] , \wColumn_47[33] , \wColumn_47[32] , 
        \wColumn_47[31] , \wColumn_47[30] , \wColumn_47[29] , \wColumn_47[28] , 
        \wColumn_47[27] , \wColumn_47[26] , \wColumn_47[25] , \wColumn_47[24] , 
        \wColumn_47[23] , \wColumn_47[22] , \wColumn_47[21] , \wColumn_47[20] , 
        \wColumn_47[19] , \wColumn_47[18] , \wColumn_47[17] , \wColumn_47[16] , 
        \wColumn_47[15] , \wColumn_47[14] , \wColumn_47[13] , \wColumn_47[12] , 
        \wColumn_47[11] , \wColumn_47[10] , \wColumn_47[9] , \wColumn_47[8] , 
        \wColumn_47[7] , \wColumn_47[6] , \wColumn_47[5] , \wColumn_47[4] , 
        \wColumn_47[3] , \wColumn_47[2] , \wColumn_47[1] , \wColumn_47[0] }), 
        .PDiagIn({\wPDiag_47[63] , \wPDiag_47[62] , \wPDiag_47[61] , 
        \wPDiag_47[60] , \wPDiag_47[59] , \wPDiag_47[58] , \wPDiag_47[57] , 
        \wPDiag_47[56] , \wPDiag_47[55] , \wPDiag_47[54] , \wPDiag_47[53] , 
        \wPDiag_47[52] , \wPDiag_47[51] , \wPDiag_47[50] , \wPDiag_47[49] , 
        \wPDiag_47[48] , \wPDiag_47[47] , \wPDiag_47[46] , \wPDiag_47[45] , 
        \wPDiag_47[44] , \wPDiag_47[43] , \wPDiag_47[42] , \wPDiag_47[41] , 
        \wPDiag_47[40] , \wPDiag_47[39] , \wPDiag_47[38] , \wPDiag_47[37] , 
        \wPDiag_47[36] , \wPDiag_47[35] , \wPDiag_47[34] , \wPDiag_47[33] , 
        \wPDiag_47[32] , \wPDiag_47[31] , \wPDiag_47[30] , \wPDiag_47[29] , 
        \wPDiag_47[28] , \wPDiag_47[27] , \wPDiag_47[26] , \wPDiag_47[25] , 
        \wPDiag_47[24] , \wPDiag_47[23] , \wPDiag_47[22] , \wPDiag_47[21] , 
        \wPDiag_47[20] , \wPDiag_47[19] , \wPDiag_47[18] , \wPDiag_47[17] , 
        \wPDiag_47[16] , \wPDiag_47[15] , \wPDiag_47[14] , \wPDiag_47[13] , 
        \wPDiag_47[12] , \wPDiag_47[11] , \wPDiag_47[10] , \wPDiag_47[9] , 
        \wPDiag_47[8] , \wPDiag_47[7] , \wPDiag_47[6] , \wPDiag_47[5] , 
        \wPDiag_47[4] , \wPDiag_47[3] , \wPDiag_47[2] , \wPDiag_47[1] , 
        \wPDiag_47[0] }), .NDiagIn({\wNDiag_47[63] , \wNDiag_47[62] , 
        \wNDiag_47[61] , \wNDiag_47[60] , \wNDiag_47[59] , \wNDiag_47[58] , 
        \wNDiag_47[57] , \wNDiag_47[56] , \wNDiag_47[55] , \wNDiag_47[54] , 
        \wNDiag_47[53] , \wNDiag_47[52] , \wNDiag_47[51] , \wNDiag_47[50] , 
        \wNDiag_47[49] , \wNDiag_47[48] , \wNDiag_47[47] , \wNDiag_47[46] , 
        \wNDiag_47[45] , \wNDiag_47[44] , \wNDiag_47[43] , \wNDiag_47[42] , 
        \wNDiag_47[41] , \wNDiag_47[40] , \wNDiag_47[39] , \wNDiag_47[38] , 
        \wNDiag_47[37] , \wNDiag_47[36] , \wNDiag_47[35] , \wNDiag_47[34] , 
        \wNDiag_47[33] , \wNDiag_47[32] , \wNDiag_47[31] , \wNDiag_47[30] , 
        \wNDiag_47[29] , \wNDiag_47[28] , \wNDiag_47[27] , \wNDiag_47[26] , 
        \wNDiag_47[25] , \wNDiag_47[24] , \wNDiag_47[23] , \wNDiag_47[22] , 
        \wNDiag_47[21] , \wNDiag_47[20] , \wNDiag_47[19] , \wNDiag_47[18] , 
        \wNDiag_47[17] , \wNDiag_47[16] , \wNDiag_47[15] , \wNDiag_47[14] , 
        \wNDiag_47[13] , \wNDiag_47[12] , \wNDiag_47[11] , \wNDiag_47[10] , 
        \wNDiag_47[9] , \wNDiag_47[8] , \wNDiag_47[7] , \wNDiag_47[6] , 
        \wNDiag_47[5] , \wNDiag_47[4] , \wNDiag_47[3] , \wNDiag_47[2] , 
        \wNDiag_47[1] , \wNDiag_47[0] }), .CallOut(\wCall_48[0] ), .ReturnOut(
        \wReturn_47[0] ), .ColOut({\wColumn_48[63] , \wColumn_48[62] , 
        \wColumn_48[61] , \wColumn_48[60] , \wColumn_48[59] , \wColumn_48[58] , 
        \wColumn_48[57] , \wColumn_48[56] , \wColumn_48[55] , \wColumn_48[54] , 
        \wColumn_48[53] , \wColumn_48[52] , \wColumn_48[51] , \wColumn_48[50] , 
        \wColumn_48[49] , \wColumn_48[48] , \wColumn_48[47] , \wColumn_48[46] , 
        \wColumn_48[45] , \wColumn_48[44] , \wColumn_48[43] , \wColumn_48[42] , 
        \wColumn_48[41] , \wColumn_48[40] , \wColumn_48[39] , \wColumn_48[38] , 
        \wColumn_48[37] , \wColumn_48[36] , \wColumn_48[35] , \wColumn_48[34] , 
        \wColumn_48[33] , \wColumn_48[32] , \wColumn_48[31] , \wColumn_48[30] , 
        \wColumn_48[29] , \wColumn_48[28] , \wColumn_48[27] , \wColumn_48[26] , 
        \wColumn_48[25] , \wColumn_48[24] , \wColumn_48[23] , \wColumn_48[22] , 
        \wColumn_48[21] , \wColumn_48[20] , \wColumn_48[19] , \wColumn_48[18] , 
        \wColumn_48[17] , \wColumn_48[16] , \wColumn_48[15] , \wColumn_48[14] , 
        \wColumn_48[13] , \wColumn_48[12] , \wColumn_48[11] , \wColumn_48[10] , 
        \wColumn_48[9] , \wColumn_48[8] , \wColumn_48[7] , \wColumn_48[6] , 
        \wColumn_48[5] , \wColumn_48[4] , \wColumn_48[3] , \wColumn_48[2] , 
        \wColumn_48[1] , \wColumn_48[0] }), .PDiagOut({\wPDiag_48[63] , 
        \wPDiag_48[62] , \wPDiag_48[61] , \wPDiag_48[60] , \wPDiag_48[59] , 
        \wPDiag_48[58] , \wPDiag_48[57] , \wPDiag_48[56] , \wPDiag_48[55] , 
        \wPDiag_48[54] , \wPDiag_48[53] , \wPDiag_48[52] , \wPDiag_48[51] , 
        \wPDiag_48[50] , \wPDiag_48[49] , \wPDiag_48[48] , \wPDiag_48[47] , 
        \wPDiag_48[46] , \wPDiag_48[45] , \wPDiag_48[44] , \wPDiag_48[43] , 
        \wPDiag_48[42] , \wPDiag_48[41] , \wPDiag_48[40] , \wPDiag_48[39] , 
        \wPDiag_48[38] , \wPDiag_48[37] , \wPDiag_48[36] , \wPDiag_48[35] , 
        \wPDiag_48[34] , \wPDiag_48[33] , \wPDiag_48[32] , \wPDiag_48[31] , 
        \wPDiag_48[30] , \wPDiag_48[29] , \wPDiag_48[28] , \wPDiag_48[27] , 
        \wPDiag_48[26] , \wPDiag_48[25] , \wPDiag_48[24] , \wPDiag_48[23] , 
        \wPDiag_48[22] , \wPDiag_48[21] , \wPDiag_48[20] , \wPDiag_48[19] , 
        \wPDiag_48[18] , \wPDiag_48[17] , \wPDiag_48[16] , \wPDiag_48[15] , 
        \wPDiag_48[14] , \wPDiag_48[13] , \wPDiag_48[12] , \wPDiag_48[11] , 
        \wPDiag_48[10] , \wPDiag_48[9] , \wPDiag_48[8] , \wPDiag_48[7] , 
        \wPDiag_48[6] , \wPDiag_48[5] , \wPDiag_48[4] , \wPDiag_48[3] , 
        \wPDiag_48[2] , \wPDiag_48[1] , \wPDiag_48[0] }), .NDiagOut({
        \wNDiag_48[63] , \wNDiag_48[62] , \wNDiag_48[61] , \wNDiag_48[60] , 
        \wNDiag_48[59] , \wNDiag_48[58] , \wNDiag_48[57] , \wNDiag_48[56] , 
        \wNDiag_48[55] , \wNDiag_48[54] , \wNDiag_48[53] , \wNDiag_48[52] , 
        \wNDiag_48[51] , \wNDiag_48[50] , \wNDiag_48[49] , \wNDiag_48[48] , 
        \wNDiag_48[47] , \wNDiag_48[46] , \wNDiag_48[45] , \wNDiag_48[44] , 
        \wNDiag_48[43] , \wNDiag_48[42] , \wNDiag_48[41] , \wNDiag_48[40] , 
        \wNDiag_48[39] , \wNDiag_48[38] , \wNDiag_48[37] , \wNDiag_48[36] , 
        \wNDiag_48[35] , \wNDiag_48[34] , \wNDiag_48[33] , \wNDiag_48[32] , 
        \wNDiag_48[31] , \wNDiag_48[30] , \wNDiag_48[29] , \wNDiag_48[28] , 
        \wNDiag_48[27] , \wNDiag_48[26] , \wNDiag_48[25] , \wNDiag_48[24] , 
        \wNDiag_48[23] , \wNDiag_48[22] , \wNDiag_48[21] , \wNDiag_48[20] , 
        \wNDiag_48[19] , \wNDiag_48[18] , \wNDiag_48[17] , \wNDiag_48[16] , 
        \wNDiag_48[15] , \wNDiag_48[14] , \wNDiag_48[13] , \wNDiag_48[12] , 
        \wNDiag_48[11] , \wNDiag_48[10] , \wNDiag_48[9] , \wNDiag_48[8] , 
        \wNDiag_48[7] , \wNDiag_48[6] , \wNDiag_48[5] , \wNDiag_48[4] , 
        \wNDiag_48[3] , \wNDiag_48[2] , \wNDiag_48[1] , \wNDiag_48[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_60 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_61[6] , \wScan_61[5] , \wScan_61[4] , 
        \wScan_61[3] , \wScan_61[2] , \wScan_61[1] , \wScan_61[0] }), 
        .ScanOut({\wScan_60[6] , \wScan_60[5] , \wScan_60[4] , \wScan_60[3] , 
        \wScan_60[2] , \wScan_60[1] , \wScan_60[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_60[0] ), .ReturnIn(\wReturn_61[0] ), .ColIn({
        \wColumn_60[63] , \wColumn_60[62] , \wColumn_60[61] , \wColumn_60[60] , 
        \wColumn_60[59] , \wColumn_60[58] , \wColumn_60[57] , \wColumn_60[56] , 
        \wColumn_60[55] , \wColumn_60[54] , \wColumn_60[53] , \wColumn_60[52] , 
        \wColumn_60[51] , \wColumn_60[50] , \wColumn_60[49] , \wColumn_60[48] , 
        \wColumn_60[47] , \wColumn_60[46] , \wColumn_60[45] , \wColumn_60[44] , 
        \wColumn_60[43] , \wColumn_60[42] , \wColumn_60[41] , \wColumn_60[40] , 
        \wColumn_60[39] , \wColumn_60[38] , \wColumn_60[37] , \wColumn_60[36] , 
        \wColumn_60[35] , \wColumn_60[34] , \wColumn_60[33] , \wColumn_60[32] , 
        \wColumn_60[31] , \wColumn_60[30] , \wColumn_60[29] , \wColumn_60[28] , 
        \wColumn_60[27] , \wColumn_60[26] , \wColumn_60[25] , \wColumn_60[24] , 
        \wColumn_60[23] , \wColumn_60[22] , \wColumn_60[21] , \wColumn_60[20] , 
        \wColumn_60[19] , \wColumn_60[18] , \wColumn_60[17] , \wColumn_60[16] , 
        \wColumn_60[15] , \wColumn_60[14] , \wColumn_60[13] , \wColumn_60[12] , 
        \wColumn_60[11] , \wColumn_60[10] , \wColumn_60[9] , \wColumn_60[8] , 
        \wColumn_60[7] , \wColumn_60[6] , \wColumn_60[5] , \wColumn_60[4] , 
        \wColumn_60[3] , \wColumn_60[2] , \wColumn_60[1] , \wColumn_60[0] }), 
        .PDiagIn({\wPDiag_60[63] , \wPDiag_60[62] , \wPDiag_60[61] , 
        \wPDiag_60[60] , \wPDiag_60[59] , \wPDiag_60[58] , \wPDiag_60[57] , 
        \wPDiag_60[56] , \wPDiag_60[55] , \wPDiag_60[54] , \wPDiag_60[53] , 
        \wPDiag_60[52] , \wPDiag_60[51] , \wPDiag_60[50] , \wPDiag_60[49] , 
        \wPDiag_60[48] , \wPDiag_60[47] , \wPDiag_60[46] , \wPDiag_60[45] , 
        \wPDiag_60[44] , \wPDiag_60[43] , \wPDiag_60[42] , \wPDiag_60[41] , 
        \wPDiag_60[40] , \wPDiag_60[39] , \wPDiag_60[38] , \wPDiag_60[37] , 
        \wPDiag_60[36] , \wPDiag_60[35] , \wPDiag_60[34] , \wPDiag_60[33] , 
        \wPDiag_60[32] , \wPDiag_60[31] , \wPDiag_60[30] , \wPDiag_60[29] , 
        \wPDiag_60[28] , \wPDiag_60[27] , \wPDiag_60[26] , \wPDiag_60[25] , 
        \wPDiag_60[24] , \wPDiag_60[23] , \wPDiag_60[22] , \wPDiag_60[21] , 
        \wPDiag_60[20] , \wPDiag_60[19] , \wPDiag_60[18] , \wPDiag_60[17] , 
        \wPDiag_60[16] , \wPDiag_60[15] , \wPDiag_60[14] , \wPDiag_60[13] , 
        \wPDiag_60[12] , \wPDiag_60[11] , \wPDiag_60[10] , \wPDiag_60[9] , 
        \wPDiag_60[8] , \wPDiag_60[7] , \wPDiag_60[6] , \wPDiag_60[5] , 
        \wPDiag_60[4] , \wPDiag_60[3] , \wPDiag_60[2] , \wPDiag_60[1] , 
        \wPDiag_60[0] }), .NDiagIn({\wNDiag_60[63] , \wNDiag_60[62] , 
        \wNDiag_60[61] , \wNDiag_60[60] , \wNDiag_60[59] , \wNDiag_60[58] , 
        \wNDiag_60[57] , \wNDiag_60[56] , \wNDiag_60[55] , \wNDiag_60[54] , 
        \wNDiag_60[53] , \wNDiag_60[52] , \wNDiag_60[51] , \wNDiag_60[50] , 
        \wNDiag_60[49] , \wNDiag_60[48] , \wNDiag_60[47] , \wNDiag_60[46] , 
        \wNDiag_60[45] , \wNDiag_60[44] , \wNDiag_60[43] , \wNDiag_60[42] , 
        \wNDiag_60[41] , \wNDiag_60[40] , \wNDiag_60[39] , \wNDiag_60[38] , 
        \wNDiag_60[37] , \wNDiag_60[36] , \wNDiag_60[35] , \wNDiag_60[34] , 
        \wNDiag_60[33] , \wNDiag_60[32] , \wNDiag_60[31] , \wNDiag_60[30] , 
        \wNDiag_60[29] , \wNDiag_60[28] , \wNDiag_60[27] , \wNDiag_60[26] , 
        \wNDiag_60[25] , \wNDiag_60[24] , \wNDiag_60[23] , \wNDiag_60[22] , 
        \wNDiag_60[21] , \wNDiag_60[20] , \wNDiag_60[19] , \wNDiag_60[18] , 
        \wNDiag_60[17] , \wNDiag_60[16] , \wNDiag_60[15] , \wNDiag_60[14] , 
        \wNDiag_60[13] , \wNDiag_60[12] , \wNDiag_60[11] , \wNDiag_60[10] , 
        \wNDiag_60[9] , \wNDiag_60[8] , \wNDiag_60[7] , \wNDiag_60[6] , 
        \wNDiag_60[5] , \wNDiag_60[4] , \wNDiag_60[3] , \wNDiag_60[2] , 
        \wNDiag_60[1] , \wNDiag_60[0] }), .CallOut(\wCall_61[0] ), .ReturnOut(
        \wReturn_60[0] ), .ColOut({\wColumn_61[63] , \wColumn_61[62] , 
        \wColumn_61[61] , \wColumn_61[60] , \wColumn_61[59] , \wColumn_61[58] , 
        \wColumn_61[57] , \wColumn_61[56] , \wColumn_61[55] , \wColumn_61[54] , 
        \wColumn_61[53] , \wColumn_61[52] , \wColumn_61[51] , \wColumn_61[50] , 
        \wColumn_61[49] , \wColumn_61[48] , \wColumn_61[47] , \wColumn_61[46] , 
        \wColumn_61[45] , \wColumn_61[44] , \wColumn_61[43] , \wColumn_61[42] , 
        \wColumn_61[41] , \wColumn_61[40] , \wColumn_61[39] , \wColumn_61[38] , 
        \wColumn_61[37] , \wColumn_61[36] , \wColumn_61[35] , \wColumn_61[34] , 
        \wColumn_61[33] , \wColumn_61[32] , \wColumn_61[31] , \wColumn_61[30] , 
        \wColumn_61[29] , \wColumn_61[28] , \wColumn_61[27] , \wColumn_61[26] , 
        \wColumn_61[25] , \wColumn_61[24] , \wColumn_61[23] , \wColumn_61[22] , 
        \wColumn_61[21] , \wColumn_61[20] , \wColumn_61[19] , \wColumn_61[18] , 
        \wColumn_61[17] , \wColumn_61[16] , \wColumn_61[15] , \wColumn_61[14] , 
        \wColumn_61[13] , \wColumn_61[12] , \wColumn_61[11] , \wColumn_61[10] , 
        \wColumn_61[9] , \wColumn_61[8] , \wColumn_61[7] , \wColumn_61[6] , 
        \wColumn_61[5] , \wColumn_61[4] , \wColumn_61[3] , \wColumn_61[2] , 
        \wColumn_61[1] , \wColumn_61[0] }), .PDiagOut({\wPDiag_61[63] , 
        \wPDiag_61[62] , \wPDiag_61[61] , \wPDiag_61[60] , \wPDiag_61[59] , 
        \wPDiag_61[58] , \wPDiag_61[57] , \wPDiag_61[56] , \wPDiag_61[55] , 
        \wPDiag_61[54] , \wPDiag_61[53] , \wPDiag_61[52] , \wPDiag_61[51] , 
        \wPDiag_61[50] , \wPDiag_61[49] , \wPDiag_61[48] , \wPDiag_61[47] , 
        \wPDiag_61[46] , \wPDiag_61[45] , \wPDiag_61[44] , \wPDiag_61[43] , 
        \wPDiag_61[42] , \wPDiag_61[41] , \wPDiag_61[40] , \wPDiag_61[39] , 
        \wPDiag_61[38] , \wPDiag_61[37] , \wPDiag_61[36] , \wPDiag_61[35] , 
        \wPDiag_61[34] , \wPDiag_61[33] , \wPDiag_61[32] , \wPDiag_61[31] , 
        \wPDiag_61[30] , \wPDiag_61[29] , \wPDiag_61[28] , \wPDiag_61[27] , 
        \wPDiag_61[26] , \wPDiag_61[25] , \wPDiag_61[24] , \wPDiag_61[23] , 
        \wPDiag_61[22] , \wPDiag_61[21] , \wPDiag_61[20] , \wPDiag_61[19] , 
        \wPDiag_61[18] , \wPDiag_61[17] , \wPDiag_61[16] , \wPDiag_61[15] , 
        \wPDiag_61[14] , \wPDiag_61[13] , \wPDiag_61[12] , \wPDiag_61[11] , 
        \wPDiag_61[10] , \wPDiag_61[9] , \wPDiag_61[8] , \wPDiag_61[7] , 
        \wPDiag_61[6] , \wPDiag_61[5] , \wPDiag_61[4] , \wPDiag_61[3] , 
        \wPDiag_61[2] , \wPDiag_61[1] , \wPDiag_61[0] }), .NDiagOut({
        \wNDiag_61[63] , \wNDiag_61[62] , \wNDiag_61[61] , \wNDiag_61[60] , 
        \wNDiag_61[59] , \wNDiag_61[58] , \wNDiag_61[57] , \wNDiag_61[56] , 
        \wNDiag_61[55] , \wNDiag_61[54] , \wNDiag_61[53] , \wNDiag_61[52] , 
        \wNDiag_61[51] , \wNDiag_61[50] , \wNDiag_61[49] , \wNDiag_61[48] , 
        \wNDiag_61[47] , \wNDiag_61[46] , \wNDiag_61[45] , \wNDiag_61[44] , 
        \wNDiag_61[43] , \wNDiag_61[42] , \wNDiag_61[41] , \wNDiag_61[40] , 
        \wNDiag_61[39] , \wNDiag_61[38] , \wNDiag_61[37] , \wNDiag_61[36] , 
        \wNDiag_61[35] , \wNDiag_61[34] , \wNDiag_61[33] , \wNDiag_61[32] , 
        \wNDiag_61[31] , \wNDiag_61[30] , \wNDiag_61[29] , \wNDiag_61[28] , 
        \wNDiag_61[27] , \wNDiag_61[26] , \wNDiag_61[25] , \wNDiag_61[24] , 
        \wNDiag_61[23] , \wNDiag_61[22] , \wNDiag_61[21] , \wNDiag_61[20] , 
        \wNDiag_61[19] , \wNDiag_61[18] , \wNDiag_61[17] , \wNDiag_61[16] , 
        \wNDiag_61[15] , \wNDiag_61[14] , \wNDiag_61[13] , \wNDiag_61[12] , 
        \wNDiag_61[11] , \wNDiag_61[10] , \wNDiag_61[9] , \wNDiag_61[8] , 
        \wNDiag_61[7] , \wNDiag_61[6] , \wNDiag_61[5] , \wNDiag_61[4] , 
        \wNDiag_61[3] , \wNDiag_61[2] , \wNDiag_61[1] , \wNDiag_61[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_13 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_14[6] , \wScan_14[5] , \wScan_14[4] , 
        \wScan_14[3] , \wScan_14[2] , \wScan_14[1] , \wScan_14[0] }), 
        .ScanOut({\wScan_13[6] , \wScan_13[5] , \wScan_13[4] , \wScan_13[3] , 
        \wScan_13[2] , \wScan_13[1] , \wScan_13[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_13[0] ), .ReturnIn(\wReturn_14[0] ), .ColIn({
        \wColumn_13[63] , \wColumn_13[62] , \wColumn_13[61] , \wColumn_13[60] , 
        \wColumn_13[59] , \wColumn_13[58] , \wColumn_13[57] , \wColumn_13[56] , 
        \wColumn_13[55] , \wColumn_13[54] , \wColumn_13[53] , \wColumn_13[52] , 
        \wColumn_13[51] , \wColumn_13[50] , \wColumn_13[49] , \wColumn_13[48] , 
        \wColumn_13[47] , \wColumn_13[46] , \wColumn_13[45] , \wColumn_13[44] , 
        \wColumn_13[43] , \wColumn_13[42] , \wColumn_13[41] , \wColumn_13[40] , 
        \wColumn_13[39] , \wColumn_13[38] , \wColumn_13[37] , \wColumn_13[36] , 
        \wColumn_13[35] , \wColumn_13[34] , \wColumn_13[33] , \wColumn_13[32] , 
        \wColumn_13[31] , \wColumn_13[30] , \wColumn_13[29] , \wColumn_13[28] , 
        \wColumn_13[27] , \wColumn_13[26] , \wColumn_13[25] , \wColumn_13[24] , 
        \wColumn_13[23] , \wColumn_13[22] , \wColumn_13[21] , \wColumn_13[20] , 
        \wColumn_13[19] , \wColumn_13[18] , \wColumn_13[17] , \wColumn_13[16] , 
        \wColumn_13[15] , \wColumn_13[14] , \wColumn_13[13] , \wColumn_13[12] , 
        \wColumn_13[11] , \wColumn_13[10] , \wColumn_13[9] , \wColumn_13[8] , 
        \wColumn_13[7] , \wColumn_13[6] , \wColumn_13[5] , \wColumn_13[4] , 
        \wColumn_13[3] , \wColumn_13[2] , \wColumn_13[1] , \wColumn_13[0] }), 
        .PDiagIn({\wPDiag_13[63] , \wPDiag_13[62] , \wPDiag_13[61] , 
        \wPDiag_13[60] , \wPDiag_13[59] , \wPDiag_13[58] , \wPDiag_13[57] , 
        \wPDiag_13[56] , \wPDiag_13[55] , \wPDiag_13[54] , \wPDiag_13[53] , 
        \wPDiag_13[52] , \wPDiag_13[51] , \wPDiag_13[50] , \wPDiag_13[49] , 
        \wPDiag_13[48] , \wPDiag_13[47] , \wPDiag_13[46] , \wPDiag_13[45] , 
        \wPDiag_13[44] , \wPDiag_13[43] , \wPDiag_13[42] , \wPDiag_13[41] , 
        \wPDiag_13[40] , \wPDiag_13[39] , \wPDiag_13[38] , \wPDiag_13[37] , 
        \wPDiag_13[36] , \wPDiag_13[35] , \wPDiag_13[34] , \wPDiag_13[33] , 
        \wPDiag_13[32] , \wPDiag_13[31] , \wPDiag_13[30] , \wPDiag_13[29] , 
        \wPDiag_13[28] , \wPDiag_13[27] , \wPDiag_13[26] , \wPDiag_13[25] , 
        \wPDiag_13[24] , \wPDiag_13[23] , \wPDiag_13[22] , \wPDiag_13[21] , 
        \wPDiag_13[20] , \wPDiag_13[19] , \wPDiag_13[18] , \wPDiag_13[17] , 
        \wPDiag_13[16] , \wPDiag_13[15] , \wPDiag_13[14] , \wPDiag_13[13] , 
        \wPDiag_13[12] , \wPDiag_13[11] , \wPDiag_13[10] , \wPDiag_13[9] , 
        \wPDiag_13[8] , \wPDiag_13[7] , \wPDiag_13[6] , \wPDiag_13[5] , 
        \wPDiag_13[4] , \wPDiag_13[3] , \wPDiag_13[2] , \wPDiag_13[1] , 
        \wPDiag_13[0] }), .NDiagIn({\wNDiag_13[63] , \wNDiag_13[62] , 
        \wNDiag_13[61] , \wNDiag_13[60] , \wNDiag_13[59] , \wNDiag_13[58] , 
        \wNDiag_13[57] , \wNDiag_13[56] , \wNDiag_13[55] , \wNDiag_13[54] , 
        \wNDiag_13[53] , \wNDiag_13[52] , \wNDiag_13[51] , \wNDiag_13[50] , 
        \wNDiag_13[49] , \wNDiag_13[48] , \wNDiag_13[47] , \wNDiag_13[46] , 
        \wNDiag_13[45] , \wNDiag_13[44] , \wNDiag_13[43] , \wNDiag_13[42] , 
        \wNDiag_13[41] , \wNDiag_13[40] , \wNDiag_13[39] , \wNDiag_13[38] , 
        \wNDiag_13[37] , \wNDiag_13[36] , \wNDiag_13[35] , \wNDiag_13[34] , 
        \wNDiag_13[33] , \wNDiag_13[32] , \wNDiag_13[31] , \wNDiag_13[30] , 
        \wNDiag_13[29] , \wNDiag_13[28] , \wNDiag_13[27] , \wNDiag_13[26] , 
        \wNDiag_13[25] , \wNDiag_13[24] , \wNDiag_13[23] , \wNDiag_13[22] , 
        \wNDiag_13[21] , \wNDiag_13[20] , \wNDiag_13[19] , \wNDiag_13[18] , 
        \wNDiag_13[17] , \wNDiag_13[16] , \wNDiag_13[15] , \wNDiag_13[14] , 
        \wNDiag_13[13] , \wNDiag_13[12] , \wNDiag_13[11] , \wNDiag_13[10] , 
        \wNDiag_13[9] , \wNDiag_13[8] , \wNDiag_13[7] , \wNDiag_13[6] , 
        \wNDiag_13[5] , \wNDiag_13[4] , \wNDiag_13[3] , \wNDiag_13[2] , 
        \wNDiag_13[1] , \wNDiag_13[0] }), .CallOut(\wCall_14[0] ), .ReturnOut(
        \wReturn_13[0] ), .ColOut({\wColumn_14[63] , \wColumn_14[62] , 
        \wColumn_14[61] , \wColumn_14[60] , \wColumn_14[59] , \wColumn_14[58] , 
        \wColumn_14[57] , \wColumn_14[56] , \wColumn_14[55] , \wColumn_14[54] , 
        \wColumn_14[53] , \wColumn_14[52] , \wColumn_14[51] , \wColumn_14[50] , 
        \wColumn_14[49] , \wColumn_14[48] , \wColumn_14[47] , \wColumn_14[46] , 
        \wColumn_14[45] , \wColumn_14[44] , \wColumn_14[43] , \wColumn_14[42] , 
        \wColumn_14[41] , \wColumn_14[40] , \wColumn_14[39] , \wColumn_14[38] , 
        \wColumn_14[37] , \wColumn_14[36] , \wColumn_14[35] , \wColumn_14[34] , 
        \wColumn_14[33] , \wColumn_14[32] , \wColumn_14[31] , \wColumn_14[30] , 
        \wColumn_14[29] , \wColumn_14[28] , \wColumn_14[27] , \wColumn_14[26] , 
        \wColumn_14[25] , \wColumn_14[24] , \wColumn_14[23] , \wColumn_14[22] , 
        \wColumn_14[21] , \wColumn_14[20] , \wColumn_14[19] , \wColumn_14[18] , 
        \wColumn_14[17] , \wColumn_14[16] , \wColumn_14[15] , \wColumn_14[14] , 
        \wColumn_14[13] , \wColumn_14[12] , \wColumn_14[11] , \wColumn_14[10] , 
        \wColumn_14[9] , \wColumn_14[8] , \wColumn_14[7] , \wColumn_14[6] , 
        \wColumn_14[5] , \wColumn_14[4] , \wColumn_14[3] , \wColumn_14[2] , 
        \wColumn_14[1] , \wColumn_14[0] }), .PDiagOut({\wPDiag_14[63] , 
        \wPDiag_14[62] , \wPDiag_14[61] , \wPDiag_14[60] , \wPDiag_14[59] , 
        \wPDiag_14[58] , \wPDiag_14[57] , \wPDiag_14[56] , \wPDiag_14[55] , 
        \wPDiag_14[54] , \wPDiag_14[53] , \wPDiag_14[52] , \wPDiag_14[51] , 
        \wPDiag_14[50] , \wPDiag_14[49] , \wPDiag_14[48] , \wPDiag_14[47] , 
        \wPDiag_14[46] , \wPDiag_14[45] , \wPDiag_14[44] , \wPDiag_14[43] , 
        \wPDiag_14[42] , \wPDiag_14[41] , \wPDiag_14[40] , \wPDiag_14[39] , 
        \wPDiag_14[38] , \wPDiag_14[37] , \wPDiag_14[36] , \wPDiag_14[35] , 
        \wPDiag_14[34] , \wPDiag_14[33] , \wPDiag_14[32] , \wPDiag_14[31] , 
        \wPDiag_14[30] , \wPDiag_14[29] , \wPDiag_14[28] , \wPDiag_14[27] , 
        \wPDiag_14[26] , \wPDiag_14[25] , \wPDiag_14[24] , \wPDiag_14[23] , 
        \wPDiag_14[22] , \wPDiag_14[21] , \wPDiag_14[20] , \wPDiag_14[19] , 
        \wPDiag_14[18] , \wPDiag_14[17] , \wPDiag_14[16] , \wPDiag_14[15] , 
        \wPDiag_14[14] , \wPDiag_14[13] , \wPDiag_14[12] , \wPDiag_14[11] , 
        \wPDiag_14[10] , \wPDiag_14[9] , \wPDiag_14[8] , \wPDiag_14[7] , 
        \wPDiag_14[6] , \wPDiag_14[5] , \wPDiag_14[4] , \wPDiag_14[3] , 
        \wPDiag_14[2] , \wPDiag_14[1] , \wPDiag_14[0] }), .NDiagOut({
        \wNDiag_14[63] , \wNDiag_14[62] , \wNDiag_14[61] , \wNDiag_14[60] , 
        \wNDiag_14[59] , \wNDiag_14[58] , \wNDiag_14[57] , \wNDiag_14[56] , 
        \wNDiag_14[55] , \wNDiag_14[54] , \wNDiag_14[53] , \wNDiag_14[52] , 
        \wNDiag_14[51] , \wNDiag_14[50] , \wNDiag_14[49] , \wNDiag_14[48] , 
        \wNDiag_14[47] , \wNDiag_14[46] , \wNDiag_14[45] , \wNDiag_14[44] , 
        \wNDiag_14[43] , \wNDiag_14[42] , \wNDiag_14[41] , \wNDiag_14[40] , 
        \wNDiag_14[39] , \wNDiag_14[38] , \wNDiag_14[37] , \wNDiag_14[36] , 
        \wNDiag_14[35] , \wNDiag_14[34] , \wNDiag_14[33] , \wNDiag_14[32] , 
        \wNDiag_14[31] , \wNDiag_14[30] , \wNDiag_14[29] , \wNDiag_14[28] , 
        \wNDiag_14[27] , \wNDiag_14[26] , \wNDiag_14[25] , \wNDiag_14[24] , 
        \wNDiag_14[23] , \wNDiag_14[22] , \wNDiag_14[21] , \wNDiag_14[20] , 
        \wNDiag_14[19] , \wNDiag_14[18] , \wNDiag_14[17] , \wNDiag_14[16] , 
        \wNDiag_14[15] , \wNDiag_14[14] , \wNDiag_14[13] , \wNDiag_14[12] , 
        \wNDiag_14[11] , \wNDiag_14[10] , \wNDiag_14[9] , \wNDiag_14[8] , 
        \wNDiag_14[7] , \wNDiag_14[6] , \wNDiag_14[5] , \wNDiag_14[4] , 
        \wNDiag_14[3] , \wNDiag_14[2] , \wNDiag_14[1] , \wNDiag_14[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_14 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_15[6] , \wScan_15[5] , \wScan_15[4] , 
        \wScan_15[3] , \wScan_15[2] , \wScan_15[1] , \wScan_15[0] }), 
        .ScanOut({\wScan_14[6] , \wScan_14[5] , \wScan_14[4] , \wScan_14[3] , 
        \wScan_14[2] , \wScan_14[1] , \wScan_14[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_14[0] ), .ReturnIn(\wReturn_15[0] ), .ColIn({
        \wColumn_14[63] , \wColumn_14[62] , \wColumn_14[61] , \wColumn_14[60] , 
        \wColumn_14[59] , \wColumn_14[58] , \wColumn_14[57] , \wColumn_14[56] , 
        \wColumn_14[55] , \wColumn_14[54] , \wColumn_14[53] , \wColumn_14[52] , 
        \wColumn_14[51] , \wColumn_14[50] , \wColumn_14[49] , \wColumn_14[48] , 
        \wColumn_14[47] , \wColumn_14[46] , \wColumn_14[45] , \wColumn_14[44] , 
        \wColumn_14[43] , \wColumn_14[42] , \wColumn_14[41] , \wColumn_14[40] , 
        \wColumn_14[39] , \wColumn_14[38] , \wColumn_14[37] , \wColumn_14[36] , 
        \wColumn_14[35] , \wColumn_14[34] , \wColumn_14[33] , \wColumn_14[32] , 
        \wColumn_14[31] , \wColumn_14[30] , \wColumn_14[29] , \wColumn_14[28] , 
        \wColumn_14[27] , \wColumn_14[26] , \wColumn_14[25] , \wColumn_14[24] , 
        \wColumn_14[23] , \wColumn_14[22] , \wColumn_14[21] , \wColumn_14[20] , 
        \wColumn_14[19] , \wColumn_14[18] , \wColumn_14[17] , \wColumn_14[16] , 
        \wColumn_14[15] , \wColumn_14[14] , \wColumn_14[13] , \wColumn_14[12] , 
        \wColumn_14[11] , \wColumn_14[10] , \wColumn_14[9] , \wColumn_14[8] , 
        \wColumn_14[7] , \wColumn_14[6] , \wColumn_14[5] , \wColumn_14[4] , 
        \wColumn_14[3] , \wColumn_14[2] , \wColumn_14[1] , \wColumn_14[0] }), 
        .PDiagIn({\wPDiag_14[63] , \wPDiag_14[62] , \wPDiag_14[61] , 
        \wPDiag_14[60] , \wPDiag_14[59] , \wPDiag_14[58] , \wPDiag_14[57] , 
        \wPDiag_14[56] , \wPDiag_14[55] , \wPDiag_14[54] , \wPDiag_14[53] , 
        \wPDiag_14[52] , \wPDiag_14[51] , \wPDiag_14[50] , \wPDiag_14[49] , 
        \wPDiag_14[48] , \wPDiag_14[47] , \wPDiag_14[46] , \wPDiag_14[45] , 
        \wPDiag_14[44] , \wPDiag_14[43] , \wPDiag_14[42] , \wPDiag_14[41] , 
        \wPDiag_14[40] , \wPDiag_14[39] , \wPDiag_14[38] , \wPDiag_14[37] , 
        \wPDiag_14[36] , \wPDiag_14[35] , \wPDiag_14[34] , \wPDiag_14[33] , 
        \wPDiag_14[32] , \wPDiag_14[31] , \wPDiag_14[30] , \wPDiag_14[29] , 
        \wPDiag_14[28] , \wPDiag_14[27] , \wPDiag_14[26] , \wPDiag_14[25] , 
        \wPDiag_14[24] , \wPDiag_14[23] , \wPDiag_14[22] , \wPDiag_14[21] , 
        \wPDiag_14[20] , \wPDiag_14[19] , \wPDiag_14[18] , \wPDiag_14[17] , 
        \wPDiag_14[16] , \wPDiag_14[15] , \wPDiag_14[14] , \wPDiag_14[13] , 
        \wPDiag_14[12] , \wPDiag_14[11] , \wPDiag_14[10] , \wPDiag_14[9] , 
        \wPDiag_14[8] , \wPDiag_14[7] , \wPDiag_14[6] , \wPDiag_14[5] , 
        \wPDiag_14[4] , \wPDiag_14[3] , \wPDiag_14[2] , \wPDiag_14[1] , 
        \wPDiag_14[0] }), .NDiagIn({\wNDiag_14[63] , \wNDiag_14[62] , 
        \wNDiag_14[61] , \wNDiag_14[60] , \wNDiag_14[59] , \wNDiag_14[58] , 
        \wNDiag_14[57] , \wNDiag_14[56] , \wNDiag_14[55] , \wNDiag_14[54] , 
        \wNDiag_14[53] , \wNDiag_14[52] , \wNDiag_14[51] , \wNDiag_14[50] , 
        \wNDiag_14[49] , \wNDiag_14[48] , \wNDiag_14[47] , \wNDiag_14[46] , 
        \wNDiag_14[45] , \wNDiag_14[44] , \wNDiag_14[43] , \wNDiag_14[42] , 
        \wNDiag_14[41] , \wNDiag_14[40] , \wNDiag_14[39] , \wNDiag_14[38] , 
        \wNDiag_14[37] , \wNDiag_14[36] , \wNDiag_14[35] , \wNDiag_14[34] , 
        \wNDiag_14[33] , \wNDiag_14[32] , \wNDiag_14[31] , \wNDiag_14[30] , 
        \wNDiag_14[29] , \wNDiag_14[28] , \wNDiag_14[27] , \wNDiag_14[26] , 
        \wNDiag_14[25] , \wNDiag_14[24] , \wNDiag_14[23] , \wNDiag_14[22] , 
        \wNDiag_14[21] , \wNDiag_14[20] , \wNDiag_14[19] , \wNDiag_14[18] , 
        \wNDiag_14[17] , \wNDiag_14[16] , \wNDiag_14[15] , \wNDiag_14[14] , 
        \wNDiag_14[13] , \wNDiag_14[12] , \wNDiag_14[11] , \wNDiag_14[10] , 
        \wNDiag_14[9] , \wNDiag_14[8] , \wNDiag_14[7] , \wNDiag_14[6] , 
        \wNDiag_14[5] , \wNDiag_14[4] , \wNDiag_14[3] , \wNDiag_14[2] , 
        \wNDiag_14[1] , \wNDiag_14[0] }), .CallOut(\wCall_15[0] ), .ReturnOut(
        \wReturn_14[0] ), .ColOut({\wColumn_15[63] , \wColumn_15[62] , 
        \wColumn_15[61] , \wColumn_15[60] , \wColumn_15[59] , \wColumn_15[58] , 
        \wColumn_15[57] , \wColumn_15[56] , \wColumn_15[55] , \wColumn_15[54] , 
        \wColumn_15[53] , \wColumn_15[52] , \wColumn_15[51] , \wColumn_15[50] , 
        \wColumn_15[49] , \wColumn_15[48] , \wColumn_15[47] , \wColumn_15[46] , 
        \wColumn_15[45] , \wColumn_15[44] , \wColumn_15[43] , \wColumn_15[42] , 
        \wColumn_15[41] , \wColumn_15[40] , \wColumn_15[39] , \wColumn_15[38] , 
        \wColumn_15[37] , \wColumn_15[36] , \wColumn_15[35] , \wColumn_15[34] , 
        \wColumn_15[33] , \wColumn_15[32] , \wColumn_15[31] , \wColumn_15[30] , 
        \wColumn_15[29] , \wColumn_15[28] , \wColumn_15[27] , \wColumn_15[26] , 
        \wColumn_15[25] , \wColumn_15[24] , \wColumn_15[23] , \wColumn_15[22] , 
        \wColumn_15[21] , \wColumn_15[20] , \wColumn_15[19] , \wColumn_15[18] , 
        \wColumn_15[17] , \wColumn_15[16] , \wColumn_15[15] , \wColumn_15[14] , 
        \wColumn_15[13] , \wColumn_15[12] , \wColumn_15[11] , \wColumn_15[10] , 
        \wColumn_15[9] , \wColumn_15[8] , \wColumn_15[7] , \wColumn_15[6] , 
        \wColumn_15[5] , \wColumn_15[4] , \wColumn_15[3] , \wColumn_15[2] , 
        \wColumn_15[1] , \wColumn_15[0] }), .PDiagOut({\wPDiag_15[63] , 
        \wPDiag_15[62] , \wPDiag_15[61] , \wPDiag_15[60] , \wPDiag_15[59] , 
        \wPDiag_15[58] , \wPDiag_15[57] , \wPDiag_15[56] , \wPDiag_15[55] , 
        \wPDiag_15[54] , \wPDiag_15[53] , \wPDiag_15[52] , \wPDiag_15[51] , 
        \wPDiag_15[50] , \wPDiag_15[49] , \wPDiag_15[48] , \wPDiag_15[47] , 
        \wPDiag_15[46] , \wPDiag_15[45] , \wPDiag_15[44] , \wPDiag_15[43] , 
        \wPDiag_15[42] , \wPDiag_15[41] , \wPDiag_15[40] , \wPDiag_15[39] , 
        \wPDiag_15[38] , \wPDiag_15[37] , \wPDiag_15[36] , \wPDiag_15[35] , 
        \wPDiag_15[34] , \wPDiag_15[33] , \wPDiag_15[32] , \wPDiag_15[31] , 
        \wPDiag_15[30] , \wPDiag_15[29] , \wPDiag_15[28] , \wPDiag_15[27] , 
        \wPDiag_15[26] , \wPDiag_15[25] , \wPDiag_15[24] , \wPDiag_15[23] , 
        \wPDiag_15[22] , \wPDiag_15[21] , \wPDiag_15[20] , \wPDiag_15[19] , 
        \wPDiag_15[18] , \wPDiag_15[17] , \wPDiag_15[16] , \wPDiag_15[15] , 
        \wPDiag_15[14] , \wPDiag_15[13] , \wPDiag_15[12] , \wPDiag_15[11] , 
        \wPDiag_15[10] , \wPDiag_15[9] , \wPDiag_15[8] , \wPDiag_15[7] , 
        \wPDiag_15[6] , \wPDiag_15[5] , \wPDiag_15[4] , \wPDiag_15[3] , 
        \wPDiag_15[2] , \wPDiag_15[1] , \wPDiag_15[0] }), .NDiagOut({
        \wNDiag_15[63] , \wNDiag_15[62] , \wNDiag_15[61] , \wNDiag_15[60] , 
        \wNDiag_15[59] , \wNDiag_15[58] , \wNDiag_15[57] , \wNDiag_15[56] , 
        \wNDiag_15[55] , \wNDiag_15[54] , \wNDiag_15[53] , \wNDiag_15[52] , 
        \wNDiag_15[51] , \wNDiag_15[50] , \wNDiag_15[49] , \wNDiag_15[48] , 
        \wNDiag_15[47] , \wNDiag_15[46] , \wNDiag_15[45] , \wNDiag_15[44] , 
        \wNDiag_15[43] , \wNDiag_15[42] , \wNDiag_15[41] , \wNDiag_15[40] , 
        \wNDiag_15[39] , \wNDiag_15[38] , \wNDiag_15[37] , \wNDiag_15[36] , 
        \wNDiag_15[35] , \wNDiag_15[34] , \wNDiag_15[33] , \wNDiag_15[32] , 
        \wNDiag_15[31] , \wNDiag_15[30] , \wNDiag_15[29] , \wNDiag_15[28] , 
        \wNDiag_15[27] , \wNDiag_15[26] , \wNDiag_15[25] , \wNDiag_15[24] , 
        \wNDiag_15[23] , \wNDiag_15[22] , \wNDiag_15[21] , \wNDiag_15[20] , 
        \wNDiag_15[19] , \wNDiag_15[18] , \wNDiag_15[17] , \wNDiag_15[16] , 
        \wNDiag_15[15] , \wNDiag_15[14] , \wNDiag_15[13] , \wNDiag_15[12] , 
        \wNDiag_15[11] , \wNDiag_15[10] , \wNDiag_15[9] , \wNDiag_15[8] , 
        \wNDiag_15[7] , \wNDiag_15[6] , \wNDiag_15[5] , \wNDiag_15[4] , 
        \wNDiag_15[3] , \wNDiag_15[2] , \wNDiag_15[1] , \wNDiag_15[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_28 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_29[6] , \wScan_29[5] , \wScan_29[4] , 
        \wScan_29[3] , \wScan_29[2] , \wScan_29[1] , \wScan_29[0] }), 
        .ScanOut({\wScan_28[6] , \wScan_28[5] , \wScan_28[4] , \wScan_28[3] , 
        \wScan_28[2] , \wScan_28[1] , \wScan_28[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_28[0] ), .ReturnIn(\wReturn_29[0] ), .ColIn({
        \wColumn_28[63] , \wColumn_28[62] , \wColumn_28[61] , \wColumn_28[60] , 
        \wColumn_28[59] , \wColumn_28[58] , \wColumn_28[57] , \wColumn_28[56] , 
        \wColumn_28[55] , \wColumn_28[54] , \wColumn_28[53] , \wColumn_28[52] , 
        \wColumn_28[51] , \wColumn_28[50] , \wColumn_28[49] , \wColumn_28[48] , 
        \wColumn_28[47] , \wColumn_28[46] , \wColumn_28[45] , \wColumn_28[44] , 
        \wColumn_28[43] , \wColumn_28[42] , \wColumn_28[41] , \wColumn_28[40] , 
        \wColumn_28[39] , \wColumn_28[38] , \wColumn_28[37] , \wColumn_28[36] , 
        \wColumn_28[35] , \wColumn_28[34] , \wColumn_28[33] , \wColumn_28[32] , 
        \wColumn_28[31] , \wColumn_28[30] , \wColumn_28[29] , \wColumn_28[28] , 
        \wColumn_28[27] , \wColumn_28[26] , \wColumn_28[25] , \wColumn_28[24] , 
        \wColumn_28[23] , \wColumn_28[22] , \wColumn_28[21] , \wColumn_28[20] , 
        \wColumn_28[19] , \wColumn_28[18] , \wColumn_28[17] , \wColumn_28[16] , 
        \wColumn_28[15] , \wColumn_28[14] , \wColumn_28[13] , \wColumn_28[12] , 
        \wColumn_28[11] , \wColumn_28[10] , \wColumn_28[9] , \wColumn_28[8] , 
        \wColumn_28[7] , \wColumn_28[6] , \wColumn_28[5] , \wColumn_28[4] , 
        \wColumn_28[3] , \wColumn_28[2] , \wColumn_28[1] , \wColumn_28[0] }), 
        .PDiagIn({\wPDiag_28[63] , \wPDiag_28[62] , \wPDiag_28[61] , 
        \wPDiag_28[60] , \wPDiag_28[59] , \wPDiag_28[58] , \wPDiag_28[57] , 
        \wPDiag_28[56] , \wPDiag_28[55] , \wPDiag_28[54] , \wPDiag_28[53] , 
        \wPDiag_28[52] , \wPDiag_28[51] , \wPDiag_28[50] , \wPDiag_28[49] , 
        \wPDiag_28[48] , \wPDiag_28[47] , \wPDiag_28[46] , \wPDiag_28[45] , 
        \wPDiag_28[44] , \wPDiag_28[43] , \wPDiag_28[42] , \wPDiag_28[41] , 
        \wPDiag_28[40] , \wPDiag_28[39] , \wPDiag_28[38] , \wPDiag_28[37] , 
        \wPDiag_28[36] , \wPDiag_28[35] , \wPDiag_28[34] , \wPDiag_28[33] , 
        \wPDiag_28[32] , \wPDiag_28[31] , \wPDiag_28[30] , \wPDiag_28[29] , 
        \wPDiag_28[28] , \wPDiag_28[27] , \wPDiag_28[26] , \wPDiag_28[25] , 
        \wPDiag_28[24] , \wPDiag_28[23] , \wPDiag_28[22] , \wPDiag_28[21] , 
        \wPDiag_28[20] , \wPDiag_28[19] , \wPDiag_28[18] , \wPDiag_28[17] , 
        \wPDiag_28[16] , \wPDiag_28[15] , \wPDiag_28[14] , \wPDiag_28[13] , 
        \wPDiag_28[12] , \wPDiag_28[11] , \wPDiag_28[10] , \wPDiag_28[9] , 
        \wPDiag_28[8] , \wPDiag_28[7] , \wPDiag_28[6] , \wPDiag_28[5] , 
        \wPDiag_28[4] , \wPDiag_28[3] , \wPDiag_28[2] , \wPDiag_28[1] , 
        \wPDiag_28[0] }), .NDiagIn({\wNDiag_28[63] , \wNDiag_28[62] , 
        \wNDiag_28[61] , \wNDiag_28[60] , \wNDiag_28[59] , \wNDiag_28[58] , 
        \wNDiag_28[57] , \wNDiag_28[56] , \wNDiag_28[55] , \wNDiag_28[54] , 
        \wNDiag_28[53] , \wNDiag_28[52] , \wNDiag_28[51] , \wNDiag_28[50] , 
        \wNDiag_28[49] , \wNDiag_28[48] , \wNDiag_28[47] , \wNDiag_28[46] , 
        \wNDiag_28[45] , \wNDiag_28[44] , \wNDiag_28[43] , \wNDiag_28[42] , 
        \wNDiag_28[41] , \wNDiag_28[40] , \wNDiag_28[39] , \wNDiag_28[38] , 
        \wNDiag_28[37] , \wNDiag_28[36] , \wNDiag_28[35] , \wNDiag_28[34] , 
        \wNDiag_28[33] , \wNDiag_28[32] , \wNDiag_28[31] , \wNDiag_28[30] , 
        \wNDiag_28[29] , \wNDiag_28[28] , \wNDiag_28[27] , \wNDiag_28[26] , 
        \wNDiag_28[25] , \wNDiag_28[24] , \wNDiag_28[23] , \wNDiag_28[22] , 
        \wNDiag_28[21] , \wNDiag_28[20] , \wNDiag_28[19] , \wNDiag_28[18] , 
        \wNDiag_28[17] , \wNDiag_28[16] , \wNDiag_28[15] , \wNDiag_28[14] , 
        \wNDiag_28[13] , \wNDiag_28[12] , \wNDiag_28[11] , \wNDiag_28[10] , 
        \wNDiag_28[9] , \wNDiag_28[8] , \wNDiag_28[7] , \wNDiag_28[6] , 
        \wNDiag_28[5] , \wNDiag_28[4] , \wNDiag_28[3] , \wNDiag_28[2] , 
        \wNDiag_28[1] , \wNDiag_28[0] }), .CallOut(\wCall_29[0] ), .ReturnOut(
        \wReturn_28[0] ), .ColOut({\wColumn_29[63] , \wColumn_29[62] , 
        \wColumn_29[61] , \wColumn_29[60] , \wColumn_29[59] , \wColumn_29[58] , 
        \wColumn_29[57] , \wColumn_29[56] , \wColumn_29[55] , \wColumn_29[54] , 
        \wColumn_29[53] , \wColumn_29[52] , \wColumn_29[51] , \wColumn_29[50] , 
        \wColumn_29[49] , \wColumn_29[48] , \wColumn_29[47] , \wColumn_29[46] , 
        \wColumn_29[45] , \wColumn_29[44] , \wColumn_29[43] , \wColumn_29[42] , 
        \wColumn_29[41] , \wColumn_29[40] , \wColumn_29[39] , \wColumn_29[38] , 
        \wColumn_29[37] , \wColumn_29[36] , \wColumn_29[35] , \wColumn_29[34] , 
        \wColumn_29[33] , \wColumn_29[32] , \wColumn_29[31] , \wColumn_29[30] , 
        \wColumn_29[29] , \wColumn_29[28] , \wColumn_29[27] , \wColumn_29[26] , 
        \wColumn_29[25] , \wColumn_29[24] , \wColumn_29[23] , \wColumn_29[22] , 
        \wColumn_29[21] , \wColumn_29[20] , \wColumn_29[19] , \wColumn_29[18] , 
        \wColumn_29[17] , \wColumn_29[16] , \wColumn_29[15] , \wColumn_29[14] , 
        \wColumn_29[13] , \wColumn_29[12] , \wColumn_29[11] , \wColumn_29[10] , 
        \wColumn_29[9] , \wColumn_29[8] , \wColumn_29[7] , \wColumn_29[6] , 
        \wColumn_29[5] , \wColumn_29[4] , \wColumn_29[3] , \wColumn_29[2] , 
        \wColumn_29[1] , \wColumn_29[0] }), .PDiagOut({\wPDiag_29[63] , 
        \wPDiag_29[62] , \wPDiag_29[61] , \wPDiag_29[60] , \wPDiag_29[59] , 
        \wPDiag_29[58] , \wPDiag_29[57] , \wPDiag_29[56] , \wPDiag_29[55] , 
        \wPDiag_29[54] , \wPDiag_29[53] , \wPDiag_29[52] , \wPDiag_29[51] , 
        \wPDiag_29[50] , \wPDiag_29[49] , \wPDiag_29[48] , \wPDiag_29[47] , 
        \wPDiag_29[46] , \wPDiag_29[45] , \wPDiag_29[44] , \wPDiag_29[43] , 
        \wPDiag_29[42] , \wPDiag_29[41] , \wPDiag_29[40] , \wPDiag_29[39] , 
        \wPDiag_29[38] , \wPDiag_29[37] , \wPDiag_29[36] , \wPDiag_29[35] , 
        \wPDiag_29[34] , \wPDiag_29[33] , \wPDiag_29[32] , \wPDiag_29[31] , 
        \wPDiag_29[30] , \wPDiag_29[29] , \wPDiag_29[28] , \wPDiag_29[27] , 
        \wPDiag_29[26] , \wPDiag_29[25] , \wPDiag_29[24] , \wPDiag_29[23] , 
        \wPDiag_29[22] , \wPDiag_29[21] , \wPDiag_29[20] , \wPDiag_29[19] , 
        \wPDiag_29[18] , \wPDiag_29[17] , \wPDiag_29[16] , \wPDiag_29[15] , 
        \wPDiag_29[14] , \wPDiag_29[13] , \wPDiag_29[12] , \wPDiag_29[11] , 
        \wPDiag_29[10] , \wPDiag_29[9] , \wPDiag_29[8] , \wPDiag_29[7] , 
        \wPDiag_29[6] , \wPDiag_29[5] , \wPDiag_29[4] , \wPDiag_29[3] , 
        \wPDiag_29[2] , \wPDiag_29[1] , \wPDiag_29[0] }), .NDiagOut({
        \wNDiag_29[63] , \wNDiag_29[62] , \wNDiag_29[61] , \wNDiag_29[60] , 
        \wNDiag_29[59] , \wNDiag_29[58] , \wNDiag_29[57] , \wNDiag_29[56] , 
        \wNDiag_29[55] , \wNDiag_29[54] , \wNDiag_29[53] , \wNDiag_29[52] , 
        \wNDiag_29[51] , \wNDiag_29[50] , \wNDiag_29[49] , \wNDiag_29[48] , 
        \wNDiag_29[47] , \wNDiag_29[46] , \wNDiag_29[45] , \wNDiag_29[44] , 
        \wNDiag_29[43] , \wNDiag_29[42] , \wNDiag_29[41] , \wNDiag_29[40] , 
        \wNDiag_29[39] , \wNDiag_29[38] , \wNDiag_29[37] , \wNDiag_29[36] , 
        \wNDiag_29[35] , \wNDiag_29[34] , \wNDiag_29[33] , \wNDiag_29[32] , 
        \wNDiag_29[31] , \wNDiag_29[30] , \wNDiag_29[29] , \wNDiag_29[28] , 
        \wNDiag_29[27] , \wNDiag_29[26] , \wNDiag_29[25] , \wNDiag_29[24] , 
        \wNDiag_29[23] , \wNDiag_29[22] , \wNDiag_29[21] , \wNDiag_29[20] , 
        \wNDiag_29[19] , \wNDiag_29[18] , \wNDiag_29[17] , \wNDiag_29[16] , 
        \wNDiag_29[15] , \wNDiag_29[14] , \wNDiag_29[13] , \wNDiag_29[12] , 
        \wNDiag_29[11] , \wNDiag_29[10] , \wNDiag_29[9] , \wNDiag_29[8] , 
        \wNDiag_29[7] , \wNDiag_29[6] , \wNDiag_29[5] , \wNDiag_29[4] , 
        \wNDiag_29[3] , \wNDiag_29[2] , \wNDiag_29[1] , \wNDiag_29[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_54 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_55[6] , \wScan_55[5] , \wScan_55[4] , 
        \wScan_55[3] , \wScan_55[2] , \wScan_55[1] , \wScan_55[0] }), 
        .ScanOut({\wScan_54[6] , \wScan_54[5] , \wScan_54[4] , \wScan_54[3] , 
        \wScan_54[2] , \wScan_54[1] , \wScan_54[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_54[0] ), .ReturnIn(\wReturn_55[0] ), .ColIn({
        \wColumn_54[63] , \wColumn_54[62] , \wColumn_54[61] , \wColumn_54[60] , 
        \wColumn_54[59] , \wColumn_54[58] , \wColumn_54[57] , \wColumn_54[56] , 
        \wColumn_54[55] , \wColumn_54[54] , \wColumn_54[53] , \wColumn_54[52] , 
        \wColumn_54[51] , \wColumn_54[50] , \wColumn_54[49] , \wColumn_54[48] , 
        \wColumn_54[47] , \wColumn_54[46] , \wColumn_54[45] , \wColumn_54[44] , 
        \wColumn_54[43] , \wColumn_54[42] , \wColumn_54[41] , \wColumn_54[40] , 
        \wColumn_54[39] , \wColumn_54[38] , \wColumn_54[37] , \wColumn_54[36] , 
        \wColumn_54[35] , \wColumn_54[34] , \wColumn_54[33] , \wColumn_54[32] , 
        \wColumn_54[31] , \wColumn_54[30] , \wColumn_54[29] , \wColumn_54[28] , 
        \wColumn_54[27] , \wColumn_54[26] , \wColumn_54[25] , \wColumn_54[24] , 
        \wColumn_54[23] , \wColumn_54[22] , \wColumn_54[21] , \wColumn_54[20] , 
        \wColumn_54[19] , \wColumn_54[18] , \wColumn_54[17] , \wColumn_54[16] , 
        \wColumn_54[15] , \wColumn_54[14] , \wColumn_54[13] , \wColumn_54[12] , 
        \wColumn_54[11] , \wColumn_54[10] , \wColumn_54[9] , \wColumn_54[8] , 
        \wColumn_54[7] , \wColumn_54[6] , \wColumn_54[5] , \wColumn_54[4] , 
        \wColumn_54[3] , \wColumn_54[2] , \wColumn_54[1] , \wColumn_54[0] }), 
        .PDiagIn({\wPDiag_54[63] , \wPDiag_54[62] , \wPDiag_54[61] , 
        \wPDiag_54[60] , \wPDiag_54[59] , \wPDiag_54[58] , \wPDiag_54[57] , 
        \wPDiag_54[56] , \wPDiag_54[55] , \wPDiag_54[54] , \wPDiag_54[53] , 
        \wPDiag_54[52] , \wPDiag_54[51] , \wPDiag_54[50] , \wPDiag_54[49] , 
        \wPDiag_54[48] , \wPDiag_54[47] , \wPDiag_54[46] , \wPDiag_54[45] , 
        \wPDiag_54[44] , \wPDiag_54[43] , \wPDiag_54[42] , \wPDiag_54[41] , 
        \wPDiag_54[40] , \wPDiag_54[39] , \wPDiag_54[38] , \wPDiag_54[37] , 
        \wPDiag_54[36] , \wPDiag_54[35] , \wPDiag_54[34] , \wPDiag_54[33] , 
        \wPDiag_54[32] , \wPDiag_54[31] , \wPDiag_54[30] , \wPDiag_54[29] , 
        \wPDiag_54[28] , \wPDiag_54[27] , \wPDiag_54[26] , \wPDiag_54[25] , 
        \wPDiag_54[24] , \wPDiag_54[23] , \wPDiag_54[22] , \wPDiag_54[21] , 
        \wPDiag_54[20] , \wPDiag_54[19] , \wPDiag_54[18] , \wPDiag_54[17] , 
        \wPDiag_54[16] , \wPDiag_54[15] , \wPDiag_54[14] , \wPDiag_54[13] , 
        \wPDiag_54[12] , \wPDiag_54[11] , \wPDiag_54[10] , \wPDiag_54[9] , 
        \wPDiag_54[8] , \wPDiag_54[7] , \wPDiag_54[6] , \wPDiag_54[5] , 
        \wPDiag_54[4] , \wPDiag_54[3] , \wPDiag_54[2] , \wPDiag_54[1] , 
        \wPDiag_54[0] }), .NDiagIn({\wNDiag_54[63] , \wNDiag_54[62] , 
        \wNDiag_54[61] , \wNDiag_54[60] , \wNDiag_54[59] , \wNDiag_54[58] , 
        \wNDiag_54[57] , \wNDiag_54[56] , \wNDiag_54[55] , \wNDiag_54[54] , 
        \wNDiag_54[53] , \wNDiag_54[52] , \wNDiag_54[51] , \wNDiag_54[50] , 
        \wNDiag_54[49] , \wNDiag_54[48] , \wNDiag_54[47] , \wNDiag_54[46] , 
        \wNDiag_54[45] , \wNDiag_54[44] , \wNDiag_54[43] , \wNDiag_54[42] , 
        \wNDiag_54[41] , \wNDiag_54[40] , \wNDiag_54[39] , \wNDiag_54[38] , 
        \wNDiag_54[37] , \wNDiag_54[36] , \wNDiag_54[35] , \wNDiag_54[34] , 
        \wNDiag_54[33] , \wNDiag_54[32] , \wNDiag_54[31] , \wNDiag_54[30] , 
        \wNDiag_54[29] , \wNDiag_54[28] , \wNDiag_54[27] , \wNDiag_54[26] , 
        \wNDiag_54[25] , \wNDiag_54[24] , \wNDiag_54[23] , \wNDiag_54[22] , 
        \wNDiag_54[21] , \wNDiag_54[20] , \wNDiag_54[19] , \wNDiag_54[18] , 
        \wNDiag_54[17] , \wNDiag_54[16] , \wNDiag_54[15] , \wNDiag_54[14] , 
        \wNDiag_54[13] , \wNDiag_54[12] , \wNDiag_54[11] , \wNDiag_54[10] , 
        \wNDiag_54[9] , \wNDiag_54[8] , \wNDiag_54[7] , \wNDiag_54[6] , 
        \wNDiag_54[5] , \wNDiag_54[4] , \wNDiag_54[3] , \wNDiag_54[2] , 
        \wNDiag_54[1] , \wNDiag_54[0] }), .CallOut(\wCall_55[0] ), .ReturnOut(
        \wReturn_54[0] ), .ColOut({\wColumn_55[63] , \wColumn_55[62] , 
        \wColumn_55[61] , \wColumn_55[60] , \wColumn_55[59] , \wColumn_55[58] , 
        \wColumn_55[57] , \wColumn_55[56] , \wColumn_55[55] , \wColumn_55[54] , 
        \wColumn_55[53] , \wColumn_55[52] , \wColumn_55[51] , \wColumn_55[50] , 
        \wColumn_55[49] , \wColumn_55[48] , \wColumn_55[47] , \wColumn_55[46] , 
        \wColumn_55[45] , \wColumn_55[44] , \wColumn_55[43] , \wColumn_55[42] , 
        \wColumn_55[41] , \wColumn_55[40] , \wColumn_55[39] , \wColumn_55[38] , 
        \wColumn_55[37] , \wColumn_55[36] , \wColumn_55[35] , \wColumn_55[34] , 
        \wColumn_55[33] , \wColumn_55[32] , \wColumn_55[31] , \wColumn_55[30] , 
        \wColumn_55[29] , \wColumn_55[28] , \wColumn_55[27] , \wColumn_55[26] , 
        \wColumn_55[25] , \wColumn_55[24] , \wColumn_55[23] , \wColumn_55[22] , 
        \wColumn_55[21] , \wColumn_55[20] , \wColumn_55[19] , \wColumn_55[18] , 
        \wColumn_55[17] , \wColumn_55[16] , \wColumn_55[15] , \wColumn_55[14] , 
        \wColumn_55[13] , \wColumn_55[12] , \wColumn_55[11] , \wColumn_55[10] , 
        \wColumn_55[9] , \wColumn_55[8] , \wColumn_55[7] , \wColumn_55[6] , 
        \wColumn_55[5] , \wColumn_55[4] , \wColumn_55[3] , \wColumn_55[2] , 
        \wColumn_55[1] , \wColumn_55[0] }), .PDiagOut({\wPDiag_55[63] , 
        \wPDiag_55[62] , \wPDiag_55[61] , \wPDiag_55[60] , \wPDiag_55[59] , 
        \wPDiag_55[58] , \wPDiag_55[57] , \wPDiag_55[56] , \wPDiag_55[55] , 
        \wPDiag_55[54] , \wPDiag_55[53] , \wPDiag_55[52] , \wPDiag_55[51] , 
        \wPDiag_55[50] , \wPDiag_55[49] , \wPDiag_55[48] , \wPDiag_55[47] , 
        \wPDiag_55[46] , \wPDiag_55[45] , \wPDiag_55[44] , \wPDiag_55[43] , 
        \wPDiag_55[42] , \wPDiag_55[41] , \wPDiag_55[40] , \wPDiag_55[39] , 
        \wPDiag_55[38] , \wPDiag_55[37] , \wPDiag_55[36] , \wPDiag_55[35] , 
        \wPDiag_55[34] , \wPDiag_55[33] , \wPDiag_55[32] , \wPDiag_55[31] , 
        \wPDiag_55[30] , \wPDiag_55[29] , \wPDiag_55[28] , \wPDiag_55[27] , 
        \wPDiag_55[26] , \wPDiag_55[25] , \wPDiag_55[24] , \wPDiag_55[23] , 
        \wPDiag_55[22] , \wPDiag_55[21] , \wPDiag_55[20] , \wPDiag_55[19] , 
        \wPDiag_55[18] , \wPDiag_55[17] , \wPDiag_55[16] , \wPDiag_55[15] , 
        \wPDiag_55[14] , \wPDiag_55[13] , \wPDiag_55[12] , \wPDiag_55[11] , 
        \wPDiag_55[10] , \wPDiag_55[9] , \wPDiag_55[8] , \wPDiag_55[7] , 
        \wPDiag_55[6] , \wPDiag_55[5] , \wPDiag_55[4] , \wPDiag_55[3] , 
        \wPDiag_55[2] , \wPDiag_55[1] , \wPDiag_55[0] }), .NDiagOut({
        \wNDiag_55[63] , \wNDiag_55[62] , \wNDiag_55[61] , \wNDiag_55[60] , 
        \wNDiag_55[59] , \wNDiag_55[58] , \wNDiag_55[57] , \wNDiag_55[56] , 
        \wNDiag_55[55] , \wNDiag_55[54] , \wNDiag_55[53] , \wNDiag_55[52] , 
        \wNDiag_55[51] , \wNDiag_55[50] , \wNDiag_55[49] , \wNDiag_55[48] , 
        \wNDiag_55[47] , \wNDiag_55[46] , \wNDiag_55[45] , \wNDiag_55[44] , 
        \wNDiag_55[43] , \wNDiag_55[42] , \wNDiag_55[41] , \wNDiag_55[40] , 
        \wNDiag_55[39] , \wNDiag_55[38] , \wNDiag_55[37] , \wNDiag_55[36] , 
        \wNDiag_55[35] , \wNDiag_55[34] , \wNDiag_55[33] , \wNDiag_55[32] , 
        \wNDiag_55[31] , \wNDiag_55[30] , \wNDiag_55[29] , \wNDiag_55[28] , 
        \wNDiag_55[27] , \wNDiag_55[26] , \wNDiag_55[25] , \wNDiag_55[24] , 
        \wNDiag_55[23] , \wNDiag_55[22] , \wNDiag_55[21] , \wNDiag_55[20] , 
        \wNDiag_55[19] , \wNDiag_55[18] , \wNDiag_55[17] , \wNDiag_55[16] , 
        \wNDiag_55[15] , \wNDiag_55[14] , \wNDiag_55[13] , \wNDiag_55[12] , 
        \wNDiag_55[11] , \wNDiag_55[10] , \wNDiag_55[9] , \wNDiag_55[8] , 
        \wNDiag_55[7] , \wNDiag_55[6] , \wNDiag_55[5] , \wNDiag_55[4] , 
        \wNDiag_55[3] , \wNDiag_55[2] , \wNDiag_55[1] , \wNDiag_55[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_46 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_47[6] , \wScan_47[5] , \wScan_47[4] , 
        \wScan_47[3] , \wScan_47[2] , \wScan_47[1] , \wScan_47[0] }), 
        .ScanOut({\wScan_46[6] , \wScan_46[5] , \wScan_46[4] , \wScan_46[3] , 
        \wScan_46[2] , \wScan_46[1] , \wScan_46[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_46[0] ), .ReturnIn(\wReturn_47[0] ), .ColIn({
        \wColumn_46[63] , \wColumn_46[62] , \wColumn_46[61] , \wColumn_46[60] , 
        \wColumn_46[59] , \wColumn_46[58] , \wColumn_46[57] , \wColumn_46[56] , 
        \wColumn_46[55] , \wColumn_46[54] , \wColumn_46[53] , \wColumn_46[52] , 
        \wColumn_46[51] , \wColumn_46[50] , \wColumn_46[49] , \wColumn_46[48] , 
        \wColumn_46[47] , \wColumn_46[46] , \wColumn_46[45] , \wColumn_46[44] , 
        \wColumn_46[43] , \wColumn_46[42] , \wColumn_46[41] , \wColumn_46[40] , 
        \wColumn_46[39] , \wColumn_46[38] , \wColumn_46[37] , \wColumn_46[36] , 
        \wColumn_46[35] , \wColumn_46[34] , \wColumn_46[33] , \wColumn_46[32] , 
        \wColumn_46[31] , \wColumn_46[30] , \wColumn_46[29] , \wColumn_46[28] , 
        \wColumn_46[27] , \wColumn_46[26] , \wColumn_46[25] , \wColumn_46[24] , 
        \wColumn_46[23] , \wColumn_46[22] , \wColumn_46[21] , \wColumn_46[20] , 
        \wColumn_46[19] , \wColumn_46[18] , \wColumn_46[17] , \wColumn_46[16] , 
        \wColumn_46[15] , \wColumn_46[14] , \wColumn_46[13] , \wColumn_46[12] , 
        \wColumn_46[11] , \wColumn_46[10] , \wColumn_46[9] , \wColumn_46[8] , 
        \wColumn_46[7] , \wColumn_46[6] , \wColumn_46[5] , \wColumn_46[4] , 
        \wColumn_46[3] , \wColumn_46[2] , \wColumn_46[1] , \wColumn_46[0] }), 
        .PDiagIn({\wPDiag_46[63] , \wPDiag_46[62] , \wPDiag_46[61] , 
        \wPDiag_46[60] , \wPDiag_46[59] , \wPDiag_46[58] , \wPDiag_46[57] , 
        \wPDiag_46[56] , \wPDiag_46[55] , \wPDiag_46[54] , \wPDiag_46[53] , 
        \wPDiag_46[52] , \wPDiag_46[51] , \wPDiag_46[50] , \wPDiag_46[49] , 
        \wPDiag_46[48] , \wPDiag_46[47] , \wPDiag_46[46] , \wPDiag_46[45] , 
        \wPDiag_46[44] , \wPDiag_46[43] , \wPDiag_46[42] , \wPDiag_46[41] , 
        \wPDiag_46[40] , \wPDiag_46[39] , \wPDiag_46[38] , \wPDiag_46[37] , 
        \wPDiag_46[36] , \wPDiag_46[35] , \wPDiag_46[34] , \wPDiag_46[33] , 
        \wPDiag_46[32] , \wPDiag_46[31] , \wPDiag_46[30] , \wPDiag_46[29] , 
        \wPDiag_46[28] , \wPDiag_46[27] , \wPDiag_46[26] , \wPDiag_46[25] , 
        \wPDiag_46[24] , \wPDiag_46[23] , \wPDiag_46[22] , \wPDiag_46[21] , 
        \wPDiag_46[20] , \wPDiag_46[19] , \wPDiag_46[18] , \wPDiag_46[17] , 
        \wPDiag_46[16] , \wPDiag_46[15] , \wPDiag_46[14] , \wPDiag_46[13] , 
        \wPDiag_46[12] , \wPDiag_46[11] , \wPDiag_46[10] , \wPDiag_46[9] , 
        \wPDiag_46[8] , \wPDiag_46[7] , \wPDiag_46[6] , \wPDiag_46[5] , 
        \wPDiag_46[4] , \wPDiag_46[3] , \wPDiag_46[2] , \wPDiag_46[1] , 
        \wPDiag_46[0] }), .NDiagIn({\wNDiag_46[63] , \wNDiag_46[62] , 
        \wNDiag_46[61] , \wNDiag_46[60] , \wNDiag_46[59] , \wNDiag_46[58] , 
        \wNDiag_46[57] , \wNDiag_46[56] , \wNDiag_46[55] , \wNDiag_46[54] , 
        \wNDiag_46[53] , \wNDiag_46[52] , \wNDiag_46[51] , \wNDiag_46[50] , 
        \wNDiag_46[49] , \wNDiag_46[48] , \wNDiag_46[47] , \wNDiag_46[46] , 
        \wNDiag_46[45] , \wNDiag_46[44] , \wNDiag_46[43] , \wNDiag_46[42] , 
        \wNDiag_46[41] , \wNDiag_46[40] , \wNDiag_46[39] , \wNDiag_46[38] , 
        \wNDiag_46[37] , \wNDiag_46[36] , \wNDiag_46[35] , \wNDiag_46[34] , 
        \wNDiag_46[33] , \wNDiag_46[32] , \wNDiag_46[31] , \wNDiag_46[30] , 
        \wNDiag_46[29] , \wNDiag_46[28] , \wNDiag_46[27] , \wNDiag_46[26] , 
        \wNDiag_46[25] , \wNDiag_46[24] , \wNDiag_46[23] , \wNDiag_46[22] , 
        \wNDiag_46[21] , \wNDiag_46[20] , \wNDiag_46[19] , \wNDiag_46[18] , 
        \wNDiag_46[17] , \wNDiag_46[16] , \wNDiag_46[15] , \wNDiag_46[14] , 
        \wNDiag_46[13] , \wNDiag_46[12] , \wNDiag_46[11] , \wNDiag_46[10] , 
        \wNDiag_46[9] , \wNDiag_46[8] , \wNDiag_46[7] , \wNDiag_46[6] , 
        \wNDiag_46[5] , \wNDiag_46[4] , \wNDiag_46[3] , \wNDiag_46[2] , 
        \wNDiag_46[1] , \wNDiag_46[0] }), .CallOut(\wCall_47[0] ), .ReturnOut(
        \wReturn_46[0] ), .ColOut({\wColumn_47[63] , \wColumn_47[62] , 
        \wColumn_47[61] , \wColumn_47[60] , \wColumn_47[59] , \wColumn_47[58] , 
        \wColumn_47[57] , \wColumn_47[56] , \wColumn_47[55] , \wColumn_47[54] , 
        \wColumn_47[53] , \wColumn_47[52] , \wColumn_47[51] , \wColumn_47[50] , 
        \wColumn_47[49] , \wColumn_47[48] , \wColumn_47[47] , \wColumn_47[46] , 
        \wColumn_47[45] , \wColumn_47[44] , \wColumn_47[43] , \wColumn_47[42] , 
        \wColumn_47[41] , \wColumn_47[40] , \wColumn_47[39] , \wColumn_47[38] , 
        \wColumn_47[37] , \wColumn_47[36] , \wColumn_47[35] , \wColumn_47[34] , 
        \wColumn_47[33] , \wColumn_47[32] , \wColumn_47[31] , \wColumn_47[30] , 
        \wColumn_47[29] , \wColumn_47[28] , \wColumn_47[27] , \wColumn_47[26] , 
        \wColumn_47[25] , \wColumn_47[24] , \wColumn_47[23] , \wColumn_47[22] , 
        \wColumn_47[21] , \wColumn_47[20] , \wColumn_47[19] , \wColumn_47[18] , 
        \wColumn_47[17] , \wColumn_47[16] , \wColumn_47[15] , \wColumn_47[14] , 
        \wColumn_47[13] , \wColumn_47[12] , \wColumn_47[11] , \wColumn_47[10] , 
        \wColumn_47[9] , \wColumn_47[8] , \wColumn_47[7] , \wColumn_47[6] , 
        \wColumn_47[5] , \wColumn_47[4] , \wColumn_47[3] , \wColumn_47[2] , 
        \wColumn_47[1] , \wColumn_47[0] }), .PDiagOut({\wPDiag_47[63] , 
        \wPDiag_47[62] , \wPDiag_47[61] , \wPDiag_47[60] , \wPDiag_47[59] , 
        \wPDiag_47[58] , \wPDiag_47[57] , \wPDiag_47[56] , \wPDiag_47[55] , 
        \wPDiag_47[54] , \wPDiag_47[53] , \wPDiag_47[52] , \wPDiag_47[51] , 
        \wPDiag_47[50] , \wPDiag_47[49] , \wPDiag_47[48] , \wPDiag_47[47] , 
        \wPDiag_47[46] , \wPDiag_47[45] , \wPDiag_47[44] , \wPDiag_47[43] , 
        \wPDiag_47[42] , \wPDiag_47[41] , \wPDiag_47[40] , \wPDiag_47[39] , 
        \wPDiag_47[38] , \wPDiag_47[37] , \wPDiag_47[36] , \wPDiag_47[35] , 
        \wPDiag_47[34] , \wPDiag_47[33] , \wPDiag_47[32] , \wPDiag_47[31] , 
        \wPDiag_47[30] , \wPDiag_47[29] , \wPDiag_47[28] , \wPDiag_47[27] , 
        \wPDiag_47[26] , \wPDiag_47[25] , \wPDiag_47[24] , \wPDiag_47[23] , 
        \wPDiag_47[22] , \wPDiag_47[21] , \wPDiag_47[20] , \wPDiag_47[19] , 
        \wPDiag_47[18] , \wPDiag_47[17] , \wPDiag_47[16] , \wPDiag_47[15] , 
        \wPDiag_47[14] , \wPDiag_47[13] , \wPDiag_47[12] , \wPDiag_47[11] , 
        \wPDiag_47[10] , \wPDiag_47[9] , \wPDiag_47[8] , \wPDiag_47[7] , 
        \wPDiag_47[6] , \wPDiag_47[5] , \wPDiag_47[4] , \wPDiag_47[3] , 
        \wPDiag_47[2] , \wPDiag_47[1] , \wPDiag_47[0] }), .NDiagOut({
        \wNDiag_47[63] , \wNDiag_47[62] , \wNDiag_47[61] , \wNDiag_47[60] , 
        \wNDiag_47[59] , \wNDiag_47[58] , \wNDiag_47[57] , \wNDiag_47[56] , 
        \wNDiag_47[55] , \wNDiag_47[54] , \wNDiag_47[53] , \wNDiag_47[52] , 
        \wNDiag_47[51] , \wNDiag_47[50] , \wNDiag_47[49] , \wNDiag_47[48] , 
        \wNDiag_47[47] , \wNDiag_47[46] , \wNDiag_47[45] , \wNDiag_47[44] , 
        \wNDiag_47[43] , \wNDiag_47[42] , \wNDiag_47[41] , \wNDiag_47[40] , 
        \wNDiag_47[39] , \wNDiag_47[38] , \wNDiag_47[37] , \wNDiag_47[36] , 
        \wNDiag_47[35] , \wNDiag_47[34] , \wNDiag_47[33] , \wNDiag_47[32] , 
        \wNDiag_47[31] , \wNDiag_47[30] , \wNDiag_47[29] , \wNDiag_47[28] , 
        \wNDiag_47[27] , \wNDiag_47[26] , \wNDiag_47[25] , \wNDiag_47[24] , 
        \wNDiag_47[23] , \wNDiag_47[22] , \wNDiag_47[21] , \wNDiag_47[20] , 
        \wNDiag_47[19] , \wNDiag_47[18] , \wNDiag_47[17] , \wNDiag_47[16] , 
        \wNDiag_47[15] , \wNDiag_47[14] , \wNDiag_47[13] , \wNDiag_47[12] , 
        \wNDiag_47[11] , \wNDiag_47[10] , \wNDiag_47[9] , \wNDiag_47[8] , 
        \wNDiag_47[7] , \wNDiag_47[6] , \wNDiag_47[5] , \wNDiag_47[4] , 
        \wNDiag_47[3] , \wNDiag_47[2] , \wNDiag_47[1] , \wNDiag_47[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_61 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_62[6] , \wScan_62[5] , \wScan_62[4] , 
        \wScan_62[3] , \wScan_62[2] , \wScan_62[1] , \wScan_62[0] }), 
        .ScanOut({\wScan_61[6] , \wScan_61[5] , \wScan_61[4] , \wScan_61[3] , 
        \wScan_61[2] , \wScan_61[1] , \wScan_61[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_61[0] ), .ReturnIn(\wReturn_62[0] ), .ColIn({
        \wColumn_61[63] , \wColumn_61[62] , \wColumn_61[61] , \wColumn_61[60] , 
        \wColumn_61[59] , \wColumn_61[58] , \wColumn_61[57] , \wColumn_61[56] , 
        \wColumn_61[55] , \wColumn_61[54] , \wColumn_61[53] , \wColumn_61[52] , 
        \wColumn_61[51] , \wColumn_61[50] , \wColumn_61[49] , \wColumn_61[48] , 
        \wColumn_61[47] , \wColumn_61[46] , \wColumn_61[45] , \wColumn_61[44] , 
        \wColumn_61[43] , \wColumn_61[42] , \wColumn_61[41] , \wColumn_61[40] , 
        \wColumn_61[39] , \wColumn_61[38] , \wColumn_61[37] , \wColumn_61[36] , 
        \wColumn_61[35] , \wColumn_61[34] , \wColumn_61[33] , \wColumn_61[32] , 
        \wColumn_61[31] , \wColumn_61[30] , \wColumn_61[29] , \wColumn_61[28] , 
        \wColumn_61[27] , \wColumn_61[26] , \wColumn_61[25] , \wColumn_61[24] , 
        \wColumn_61[23] , \wColumn_61[22] , \wColumn_61[21] , \wColumn_61[20] , 
        \wColumn_61[19] , \wColumn_61[18] , \wColumn_61[17] , \wColumn_61[16] , 
        \wColumn_61[15] , \wColumn_61[14] , \wColumn_61[13] , \wColumn_61[12] , 
        \wColumn_61[11] , \wColumn_61[10] , \wColumn_61[9] , \wColumn_61[8] , 
        \wColumn_61[7] , \wColumn_61[6] , \wColumn_61[5] , \wColumn_61[4] , 
        \wColumn_61[3] , \wColumn_61[2] , \wColumn_61[1] , \wColumn_61[0] }), 
        .PDiagIn({\wPDiag_61[63] , \wPDiag_61[62] , \wPDiag_61[61] , 
        \wPDiag_61[60] , \wPDiag_61[59] , \wPDiag_61[58] , \wPDiag_61[57] , 
        \wPDiag_61[56] , \wPDiag_61[55] , \wPDiag_61[54] , \wPDiag_61[53] , 
        \wPDiag_61[52] , \wPDiag_61[51] , \wPDiag_61[50] , \wPDiag_61[49] , 
        \wPDiag_61[48] , \wPDiag_61[47] , \wPDiag_61[46] , \wPDiag_61[45] , 
        \wPDiag_61[44] , \wPDiag_61[43] , \wPDiag_61[42] , \wPDiag_61[41] , 
        \wPDiag_61[40] , \wPDiag_61[39] , \wPDiag_61[38] , \wPDiag_61[37] , 
        \wPDiag_61[36] , \wPDiag_61[35] , \wPDiag_61[34] , \wPDiag_61[33] , 
        \wPDiag_61[32] , \wPDiag_61[31] , \wPDiag_61[30] , \wPDiag_61[29] , 
        \wPDiag_61[28] , \wPDiag_61[27] , \wPDiag_61[26] , \wPDiag_61[25] , 
        \wPDiag_61[24] , \wPDiag_61[23] , \wPDiag_61[22] , \wPDiag_61[21] , 
        \wPDiag_61[20] , \wPDiag_61[19] , \wPDiag_61[18] , \wPDiag_61[17] , 
        \wPDiag_61[16] , \wPDiag_61[15] , \wPDiag_61[14] , \wPDiag_61[13] , 
        \wPDiag_61[12] , \wPDiag_61[11] , \wPDiag_61[10] , \wPDiag_61[9] , 
        \wPDiag_61[8] , \wPDiag_61[7] , \wPDiag_61[6] , \wPDiag_61[5] , 
        \wPDiag_61[4] , \wPDiag_61[3] , \wPDiag_61[2] , \wPDiag_61[1] , 
        \wPDiag_61[0] }), .NDiagIn({\wNDiag_61[63] , \wNDiag_61[62] , 
        \wNDiag_61[61] , \wNDiag_61[60] , \wNDiag_61[59] , \wNDiag_61[58] , 
        \wNDiag_61[57] , \wNDiag_61[56] , \wNDiag_61[55] , \wNDiag_61[54] , 
        \wNDiag_61[53] , \wNDiag_61[52] , \wNDiag_61[51] , \wNDiag_61[50] , 
        \wNDiag_61[49] , \wNDiag_61[48] , \wNDiag_61[47] , \wNDiag_61[46] , 
        \wNDiag_61[45] , \wNDiag_61[44] , \wNDiag_61[43] , \wNDiag_61[42] , 
        \wNDiag_61[41] , \wNDiag_61[40] , \wNDiag_61[39] , \wNDiag_61[38] , 
        \wNDiag_61[37] , \wNDiag_61[36] , \wNDiag_61[35] , \wNDiag_61[34] , 
        \wNDiag_61[33] , \wNDiag_61[32] , \wNDiag_61[31] , \wNDiag_61[30] , 
        \wNDiag_61[29] , \wNDiag_61[28] , \wNDiag_61[27] , \wNDiag_61[26] , 
        \wNDiag_61[25] , \wNDiag_61[24] , \wNDiag_61[23] , \wNDiag_61[22] , 
        \wNDiag_61[21] , \wNDiag_61[20] , \wNDiag_61[19] , \wNDiag_61[18] , 
        \wNDiag_61[17] , \wNDiag_61[16] , \wNDiag_61[15] , \wNDiag_61[14] , 
        \wNDiag_61[13] , \wNDiag_61[12] , \wNDiag_61[11] , \wNDiag_61[10] , 
        \wNDiag_61[9] , \wNDiag_61[8] , \wNDiag_61[7] , \wNDiag_61[6] , 
        \wNDiag_61[5] , \wNDiag_61[4] , \wNDiag_61[3] , \wNDiag_61[2] , 
        \wNDiag_61[1] , \wNDiag_61[0] }), .CallOut(\wCall_62[0] ), .ReturnOut(
        \wReturn_61[0] ), .ColOut({\wColumn_62[63] , \wColumn_62[62] , 
        \wColumn_62[61] , \wColumn_62[60] , \wColumn_62[59] , \wColumn_62[58] , 
        \wColumn_62[57] , \wColumn_62[56] , \wColumn_62[55] , \wColumn_62[54] , 
        \wColumn_62[53] , \wColumn_62[52] , \wColumn_62[51] , \wColumn_62[50] , 
        \wColumn_62[49] , \wColumn_62[48] , \wColumn_62[47] , \wColumn_62[46] , 
        \wColumn_62[45] , \wColumn_62[44] , \wColumn_62[43] , \wColumn_62[42] , 
        \wColumn_62[41] , \wColumn_62[40] , \wColumn_62[39] , \wColumn_62[38] , 
        \wColumn_62[37] , \wColumn_62[36] , \wColumn_62[35] , \wColumn_62[34] , 
        \wColumn_62[33] , \wColumn_62[32] , \wColumn_62[31] , \wColumn_62[30] , 
        \wColumn_62[29] , \wColumn_62[28] , \wColumn_62[27] , \wColumn_62[26] , 
        \wColumn_62[25] , \wColumn_62[24] , \wColumn_62[23] , \wColumn_62[22] , 
        \wColumn_62[21] , \wColumn_62[20] , \wColumn_62[19] , \wColumn_62[18] , 
        \wColumn_62[17] , \wColumn_62[16] , \wColumn_62[15] , \wColumn_62[14] , 
        \wColumn_62[13] , \wColumn_62[12] , \wColumn_62[11] , \wColumn_62[10] , 
        \wColumn_62[9] , \wColumn_62[8] , \wColumn_62[7] , \wColumn_62[6] , 
        \wColumn_62[5] , \wColumn_62[4] , \wColumn_62[3] , \wColumn_62[2] , 
        \wColumn_62[1] , \wColumn_62[0] }), .PDiagOut({\wPDiag_62[63] , 
        \wPDiag_62[62] , \wPDiag_62[61] , \wPDiag_62[60] , \wPDiag_62[59] , 
        \wPDiag_62[58] , \wPDiag_62[57] , \wPDiag_62[56] , \wPDiag_62[55] , 
        \wPDiag_62[54] , \wPDiag_62[53] , \wPDiag_62[52] , \wPDiag_62[51] , 
        \wPDiag_62[50] , \wPDiag_62[49] , \wPDiag_62[48] , \wPDiag_62[47] , 
        \wPDiag_62[46] , \wPDiag_62[45] , \wPDiag_62[44] , \wPDiag_62[43] , 
        \wPDiag_62[42] , \wPDiag_62[41] , \wPDiag_62[40] , \wPDiag_62[39] , 
        \wPDiag_62[38] , \wPDiag_62[37] , \wPDiag_62[36] , \wPDiag_62[35] , 
        \wPDiag_62[34] , \wPDiag_62[33] , \wPDiag_62[32] , \wPDiag_62[31] , 
        \wPDiag_62[30] , \wPDiag_62[29] , \wPDiag_62[28] , \wPDiag_62[27] , 
        \wPDiag_62[26] , \wPDiag_62[25] , \wPDiag_62[24] , \wPDiag_62[23] , 
        \wPDiag_62[22] , \wPDiag_62[21] , \wPDiag_62[20] , \wPDiag_62[19] , 
        \wPDiag_62[18] , \wPDiag_62[17] , \wPDiag_62[16] , \wPDiag_62[15] , 
        \wPDiag_62[14] , \wPDiag_62[13] , \wPDiag_62[12] , \wPDiag_62[11] , 
        \wPDiag_62[10] , \wPDiag_62[9] , \wPDiag_62[8] , \wPDiag_62[7] , 
        \wPDiag_62[6] , \wPDiag_62[5] , \wPDiag_62[4] , \wPDiag_62[3] , 
        \wPDiag_62[2] , \wPDiag_62[1] , \wPDiag_62[0] }), .NDiagOut({
        \wNDiag_62[63] , \wNDiag_62[62] , \wNDiag_62[61] , \wNDiag_62[60] , 
        \wNDiag_62[59] , \wNDiag_62[58] , \wNDiag_62[57] , \wNDiag_62[56] , 
        \wNDiag_62[55] , \wNDiag_62[54] , \wNDiag_62[53] , \wNDiag_62[52] , 
        \wNDiag_62[51] , \wNDiag_62[50] , \wNDiag_62[49] , \wNDiag_62[48] , 
        \wNDiag_62[47] , \wNDiag_62[46] , \wNDiag_62[45] , \wNDiag_62[44] , 
        \wNDiag_62[43] , \wNDiag_62[42] , \wNDiag_62[41] , \wNDiag_62[40] , 
        \wNDiag_62[39] , \wNDiag_62[38] , \wNDiag_62[37] , \wNDiag_62[36] , 
        \wNDiag_62[35] , \wNDiag_62[34] , \wNDiag_62[33] , \wNDiag_62[32] , 
        \wNDiag_62[31] , \wNDiag_62[30] , \wNDiag_62[29] , \wNDiag_62[28] , 
        \wNDiag_62[27] , \wNDiag_62[26] , \wNDiag_62[25] , \wNDiag_62[24] , 
        \wNDiag_62[23] , \wNDiag_62[22] , \wNDiag_62[21] , \wNDiag_62[20] , 
        \wNDiag_62[19] , \wNDiag_62[18] , \wNDiag_62[17] , \wNDiag_62[16] , 
        \wNDiag_62[15] , \wNDiag_62[14] , \wNDiag_62[13] , \wNDiag_62[12] , 
        \wNDiag_62[11] , \wNDiag_62[10] , \wNDiag_62[9] , \wNDiag_62[8] , 
        \wNDiag_62[7] , \wNDiag_62[6] , \wNDiag_62[5] , \wNDiag_62[4] , 
        \wNDiag_62[3] , \wNDiag_62[2] , \wNDiag_62[1] , \wNDiag_62[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_33 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_34[6] , \wScan_34[5] , \wScan_34[4] , 
        \wScan_34[3] , \wScan_34[2] , \wScan_34[1] , \wScan_34[0] }), 
        .ScanOut({\wScan_33[6] , \wScan_33[5] , \wScan_33[4] , \wScan_33[3] , 
        \wScan_33[2] , \wScan_33[1] , \wScan_33[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_33[0] ), .ReturnIn(\wReturn_34[0] ), .ColIn({
        \wColumn_33[63] , \wColumn_33[62] , \wColumn_33[61] , \wColumn_33[60] , 
        \wColumn_33[59] , \wColumn_33[58] , \wColumn_33[57] , \wColumn_33[56] , 
        \wColumn_33[55] , \wColumn_33[54] , \wColumn_33[53] , \wColumn_33[52] , 
        \wColumn_33[51] , \wColumn_33[50] , \wColumn_33[49] , \wColumn_33[48] , 
        \wColumn_33[47] , \wColumn_33[46] , \wColumn_33[45] , \wColumn_33[44] , 
        \wColumn_33[43] , \wColumn_33[42] , \wColumn_33[41] , \wColumn_33[40] , 
        \wColumn_33[39] , \wColumn_33[38] , \wColumn_33[37] , \wColumn_33[36] , 
        \wColumn_33[35] , \wColumn_33[34] , \wColumn_33[33] , \wColumn_33[32] , 
        \wColumn_33[31] , \wColumn_33[30] , \wColumn_33[29] , \wColumn_33[28] , 
        \wColumn_33[27] , \wColumn_33[26] , \wColumn_33[25] , \wColumn_33[24] , 
        \wColumn_33[23] , \wColumn_33[22] , \wColumn_33[21] , \wColumn_33[20] , 
        \wColumn_33[19] , \wColumn_33[18] , \wColumn_33[17] , \wColumn_33[16] , 
        \wColumn_33[15] , \wColumn_33[14] , \wColumn_33[13] , \wColumn_33[12] , 
        \wColumn_33[11] , \wColumn_33[10] , \wColumn_33[9] , \wColumn_33[8] , 
        \wColumn_33[7] , \wColumn_33[6] , \wColumn_33[5] , \wColumn_33[4] , 
        \wColumn_33[3] , \wColumn_33[2] , \wColumn_33[1] , \wColumn_33[0] }), 
        .PDiagIn({\wPDiag_33[63] , \wPDiag_33[62] , \wPDiag_33[61] , 
        \wPDiag_33[60] , \wPDiag_33[59] , \wPDiag_33[58] , \wPDiag_33[57] , 
        \wPDiag_33[56] , \wPDiag_33[55] , \wPDiag_33[54] , \wPDiag_33[53] , 
        \wPDiag_33[52] , \wPDiag_33[51] , \wPDiag_33[50] , \wPDiag_33[49] , 
        \wPDiag_33[48] , \wPDiag_33[47] , \wPDiag_33[46] , \wPDiag_33[45] , 
        \wPDiag_33[44] , \wPDiag_33[43] , \wPDiag_33[42] , \wPDiag_33[41] , 
        \wPDiag_33[40] , \wPDiag_33[39] , \wPDiag_33[38] , \wPDiag_33[37] , 
        \wPDiag_33[36] , \wPDiag_33[35] , \wPDiag_33[34] , \wPDiag_33[33] , 
        \wPDiag_33[32] , \wPDiag_33[31] , \wPDiag_33[30] , \wPDiag_33[29] , 
        \wPDiag_33[28] , \wPDiag_33[27] , \wPDiag_33[26] , \wPDiag_33[25] , 
        \wPDiag_33[24] , \wPDiag_33[23] , \wPDiag_33[22] , \wPDiag_33[21] , 
        \wPDiag_33[20] , \wPDiag_33[19] , \wPDiag_33[18] , \wPDiag_33[17] , 
        \wPDiag_33[16] , \wPDiag_33[15] , \wPDiag_33[14] , \wPDiag_33[13] , 
        \wPDiag_33[12] , \wPDiag_33[11] , \wPDiag_33[10] , \wPDiag_33[9] , 
        \wPDiag_33[8] , \wPDiag_33[7] , \wPDiag_33[6] , \wPDiag_33[5] , 
        \wPDiag_33[4] , \wPDiag_33[3] , \wPDiag_33[2] , \wPDiag_33[1] , 
        \wPDiag_33[0] }), .NDiagIn({\wNDiag_33[63] , \wNDiag_33[62] , 
        \wNDiag_33[61] , \wNDiag_33[60] , \wNDiag_33[59] , \wNDiag_33[58] , 
        \wNDiag_33[57] , \wNDiag_33[56] , \wNDiag_33[55] , \wNDiag_33[54] , 
        \wNDiag_33[53] , \wNDiag_33[52] , \wNDiag_33[51] , \wNDiag_33[50] , 
        \wNDiag_33[49] , \wNDiag_33[48] , \wNDiag_33[47] , \wNDiag_33[46] , 
        \wNDiag_33[45] , \wNDiag_33[44] , \wNDiag_33[43] , \wNDiag_33[42] , 
        \wNDiag_33[41] , \wNDiag_33[40] , \wNDiag_33[39] , \wNDiag_33[38] , 
        \wNDiag_33[37] , \wNDiag_33[36] , \wNDiag_33[35] , \wNDiag_33[34] , 
        \wNDiag_33[33] , \wNDiag_33[32] , \wNDiag_33[31] , \wNDiag_33[30] , 
        \wNDiag_33[29] , \wNDiag_33[28] , \wNDiag_33[27] , \wNDiag_33[26] , 
        \wNDiag_33[25] , \wNDiag_33[24] , \wNDiag_33[23] , \wNDiag_33[22] , 
        \wNDiag_33[21] , \wNDiag_33[20] , \wNDiag_33[19] , \wNDiag_33[18] , 
        \wNDiag_33[17] , \wNDiag_33[16] , \wNDiag_33[15] , \wNDiag_33[14] , 
        \wNDiag_33[13] , \wNDiag_33[12] , \wNDiag_33[11] , \wNDiag_33[10] , 
        \wNDiag_33[9] , \wNDiag_33[8] , \wNDiag_33[7] , \wNDiag_33[6] , 
        \wNDiag_33[5] , \wNDiag_33[4] , \wNDiag_33[3] , \wNDiag_33[2] , 
        \wNDiag_33[1] , \wNDiag_33[0] }), .CallOut(\wCall_34[0] ), .ReturnOut(
        \wReturn_33[0] ), .ColOut({\wColumn_34[63] , \wColumn_34[62] , 
        \wColumn_34[61] , \wColumn_34[60] , \wColumn_34[59] , \wColumn_34[58] , 
        \wColumn_34[57] , \wColumn_34[56] , \wColumn_34[55] , \wColumn_34[54] , 
        \wColumn_34[53] , \wColumn_34[52] , \wColumn_34[51] , \wColumn_34[50] , 
        \wColumn_34[49] , \wColumn_34[48] , \wColumn_34[47] , \wColumn_34[46] , 
        \wColumn_34[45] , \wColumn_34[44] , \wColumn_34[43] , \wColumn_34[42] , 
        \wColumn_34[41] , \wColumn_34[40] , \wColumn_34[39] , \wColumn_34[38] , 
        \wColumn_34[37] , \wColumn_34[36] , \wColumn_34[35] , \wColumn_34[34] , 
        \wColumn_34[33] , \wColumn_34[32] , \wColumn_34[31] , \wColumn_34[30] , 
        \wColumn_34[29] , \wColumn_34[28] , \wColumn_34[27] , \wColumn_34[26] , 
        \wColumn_34[25] , \wColumn_34[24] , \wColumn_34[23] , \wColumn_34[22] , 
        \wColumn_34[21] , \wColumn_34[20] , \wColumn_34[19] , \wColumn_34[18] , 
        \wColumn_34[17] , \wColumn_34[16] , \wColumn_34[15] , \wColumn_34[14] , 
        \wColumn_34[13] , \wColumn_34[12] , \wColumn_34[11] , \wColumn_34[10] , 
        \wColumn_34[9] , \wColumn_34[8] , \wColumn_34[7] , \wColumn_34[6] , 
        \wColumn_34[5] , \wColumn_34[4] , \wColumn_34[3] , \wColumn_34[2] , 
        \wColumn_34[1] , \wColumn_34[0] }), .PDiagOut({\wPDiag_34[63] , 
        \wPDiag_34[62] , \wPDiag_34[61] , \wPDiag_34[60] , \wPDiag_34[59] , 
        \wPDiag_34[58] , \wPDiag_34[57] , \wPDiag_34[56] , \wPDiag_34[55] , 
        \wPDiag_34[54] , \wPDiag_34[53] , \wPDiag_34[52] , \wPDiag_34[51] , 
        \wPDiag_34[50] , \wPDiag_34[49] , \wPDiag_34[48] , \wPDiag_34[47] , 
        \wPDiag_34[46] , \wPDiag_34[45] , \wPDiag_34[44] , \wPDiag_34[43] , 
        \wPDiag_34[42] , \wPDiag_34[41] , \wPDiag_34[40] , \wPDiag_34[39] , 
        \wPDiag_34[38] , \wPDiag_34[37] , \wPDiag_34[36] , \wPDiag_34[35] , 
        \wPDiag_34[34] , \wPDiag_34[33] , \wPDiag_34[32] , \wPDiag_34[31] , 
        \wPDiag_34[30] , \wPDiag_34[29] , \wPDiag_34[28] , \wPDiag_34[27] , 
        \wPDiag_34[26] , \wPDiag_34[25] , \wPDiag_34[24] , \wPDiag_34[23] , 
        \wPDiag_34[22] , \wPDiag_34[21] , \wPDiag_34[20] , \wPDiag_34[19] , 
        \wPDiag_34[18] , \wPDiag_34[17] , \wPDiag_34[16] , \wPDiag_34[15] , 
        \wPDiag_34[14] , \wPDiag_34[13] , \wPDiag_34[12] , \wPDiag_34[11] , 
        \wPDiag_34[10] , \wPDiag_34[9] , \wPDiag_34[8] , \wPDiag_34[7] , 
        \wPDiag_34[6] , \wPDiag_34[5] , \wPDiag_34[4] , \wPDiag_34[3] , 
        \wPDiag_34[2] , \wPDiag_34[1] , \wPDiag_34[0] }), .NDiagOut({
        \wNDiag_34[63] , \wNDiag_34[62] , \wNDiag_34[61] , \wNDiag_34[60] , 
        \wNDiag_34[59] , \wNDiag_34[58] , \wNDiag_34[57] , \wNDiag_34[56] , 
        \wNDiag_34[55] , \wNDiag_34[54] , \wNDiag_34[53] , \wNDiag_34[52] , 
        \wNDiag_34[51] , \wNDiag_34[50] , \wNDiag_34[49] , \wNDiag_34[48] , 
        \wNDiag_34[47] , \wNDiag_34[46] , \wNDiag_34[45] , \wNDiag_34[44] , 
        \wNDiag_34[43] , \wNDiag_34[42] , \wNDiag_34[41] , \wNDiag_34[40] , 
        \wNDiag_34[39] , \wNDiag_34[38] , \wNDiag_34[37] , \wNDiag_34[36] , 
        \wNDiag_34[35] , \wNDiag_34[34] , \wNDiag_34[33] , \wNDiag_34[32] , 
        \wNDiag_34[31] , \wNDiag_34[30] , \wNDiag_34[29] , \wNDiag_34[28] , 
        \wNDiag_34[27] , \wNDiag_34[26] , \wNDiag_34[25] , \wNDiag_34[24] , 
        \wNDiag_34[23] , \wNDiag_34[22] , \wNDiag_34[21] , \wNDiag_34[20] , 
        \wNDiag_34[19] , \wNDiag_34[18] , \wNDiag_34[17] , \wNDiag_34[16] , 
        \wNDiag_34[15] , \wNDiag_34[14] , \wNDiag_34[13] , \wNDiag_34[12] , 
        \wNDiag_34[11] , \wNDiag_34[10] , \wNDiag_34[9] , \wNDiag_34[8] , 
        \wNDiag_34[7] , \wNDiag_34[6] , \wNDiag_34[5] , \wNDiag_34[4] , 
        \wNDiag_34[3] , \wNDiag_34[2] , \wNDiag_34[1] , \wNDiag_34[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_34 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_35[6] , \wScan_35[5] , \wScan_35[4] , 
        \wScan_35[3] , \wScan_35[2] , \wScan_35[1] , \wScan_35[0] }), 
        .ScanOut({\wScan_34[6] , \wScan_34[5] , \wScan_34[4] , \wScan_34[3] , 
        \wScan_34[2] , \wScan_34[1] , \wScan_34[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_34[0] ), .ReturnIn(\wReturn_35[0] ), .ColIn({
        \wColumn_34[63] , \wColumn_34[62] , \wColumn_34[61] , \wColumn_34[60] , 
        \wColumn_34[59] , \wColumn_34[58] , \wColumn_34[57] , \wColumn_34[56] , 
        \wColumn_34[55] , \wColumn_34[54] , \wColumn_34[53] , \wColumn_34[52] , 
        \wColumn_34[51] , \wColumn_34[50] , \wColumn_34[49] , \wColumn_34[48] , 
        \wColumn_34[47] , \wColumn_34[46] , \wColumn_34[45] , \wColumn_34[44] , 
        \wColumn_34[43] , \wColumn_34[42] , \wColumn_34[41] , \wColumn_34[40] , 
        \wColumn_34[39] , \wColumn_34[38] , \wColumn_34[37] , \wColumn_34[36] , 
        \wColumn_34[35] , \wColumn_34[34] , \wColumn_34[33] , \wColumn_34[32] , 
        \wColumn_34[31] , \wColumn_34[30] , \wColumn_34[29] , \wColumn_34[28] , 
        \wColumn_34[27] , \wColumn_34[26] , \wColumn_34[25] , \wColumn_34[24] , 
        \wColumn_34[23] , \wColumn_34[22] , \wColumn_34[21] , \wColumn_34[20] , 
        \wColumn_34[19] , \wColumn_34[18] , \wColumn_34[17] , \wColumn_34[16] , 
        \wColumn_34[15] , \wColumn_34[14] , \wColumn_34[13] , \wColumn_34[12] , 
        \wColumn_34[11] , \wColumn_34[10] , \wColumn_34[9] , \wColumn_34[8] , 
        \wColumn_34[7] , \wColumn_34[6] , \wColumn_34[5] , \wColumn_34[4] , 
        \wColumn_34[3] , \wColumn_34[2] , \wColumn_34[1] , \wColumn_34[0] }), 
        .PDiagIn({\wPDiag_34[63] , \wPDiag_34[62] , \wPDiag_34[61] , 
        \wPDiag_34[60] , \wPDiag_34[59] , \wPDiag_34[58] , \wPDiag_34[57] , 
        \wPDiag_34[56] , \wPDiag_34[55] , \wPDiag_34[54] , \wPDiag_34[53] , 
        \wPDiag_34[52] , \wPDiag_34[51] , \wPDiag_34[50] , \wPDiag_34[49] , 
        \wPDiag_34[48] , \wPDiag_34[47] , \wPDiag_34[46] , \wPDiag_34[45] , 
        \wPDiag_34[44] , \wPDiag_34[43] , \wPDiag_34[42] , \wPDiag_34[41] , 
        \wPDiag_34[40] , \wPDiag_34[39] , \wPDiag_34[38] , \wPDiag_34[37] , 
        \wPDiag_34[36] , \wPDiag_34[35] , \wPDiag_34[34] , \wPDiag_34[33] , 
        \wPDiag_34[32] , \wPDiag_34[31] , \wPDiag_34[30] , \wPDiag_34[29] , 
        \wPDiag_34[28] , \wPDiag_34[27] , \wPDiag_34[26] , \wPDiag_34[25] , 
        \wPDiag_34[24] , \wPDiag_34[23] , \wPDiag_34[22] , \wPDiag_34[21] , 
        \wPDiag_34[20] , \wPDiag_34[19] , \wPDiag_34[18] , \wPDiag_34[17] , 
        \wPDiag_34[16] , \wPDiag_34[15] , \wPDiag_34[14] , \wPDiag_34[13] , 
        \wPDiag_34[12] , \wPDiag_34[11] , \wPDiag_34[10] , \wPDiag_34[9] , 
        \wPDiag_34[8] , \wPDiag_34[7] , \wPDiag_34[6] , \wPDiag_34[5] , 
        \wPDiag_34[4] , \wPDiag_34[3] , \wPDiag_34[2] , \wPDiag_34[1] , 
        \wPDiag_34[0] }), .NDiagIn({\wNDiag_34[63] , \wNDiag_34[62] , 
        \wNDiag_34[61] , \wNDiag_34[60] , \wNDiag_34[59] , \wNDiag_34[58] , 
        \wNDiag_34[57] , \wNDiag_34[56] , \wNDiag_34[55] , \wNDiag_34[54] , 
        \wNDiag_34[53] , \wNDiag_34[52] , \wNDiag_34[51] , \wNDiag_34[50] , 
        \wNDiag_34[49] , \wNDiag_34[48] , \wNDiag_34[47] , \wNDiag_34[46] , 
        \wNDiag_34[45] , \wNDiag_34[44] , \wNDiag_34[43] , \wNDiag_34[42] , 
        \wNDiag_34[41] , \wNDiag_34[40] , \wNDiag_34[39] , \wNDiag_34[38] , 
        \wNDiag_34[37] , \wNDiag_34[36] , \wNDiag_34[35] , \wNDiag_34[34] , 
        \wNDiag_34[33] , \wNDiag_34[32] , \wNDiag_34[31] , \wNDiag_34[30] , 
        \wNDiag_34[29] , \wNDiag_34[28] , \wNDiag_34[27] , \wNDiag_34[26] , 
        \wNDiag_34[25] , \wNDiag_34[24] , \wNDiag_34[23] , \wNDiag_34[22] , 
        \wNDiag_34[21] , \wNDiag_34[20] , \wNDiag_34[19] , \wNDiag_34[18] , 
        \wNDiag_34[17] , \wNDiag_34[16] , \wNDiag_34[15] , \wNDiag_34[14] , 
        \wNDiag_34[13] , \wNDiag_34[12] , \wNDiag_34[11] , \wNDiag_34[10] , 
        \wNDiag_34[9] , \wNDiag_34[8] , \wNDiag_34[7] , \wNDiag_34[6] , 
        \wNDiag_34[5] , \wNDiag_34[4] , \wNDiag_34[3] , \wNDiag_34[2] , 
        \wNDiag_34[1] , \wNDiag_34[0] }), .CallOut(\wCall_35[0] ), .ReturnOut(
        \wReturn_34[0] ), .ColOut({\wColumn_35[63] , \wColumn_35[62] , 
        \wColumn_35[61] , \wColumn_35[60] , \wColumn_35[59] , \wColumn_35[58] , 
        \wColumn_35[57] , \wColumn_35[56] , \wColumn_35[55] , \wColumn_35[54] , 
        \wColumn_35[53] , \wColumn_35[52] , \wColumn_35[51] , \wColumn_35[50] , 
        \wColumn_35[49] , \wColumn_35[48] , \wColumn_35[47] , \wColumn_35[46] , 
        \wColumn_35[45] , \wColumn_35[44] , \wColumn_35[43] , \wColumn_35[42] , 
        \wColumn_35[41] , \wColumn_35[40] , \wColumn_35[39] , \wColumn_35[38] , 
        \wColumn_35[37] , \wColumn_35[36] , \wColumn_35[35] , \wColumn_35[34] , 
        \wColumn_35[33] , \wColumn_35[32] , \wColumn_35[31] , \wColumn_35[30] , 
        \wColumn_35[29] , \wColumn_35[28] , \wColumn_35[27] , \wColumn_35[26] , 
        \wColumn_35[25] , \wColumn_35[24] , \wColumn_35[23] , \wColumn_35[22] , 
        \wColumn_35[21] , \wColumn_35[20] , \wColumn_35[19] , \wColumn_35[18] , 
        \wColumn_35[17] , \wColumn_35[16] , \wColumn_35[15] , \wColumn_35[14] , 
        \wColumn_35[13] , \wColumn_35[12] , \wColumn_35[11] , \wColumn_35[10] , 
        \wColumn_35[9] , \wColumn_35[8] , \wColumn_35[7] , \wColumn_35[6] , 
        \wColumn_35[5] , \wColumn_35[4] , \wColumn_35[3] , \wColumn_35[2] , 
        \wColumn_35[1] , \wColumn_35[0] }), .PDiagOut({\wPDiag_35[63] , 
        \wPDiag_35[62] , \wPDiag_35[61] , \wPDiag_35[60] , \wPDiag_35[59] , 
        \wPDiag_35[58] , \wPDiag_35[57] , \wPDiag_35[56] , \wPDiag_35[55] , 
        \wPDiag_35[54] , \wPDiag_35[53] , \wPDiag_35[52] , \wPDiag_35[51] , 
        \wPDiag_35[50] , \wPDiag_35[49] , \wPDiag_35[48] , \wPDiag_35[47] , 
        \wPDiag_35[46] , \wPDiag_35[45] , \wPDiag_35[44] , \wPDiag_35[43] , 
        \wPDiag_35[42] , \wPDiag_35[41] , \wPDiag_35[40] , \wPDiag_35[39] , 
        \wPDiag_35[38] , \wPDiag_35[37] , \wPDiag_35[36] , \wPDiag_35[35] , 
        \wPDiag_35[34] , \wPDiag_35[33] , \wPDiag_35[32] , \wPDiag_35[31] , 
        \wPDiag_35[30] , \wPDiag_35[29] , \wPDiag_35[28] , \wPDiag_35[27] , 
        \wPDiag_35[26] , \wPDiag_35[25] , \wPDiag_35[24] , \wPDiag_35[23] , 
        \wPDiag_35[22] , \wPDiag_35[21] , \wPDiag_35[20] , \wPDiag_35[19] , 
        \wPDiag_35[18] , \wPDiag_35[17] , \wPDiag_35[16] , \wPDiag_35[15] , 
        \wPDiag_35[14] , \wPDiag_35[13] , \wPDiag_35[12] , \wPDiag_35[11] , 
        \wPDiag_35[10] , \wPDiag_35[9] , \wPDiag_35[8] , \wPDiag_35[7] , 
        \wPDiag_35[6] , \wPDiag_35[5] , \wPDiag_35[4] , \wPDiag_35[3] , 
        \wPDiag_35[2] , \wPDiag_35[1] , \wPDiag_35[0] }), .NDiagOut({
        \wNDiag_35[63] , \wNDiag_35[62] , \wNDiag_35[61] , \wNDiag_35[60] , 
        \wNDiag_35[59] , \wNDiag_35[58] , \wNDiag_35[57] , \wNDiag_35[56] , 
        \wNDiag_35[55] , \wNDiag_35[54] , \wNDiag_35[53] , \wNDiag_35[52] , 
        \wNDiag_35[51] , \wNDiag_35[50] , \wNDiag_35[49] , \wNDiag_35[48] , 
        \wNDiag_35[47] , \wNDiag_35[46] , \wNDiag_35[45] , \wNDiag_35[44] , 
        \wNDiag_35[43] , \wNDiag_35[42] , \wNDiag_35[41] , \wNDiag_35[40] , 
        \wNDiag_35[39] , \wNDiag_35[38] , \wNDiag_35[37] , \wNDiag_35[36] , 
        \wNDiag_35[35] , \wNDiag_35[34] , \wNDiag_35[33] , \wNDiag_35[32] , 
        \wNDiag_35[31] , \wNDiag_35[30] , \wNDiag_35[29] , \wNDiag_35[28] , 
        \wNDiag_35[27] , \wNDiag_35[26] , \wNDiag_35[25] , \wNDiag_35[24] , 
        \wNDiag_35[23] , \wNDiag_35[22] , \wNDiag_35[21] , \wNDiag_35[20] , 
        \wNDiag_35[19] , \wNDiag_35[18] , \wNDiag_35[17] , \wNDiag_35[16] , 
        \wNDiag_35[15] , \wNDiag_35[14] , \wNDiag_35[13] , \wNDiag_35[12] , 
        \wNDiag_35[11] , \wNDiag_35[10] , \wNDiag_35[9] , \wNDiag_35[8] , 
        \wNDiag_35[7] , \wNDiag_35[6] , \wNDiag_35[5] , \wNDiag_35[4] , 
        \wNDiag_35[3] , \wNDiag_35[2] , \wNDiag_35[1] , \wNDiag_35[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_41 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_42[6] , \wScan_42[5] , \wScan_42[4] , 
        \wScan_42[3] , \wScan_42[2] , \wScan_42[1] , \wScan_42[0] }), 
        .ScanOut({\wScan_41[6] , \wScan_41[5] , \wScan_41[4] , \wScan_41[3] , 
        \wScan_41[2] , \wScan_41[1] , \wScan_41[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_41[0] ), .ReturnIn(\wReturn_42[0] ), .ColIn({
        \wColumn_41[63] , \wColumn_41[62] , \wColumn_41[61] , \wColumn_41[60] , 
        \wColumn_41[59] , \wColumn_41[58] , \wColumn_41[57] , \wColumn_41[56] , 
        \wColumn_41[55] , \wColumn_41[54] , \wColumn_41[53] , \wColumn_41[52] , 
        \wColumn_41[51] , \wColumn_41[50] , \wColumn_41[49] , \wColumn_41[48] , 
        \wColumn_41[47] , \wColumn_41[46] , \wColumn_41[45] , \wColumn_41[44] , 
        \wColumn_41[43] , \wColumn_41[42] , \wColumn_41[41] , \wColumn_41[40] , 
        \wColumn_41[39] , \wColumn_41[38] , \wColumn_41[37] , \wColumn_41[36] , 
        \wColumn_41[35] , \wColumn_41[34] , \wColumn_41[33] , \wColumn_41[32] , 
        \wColumn_41[31] , \wColumn_41[30] , \wColumn_41[29] , \wColumn_41[28] , 
        \wColumn_41[27] , \wColumn_41[26] , \wColumn_41[25] , \wColumn_41[24] , 
        \wColumn_41[23] , \wColumn_41[22] , \wColumn_41[21] , \wColumn_41[20] , 
        \wColumn_41[19] , \wColumn_41[18] , \wColumn_41[17] , \wColumn_41[16] , 
        \wColumn_41[15] , \wColumn_41[14] , \wColumn_41[13] , \wColumn_41[12] , 
        \wColumn_41[11] , \wColumn_41[10] , \wColumn_41[9] , \wColumn_41[8] , 
        \wColumn_41[7] , \wColumn_41[6] , \wColumn_41[5] , \wColumn_41[4] , 
        \wColumn_41[3] , \wColumn_41[2] , \wColumn_41[1] , \wColumn_41[0] }), 
        .PDiagIn({\wPDiag_41[63] , \wPDiag_41[62] , \wPDiag_41[61] , 
        \wPDiag_41[60] , \wPDiag_41[59] , \wPDiag_41[58] , \wPDiag_41[57] , 
        \wPDiag_41[56] , \wPDiag_41[55] , \wPDiag_41[54] , \wPDiag_41[53] , 
        \wPDiag_41[52] , \wPDiag_41[51] , \wPDiag_41[50] , \wPDiag_41[49] , 
        \wPDiag_41[48] , \wPDiag_41[47] , \wPDiag_41[46] , \wPDiag_41[45] , 
        \wPDiag_41[44] , \wPDiag_41[43] , \wPDiag_41[42] , \wPDiag_41[41] , 
        \wPDiag_41[40] , \wPDiag_41[39] , \wPDiag_41[38] , \wPDiag_41[37] , 
        \wPDiag_41[36] , \wPDiag_41[35] , \wPDiag_41[34] , \wPDiag_41[33] , 
        \wPDiag_41[32] , \wPDiag_41[31] , \wPDiag_41[30] , \wPDiag_41[29] , 
        \wPDiag_41[28] , \wPDiag_41[27] , \wPDiag_41[26] , \wPDiag_41[25] , 
        \wPDiag_41[24] , \wPDiag_41[23] , \wPDiag_41[22] , \wPDiag_41[21] , 
        \wPDiag_41[20] , \wPDiag_41[19] , \wPDiag_41[18] , \wPDiag_41[17] , 
        \wPDiag_41[16] , \wPDiag_41[15] , \wPDiag_41[14] , \wPDiag_41[13] , 
        \wPDiag_41[12] , \wPDiag_41[11] , \wPDiag_41[10] , \wPDiag_41[9] , 
        \wPDiag_41[8] , \wPDiag_41[7] , \wPDiag_41[6] , \wPDiag_41[5] , 
        \wPDiag_41[4] , \wPDiag_41[3] , \wPDiag_41[2] , \wPDiag_41[1] , 
        \wPDiag_41[0] }), .NDiagIn({\wNDiag_41[63] , \wNDiag_41[62] , 
        \wNDiag_41[61] , \wNDiag_41[60] , \wNDiag_41[59] , \wNDiag_41[58] , 
        \wNDiag_41[57] , \wNDiag_41[56] , \wNDiag_41[55] , \wNDiag_41[54] , 
        \wNDiag_41[53] , \wNDiag_41[52] , \wNDiag_41[51] , \wNDiag_41[50] , 
        \wNDiag_41[49] , \wNDiag_41[48] , \wNDiag_41[47] , \wNDiag_41[46] , 
        \wNDiag_41[45] , \wNDiag_41[44] , \wNDiag_41[43] , \wNDiag_41[42] , 
        \wNDiag_41[41] , \wNDiag_41[40] , \wNDiag_41[39] , \wNDiag_41[38] , 
        \wNDiag_41[37] , \wNDiag_41[36] , \wNDiag_41[35] , \wNDiag_41[34] , 
        \wNDiag_41[33] , \wNDiag_41[32] , \wNDiag_41[31] , \wNDiag_41[30] , 
        \wNDiag_41[29] , \wNDiag_41[28] , \wNDiag_41[27] , \wNDiag_41[26] , 
        \wNDiag_41[25] , \wNDiag_41[24] , \wNDiag_41[23] , \wNDiag_41[22] , 
        \wNDiag_41[21] , \wNDiag_41[20] , \wNDiag_41[19] , \wNDiag_41[18] , 
        \wNDiag_41[17] , \wNDiag_41[16] , \wNDiag_41[15] , \wNDiag_41[14] , 
        \wNDiag_41[13] , \wNDiag_41[12] , \wNDiag_41[11] , \wNDiag_41[10] , 
        \wNDiag_41[9] , \wNDiag_41[8] , \wNDiag_41[7] , \wNDiag_41[6] , 
        \wNDiag_41[5] , \wNDiag_41[4] , \wNDiag_41[3] , \wNDiag_41[2] , 
        \wNDiag_41[1] , \wNDiag_41[0] }), .CallOut(\wCall_42[0] ), .ReturnOut(
        \wReturn_41[0] ), .ColOut({\wColumn_42[63] , \wColumn_42[62] , 
        \wColumn_42[61] , \wColumn_42[60] , \wColumn_42[59] , \wColumn_42[58] , 
        \wColumn_42[57] , \wColumn_42[56] , \wColumn_42[55] , \wColumn_42[54] , 
        \wColumn_42[53] , \wColumn_42[52] , \wColumn_42[51] , \wColumn_42[50] , 
        \wColumn_42[49] , \wColumn_42[48] , \wColumn_42[47] , \wColumn_42[46] , 
        \wColumn_42[45] , \wColumn_42[44] , \wColumn_42[43] , \wColumn_42[42] , 
        \wColumn_42[41] , \wColumn_42[40] , \wColumn_42[39] , \wColumn_42[38] , 
        \wColumn_42[37] , \wColumn_42[36] , \wColumn_42[35] , \wColumn_42[34] , 
        \wColumn_42[33] , \wColumn_42[32] , \wColumn_42[31] , \wColumn_42[30] , 
        \wColumn_42[29] , \wColumn_42[28] , \wColumn_42[27] , \wColumn_42[26] , 
        \wColumn_42[25] , \wColumn_42[24] , \wColumn_42[23] , \wColumn_42[22] , 
        \wColumn_42[21] , \wColumn_42[20] , \wColumn_42[19] , \wColumn_42[18] , 
        \wColumn_42[17] , \wColumn_42[16] , \wColumn_42[15] , \wColumn_42[14] , 
        \wColumn_42[13] , \wColumn_42[12] , \wColumn_42[11] , \wColumn_42[10] , 
        \wColumn_42[9] , \wColumn_42[8] , \wColumn_42[7] , \wColumn_42[6] , 
        \wColumn_42[5] , \wColumn_42[4] , \wColumn_42[3] , \wColumn_42[2] , 
        \wColumn_42[1] , \wColumn_42[0] }), .PDiagOut({\wPDiag_42[63] , 
        \wPDiag_42[62] , \wPDiag_42[61] , \wPDiag_42[60] , \wPDiag_42[59] , 
        \wPDiag_42[58] , \wPDiag_42[57] , \wPDiag_42[56] , \wPDiag_42[55] , 
        \wPDiag_42[54] , \wPDiag_42[53] , \wPDiag_42[52] , \wPDiag_42[51] , 
        \wPDiag_42[50] , \wPDiag_42[49] , \wPDiag_42[48] , \wPDiag_42[47] , 
        \wPDiag_42[46] , \wPDiag_42[45] , \wPDiag_42[44] , \wPDiag_42[43] , 
        \wPDiag_42[42] , \wPDiag_42[41] , \wPDiag_42[40] , \wPDiag_42[39] , 
        \wPDiag_42[38] , \wPDiag_42[37] , \wPDiag_42[36] , \wPDiag_42[35] , 
        \wPDiag_42[34] , \wPDiag_42[33] , \wPDiag_42[32] , \wPDiag_42[31] , 
        \wPDiag_42[30] , \wPDiag_42[29] , \wPDiag_42[28] , \wPDiag_42[27] , 
        \wPDiag_42[26] , \wPDiag_42[25] , \wPDiag_42[24] , \wPDiag_42[23] , 
        \wPDiag_42[22] , \wPDiag_42[21] , \wPDiag_42[20] , \wPDiag_42[19] , 
        \wPDiag_42[18] , \wPDiag_42[17] , \wPDiag_42[16] , \wPDiag_42[15] , 
        \wPDiag_42[14] , \wPDiag_42[13] , \wPDiag_42[12] , \wPDiag_42[11] , 
        \wPDiag_42[10] , \wPDiag_42[9] , \wPDiag_42[8] , \wPDiag_42[7] , 
        \wPDiag_42[6] , \wPDiag_42[5] , \wPDiag_42[4] , \wPDiag_42[3] , 
        \wPDiag_42[2] , \wPDiag_42[1] , \wPDiag_42[0] }), .NDiagOut({
        \wNDiag_42[63] , \wNDiag_42[62] , \wNDiag_42[61] , \wNDiag_42[60] , 
        \wNDiag_42[59] , \wNDiag_42[58] , \wNDiag_42[57] , \wNDiag_42[56] , 
        \wNDiag_42[55] , \wNDiag_42[54] , \wNDiag_42[53] , \wNDiag_42[52] , 
        \wNDiag_42[51] , \wNDiag_42[50] , \wNDiag_42[49] , \wNDiag_42[48] , 
        \wNDiag_42[47] , \wNDiag_42[46] , \wNDiag_42[45] , \wNDiag_42[44] , 
        \wNDiag_42[43] , \wNDiag_42[42] , \wNDiag_42[41] , \wNDiag_42[40] , 
        \wNDiag_42[39] , \wNDiag_42[38] , \wNDiag_42[37] , \wNDiag_42[36] , 
        \wNDiag_42[35] , \wNDiag_42[34] , \wNDiag_42[33] , \wNDiag_42[32] , 
        \wNDiag_42[31] , \wNDiag_42[30] , \wNDiag_42[29] , \wNDiag_42[28] , 
        \wNDiag_42[27] , \wNDiag_42[26] , \wNDiag_42[25] , \wNDiag_42[24] , 
        \wNDiag_42[23] , \wNDiag_42[22] , \wNDiag_42[21] , \wNDiag_42[20] , 
        \wNDiag_42[19] , \wNDiag_42[18] , \wNDiag_42[17] , \wNDiag_42[16] , 
        \wNDiag_42[15] , \wNDiag_42[14] , \wNDiag_42[13] , \wNDiag_42[12] , 
        \wNDiag_42[11] , \wNDiag_42[10] , \wNDiag_42[9] , \wNDiag_42[8] , 
        \wNDiag_42[7] , \wNDiag_42[6] , \wNDiag_42[5] , \wNDiag_42[4] , 
        \wNDiag_42[3] , \wNDiag_42[2] , \wNDiag_42[1] , \wNDiag_42[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_53 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_54[6] , \wScan_54[5] , \wScan_54[4] , 
        \wScan_54[3] , \wScan_54[2] , \wScan_54[1] , \wScan_54[0] }), 
        .ScanOut({\wScan_53[6] , \wScan_53[5] , \wScan_53[4] , \wScan_53[3] , 
        \wScan_53[2] , \wScan_53[1] , \wScan_53[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_53[0] ), .ReturnIn(\wReturn_54[0] ), .ColIn({
        \wColumn_53[63] , \wColumn_53[62] , \wColumn_53[61] , \wColumn_53[60] , 
        \wColumn_53[59] , \wColumn_53[58] , \wColumn_53[57] , \wColumn_53[56] , 
        \wColumn_53[55] , \wColumn_53[54] , \wColumn_53[53] , \wColumn_53[52] , 
        \wColumn_53[51] , \wColumn_53[50] , \wColumn_53[49] , \wColumn_53[48] , 
        \wColumn_53[47] , \wColumn_53[46] , \wColumn_53[45] , \wColumn_53[44] , 
        \wColumn_53[43] , \wColumn_53[42] , \wColumn_53[41] , \wColumn_53[40] , 
        \wColumn_53[39] , \wColumn_53[38] , \wColumn_53[37] , \wColumn_53[36] , 
        \wColumn_53[35] , \wColumn_53[34] , \wColumn_53[33] , \wColumn_53[32] , 
        \wColumn_53[31] , \wColumn_53[30] , \wColumn_53[29] , \wColumn_53[28] , 
        \wColumn_53[27] , \wColumn_53[26] , \wColumn_53[25] , \wColumn_53[24] , 
        \wColumn_53[23] , \wColumn_53[22] , \wColumn_53[21] , \wColumn_53[20] , 
        \wColumn_53[19] , \wColumn_53[18] , \wColumn_53[17] , \wColumn_53[16] , 
        \wColumn_53[15] , \wColumn_53[14] , \wColumn_53[13] , \wColumn_53[12] , 
        \wColumn_53[11] , \wColumn_53[10] , \wColumn_53[9] , \wColumn_53[8] , 
        \wColumn_53[7] , \wColumn_53[6] , \wColumn_53[5] , \wColumn_53[4] , 
        \wColumn_53[3] , \wColumn_53[2] , \wColumn_53[1] , \wColumn_53[0] }), 
        .PDiagIn({\wPDiag_53[63] , \wPDiag_53[62] , \wPDiag_53[61] , 
        \wPDiag_53[60] , \wPDiag_53[59] , \wPDiag_53[58] , \wPDiag_53[57] , 
        \wPDiag_53[56] , \wPDiag_53[55] , \wPDiag_53[54] , \wPDiag_53[53] , 
        \wPDiag_53[52] , \wPDiag_53[51] , \wPDiag_53[50] , \wPDiag_53[49] , 
        \wPDiag_53[48] , \wPDiag_53[47] , \wPDiag_53[46] , \wPDiag_53[45] , 
        \wPDiag_53[44] , \wPDiag_53[43] , \wPDiag_53[42] , \wPDiag_53[41] , 
        \wPDiag_53[40] , \wPDiag_53[39] , \wPDiag_53[38] , \wPDiag_53[37] , 
        \wPDiag_53[36] , \wPDiag_53[35] , \wPDiag_53[34] , \wPDiag_53[33] , 
        \wPDiag_53[32] , \wPDiag_53[31] , \wPDiag_53[30] , \wPDiag_53[29] , 
        \wPDiag_53[28] , \wPDiag_53[27] , \wPDiag_53[26] , \wPDiag_53[25] , 
        \wPDiag_53[24] , \wPDiag_53[23] , \wPDiag_53[22] , \wPDiag_53[21] , 
        \wPDiag_53[20] , \wPDiag_53[19] , \wPDiag_53[18] , \wPDiag_53[17] , 
        \wPDiag_53[16] , \wPDiag_53[15] , \wPDiag_53[14] , \wPDiag_53[13] , 
        \wPDiag_53[12] , \wPDiag_53[11] , \wPDiag_53[10] , \wPDiag_53[9] , 
        \wPDiag_53[8] , \wPDiag_53[7] , \wPDiag_53[6] , \wPDiag_53[5] , 
        \wPDiag_53[4] , \wPDiag_53[3] , \wPDiag_53[2] , \wPDiag_53[1] , 
        \wPDiag_53[0] }), .NDiagIn({\wNDiag_53[63] , \wNDiag_53[62] , 
        \wNDiag_53[61] , \wNDiag_53[60] , \wNDiag_53[59] , \wNDiag_53[58] , 
        \wNDiag_53[57] , \wNDiag_53[56] , \wNDiag_53[55] , \wNDiag_53[54] , 
        \wNDiag_53[53] , \wNDiag_53[52] , \wNDiag_53[51] , \wNDiag_53[50] , 
        \wNDiag_53[49] , \wNDiag_53[48] , \wNDiag_53[47] , \wNDiag_53[46] , 
        \wNDiag_53[45] , \wNDiag_53[44] , \wNDiag_53[43] , \wNDiag_53[42] , 
        \wNDiag_53[41] , \wNDiag_53[40] , \wNDiag_53[39] , \wNDiag_53[38] , 
        \wNDiag_53[37] , \wNDiag_53[36] , \wNDiag_53[35] , \wNDiag_53[34] , 
        \wNDiag_53[33] , \wNDiag_53[32] , \wNDiag_53[31] , \wNDiag_53[30] , 
        \wNDiag_53[29] , \wNDiag_53[28] , \wNDiag_53[27] , \wNDiag_53[26] , 
        \wNDiag_53[25] , \wNDiag_53[24] , \wNDiag_53[23] , \wNDiag_53[22] , 
        \wNDiag_53[21] , \wNDiag_53[20] , \wNDiag_53[19] , \wNDiag_53[18] , 
        \wNDiag_53[17] , \wNDiag_53[16] , \wNDiag_53[15] , \wNDiag_53[14] , 
        \wNDiag_53[13] , \wNDiag_53[12] , \wNDiag_53[11] , \wNDiag_53[10] , 
        \wNDiag_53[9] , \wNDiag_53[8] , \wNDiag_53[7] , \wNDiag_53[6] , 
        \wNDiag_53[5] , \wNDiag_53[4] , \wNDiag_53[3] , \wNDiag_53[2] , 
        \wNDiag_53[1] , \wNDiag_53[0] }), .CallOut(\wCall_54[0] ), .ReturnOut(
        \wReturn_53[0] ), .ColOut({\wColumn_54[63] , \wColumn_54[62] , 
        \wColumn_54[61] , \wColumn_54[60] , \wColumn_54[59] , \wColumn_54[58] , 
        \wColumn_54[57] , \wColumn_54[56] , \wColumn_54[55] , \wColumn_54[54] , 
        \wColumn_54[53] , \wColumn_54[52] , \wColumn_54[51] , \wColumn_54[50] , 
        \wColumn_54[49] , \wColumn_54[48] , \wColumn_54[47] , \wColumn_54[46] , 
        \wColumn_54[45] , \wColumn_54[44] , \wColumn_54[43] , \wColumn_54[42] , 
        \wColumn_54[41] , \wColumn_54[40] , \wColumn_54[39] , \wColumn_54[38] , 
        \wColumn_54[37] , \wColumn_54[36] , \wColumn_54[35] , \wColumn_54[34] , 
        \wColumn_54[33] , \wColumn_54[32] , \wColumn_54[31] , \wColumn_54[30] , 
        \wColumn_54[29] , \wColumn_54[28] , \wColumn_54[27] , \wColumn_54[26] , 
        \wColumn_54[25] , \wColumn_54[24] , \wColumn_54[23] , \wColumn_54[22] , 
        \wColumn_54[21] , \wColumn_54[20] , \wColumn_54[19] , \wColumn_54[18] , 
        \wColumn_54[17] , \wColumn_54[16] , \wColumn_54[15] , \wColumn_54[14] , 
        \wColumn_54[13] , \wColumn_54[12] , \wColumn_54[11] , \wColumn_54[10] , 
        \wColumn_54[9] , \wColumn_54[8] , \wColumn_54[7] , \wColumn_54[6] , 
        \wColumn_54[5] , \wColumn_54[4] , \wColumn_54[3] , \wColumn_54[2] , 
        \wColumn_54[1] , \wColumn_54[0] }), .PDiagOut({\wPDiag_54[63] , 
        \wPDiag_54[62] , \wPDiag_54[61] , \wPDiag_54[60] , \wPDiag_54[59] , 
        \wPDiag_54[58] , \wPDiag_54[57] , \wPDiag_54[56] , \wPDiag_54[55] , 
        \wPDiag_54[54] , \wPDiag_54[53] , \wPDiag_54[52] , \wPDiag_54[51] , 
        \wPDiag_54[50] , \wPDiag_54[49] , \wPDiag_54[48] , \wPDiag_54[47] , 
        \wPDiag_54[46] , \wPDiag_54[45] , \wPDiag_54[44] , \wPDiag_54[43] , 
        \wPDiag_54[42] , \wPDiag_54[41] , \wPDiag_54[40] , \wPDiag_54[39] , 
        \wPDiag_54[38] , \wPDiag_54[37] , \wPDiag_54[36] , \wPDiag_54[35] , 
        \wPDiag_54[34] , \wPDiag_54[33] , \wPDiag_54[32] , \wPDiag_54[31] , 
        \wPDiag_54[30] , \wPDiag_54[29] , \wPDiag_54[28] , \wPDiag_54[27] , 
        \wPDiag_54[26] , \wPDiag_54[25] , \wPDiag_54[24] , \wPDiag_54[23] , 
        \wPDiag_54[22] , \wPDiag_54[21] , \wPDiag_54[20] , \wPDiag_54[19] , 
        \wPDiag_54[18] , \wPDiag_54[17] , \wPDiag_54[16] , \wPDiag_54[15] , 
        \wPDiag_54[14] , \wPDiag_54[13] , \wPDiag_54[12] , \wPDiag_54[11] , 
        \wPDiag_54[10] , \wPDiag_54[9] , \wPDiag_54[8] , \wPDiag_54[7] , 
        \wPDiag_54[6] , \wPDiag_54[5] , \wPDiag_54[4] , \wPDiag_54[3] , 
        \wPDiag_54[2] , \wPDiag_54[1] , \wPDiag_54[0] }), .NDiagOut({
        \wNDiag_54[63] , \wNDiag_54[62] , \wNDiag_54[61] , \wNDiag_54[60] , 
        \wNDiag_54[59] , \wNDiag_54[58] , \wNDiag_54[57] , \wNDiag_54[56] , 
        \wNDiag_54[55] , \wNDiag_54[54] , \wNDiag_54[53] , \wNDiag_54[52] , 
        \wNDiag_54[51] , \wNDiag_54[50] , \wNDiag_54[49] , \wNDiag_54[48] , 
        \wNDiag_54[47] , \wNDiag_54[46] , \wNDiag_54[45] , \wNDiag_54[44] , 
        \wNDiag_54[43] , \wNDiag_54[42] , \wNDiag_54[41] , \wNDiag_54[40] , 
        \wNDiag_54[39] , \wNDiag_54[38] , \wNDiag_54[37] , \wNDiag_54[36] , 
        \wNDiag_54[35] , \wNDiag_54[34] , \wNDiag_54[33] , \wNDiag_54[32] , 
        \wNDiag_54[31] , \wNDiag_54[30] , \wNDiag_54[29] , \wNDiag_54[28] , 
        \wNDiag_54[27] , \wNDiag_54[26] , \wNDiag_54[25] , \wNDiag_54[24] , 
        \wNDiag_54[23] , \wNDiag_54[22] , \wNDiag_54[21] , \wNDiag_54[20] , 
        \wNDiag_54[19] , \wNDiag_54[18] , \wNDiag_54[17] , \wNDiag_54[16] , 
        \wNDiag_54[15] , \wNDiag_54[14] , \wNDiag_54[13] , \wNDiag_54[12] , 
        \wNDiag_54[11] , \wNDiag_54[10] , \wNDiag_54[9] , \wNDiag_54[8] , 
        \wNDiag_54[7] , \wNDiag_54[6] , \wNDiag_54[5] , \wNDiag_54[4] , 
        \wNDiag_54[3] , \wNDiag_54[2] , \wNDiag_54[1] , \wNDiag_54[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_9 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_10[6] , \wScan_10[5] , \wScan_10[4] , 
        \wScan_10[3] , \wScan_10[2] , \wScan_10[1] , \wScan_10[0] }), 
        .ScanOut({\wScan_9[6] , \wScan_9[5] , \wScan_9[4] , \wScan_9[3] , 
        \wScan_9[2] , \wScan_9[1] , \wScan_9[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_9[0] ), .ReturnIn(\wReturn_10[0] ), .ColIn({
        \wColumn_9[63] , \wColumn_9[62] , \wColumn_9[61] , \wColumn_9[60] , 
        \wColumn_9[59] , \wColumn_9[58] , \wColumn_9[57] , \wColumn_9[56] , 
        \wColumn_9[55] , \wColumn_9[54] , \wColumn_9[53] , \wColumn_9[52] , 
        \wColumn_9[51] , \wColumn_9[50] , \wColumn_9[49] , \wColumn_9[48] , 
        \wColumn_9[47] , \wColumn_9[46] , \wColumn_9[45] , \wColumn_9[44] , 
        \wColumn_9[43] , \wColumn_9[42] , \wColumn_9[41] , \wColumn_9[40] , 
        \wColumn_9[39] , \wColumn_9[38] , \wColumn_9[37] , \wColumn_9[36] , 
        \wColumn_9[35] , \wColumn_9[34] , \wColumn_9[33] , \wColumn_9[32] , 
        \wColumn_9[31] , \wColumn_9[30] , \wColumn_9[29] , \wColumn_9[28] , 
        \wColumn_9[27] , \wColumn_9[26] , \wColumn_9[25] , \wColumn_9[24] , 
        \wColumn_9[23] , \wColumn_9[22] , \wColumn_9[21] , \wColumn_9[20] , 
        \wColumn_9[19] , \wColumn_9[18] , \wColumn_9[17] , \wColumn_9[16] , 
        \wColumn_9[15] , \wColumn_9[14] , \wColumn_9[13] , \wColumn_9[12] , 
        \wColumn_9[11] , \wColumn_9[10] , \wColumn_9[9] , \wColumn_9[8] , 
        \wColumn_9[7] , \wColumn_9[6] , \wColumn_9[5] , \wColumn_9[4] , 
        \wColumn_9[3] , \wColumn_9[2] , \wColumn_9[1] , \wColumn_9[0] }), 
        .PDiagIn({\wPDiag_9[63] , \wPDiag_9[62] , \wPDiag_9[61] , 
        \wPDiag_9[60] , \wPDiag_9[59] , \wPDiag_9[58] , \wPDiag_9[57] , 
        \wPDiag_9[56] , \wPDiag_9[55] , \wPDiag_9[54] , \wPDiag_9[53] , 
        \wPDiag_9[52] , \wPDiag_9[51] , \wPDiag_9[50] , \wPDiag_9[49] , 
        \wPDiag_9[48] , \wPDiag_9[47] , \wPDiag_9[46] , \wPDiag_9[45] , 
        \wPDiag_9[44] , \wPDiag_9[43] , \wPDiag_9[42] , \wPDiag_9[41] , 
        \wPDiag_9[40] , \wPDiag_9[39] , \wPDiag_9[38] , \wPDiag_9[37] , 
        \wPDiag_9[36] , \wPDiag_9[35] , \wPDiag_9[34] , \wPDiag_9[33] , 
        \wPDiag_9[32] , \wPDiag_9[31] , \wPDiag_9[30] , \wPDiag_9[29] , 
        \wPDiag_9[28] , \wPDiag_9[27] , \wPDiag_9[26] , \wPDiag_9[25] , 
        \wPDiag_9[24] , \wPDiag_9[23] , \wPDiag_9[22] , \wPDiag_9[21] , 
        \wPDiag_9[20] , \wPDiag_9[19] , \wPDiag_9[18] , \wPDiag_9[17] , 
        \wPDiag_9[16] , \wPDiag_9[15] , \wPDiag_9[14] , \wPDiag_9[13] , 
        \wPDiag_9[12] , \wPDiag_9[11] , \wPDiag_9[10] , \wPDiag_9[9] , 
        \wPDiag_9[8] , \wPDiag_9[7] , \wPDiag_9[6] , \wPDiag_9[5] , 
        \wPDiag_9[4] , \wPDiag_9[3] , \wPDiag_9[2] , \wPDiag_9[1] , 
        \wPDiag_9[0] }), .NDiagIn({\wNDiag_9[63] , \wNDiag_9[62] , 
        \wNDiag_9[61] , \wNDiag_9[60] , \wNDiag_9[59] , \wNDiag_9[58] , 
        \wNDiag_9[57] , \wNDiag_9[56] , \wNDiag_9[55] , \wNDiag_9[54] , 
        \wNDiag_9[53] , \wNDiag_9[52] , \wNDiag_9[51] , \wNDiag_9[50] , 
        \wNDiag_9[49] , \wNDiag_9[48] , \wNDiag_9[47] , \wNDiag_9[46] , 
        \wNDiag_9[45] , \wNDiag_9[44] , \wNDiag_9[43] , \wNDiag_9[42] , 
        \wNDiag_9[41] , \wNDiag_9[40] , \wNDiag_9[39] , \wNDiag_9[38] , 
        \wNDiag_9[37] , \wNDiag_9[36] , \wNDiag_9[35] , \wNDiag_9[34] , 
        \wNDiag_9[33] , \wNDiag_9[32] , \wNDiag_9[31] , \wNDiag_9[30] , 
        \wNDiag_9[29] , \wNDiag_9[28] , \wNDiag_9[27] , \wNDiag_9[26] , 
        \wNDiag_9[25] , \wNDiag_9[24] , \wNDiag_9[23] , \wNDiag_9[22] , 
        \wNDiag_9[21] , \wNDiag_9[20] , \wNDiag_9[19] , \wNDiag_9[18] , 
        \wNDiag_9[17] , \wNDiag_9[16] , \wNDiag_9[15] , \wNDiag_9[14] , 
        \wNDiag_9[13] , \wNDiag_9[12] , \wNDiag_9[11] , \wNDiag_9[10] , 
        \wNDiag_9[9] , \wNDiag_9[8] , \wNDiag_9[7] , \wNDiag_9[6] , 
        \wNDiag_9[5] , \wNDiag_9[4] , \wNDiag_9[3] , \wNDiag_9[2] , 
        \wNDiag_9[1] , \wNDiag_9[0] }), .CallOut(\wCall_10[0] ), .ReturnOut(
        \wReturn_9[0] ), .ColOut({\wColumn_10[63] , \wColumn_10[62] , 
        \wColumn_10[61] , \wColumn_10[60] , \wColumn_10[59] , \wColumn_10[58] , 
        \wColumn_10[57] , \wColumn_10[56] , \wColumn_10[55] , \wColumn_10[54] , 
        \wColumn_10[53] , \wColumn_10[52] , \wColumn_10[51] , \wColumn_10[50] , 
        \wColumn_10[49] , \wColumn_10[48] , \wColumn_10[47] , \wColumn_10[46] , 
        \wColumn_10[45] , \wColumn_10[44] , \wColumn_10[43] , \wColumn_10[42] , 
        \wColumn_10[41] , \wColumn_10[40] , \wColumn_10[39] , \wColumn_10[38] , 
        \wColumn_10[37] , \wColumn_10[36] , \wColumn_10[35] , \wColumn_10[34] , 
        \wColumn_10[33] , \wColumn_10[32] , \wColumn_10[31] , \wColumn_10[30] , 
        \wColumn_10[29] , \wColumn_10[28] , \wColumn_10[27] , \wColumn_10[26] , 
        \wColumn_10[25] , \wColumn_10[24] , \wColumn_10[23] , \wColumn_10[22] , 
        \wColumn_10[21] , \wColumn_10[20] , \wColumn_10[19] , \wColumn_10[18] , 
        \wColumn_10[17] , \wColumn_10[16] , \wColumn_10[15] , \wColumn_10[14] , 
        \wColumn_10[13] , \wColumn_10[12] , \wColumn_10[11] , \wColumn_10[10] , 
        \wColumn_10[9] , \wColumn_10[8] , \wColumn_10[7] , \wColumn_10[6] , 
        \wColumn_10[5] , \wColumn_10[4] , \wColumn_10[3] , \wColumn_10[2] , 
        \wColumn_10[1] , \wColumn_10[0] }), .PDiagOut({\wPDiag_10[63] , 
        \wPDiag_10[62] , \wPDiag_10[61] , \wPDiag_10[60] , \wPDiag_10[59] , 
        \wPDiag_10[58] , \wPDiag_10[57] , \wPDiag_10[56] , \wPDiag_10[55] , 
        \wPDiag_10[54] , \wPDiag_10[53] , \wPDiag_10[52] , \wPDiag_10[51] , 
        \wPDiag_10[50] , \wPDiag_10[49] , \wPDiag_10[48] , \wPDiag_10[47] , 
        \wPDiag_10[46] , \wPDiag_10[45] , \wPDiag_10[44] , \wPDiag_10[43] , 
        \wPDiag_10[42] , \wPDiag_10[41] , \wPDiag_10[40] , \wPDiag_10[39] , 
        \wPDiag_10[38] , \wPDiag_10[37] , \wPDiag_10[36] , \wPDiag_10[35] , 
        \wPDiag_10[34] , \wPDiag_10[33] , \wPDiag_10[32] , \wPDiag_10[31] , 
        \wPDiag_10[30] , \wPDiag_10[29] , \wPDiag_10[28] , \wPDiag_10[27] , 
        \wPDiag_10[26] , \wPDiag_10[25] , \wPDiag_10[24] , \wPDiag_10[23] , 
        \wPDiag_10[22] , \wPDiag_10[21] , \wPDiag_10[20] , \wPDiag_10[19] , 
        \wPDiag_10[18] , \wPDiag_10[17] , \wPDiag_10[16] , \wPDiag_10[15] , 
        \wPDiag_10[14] , \wPDiag_10[13] , \wPDiag_10[12] , \wPDiag_10[11] , 
        \wPDiag_10[10] , \wPDiag_10[9] , \wPDiag_10[8] , \wPDiag_10[7] , 
        \wPDiag_10[6] , \wPDiag_10[5] , \wPDiag_10[4] , \wPDiag_10[3] , 
        \wPDiag_10[2] , \wPDiag_10[1] , \wPDiag_10[0] }), .NDiagOut({
        \wNDiag_10[63] , \wNDiag_10[62] , \wNDiag_10[61] , \wNDiag_10[60] , 
        \wNDiag_10[59] , \wNDiag_10[58] , \wNDiag_10[57] , \wNDiag_10[56] , 
        \wNDiag_10[55] , \wNDiag_10[54] , \wNDiag_10[53] , \wNDiag_10[52] , 
        \wNDiag_10[51] , \wNDiag_10[50] , \wNDiag_10[49] , \wNDiag_10[48] , 
        \wNDiag_10[47] , \wNDiag_10[46] , \wNDiag_10[45] , \wNDiag_10[44] , 
        \wNDiag_10[43] , \wNDiag_10[42] , \wNDiag_10[41] , \wNDiag_10[40] , 
        \wNDiag_10[39] , \wNDiag_10[38] , \wNDiag_10[37] , \wNDiag_10[36] , 
        \wNDiag_10[35] , \wNDiag_10[34] , \wNDiag_10[33] , \wNDiag_10[32] , 
        \wNDiag_10[31] , \wNDiag_10[30] , \wNDiag_10[29] , \wNDiag_10[28] , 
        \wNDiag_10[27] , \wNDiag_10[26] , \wNDiag_10[25] , \wNDiag_10[24] , 
        \wNDiag_10[23] , \wNDiag_10[22] , \wNDiag_10[21] , \wNDiag_10[20] , 
        \wNDiag_10[19] , \wNDiag_10[18] , \wNDiag_10[17] , \wNDiag_10[16] , 
        \wNDiag_10[15] , \wNDiag_10[14] , \wNDiag_10[13] , \wNDiag_10[12] , 
        \wNDiag_10[11] , \wNDiag_10[10] , \wNDiag_10[9] , \wNDiag_10[8] , 
        \wNDiag_10[7] , \wNDiag_10[6] , \wNDiag_10[5] , \wNDiag_10[4] , 
        \wNDiag_10[3] , \wNDiag_10[2] , \wNDiag_10[1] , \wNDiag_10[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_26 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_27[6] , \wScan_27[5] , \wScan_27[4] , 
        \wScan_27[3] , \wScan_27[2] , \wScan_27[1] , \wScan_27[0] }), 
        .ScanOut({\wScan_26[6] , \wScan_26[5] , \wScan_26[4] , \wScan_26[3] , 
        \wScan_26[2] , \wScan_26[1] , \wScan_26[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_26[0] ), .ReturnIn(\wReturn_27[0] ), .ColIn({
        \wColumn_26[63] , \wColumn_26[62] , \wColumn_26[61] , \wColumn_26[60] , 
        \wColumn_26[59] , \wColumn_26[58] , \wColumn_26[57] , \wColumn_26[56] , 
        \wColumn_26[55] , \wColumn_26[54] , \wColumn_26[53] , \wColumn_26[52] , 
        \wColumn_26[51] , \wColumn_26[50] , \wColumn_26[49] , \wColumn_26[48] , 
        \wColumn_26[47] , \wColumn_26[46] , \wColumn_26[45] , \wColumn_26[44] , 
        \wColumn_26[43] , \wColumn_26[42] , \wColumn_26[41] , \wColumn_26[40] , 
        \wColumn_26[39] , \wColumn_26[38] , \wColumn_26[37] , \wColumn_26[36] , 
        \wColumn_26[35] , \wColumn_26[34] , \wColumn_26[33] , \wColumn_26[32] , 
        \wColumn_26[31] , \wColumn_26[30] , \wColumn_26[29] , \wColumn_26[28] , 
        \wColumn_26[27] , \wColumn_26[26] , \wColumn_26[25] , \wColumn_26[24] , 
        \wColumn_26[23] , \wColumn_26[22] , \wColumn_26[21] , \wColumn_26[20] , 
        \wColumn_26[19] , \wColumn_26[18] , \wColumn_26[17] , \wColumn_26[16] , 
        \wColumn_26[15] , \wColumn_26[14] , \wColumn_26[13] , \wColumn_26[12] , 
        \wColumn_26[11] , \wColumn_26[10] , \wColumn_26[9] , \wColumn_26[8] , 
        \wColumn_26[7] , \wColumn_26[6] , \wColumn_26[5] , \wColumn_26[4] , 
        \wColumn_26[3] , \wColumn_26[2] , \wColumn_26[1] , \wColumn_26[0] }), 
        .PDiagIn({\wPDiag_26[63] , \wPDiag_26[62] , \wPDiag_26[61] , 
        \wPDiag_26[60] , \wPDiag_26[59] , \wPDiag_26[58] , \wPDiag_26[57] , 
        \wPDiag_26[56] , \wPDiag_26[55] , \wPDiag_26[54] , \wPDiag_26[53] , 
        \wPDiag_26[52] , \wPDiag_26[51] , \wPDiag_26[50] , \wPDiag_26[49] , 
        \wPDiag_26[48] , \wPDiag_26[47] , \wPDiag_26[46] , \wPDiag_26[45] , 
        \wPDiag_26[44] , \wPDiag_26[43] , \wPDiag_26[42] , \wPDiag_26[41] , 
        \wPDiag_26[40] , \wPDiag_26[39] , \wPDiag_26[38] , \wPDiag_26[37] , 
        \wPDiag_26[36] , \wPDiag_26[35] , \wPDiag_26[34] , \wPDiag_26[33] , 
        \wPDiag_26[32] , \wPDiag_26[31] , \wPDiag_26[30] , \wPDiag_26[29] , 
        \wPDiag_26[28] , \wPDiag_26[27] , \wPDiag_26[26] , \wPDiag_26[25] , 
        \wPDiag_26[24] , \wPDiag_26[23] , \wPDiag_26[22] , \wPDiag_26[21] , 
        \wPDiag_26[20] , \wPDiag_26[19] , \wPDiag_26[18] , \wPDiag_26[17] , 
        \wPDiag_26[16] , \wPDiag_26[15] , \wPDiag_26[14] , \wPDiag_26[13] , 
        \wPDiag_26[12] , \wPDiag_26[11] , \wPDiag_26[10] , \wPDiag_26[9] , 
        \wPDiag_26[8] , \wPDiag_26[7] , \wPDiag_26[6] , \wPDiag_26[5] , 
        \wPDiag_26[4] , \wPDiag_26[3] , \wPDiag_26[2] , \wPDiag_26[1] , 
        \wPDiag_26[0] }), .NDiagIn({\wNDiag_26[63] , \wNDiag_26[62] , 
        \wNDiag_26[61] , \wNDiag_26[60] , \wNDiag_26[59] , \wNDiag_26[58] , 
        \wNDiag_26[57] , \wNDiag_26[56] , \wNDiag_26[55] , \wNDiag_26[54] , 
        \wNDiag_26[53] , \wNDiag_26[52] , \wNDiag_26[51] , \wNDiag_26[50] , 
        \wNDiag_26[49] , \wNDiag_26[48] , \wNDiag_26[47] , \wNDiag_26[46] , 
        \wNDiag_26[45] , \wNDiag_26[44] , \wNDiag_26[43] , \wNDiag_26[42] , 
        \wNDiag_26[41] , \wNDiag_26[40] , \wNDiag_26[39] , \wNDiag_26[38] , 
        \wNDiag_26[37] , \wNDiag_26[36] , \wNDiag_26[35] , \wNDiag_26[34] , 
        \wNDiag_26[33] , \wNDiag_26[32] , \wNDiag_26[31] , \wNDiag_26[30] , 
        \wNDiag_26[29] , \wNDiag_26[28] , \wNDiag_26[27] , \wNDiag_26[26] , 
        \wNDiag_26[25] , \wNDiag_26[24] , \wNDiag_26[23] , \wNDiag_26[22] , 
        \wNDiag_26[21] , \wNDiag_26[20] , \wNDiag_26[19] , \wNDiag_26[18] , 
        \wNDiag_26[17] , \wNDiag_26[16] , \wNDiag_26[15] , \wNDiag_26[14] , 
        \wNDiag_26[13] , \wNDiag_26[12] , \wNDiag_26[11] , \wNDiag_26[10] , 
        \wNDiag_26[9] , \wNDiag_26[8] , \wNDiag_26[7] , \wNDiag_26[6] , 
        \wNDiag_26[5] , \wNDiag_26[4] , \wNDiag_26[3] , \wNDiag_26[2] , 
        \wNDiag_26[1] , \wNDiag_26[0] }), .CallOut(\wCall_27[0] ), .ReturnOut(
        \wReturn_26[0] ), .ColOut({\wColumn_27[63] , \wColumn_27[62] , 
        \wColumn_27[61] , \wColumn_27[60] , \wColumn_27[59] , \wColumn_27[58] , 
        \wColumn_27[57] , \wColumn_27[56] , \wColumn_27[55] , \wColumn_27[54] , 
        \wColumn_27[53] , \wColumn_27[52] , \wColumn_27[51] , \wColumn_27[50] , 
        \wColumn_27[49] , \wColumn_27[48] , \wColumn_27[47] , \wColumn_27[46] , 
        \wColumn_27[45] , \wColumn_27[44] , \wColumn_27[43] , \wColumn_27[42] , 
        \wColumn_27[41] , \wColumn_27[40] , \wColumn_27[39] , \wColumn_27[38] , 
        \wColumn_27[37] , \wColumn_27[36] , \wColumn_27[35] , \wColumn_27[34] , 
        \wColumn_27[33] , \wColumn_27[32] , \wColumn_27[31] , \wColumn_27[30] , 
        \wColumn_27[29] , \wColumn_27[28] , \wColumn_27[27] , \wColumn_27[26] , 
        \wColumn_27[25] , \wColumn_27[24] , \wColumn_27[23] , \wColumn_27[22] , 
        \wColumn_27[21] , \wColumn_27[20] , \wColumn_27[19] , \wColumn_27[18] , 
        \wColumn_27[17] , \wColumn_27[16] , \wColumn_27[15] , \wColumn_27[14] , 
        \wColumn_27[13] , \wColumn_27[12] , \wColumn_27[11] , \wColumn_27[10] , 
        \wColumn_27[9] , \wColumn_27[8] , \wColumn_27[7] , \wColumn_27[6] , 
        \wColumn_27[5] , \wColumn_27[4] , \wColumn_27[3] , \wColumn_27[2] , 
        \wColumn_27[1] , \wColumn_27[0] }), .PDiagOut({\wPDiag_27[63] , 
        \wPDiag_27[62] , \wPDiag_27[61] , \wPDiag_27[60] , \wPDiag_27[59] , 
        \wPDiag_27[58] , \wPDiag_27[57] , \wPDiag_27[56] , \wPDiag_27[55] , 
        \wPDiag_27[54] , \wPDiag_27[53] , \wPDiag_27[52] , \wPDiag_27[51] , 
        \wPDiag_27[50] , \wPDiag_27[49] , \wPDiag_27[48] , \wPDiag_27[47] , 
        \wPDiag_27[46] , \wPDiag_27[45] , \wPDiag_27[44] , \wPDiag_27[43] , 
        \wPDiag_27[42] , \wPDiag_27[41] , \wPDiag_27[40] , \wPDiag_27[39] , 
        \wPDiag_27[38] , \wPDiag_27[37] , \wPDiag_27[36] , \wPDiag_27[35] , 
        \wPDiag_27[34] , \wPDiag_27[33] , \wPDiag_27[32] , \wPDiag_27[31] , 
        \wPDiag_27[30] , \wPDiag_27[29] , \wPDiag_27[28] , \wPDiag_27[27] , 
        \wPDiag_27[26] , \wPDiag_27[25] , \wPDiag_27[24] , \wPDiag_27[23] , 
        \wPDiag_27[22] , \wPDiag_27[21] , \wPDiag_27[20] , \wPDiag_27[19] , 
        \wPDiag_27[18] , \wPDiag_27[17] , \wPDiag_27[16] , \wPDiag_27[15] , 
        \wPDiag_27[14] , \wPDiag_27[13] , \wPDiag_27[12] , \wPDiag_27[11] , 
        \wPDiag_27[10] , \wPDiag_27[9] , \wPDiag_27[8] , \wPDiag_27[7] , 
        \wPDiag_27[6] , \wPDiag_27[5] , \wPDiag_27[4] , \wPDiag_27[3] , 
        \wPDiag_27[2] , \wPDiag_27[1] , \wPDiag_27[0] }), .NDiagOut({
        \wNDiag_27[63] , \wNDiag_27[62] , \wNDiag_27[61] , \wNDiag_27[60] , 
        \wNDiag_27[59] , \wNDiag_27[58] , \wNDiag_27[57] , \wNDiag_27[56] , 
        \wNDiag_27[55] , \wNDiag_27[54] , \wNDiag_27[53] , \wNDiag_27[52] , 
        \wNDiag_27[51] , \wNDiag_27[50] , \wNDiag_27[49] , \wNDiag_27[48] , 
        \wNDiag_27[47] , \wNDiag_27[46] , \wNDiag_27[45] , \wNDiag_27[44] , 
        \wNDiag_27[43] , \wNDiag_27[42] , \wNDiag_27[41] , \wNDiag_27[40] , 
        \wNDiag_27[39] , \wNDiag_27[38] , \wNDiag_27[37] , \wNDiag_27[36] , 
        \wNDiag_27[35] , \wNDiag_27[34] , \wNDiag_27[33] , \wNDiag_27[32] , 
        \wNDiag_27[31] , \wNDiag_27[30] , \wNDiag_27[29] , \wNDiag_27[28] , 
        \wNDiag_27[27] , \wNDiag_27[26] , \wNDiag_27[25] , \wNDiag_27[24] , 
        \wNDiag_27[23] , \wNDiag_27[22] , \wNDiag_27[21] , \wNDiag_27[20] , 
        \wNDiag_27[19] , \wNDiag_27[18] , \wNDiag_27[17] , \wNDiag_27[16] , 
        \wNDiag_27[15] , \wNDiag_27[14] , \wNDiag_27[13] , \wNDiag_27[12] , 
        \wNDiag_27[11] , \wNDiag_27[10] , \wNDiag_27[9] , \wNDiag_27[8] , 
        \wNDiag_27[7] , \wNDiag_27[6] , \wNDiag_27[5] , \wNDiag_27[4] , 
        \wNDiag_27[3] , \wNDiag_27[2] , \wNDiag_27[1] , \wNDiag_27[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_48 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_49[6] , \wScan_49[5] , \wScan_49[4] , 
        \wScan_49[3] , \wScan_49[2] , \wScan_49[1] , \wScan_49[0] }), 
        .ScanOut({\wScan_48[6] , \wScan_48[5] , \wScan_48[4] , \wScan_48[3] , 
        \wScan_48[2] , \wScan_48[1] , \wScan_48[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_48[0] ), .ReturnIn(\wReturn_49[0] ), .ColIn({
        \wColumn_48[63] , \wColumn_48[62] , \wColumn_48[61] , \wColumn_48[60] , 
        \wColumn_48[59] , \wColumn_48[58] , \wColumn_48[57] , \wColumn_48[56] , 
        \wColumn_48[55] , \wColumn_48[54] , \wColumn_48[53] , \wColumn_48[52] , 
        \wColumn_48[51] , \wColumn_48[50] , \wColumn_48[49] , \wColumn_48[48] , 
        \wColumn_48[47] , \wColumn_48[46] , \wColumn_48[45] , \wColumn_48[44] , 
        \wColumn_48[43] , \wColumn_48[42] , \wColumn_48[41] , \wColumn_48[40] , 
        \wColumn_48[39] , \wColumn_48[38] , \wColumn_48[37] , \wColumn_48[36] , 
        \wColumn_48[35] , \wColumn_48[34] , \wColumn_48[33] , \wColumn_48[32] , 
        \wColumn_48[31] , \wColumn_48[30] , \wColumn_48[29] , \wColumn_48[28] , 
        \wColumn_48[27] , \wColumn_48[26] , \wColumn_48[25] , \wColumn_48[24] , 
        \wColumn_48[23] , \wColumn_48[22] , \wColumn_48[21] , \wColumn_48[20] , 
        \wColumn_48[19] , \wColumn_48[18] , \wColumn_48[17] , \wColumn_48[16] , 
        \wColumn_48[15] , \wColumn_48[14] , \wColumn_48[13] , \wColumn_48[12] , 
        \wColumn_48[11] , \wColumn_48[10] , \wColumn_48[9] , \wColumn_48[8] , 
        \wColumn_48[7] , \wColumn_48[6] , \wColumn_48[5] , \wColumn_48[4] , 
        \wColumn_48[3] , \wColumn_48[2] , \wColumn_48[1] , \wColumn_48[0] }), 
        .PDiagIn({\wPDiag_48[63] , \wPDiag_48[62] , \wPDiag_48[61] , 
        \wPDiag_48[60] , \wPDiag_48[59] , \wPDiag_48[58] , \wPDiag_48[57] , 
        \wPDiag_48[56] , \wPDiag_48[55] , \wPDiag_48[54] , \wPDiag_48[53] , 
        \wPDiag_48[52] , \wPDiag_48[51] , \wPDiag_48[50] , \wPDiag_48[49] , 
        \wPDiag_48[48] , \wPDiag_48[47] , \wPDiag_48[46] , \wPDiag_48[45] , 
        \wPDiag_48[44] , \wPDiag_48[43] , \wPDiag_48[42] , \wPDiag_48[41] , 
        \wPDiag_48[40] , \wPDiag_48[39] , \wPDiag_48[38] , \wPDiag_48[37] , 
        \wPDiag_48[36] , \wPDiag_48[35] , \wPDiag_48[34] , \wPDiag_48[33] , 
        \wPDiag_48[32] , \wPDiag_48[31] , \wPDiag_48[30] , \wPDiag_48[29] , 
        \wPDiag_48[28] , \wPDiag_48[27] , \wPDiag_48[26] , \wPDiag_48[25] , 
        \wPDiag_48[24] , \wPDiag_48[23] , \wPDiag_48[22] , \wPDiag_48[21] , 
        \wPDiag_48[20] , \wPDiag_48[19] , \wPDiag_48[18] , \wPDiag_48[17] , 
        \wPDiag_48[16] , \wPDiag_48[15] , \wPDiag_48[14] , \wPDiag_48[13] , 
        \wPDiag_48[12] , \wPDiag_48[11] , \wPDiag_48[10] , \wPDiag_48[9] , 
        \wPDiag_48[8] , \wPDiag_48[7] , \wPDiag_48[6] , \wPDiag_48[5] , 
        \wPDiag_48[4] , \wPDiag_48[3] , \wPDiag_48[2] , \wPDiag_48[1] , 
        \wPDiag_48[0] }), .NDiagIn({\wNDiag_48[63] , \wNDiag_48[62] , 
        \wNDiag_48[61] , \wNDiag_48[60] , \wNDiag_48[59] , \wNDiag_48[58] , 
        \wNDiag_48[57] , \wNDiag_48[56] , \wNDiag_48[55] , \wNDiag_48[54] , 
        \wNDiag_48[53] , \wNDiag_48[52] , \wNDiag_48[51] , \wNDiag_48[50] , 
        \wNDiag_48[49] , \wNDiag_48[48] , \wNDiag_48[47] , \wNDiag_48[46] , 
        \wNDiag_48[45] , \wNDiag_48[44] , \wNDiag_48[43] , \wNDiag_48[42] , 
        \wNDiag_48[41] , \wNDiag_48[40] , \wNDiag_48[39] , \wNDiag_48[38] , 
        \wNDiag_48[37] , \wNDiag_48[36] , \wNDiag_48[35] , \wNDiag_48[34] , 
        \wNDiag_48[33] , \wNDiag_48[32] , \wNDiag_48[31] , \wNDiag_48[30] , 
        \wNDiag_48[29] , \wNDiag_48[28] , \wNDiag_48[27] , \wNDiag_48[26] , 
        \wNDiag_48[25] , \wNDiag_48[24] , \wNDiag_48[23] , \wNDiag_48[22] , 
        \wNDiag_48[21] , \wNDiag_48[20] , \wNDiag_48[19] , \wNDiag_48[18] , 
        \wNDiag_48[17] , \wNDiag_48[16] , \wNDiag_48[15] , \wNDiag_48[14] , 
        \wNDiag_48[13] , \wNDiag_48[12] , \wNDiag_48[11] , \wNDiag_48[10] , 
        \wNDiag_48[9] , \wNDiag_48[8] , \wNDiag_48[7] , \wNDiag_48[6] , 
        \wNDiag_48[5] , \wNDiag_48[4] , \wNDiag_48[3] , \wNDiag_48[2] , 
        \wNDiag_48[1] , \wNDiag_48[0] }), .CallOut(\wCall_49[0] ), .ReturnOut(
        \wReturn_48[0] ), .ColOut({\wColumn_49[63] , \wColumn_49[62] , 
        \wColumn_49[61] , \wColumn_49[60] , \wColumn_49[59] , \wColumn_49[58] , 
        \wColumn_49[57] , \wColumn_49[56] , \wColumn_49[55] , \wColumn_49[54] , 
        \wColumn_49[53] , \wColumn_49[52] , \wColumn_49[51] , \wColumn_49[50] , 
        \wColumn_49[49] , \wColumn_49[48] , \wColumn_49[47] , \wColumn_49[46] , 
        \wColumn_49[45] , \wColumn_49[44] , \wColumn_49[43] , \wColumn_49[42] , 
        \wColumn_49[41] , \wColumn_49[40] , \wColumn_49[39] , \wColumn_49[38] , 
        \wColumn_49[37] , \wColumn_49[36] , \wColumn_49[35] , \wColumn_49[34] , 
        \wColumn_49[33] , \wColumn_49[32] , \wColumn_49[31] , \wColumn_49[30] , 
        \wColumn_49[29] , \wColumn_49[28] , \wColumn_49[27] , \wColumn_49[26] , 
        \wColumn_49[25] , \wColumn_49[24] , \wColumn_49[23] , \wColumn_49[22] , 
        \wColumn_49[21] , \wColumn_49[20] , \wColumn_49[19] , \wColumn_49[18] , 
        \wColumn_49[17] , \wColumn_49[16] , \wColumn_49[15] , \wColumn_49[14] , 
        \wColumn_49[13] , \wColumn_49[12] , \wColumn_49[11] , \wColumn_49[10] , 
        \wColumn_49[9] , \wColumn_49[8] , \wColumn_49[7] , \wColumn_49[6] , 
        \wColumn_49[5] , \wColumn_49[4] , \wColumn_49[3] , \wColumn_49[2] , 
        \wColumn_49[1] , \wColumn_49[0] }), .PDiagOut({\wPDiag_49[63] , 
        \wPDiag_49[62] , \wPDiag_49[61] , \wPDiag_49[60] , \wPDiag_49[59] , 
        \wPDiag_49[58] , \wPDiag_49[57] , \wPDiag_49[56] , \wPDiag_49[55] , 
        \wPDiag_49[54] , \wPDiag_49[53] , \wPDiag_49[52] , \wPDiag_49[51] , 
        \wPDiag_49[50] , \wPDiag_49[49] , \wPDiag_49[48] , \wPDiag_49[47] , 
        \wPDiag_49[46] , \wPDiag_49[45] , \wPDiag_49[44] , \wPDiag_49[43] , 
        \wPDiag_49[42] , \wPDiag_49[41] , \wPDiag_49[40] , \wPDiag_49[39] , 
        \wPDiag_49[38] , \wPDiag_49[37] , \wPDiag_49[36] , \wPDiag_49[35] , 
        \wPDiag_49[34] , \wPDiag_49[33] , \wPDiag_49[32] , \wPDiag_49[31] , 
        \wPDiag_49[30] , \wPDiag_49[29] , \wPDiag_49[28] , \wPDiag_49[27] , 
        \wPDiag_49[26] , \wPDiag_49[25] , \wPDiag_49[24] , \wPDiag_49[23] , 
        \wPDiag_49[22] , \wPDiag_49[21] , \wPDiag_49[20] , \wPDiag_49[19] , 
        \wPDiag_49[18] , \wPDiag_49[17] , \wPDiag_49[16] , \wPDiag_49[15] , 
        \wPDiag_49[14] , \wPDiag_49[13] , \wPDiag_49[12] , \wPDiag_49[11] , 
        \wPDiag_49[10] , \wPDiag_49[9] , \wPDiag_49[8] , \wPDiag_49[7] , 
        \wPDiag_49[6] , \wPDiag_49[5] , \wPDiag_49[4] , \wPDiag_49[3] , 
        \wPDiag_49[2] , \wPDiag_49[1] , \wPDiag_49[0] }), .NDiagOut({
        \wNDiag_49[63] , \wNDiag_49[62] , \wNDiag_49[61] , \wNDiag_49[60] , 
        \wNDiag_49[59] , \wNDiag_49[58] , \wNDiag_49[57] , \wNDiag_49[56] , 
        \wNDiag_49[55] , \wNDiag_49[54] , \wNDiag_49[53] , \wNDiag_49[52] , 
        \wNDiag_49[51] , \wNDiag_49[50] , \wNDiag_49[49] , \wNDiag_49[48] , 
        \wNDiag_49[47] , \wNDiag_49[46] , \wNDiag_49[45] , \wNDiag_49[44] , 
        \wNDiag_49[43] , \wNDiag_49[42] , \wNDiag_49[41] , \wNDiag_49[40] , 
        \wNDiag_49[39] , \wNDiag_49[38] , \wNDiag_49[37] , \wNDiag_49[36] , 
        \wNDiag_49[35] , \wNDiag_49[34] , \wNDiag_49[33] , \wNDiag_49[32] , 
        \wNDiag_49[31] , \wNDiag_49[30] , \wNDiag_49[29] , \wNDiag_49[28] , 
        \wNDiag_49[27] , \wNDiag_49[26] , \wNDiag_49[25] , \wNDiag_49[24] , 
        \wNDiag_49[23] , \wNDiag_49[22] , \wNDiag_49[21] , \wNDiag_49[20] , 
        \wNDiag_49[19] , \wNDiag_49[18] , \wNDiag_49[17] , \wNDiag_49[16] , 
        \wNDiag_49[15] , \wNDiag_49[14] , \wNDiag_49[13] , \wNDiag_49[12] , 
        \wNDiag_49[11] , \wNDiag_49[10] , \wNDiag_49[9] , \wNDiag_49[8] , 
        \wNDiag_49[7] , \wNDiag_49[6] , \wNDiag_49[5] , \wNDiag_49[4] , 
        \wNDiag_49[3] , \wNDiag_49[2] , \wNDiag_49[1] , \wNDiag_49[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_43 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_44[6] , \wScan_44[5] , \wScan_44[4] , 
        \wScan_44[3] , \wScan_44[2] , \wScan_44[1] , \wScan_44[0] }), 
        .ScanOut({\wScan_43[6] , \wScan_43[5] , \wScan_43[4] , \wScan_43[3] , 
        \wScan_43[2] , \wScan_43[1] , \wScan_43[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_43[0] ), .ReturnIn(\wReturn_44[0] ), .ColIn({
        \wColumn_43[63] , \wColumn_43[62] , \wColumn_43[61] , \wColumn_43[60] , 
        \wColumn_43[59] , \wColumn_43[58] , \wColumn_43[57] , \wColumn_43[56] , 
        \wColumn_43[55] , \wColumn_43[54] , \wColumn_43[53] , \wColumn_43[52] , 
        \wColumn_43[51] , \wColumn_43[50] , \wColumn_43[49] , \wColumn_43[48] , 
        \wColumn_43[47] , \wColumn_43[46] , \wColumn_43[45] , \wColumn_43[44] , 
        \wColumn_43[43] , \wColumn_43[42] , \wColumn_43[41] , \wColumn_43[40] , 
        \wColumn_43[39] , \wColumn_43[38] , \wColumn_43[37] , \wColumn_43[36] , 
        \wColumn_43[35] , \wColumn_43[34] , \wColumn_43[33] , \wColumn_43[32] , 
        \wColumn_43[31] , \wColumn_43[30] , \wColumn_43[29] , \wColumn_43[28] , 
        \wColumn_43[27] , \wColumn_43[26] , \wColumn_43[25] , \wColumn_43[24] , 
        \wColumn_43[23] , \wColumn_43[22] , \wColumn_43[21] , \wColumn_43[20] , 
        \wColumn_43[19] , \wColumn_43[18] , \wColumn_43[17] , \wColumn_43[16] , 
        \wColumn_43[15] , \wColumn_43[14] , \wColumn_43[13] , \wColumn_43[12] , 
        \wColumn_43[11] , \wColumn_43[10] , \wColumn_43[9] , \wColumn_43[8] , 
        \wColumn_43[7] , \wColumn_43[6] , \wColumn_43[5] , \wColumn_43[4] , 
        \wColumn_43[3] , \wColumn_43[2] , \wColumn_43[1] , \wColumn_43[0] }), 
        .PDiagIn({\wPDiag_43[63] , \wPDiag_43[62] , \wPDiag_43[61] , 
        \wPDiag_43[60] , \wPDiag_43[59] , \wPDiag_43[58] , \wPDiag_43[57] , 
        \wPDiag_43[56] , \wPDiag_43[55] , \wPDiag_43[54] , \wPDiag_43[53] , 
        \wPDiag_43[52] , \wPDiag_43[51] , \wPDiag_43[50] , \wPDiag_43[49] , 
        \wPDiag_43[48] , \wPDiag_43[47] , \wPDiag_43[46] , \wPDiag_43[45] , 
        \wPDiag_43[44] , \wPDiag_43[43] , \wPDiag_43[42] , \wPDiag_43[41] , 
        \wPDiag_43[40] , \wPDiag_43[39] , \wPDiag_43[38] , \wPDiag_43[37] , 
        \wPDiag_43[36] , \wPDiag_43[35] , \wPDiag_43[34] , \wPDiag_43[33] , 
        \wPDiag_43[32] , \wPDiag_43[31] , \wPDiag_43[30] , \wPDiag_43[29] , 
        \wPDiag_43[28] , \wPDiag_43[27] , \wPDiag_43[26] , \wPDiag_43[25] , 
        \wPDiag_43[24] , \wPDiag_43[23] , \wPDiag_43[22] , \wPDiag_43[21] , 
        \wPDiag_43[20] , \wPDiag_43[19] , \wPDiag_43[18] , \wPDiag_43[17] , 
        \wPDiag_43[16] , \wPDiag_43[15] , \wPDiag_43[14] , \wPDiag_43[13] , 
        \wPDiag_43[12] , \wPDiag_43[11] , \wPDiag_43[10] , \wPDiag_43[9] , 
        \wPDiag_43[8] , \wPDiag_43[7] , \wPDiag_43[6] , \wPDiag_43[5] , 
        \wPDiag_43[4] , \wPDiag_43[3] , \wPDiag_43[2] , \wPDiag_43[1] , 
        \wPDiag_43[0] }), .NDiagIn({\wNDiag_43[63] , \wNDiag_43[62] , 
        \wNDiag_43[61] , \wNDiag_43[60] , \wNDiag_43[59] , \wNDiag_43[58] , 
        \wNDiag_43[57] , \wNDiag_43[56] , \wNDiag_43[55] , \wNDiag_43[54] , 
        \wNDiag_43[53] , \wNDiag_43[52] , \wNDiag_43[51] , \wNDiag_43[50] , 
        \wNDiag_43[49] , \wNDiag_43[48] , \wNDiag_43[47] , \wNDiag_43[46] , 
        \wNDiag_43[45] , \wNDiag_43[44] , \wNDiag_43[43] , \wNDiag_43[42] , 
        \wNDiag_43[41] , \wNDiag_43[40] , \wNDiag_43[39] , \wNDiag_43[38] , 
        \wNDiag_43[37] , \wNDiag_43[36] , \wNDiag_43[35] , \wNDiag_43[34] , 
        \wNDiag_43[33] , \wNDiag_43[32] , \wNDiag_43[31] , \wNDiag_43[30] , 
        \wNDiag_43[29] , \wNDiag_43[28] , \wNDiag_43[27] , \wNDiag_43[26] , 
        \wNDiag_43[25] , \wNDiag_43[24] , \wNDiag_43[23] , \wNDiag_43[22] , 
        \wNDiag_43[21] , \wNDiag_43[20] , \wNDiag_43[19] , \wNDiag_43[18] , 
        \wNDiag_43[17] , \wNDiag_43[16] , \wNDiag_43[15] , \wNDiag_43[14] , 
        \wNDiag_43[13] , \wNDiag_43[12] , \wNDiag_43[11] , \wNDiag_43[10] , 
        \wNDiag_43[9] , \wNDiag_43[8] , \wNDiag_43[7] , \wNDiag_43[6] , 
        \wNDiag_43[5] , \wNDiag_43[4] , \wNDiag_43[3] , \wNDiag_43[2] , 
        \wNDiag_43[1] , \wNDiag_43[0] }), .CallOut(\wCall_44[0] ), .ReturnOut(
        \wReturn_43[0] ), .ColOut({\wColumn_44[63] , \wColumn_44[62] , 
        \wColumn_44[61] , \wColumn_44[60] , \wColumn_44[59] , \wColumn_44[58] , 
        \wColumn_44[57] , \wColumn_44[56] , \wColumn_44[55] , \wColumn_44[54] , 
        \wColumn_44[53] , \wColumn_44[52] , \wColumn_44[51] , \wColumn_44[50] , 
        \wColumn_44[49] , \wColumn_44[48] , \wColumn_44[47] , \wColumn_44[46] , 
        \wColumn_44[45] , \wColumn_44[44] , \wColumn_44[43] , \wColumn_44[42] , 
        \wColumn_44[41] , \wColumn_44[40] , \wColumn_44[39] , \wColumn_44[38] , 
        \wColumn_44[37] , \wColumn_44[36] , \wColumn_44[35] , \wColumn_44[34] , 
        \wColumn_44[33] , \wColumn_44[32] , \wColumn_44[31] , \wColumn_44[30] , 
        \wColumn_44[29] , \wColumn_44[28] , \wColumn_44[27] , \wColumn_44[26] , 
        \wColumn_44[25] , \wColumn_44[24] , \wColumn_44[23] , \wColumn_44[22] , 
        \wColumn_44[21] , \wColumn_44[20] , \wColumn_44[19] , \wColumn_44[18] , 
        \wColumn_44[17] , \wColumn_44[16] , \wColumn_44[15] , \wColumn_44[14] , 
        \wColumn_44[13] , \wColumn_44[12] , \wColumn_44[11] , \wColumn_44[10] , 
        \wColumn_44[9] , \wColumn_44[8] , \wColumn_44[7] , \wColumn_44[6] , 
        \wColumn_44[5] , \wColumn_44[4] , \wColumn_44[3] , \wColumn_44[2] , 
        \wColumn_44[1] , \wColumn_44[0] }), .PDiagOut({\wPDiag_44[63] , 
        \wPDiag_44[62] , \wPDiag_44[61] , \wPDiag_44[60] , \wPDiag_44[59] , 
        \wPDiag_44[58] , \wPDiag_44[57] , \wPDiag_44[56] , \wPDiag_44[55] , 
        \wPDiag_44[54] , \wPDiag_44[53] , \wPDiag_44[52] , \wPDiag_44[51] , 
        \wPDiag_44[50] , \wPDiag_44[49] , \wPDiag_44[48] , \wPDiag_44[47] , 
        \wPDiag_44[46] , \wPDiag_44[45] , \wPDiag_44[44] , \wPDiag_44[43] , 
        \wPDiag_44[42] , \wPDiag_44[41] , \wPDiag_44[40] , \wPDiag_44[39] , 
        \wPDiag_44[38] , \wPDiag_44[37] , \wPDiag_44[36] , \wPDiag_44[35] , 
        \wPDiag_44[34] , \wPDiag_44[33] , \wPDiag_44[32] , \wPDiag_44[31] , 
        \wPDiag_44[30] , \wPDiag_44[29] , \wPDiag_44[28] , \wPDiag_44[27] , 
        \wPDiag_44[26] , \wPDiag_44[25] , \wPDiag_44[24] , \wPDiag_44[23] , 
        \wPDiag_44[22] , \wPDiag_44[21] , \wPDiag_44[20] , \wPDiag_44[19] , 
        \wPDiag_44[18] , \wPDiag_44[17] , \wPDiag_44[16] , \wPDiag_44[15] , 
        \wPDiag_44[14] , \wPDiag_44[13] , \wPDiag_44[12] , \wPDiag_44[11] , 
        \wPDiag_44[10] , \wPDiag_44[9] , \wPDiag_44[8] , \wPDiag_44[7] , 
        \wPDiag_44[6] , \wPDiag_44[5] , \wPDiag_44[4] , \wPDiag_44[3] , 
        \wPDiag_44[2] , \wPDiag_44[1] , \wPDiag_44[0] }), .NDiagOut({
        \wNDiag_44[63] , \wNDiag_44[62] , \wNDiag_44[61] , \wNDiag_44[60] , 
        \wNDiag_44[59] , \wNDiag_44[58] , \wNDiag_44[57] , \wNDiag_44[56] , 
        \wNDiag_44[55] , \wNDiag_44[54] , \wNDiag_44[53] , \wNDiag_44[52] , 
        \wNDiag_44[51] , \wNDiag_44[50] , \wNDiag_44[49] , \wNDiag_44[48] , 
        \wNDiag_44[47] , \wNDiag_44[46] , \wNDiag_44[45] , \wNDiag_44[44] , 
        \wNDiag_44[43] , \wNDiag_44[42] , \wNDiag_44[41] , \wNDiag_44[40] , 
        \wNDiag_44[39] , \wNDiag_44[38] , \wNDiag_44[37] , \wNDiag_44[36] , 
        \wNDiag_44[35] , \wNDiag_44[34] , \wNDiag_44[33] , \wNDiag_44[32] , 
        \wNDiag_44[31] , \wNDiag_44[30] , \wNDiag_44[29] , \wNDiag_44[28] , 
        \wNDiag_44[27] , \wNDiag_44[26] , \wNDiag_44[25] , \wNDiag_44[24] , 
        \wNDiag_44[23] , \wNDiag_44[22] , \wNDiag_44[21] , \wNDiag_44[20] , 
        \wNDiag_44[19] , \wNDiag_44[18] , \wNDiag_44[17] , \wNDiag_44[16] , 
        \wNDiag_44[15] , \wNDiag_44[14] , \wNDiag_44[13] , \wNDiag_44[12] , 
        \wNDiag_44[11] , \wNDiag_44[10] , \wNDiag_44[9] , \wNDiag_44[8] , 
        \wNDiag_44[7] , \wNDiag_44[6] , \wNDiag_44[5] , \wNDiag_44[4] , 
        \wNDiag_44[3] , \wNDiag_44[2] , \wNDiag_44[1] , \wNDiag_44[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_58 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_59[6] , \wScan_59[5] , \wScan_59[4] , 
        \wScan_59[3] , \wScan_59[2] , \wScan_59[1] , \wScan_59[0] }), 
        .ScanOut({\wScan_58[6] , \wScan_58[5] , \wScan_58[4] , \wScan_58[3] , 
        \wScan_58[2] , \wScan_58[1] , \wScan_58[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_58[0] ), .ReturnIn(\wReturn_59[0] ), .ColIn({
        \wColumn_58[63] , \wColumn_58[62] , \wColumn_58[61] , \wColumn_58[60] , 
        \wColumn_58[59] , \wColumn_58[58] , \wColumn_58[57] , \wColumn_58[56] , 
        \wColumn_58[55] , \wColumn_58[54] , \wColumn_58[53] , \wColumn_58[52] , 
        \wColumn_58[51] , \wColumn_58[50] , \wColumn_58[49] , \wColumn_58[48] , 
        \wColumn_58[47] , \wColumn_58[46] , \wColumn_58[45] , \wColumn_58[44] , 
        \wColumn_58[43] , \wColumn_58[42] , \wColumn_58[41] , \wColumn_58[40] , 
        \wColumn_58[39] , \wColumn_58[38] , \wColumn_58[37] , \wColumn_58[36] , 
        \wColumn_58[35] , \wColumn_58[34] , \wColumn_58[33] , \wColumn_58[32] , 
        \wColumn_58[31] , \wColumn_58[30] , \wColumn_58[29] , \wColumn_58[28] , 
        \wColumn_58[27] , \wColumn_58[26] , \wColumn_58[25] , \wColumn_58[24] , 
        \wColumn_58[23] , \wColumn_58[22] , \wColumn_58[21] , \wColumn_58[20] , 
        \wColumn_58[19] , \wColumn_58[18] , \wColumn_58[17] , \wColumn_58[16] , 
        \wColumn_58[15] , \wColumn_58[14] , \wColumn_58[13] , \wColumn_58[12] , 
        \wColumn_58[11] , \wColumn_58[10] , \wColumn_58[9] , \wColumn_58[8] , 
        \wColumn_58[7] , \wColumn_58[6] , \wColumn_58[5] , \wColumn_58[4] , 
        \wColumn_58[3] , \wColumn_58[2] , \wColumn_58[1] , \wColumn_58[0] }), 
        .PDiagIn({\wPDiag_58[63] , \wPDiag_58[62] , \wPDiag_58[61] , 
        \wPDiag_58[60] , \wPDiag_58[59] , \wPDiag_58[58] , \wPDiag_58[57] , 
        \wPDiag_58[56] , \wPDiag_58[55] , \wPDiag_58[54] , \wPDiag_58[53] , 
        \wPDiag_58[52] , \wPDiag_58[51] , \wPDiag_58[50] , \wPDiag_58[49] , 
        \wPDiag_58[48] , \wPDiag_58[47] , \wPDiag_58[46] , \wPDiag_58[45] , 
        \wPDiag_58[44] , \wPDiag_58[43] , \wPDiag_58[42] , \wPDiag_58[41] , 
        \wPDiag_58[40] , \wPDiag_58[39] , \wPDiag_58[38] , \wPDiag_58[37] , 
        \wPDiag_58[36] , \wPDiag_58[35] , \wPDiag_58[34] , \wPDiag_58[33] , 
        \wPDiag_58[32] , \wPDiag_58[31] , \wPDiag_58[30] , \wPDiag_58[29] , 
        \wPDiag_58[28] , \wPDiag_58[27] , \wPDiag_58[26] , \wPDiag_58[25] , 
        \wPDiag_58[24] , \wPDiag_58[23] , \wPDiag_58[22] , \wPDiag_58[21] , 
        \wPDiag_58[20] , \wPDiag_58[19] , \wPDiag_58[18] , \wPDiag_58[17] , 
        \wPDiag_58[16] , \wPDiag_58[15] , \wPDiag_58[14] , \wPDiag_58[13] , 
        \wPDiag_58[12] , \wPDiag_58[11] , \wPDiag_58[10] , \wPDiag_58[9] , 
        \wPDiag_58[8] , \wPDiag_58[7] , \wPDiag_58[6] , \wPDiag_58[5] , 
        \wPDiag_58[4] , \wPDiag_58[3] , \wPDiag_58[2] , \wPDiag_58[1] , 
        \wPDiag_58[0] }), .NDiagIn({\wNDiag_58[63] , \wNDiag_58[62] , 
        \wNDiag_58[61] , \wNDiag_58[60] , \wNDiag_58[59] , \wNDiag_58[58] , 
        \wNDiag_58[57] , \wNDiag_58[56] , \wNDiag_58[55] , \wNDiag_58[54] , 
        \wNDiag_58[53] , \wNDiag_58[52] , \wNDiag_58[51] , \wNDiag_58[50] , 
        \wNDiag_58[49] , \wNDiag_58[48] , \wNDiag_58[47] , \wNDiag_58[46] , 
        \wNDiag_58[45] , \wNDiag_58[44] , \wNDiag_58[43] , \wNDiag_58[42] , 
        \wNDiag_58[41] , \wNDiag_58[40] , \wNDiag_58[39] , \wNDiag_58[38] , 
        \wNDiag_58[37] , \wNDiag_58[36] , \wNDiag_58[35] , \wNDiag_58[34] , 
        \wNDiag_58[33] , \wNDiag_58[32] , \wNDiag_58[31] , \wNDiag_58[30] , 
        \wNDiag_58[29] , \wNDiag_58[28] , \wNDiag_58[27] , \wNDiag_58[26] , 
        \wNDiag_58[25] , \wNDiag_58[24] , \wNDiag_58[23] , \wNDiag_58[22] , 
        \wNDiag_58[21] , \wNDiag_58[20] , \wNDiag_58[19] , \wNDiag_58[18] , 
        \wNDiag_58[17] , \wNDiag_58[16] , \wNDiag_58[15] , \wNDiag_58[14] , 
        \wNDiag_58[13] , \wNDiag_58[12] , \wNDiag_58[11] , \wNDiag_58[10] , 
        \wNDiag_58[9] , \wNDiag_58[8] , \wNDiag_58[7] , \wNDiag_58[6] , 
        \wNDiag_58[5] , \wNDiag_58[4] , \wNDiag_58[3] , \wNDiag_58[2] , 
        \wNDiag_58[1] , \wNDiag_58[0] }), .CallOut(\wCall_59[0] ), .ReturnOut(
        \wReturn_58[0] ), .ColOut({\wColumn_59[63] , \wColumn_59[62] , 
        \wColumn_59[61] , \wColumn_59[60] , \wColumn_59[59] , \wColumn_59[58] , 
        \wColumn_59[57] , \wColumn_59[56] , \wColumn_59[55] , \wColumn_59[54] , 
        \wColumn_59[53] , \wColumn_59[52] , \wColumn_59[51] , \wColumn_59[50] , 
        \wColumn_59[49] , \wColumn_59[48] , \wColumn_59[47] , \wColumn_59[46] , 
        \wColumn_59[45] , \wColumn_59[44] , \wColumn_59[43] , \wColumn_59[42] , 
        \wColumn_59[41] , \wColumn_59[40] , \wColumn_59[39] , \wColumn_59[38] , 
        \wColumn_59[37] , \wColumn_59[36] , \wColumn_59[35] , \wColumn_59[34] , 
        \wColumn_59[33] , \wColumn_59[32] , \wColumn_59[31] , \wColumn_59[30] , 
        \wColumn_59[29] , \wColumn_59[28] , \wColumn_59[27] , \wColumn_59[26] , 
        \wColumn_59[25] , \wColumn_59[24] , \wColumn_59[23] , \wColumn_59[22] , 
        \wColumn_59[21] , \wColumn_59[20] , \wColumn_59[19] , \wColumn_59[18] , 
        \wColumn_59[17] , \wColumn_59[16] , \wColumn_59[15] , \wColumn_59[14] , 
        \wColumn_59[13] , \wColumn_59[12] , \wColumn_59[11] , \wColumn_59[10] , 
        \wColumn_59[9] , \wColumn_59[8] , \wColumn_59[7] , \wColumn_59[6] , 
        \wColumn_59[5] , \wColumn_59[4] , \wColumn_59[3] , \wColumn_59[2] , 
        \wColumn_59[1] , \wColumn_59[0] }), .PDiagOut({\wPDiag_59[63] , 
        \wPDiag_59[62] , \wPDiag_59[61] , \wPDiag_59[60] , \wPDiag_59[59] , 
        \wPDiag_59[58] , \wPDiag_59[57] , \wPDiag_59[56] , \wPDiag_59[55] , 
        \wPDiag_59[54] , \wPDiag_59[53] , \wPDiag_59[52] , \wPDiag_59[51] , 
        \wPDiag_59[50] , \wPDiag_59[49] , \wPDiag_59[48] , \wPDiag_59[47] , 
        \wPDiag_59[46] , \wPDiag_59[45] , \wPDiag_59[44] , \wPDiag_59[43] , 
        \wPDiag_59[42] , \wPDiag_59[41] , \wPDiag_59[40] , \wPDiag_59[39] , 
        \wPDiag_59[38] , \wPDiag_59[37] , \wPDiag_59[36] , \wPDiag_59[35] , 
        \wPDiag_59[34] , \wPDiag_59[33] , \wPDiag_59[32] , \wPDiag_59[31] , 
        \wPDiag_59[30] , \wPDiag_59[29] , \wPDiag_59[28] , \wPDiag_59[27] , 
        \wPDiag_59[26] , \wPDiag_59[25] , \wPDiag_59[24] , \wPDiag_59[23] , 
        \wPDiag_59[22] , \wPDiag_59[21] , \wPDiag_59[20] , \wPDiag_59[19] , 
        \wPDiag_59[18] , \wPDiag_59[17] , \wPDiag_59[16] , \wPDiag_59[15] , 
        \wPDiag_59[14] , \wPDiag_59[13] , \wPDiag_59[12] , \wPDiag_59[11] , 
        \wPDiag_59[10] , \wPDiag_59[9] , \wPDiag_59[8] , \wPDiag_59[7] , 
        \wPDiag_59[6] , \wPDiag_59[5] , \wPDiag_59[4] , \wPDiag_59[3] , 
        \wPDiag_59[2] , \wPDiag_59[1] , \wPDiag_59[0] }), .NDiagOut({
        \wNDiag_59[63] , \wNDiag_59[62] , \wNDiag_59[61] , \wNDiag_59[60] , 
        \wNDiag_59[59] , \wNDiag_59[58] , \wNDiag_59[57] , \wNDiag_59[56] , 
        \wNDiag_59[55] , \wNDiag_59[54] , \wNDiag_59[53] , \wNDiag_59[52] , 
        \wNDiag_59[51] , \wNDiag_59[50] , \wNDiag_59[49] , \wNDiag_59[48] , 
        \wNDiag_59[47] , \wNDiag_59[46] , \wNDiag_59[45] , \wNDiag_59[44] , 
        \wNDiag_59[43] , \wNDiag_59[42] , \wNDiag_59[41] , \wNDiag_59[40] , 
        \wNDiag_59[39] , \wNDiag_59[38] , \wNDiag_59[37] , \wNDiag_59[36] , 
        \wNDiag_59[35] , \wNDiag_59[34] , \wNDiag_59[33] , \wNDiag_59[32] , 
        \wNDiag_59[31] , \wNDiag_59[30] , \wNDiag_59[29] , \wNDiag_59[28] , 
        \wNDiag_59[27] , \wNDiag_59[26] , \wNDiag_59[25] , \wNDiag_59[24] , 
        \wNDiag_59[23] , \wNDiag_59[22] , \wNDiag_59[21] , \wNDiag_59[20] , 
        \wNDiag_59[19] , \wNDiag_59[18] , \wNDiag_59[17] , \wNDiag_59[16] , 
        \wNDiag_59[15] , \wNDiag_59[14] , \wNDiag_59[13] , \wNDiag_59[12] , 
        \wNDiag_59[11] , \wNDiag_59[10] , \wNDiag_59[9] , \wNDiag_59[8] , 
        \wNDiag_59[7] , \wNDiag_59[6] , \wNDiag_59[5] , \wNDiag_59[4] , 
        \wNDiag_59[3] , \wNDiag_59[2] , \wNDiag_59[1] , \wNDiag_59[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_11 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_12[6] , \wScan_12[5] , \wScan_12[4] , 
        \wScan_12[3] , \wScan_12[2] , \wScan_12[1] , \wScan_12[0] }), 
        .ScanOut({\wScan_11[6] , \wScan_11[5] , \wScan_11[4] , \wScan_11[3] , 
        \wScan_11[2] , \wScan_11[1] , \wScan_11[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_11[0] ), .ReturnIn(\wReturn_12[0] ), .ColIn({
        \wColumn_11[63] , \wColumn_11[62] , \wColumn_11[61] , \wColumn_11[60] , 
        \wColumn_11[59] , \wColumn_11[58] , \wColumn_11[57] , \wColumn_11[56] , 
        \wColumn_11[55] , \wColumn_11[54] , \wColumn_11[53] , \wColumn_11[52] , 
        \wColumn_11[51] , \wColumn_11[50] , \wColumn_11[49] , \wColumn_11[48] , 
        \wColumn_11[47] , \wColumn_11[46] , \wColumn_11[45] , \wColumn_11[44] , 
        \wColumn_11[43] , \wColumn_11[42] , \wColumn_11[41] , \wColumn_11[40] , 
        \wColumn_11[39] , \wColumn_11[38] , \wColumn_11[37] , \wColumn_11[36] , 
        \wColumn_11[35] , \wColumn_11[34] , \wColumn_11[33] , \wColumn_11[32] , 
        \wColumn_11[31] , \wColumn_11[30] , \wColumn_11[29] , \wColumn_11[28] , 
        \wColumn_11[27] , \wColumn_11[26] , \wColumn_11[25] , \wColumn_11[24] , 
        \wColumn_11[23] , \wColumn_11[22] , \wColumn_11[21] , \wColumn_11[20] , 
        \wColumn_11[19] , \wColumn_11[18] , \wColumn_11[17] , \wColumn_11[16] , 
        \wColumn_11[15] , \wColumn_11[14] , \wColumn_11[13] , \wColumn_11[12] , 
        \wColumn_11[11] , \wColumn_11[10] , \wColumn_11[9] , \wColumn_11[8] , 
        \wColumn_11[7] , \wColumn_11[6] , \wColumn_11[5] , \wColumn_11[4] , 
        \wColumn_11[3] , \wColumn_11[2] , \wColumn_11[1] , \wColumn_11[0] }), 
        .PDiagIn({\wPDiag_11[63] , \wPDiag_11[62] , \wPDiag_11[61] , 
        \wPDiag_11[60] , \wPDiag_11[59] , \wPDiag_11[58] , \wPDiag_11[57] , 
        \wPDiag_11[56] , \wPDiag_11[55] , \wPDiag_11[54] , \wPDiag_11[53] , 
        \wPDiag_11[52] , \wPDiag_11[51] , \wPDiag_11[50] , \wPDiag_11[49] , 
        \wPDiag_11[48] , \wPDiag_11[47] , \wPDiag_11[46] , \wPDiag_11[45] , 
        \wPDiag_11[44] , \wPDiag_11[43] , \wPDiag_11[42] , \wPDiag_11[41] , 
        \wPDiag_11[40] , \wPDiag_11[39] , \wPDiag_11[38] , \wPDiag_11[37] , 
        \wPDiag_11[36] , \wPDiag_11[35] , \wPDiag_11[34] , \wPDiag_11[33] , 
        \wPDiag_11[32] , \wPDiag_11[31] , \wPDiag_11[30] , \wPDiag_11[29] , 
        \wPDiag_11[28] , \wPDiag_11[27] , \wPDiag_11[26] , \wPDiag_11[25] , 
        \wPDiag_11[24] , \wPDiag_11[23] , \wPDiag_11[22] , \wPDiag_11[21] , 
        \wPDiag_11[20] , \wPDiag_11[19] , \wPDiag_11[18] , \wPDiag_11[17] , 
        \wPDiag_11[16] , \wPDiag_11[15] , \wPDiag_11[14] , \wPDiag_11[13] , 
        \wPDiag_11[12] , \wPDiag_11[11] , \wPDiag_11[10] , \wPDiag_11[9] , 
        \wPDiag_11[8] , \wPDiag_11[7] , \wPDiag_11[6] , \wPDiag_11[5] , 
        \wPDiag_11[4] , \wPDiag_11[3] , \wPDiag_11[2] , \wPDiag_11[1] , 
        \wPDiag_11[0] }), .NDiagIn({\wNDiag_11[63] , \wNDiag_11[62] , 
        \wNDiag_11[61] , \wNDiag_11[60] , \wNDiag_11[59] , \wNDiag_11[58] , 
        \wNDiag_11[57] , \wNDiag_11[56] , \wNDiag_11[55] , \wNDiag_11[54] , 
        \wNDiag_11[53] , \wNDiag_11[52] , \wNDiag_11[51] , \wNDiag_11[50] , 
        \wNDiag_11[49] , \wNDiag_11[48] , \wNDiag_11[47] , \wNDiag_11[46] , 
        \wNDiag_11[45] , \wNDiag_11[44] , \wNDiag_11[43] , \wNDiag_11[42] , 
        \wNDiag_11[41] , \wNDiag_11[40] , \wNDiag_11[39] , \wNDiag_11[38] , 
        \wNDiag_11[37] , \wNDiag_11[36] , \wNDiag_11[35] , \wNDiag_11[34] , 
        \wNDiag_11[33] , \wNDiag_11[32] , \wNDiag_11[31] , \wNDiag_11[30] , 
        \wNDiag_11[29] , \wNDiag_11[28] , \wNDiag_11[27] , \wNDiag_11[26] , 
        \wNDiag_11[25] , \wNDiag_11[24] , \wNDiag_11[23] , \wNDiag_11[22] , 
        \wNDiag_11[21] , \wNDiag_11[20] , \wNDiag_11[19] , \wNDiag_11[18] , 
        \wNDiag_11[17] , \wNDiag_11[16] , \wNDiag_11[15] , \wNDiag_11[14] , 
        \wNDiag_11[13] , \wNDiag_11[12] , \wNDiag_11[11] , \wNDiag_11[10] , 
        \wNDiag_11[9] , \wNDiag_11[8] , \wNDiag_11[7] , \wNDiag_11[6] , 
        \wNDiag_11[5] , \wNDiag_11[4] , \wNDiag_11[3] , \wNDiag_11[2] , 
        \wNDiag_11[1] , \wNDiag_11[0] }), .CallOut(\wCall_12[0] ), .ReturnOut(
        \wReturn_11[0] ), .ColOut({\wColumn_12[63] , \wColumn_12[62] , 
        \wColumn_12[61] , \wColumn_12[60] , \wColumn_12[59] , \wColumn_12[58] , 
        \wColumn_12[57] , \wColumn_12[56] , \wColumn_12[55] , \wColumn_12[54] , 
        \wColumn_12[53] , \wColumn_12[52] , \wColumn_12[51] , \wColumn_12[50] , 
        \wColumn_12[49] , \wColumn_12[48] , \wColumn_12[47] , \wColumn_12[46] , 
        \wColumn_12[45] , \wColumn_12[44] , \wColumn_12[43] , \wColumn_12[42] , 
        \wColumn_12[41] , \wColumn_12[40] , \wColumn_12[39] , \wColumn_12[38] , 
        \wColumn_12[37] , \wColumn_12[36] , \wColumn_12[35] , \wColumn_12[34] , 
        \wColumn_12[33] , \wColumn_12[32] , \wColumn_12[31] , \wColumn_12[30] , 
        \wColumn_12[29] , \wColumn_12[28] , \wColumn_12[27] , \wColumn_12[26] , 
        \wColumn_12[25] , \wColumn_12[24] , \wColumn_12[23] , \wColumn_12[22] , 
        \wColumn_12[21] , \wColumn_12[20] , \wColumn_12[19] , \wColumn_12[18] , 
        \wColumn_12[17] , \wColumn_12[16] , \wColumn_12[15] , \wColumn_12[14] , 
        \wColumn_12[13] , \wColumn_12[12] , \wColumn_12[11] , \wColumn_12[10] , 
        \wColumn_12[9] , \wColumn_12[8] , \wColumn_12[7] , \wColumn_12[6] , 
        \wColumn_12[5] , \wColumn_12[4] , \wColumn_12[3] , \wColumn_12[2] , 
        \wColumn_12[1] , \wColumn_12[0] }), .PDiagOut({\wPDiag_12[63] , 
        \wPDiag_12[62] , \wPDiag_12[61] , \wPDiag_12[60] , \wPDiag_12[59] , 
        \wPDiag_12[58] , \wPDiag_12[57] , \wPDiag_12[56] , \wPDiag_12[55] , 
        \wPDiag_12[54] , \wPDiag_12[53] , \wPDiag_12[52] , \wPDiag_12[51] , 
        \wPDiag_12[50] , \wPDiag_12[49] , \wPDiag_12[48] , \wPDiag_12[47] , 
        \wPDiag_12[46] , \wPDiag_12[45] , \wPDiag_12[44] , \wPDiag_12[43] , 
        \wPDiag_12[42] , \wPDiag_12[41] , \wPDiag_12[40] , \wPDiag_12[39] , 
        \wPDiag_12[38] , \wPDiag_12[37] , \wPDiag_12[36] , \wPDiag_12[35] , 
        \wPDiag_12[34] , \wPDiag_12[33] , \wPDiag_12[32] , \wPDiag_12[31] , 
        \wPDiag_12[30] , \wPDiag_12[29] , \wPDiag_12[28] , \wPDiag_12[27] , 
        \wPDiag_12[26] , \wPDiag_12[25] , \wPDiag_12[24] , \wPDiag_12[23] , 
        \wPDiag_12[22] , \wPDiag_12[21] , \wPDiag_12[20] , \wPDiag_12[19] , 
        \wPDiag_12[18] , \wPDiag_12[17] , \wPDiag_12[16] , \wPDiag_12[15] , 
        \wPDiag_12[14] , \wPDiag_12[13] , \wPDiag_12[12] , \wPDiag_12[11] , 
        \wPDiag_12[10] , \wPDiag_12[9] , \wPDiag_12[8] , \wPDiag_12[7] , 
        \wPDiag_12[6] , \wPDiag_12[5] , \wPDiag_12[4] , \wPDiag_12[3] , 
        \wPDiag_12[2] , \wPDiag_12[1] , \wPDiag_12[0] }), .NDiagOut({
        \wNDiag_12[63] , \wNDiag_12[62] , \wNDiag_12[61] , \wNDiag_12[60] , 
        \wNDiag_12[59] , \wNDiag_12[58] , \wNDiag_12[57] , \wNDiag_12[56] , 
        \wNDiag_12[55] , \wNDiag_12[54] , \wNDiag_12[53] , \wNDiag_12[52] , 
        \wNDiag_12[51] , \wNDiag_12[50] , \wNDiag_12[49] , \wNDiag_12[48] , 
        \wNDiag_12[47] , \wNDiag_12[46] , \wNDiag_12[45] , \wNDiag_12[44] , 
        \wNDiag_12[43] , \wNDiag_12[42] , \wNDiag_12[41] , \wNDiag_12[40] , 
        \wNDiag_12[39] , \wNDiag_12[38] , \wNDiag_12[37] , \wNDiag_12[36] , 
        \wNDiag_12[35] , \wNDiag_12[34] , \wNDiag_12[33] , \wNDiag_12[32] , 
        \wNDiag_12[31] , \wNDiag_12[30] , \wNDiag_12[29] , \wNDiag_12[28] , 
        \wNDiag_12[27] , \wNDiag_12[26] , \wNDiag_12[25] , \wNDiag_12[24] , 
        \wNDiag_12[23] , \wNDiag_12[22] , \wNDiag_12[21] , \wNDiag_12[20] , 
        \wNDiag_12[19] , \wNDiag_12[18] , \wNDiag_12[17] , \wNDiag_12[16] , 
        \wNDiag_12[15] , \wNDiag_12[14] , \wNDiag_12[13] , \wNDiag_12[12] , 
        \wNDiag_12[11] , \wNDiag_12[10] , \wNDiag_12[9] , \wNDiag_12[8] , 
        \wNDiag_12[7] , \wNDiag_12[6] , \wNDiag_12[5] , \wNDiag_12[4] , 
        \wNDiag_12[3] , \wNDiag_12[2] , \wNDiag_12[1] , \wNDiag_12[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_24 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_25[6] , \wScan_25[5] , \wScan_25[4] , 
        \wScan_25[3] , \wScan_25[2] , \wScan_25[1] , \wScan_25[0] }), 
        .ScanOut({\wScan_24[6] , \wScan_24[5] , \wScan_24[4] , \wScan_24[3] , 
        \wScan_24[2] , \wScan_24[1] , \wScan_24[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_24[0] ), .ReturnIn(\wReturn_25[0] ), .ColIn({
        \wColumn_24[63] , \wColumn_24[62] , \wColumn_24[61] , \wColumn_24[60] , 
        \wColumn_24[59] , \wColumn_24[58] , \wColumn_24[57] , \wColumn_24[56] , 
        \wColumn_24[55] , \wColumn_24[54] , \wColumn_24[53] , \wColumn_24[52] , 
        \wColumn_24[51] , \wColumn_24[50] , \wColumn_24[49] , \wColumn_24[48] , 
        \wColumn_24[47] , \wColumn_24[46] , \wColumn_24[45] , \wColumn_24[44] , 
        \wColumn_24[43] , \wColumn_24[42] , \wColumn_24[41] , \wColumn_24[40] , 
        \wColumn_24[39] , \wColumn_24[38] , \wColumn_24[37] , \wColumn_24[36] , 
        \wColumn_24[35] , \wColumn_24[34] , \wColumn_24[33] , \wColumn_24[32] , 
        \wColumn_24[31] , \wColumn_24[30] , \wColumn_24[29] , \wColumn_24[28] , 
        \wColumn_24[27] , \wColumn_24[26] , \wColumn_24[25] , \wColumn_24[24] , 
        \wColumn_24[23] , \wColumn_24[22] , \wColumn_24[21] , \wColumn_24[20] , 
        \wColumn_24[19] , \wColumn_24[18] , \wColumn_24[17] , \wColumn_24[16] , 
        \wColumn_24[15] , \wColumn_24[14] , \wColumn_24[13] , \wColumn_24[12] , 
        \wColumn_24[11] , \wColumn_24[10] , \wColumn_24[9] , \wColumn_24[8] , 
        \wColumn_24[7] , \wColumn_24[6] , \wColumn_24[5] , \wColumn_24[4] , 
        \wColumn_24[3] , \wColumn_24[2] , \wColumn_24[1] , \wColumn_24[0] }), 
        .PDiagIn({\wPDiag_24[63] , \wPDiag_24[62] , \wPDiag_24[61] , 
        \wPDiag_24[60] , \wPDiag_24[59] , \wPDiag_24[58] , \wPDiag_24[57] , 
        \wPDiag_24[56] , \wPDiag_24[55] , \wPDiag_24[54] , \wPDiag_24[53] , 
        \wPDiag_24[52] , \wPDiag_24[51] , \wPDiag_24[50] , \wPDiag_24[49] , 
        \wPDiag_24[48] , \wPDiag_24[47] , \wPDiag_24[46] , \wPDiag_24[45] , 
        \wPDiag_24[44] , \wPDiag_24[43] , \wPDiag_24[42] , \wPDiag_24[41] , 
        \wPDiag_24[40] , \wPDiag_24[39] , \wPDiag_24[38] , \wPDiag_24[37] , 
        \wPDiag_24[36] , \wPDiag_24[35] , \wPDiag_24[34] , \wPDiag_24[33] , 
        \wPDiag_24[32] , \wPDiag_24[31] , \wPDiag_24[30] , \wPDiag_24[29] , 
        \wPDiag_24[28] , \wPDiag_24[27] , \wPDiag_24[26] , \wPDiag_24[25] , 
        \wPDiag_24[24] , \wPDiag_24[23] , \wPDiag_24[22] , \wPDiag_24[21] , 
        \wPDiag_24[20] , \wPDiag_24[19] , \wPDiag_24[18] , \wPDiag_24[17] , 
        \wPDiag_24[16] , \wPDiag_24[15] , \wPDiag_24[14] , \wPDiag_24[13] , 
        \wPDiag_24[12] , \wPDiag_24[11] , \wPDiag_24[10] , \wPDiag_24[9] , 
        \wPDiag_24[8] , \wPDiag_24[7] , \wPDiag_24[6] , \wPDiag_24[5] , 
        \wPDiag_24[4] , \wPDiag_24[3] , \wPDiag_24[2] , \wPDiag_24[1] , 
        \wPDiag_24[0] }), .NDiagIn({\wNDiag_24[63] , \wNDiag_24[62] , 
        \wNDiag_24[61] , \wNDiag_24[60] , \wNDiag_24[59] , \wNDiag_24[58] , 
        \wNDiag_24[57] , \wNDiag_24[56] , \wNDiag_24[55] , \wNDiag_24[54] , 
        \wNDiag_24[53] , \wNDiag_24[52] , \wNDiag_24[51] , \wNDiag_24[50] , 
        \wNDiag_24[49] , \wNDiag_24[48] , \wNDiag_24[47] , \wNDiag_24[46] , 
        \wNDiag_24[45] , \wNDiag_24[44] , \wNDiag_24[43] , \wNDiag_24[42] , 
        \wNDiag_24[41] , \wNDiag_24[40] , \wNDiag_24[39] , \wNDiag_24[38] , 
        \wNDiag_24[37] , \wNDiag_24[36] , \wNDiag_24[35] , \wNDiag_24[34] , 
        \wNDiag_24[33] , \wNDiag_24[32] , \wNDiag_24[31] , \wNDiag_24[30] , 
        \wNDiag_24[29] , \wNDiag_24[28] , \wNDiag_24[27] , \wNDiag_24[26] , 
        \wNDiag_24[25] , \wNDiag_24[24] , \wNDiag_24[23] , \wNDiag_24[22] , 
        \wNDiag_24[21] , \wNDiag_24[20] , \wNDiag_24[19] , \wNDiag_24[18] , 
        \wNDiag_24[17] , \wNDiag_24[16] , \wNDiag_24[15] , \wNDiag_24[14] , 
        \wNDiag_24[13] , \wNDiag_24[12] , \wNDiag_24[11] , \wNDiag_24[10] , 
        \wNDiag_24[9] , \wNDiag_24[8] , \wNDiag_24[7] , \wNDiag_24[6] , 
        \wNDiag_24[5] , \wNDiag_24[4] , \wNDiag_24[3] , \wNDiag_24[2] , 
        \wNDiag_24[1] , \wNDiag_24[0] }), .CallOut(\wCall_25[0] ), .ReturnOut(
        \wReturn_24[0] ), .ColOut({\wColumn_25[63] , \wColumn_25[62] , 
        \wColumn_25[61] , \wColumn_25[60] , \wColumn_25[59] , \wColumn_25[58] , 
        \wColumn_25[57] , \wColumn_25[56] , \wColumn_25[55] , \wColumn_25[54] , 
        \wColumn_25[53] , \wColumn_25[52] , \wColumn_25[51] , \wColumn_25[50] , 
        \wColumn_25[49] , \wColumn_25[48] , \wColumn_25[47] , \wColumn_25[46] , 
        \wColumn_25[45] , \wColumn_25[44] , \wColumn_25[43] , \wColumn_25[42] , 
        \wColumn_25[41] , \wColumn_25[40] , \wColumn_25[39] , \wColumn_25[38] , 
        \wColumn_25[37] , \wColumn_25[36] , \wColumn_25[35] , \wColumn_25[34] , 
        \wColumn_25[33] , \wColumn_25[32] , \wColumn_25[31] , \wColumn_25[30] , 
        \wColumn_25[29] , \wColumn_25[28] , \wColumn_25[27] , \wColumn_25[26] , 
        \wColumn_25[25] , \wColumn_25[24] , \wColumn_25[23] , \wColumn_25[22] , 
        \wColumn_25[21] , \wColumn_25[20] , \wColumn_25[19] , \wColumn_25[18] , 
        \wColumn_25[17] , \wColumn_25[16] , \wColumn_25[15] , \wColumn_25[14] , 
        \wColumn_25[13] , \wColumn_25[12] , \wColumn_25[11] , \wColumn_25[10] , 
        \wColumn_25[9] , \wColumn_25[8] , \wColumn_25[7] , \wColumn_25[6] , 
        \wColumn_25[5] , \wColumn_25[4] , \wColumn_25[3] , \wColumn_25[2] , 
        \wColumn_25[1] , \wColumn_25[0] }), .PDiagOut({\wPDiag_25[63] , 
        \wPDiag_25[62] , \wPDiag_25[61] , \wPDiag_25[60] , \wPDiag_25[59] , 
        \wPDiag_25[58] , \wPDiag_25[57] , \wPDiag_25[56] , \wPDiag_25[55] , 
        \wPDiag_25[54] , \wPDiag_25[53] , \wPDiag_25[52] , \wPDiag_25[51] , 
        \wPDiag_25[50] , \wPDiag_25[49] , \wPDiag_25[48] , \wPDiag_25[47] , 
        \wPDiag_25[46] , \wPDiag_25[45] , \wPDiag_25[44] , \wPDiag_25[43] , 
        \wPDiag_25[42] , \wPDiag_25[41] , \wPDiag_25[40] , \wPDiag_25[39] , 
        \wPDiag_25[38] , \wPDiag_25[37] , \wPDiag_25[36] , \wPDiag_25[35] , 
        \wPDiag_25[34] , \wPDiag_25[33] , \wPDiag_25[32] , \wPDiag_25[31] , 
        \wPDiag_25[30] , \wPDiag_25[29] , \wPDiag_25[28] , \wPDiag_25[27] , 
        \wPDiag_25[26] , \wPDiag_25[25] , \wPDiag_25[24] , \wPDiag_25[23] , 
        \wPDiag_25[22] , \wPDiag_25[21] , \wPDiag_25[20] , \wPDiag_25[19] , 
        \wPDiag_25[18] , \wPDiag_25[17] , \wPDiag_25[16] , \wPDiag_25[15] , 
        \wPDiag_25[14] , \wPDiag_25[13] , \wPDiag_25[12] , \wPDiag_25[11] , 
        \wPDiag_25[10] , \wPDiag_25[9] , \wPDiag_25[8] , \wPDiag_25[7] , 
        \wPDiag_25[6] , \wPDiag_25[5] , \wPDiag_25[4] , \wPDiag_25[3] , 
        \wPDiag_25[2] , \wPDiag_25[1] , \wPDiag_25[0] }), .NDiagOut({
        \wNDiag_25[63] , \wNDiag_25[62] , \wNDiag_25[61] , \wNDiag_25[60] , 
        \wNDiag_25[59] , \wNDiag_25[58] , \wNDiag_25[57] , \wNDiag_25[56] , 
        \wNDiag_25[55] , \wNDiag_25[54] , \wNDiag_25[53] , \wNDiag_25[52] , 
        \wNDiag_25[51] , \wNDiag_25[50] , \wNDiag_25[49] , \wNDiag_25[48] , 
        \wNDiag_25[47] , \wNDiag_25[46] , \wNDiag_25[45] , \wNDiag_25[44] , 
        \wNDiag_25[43] , \wNDiag_25[42] , \wNDiag_25[41] , \wNDiag_25[40] , 
        \wNDiag_25[39] , \wNDiag_25[38] , \wNDiag_25[37] , \wNDiag_25[36] , 
        \wNDiag_25[35] , \wNDiag_25[34] , \wNDiag_25[33] , \wNDiag_25[32] , 
        \wNDiag_25[31] , \wNDiag_25[30] , \wNDiag_25[29] , \wNDiag_25[28] , 
        \wNDiag_25[27] , \wNDiag_25[26] , \wNDiag_25[25] , \wNDiag_25[24] , 
        \wNDiag_25[23] , \wNDiag_25[22] , \wNDiag_25[21] , \wNDiag_25[20] , 
        \wNDiag_25[19] , \wNDiag_25[18] , \wNDiag_25[17] , \wNDiag_25[16] , 
        \wNDiag_25[15] , \wNDiag_25[14] , \wNDiag_25[13] , \wNDiag_25[12] , 
        \wNDiag_25[11] , \wNDiag_25[10] , \wNDiag_25[9] , \wNDiag_25[8] , 
        \wNDiag_25[7] , \wNDiag_25[6] , \wNDiag_25[5] , \wNDiag_25[4] , 
        \wNDiag_25[3] , \wNDiag_25[2] , \wNDiag_25[1] , \wNDiag_25[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_36 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_37[6] , \wScan_37[5] , \wScan_37[4] , 
        \wScan_37[3] , \wScan_37[2] , \wScan_37[1] , \wScan_37[0] }), 
        .ScanOut({\wScan_36[6] , \wScan_36[5] , \wScan_36[4] , \wScan_36[3] , 
        \wScan_36[2] , \wScan_36[1] , \wScan_36[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_36[0] ), .ReturnIn(\wReturn_37[0] ), .ColIn({
        \wColumn_36[63] , \wColumn_36[62] , \wColumn_36[61] , \wColumn_36[60] , 
        \wColumn_36[59] , \wColumn_36[58] , \wColumn_36[57] , \wColumn_36[56] , 
        \wColumn_36[55] , \wColumn_36[54] , \wColumn_36[53] , \wColumn_36[52] , 
        \wColumn_36[51] , \wColumn_36[50] , \wColumn_36[49] , \wColumn_36[48] , 
        \wColumn_36[47] , \wColumn_36[46] , \wColumn_36[45] , \wColumn_36[44] , 
        \wColumn_36[43] , \wColumn_36[42] , \wColumn_36[41] , \wColumn_36[40] , 
        \wColumn_36[39] , \wColumn_36[38] , \wColumn_36[37] , \wColumn_36[36] , 
        \wColumn_36[35] , \wColumn_36[34] , \wColumn_36[33] , \wColumn_36[32] , 
        \wColumn_36[31] , \wColumn_36[30] , \wColumn_36[29] , \wColumn_36[28] , 
        \wColumn_36[27] , \wColumn_36[26] , \wColumn_36[25] , \wColumn_36[24] , 
        \wColumn_36[23] , \wColumn_36[22] , \wColumn_36[21] , \wColumn_36[20] , 
        \wColumn_36[19] , \wColumn_36[18] , \wColumn_36[17] , \wColumn_36[16] , 
        \wColumn_36[15] , \wColumn_36[14] , \wColumn_36[13] , \wColumn_36[12] , 
        \wColumn_36[11] , \wColumn_36[10] , \wColumn_36[9] , \wColumn_36[8] , 
        \wColumn_36[7] , \wColumn_36[6] , \wColumn_36[5] , \wColumn_36[4] , 
        \wColumn_36[3] , \wColumn_36[2] , \wColumn_36[1] , \wColumn_36[0] }), 
        .PDiagIn({\wPDiag_36[63] , \wPDiag_36[62] , \wPDiag_36[61] , 
        \wPDiag_36[60] , \wPDiag_36[59] , \wPDiag_36[58] , \wPDiag_36[57] , 
        \wPDiag_36[56] , \wPDiag_36[55] , \wPDiag_36[54] , \wPDiag_36[53] , 
        \wPDiag_36[52] , \wPDiag_36[51] , \wPDiag_36[50] , \wPDiag_36[49] , 
        \wPDiag_36[48] , \wPDiag_36[47] , \wPDiag_36[46] , \wPDiag_36[45] , 
        \wPDiag_36[44] , \wPDiag_36[43] , \wPDiag_36[42] , \wPDiag_36[41] , 
        \wPDiag_36[40] , \wPDiag_36[39] , \wPDiag_36[38] , \wPDiag_36[37] , 
        \wPDiag_36[36] , \wPDiag_36[35] , \wPDiag_36[34] , \wPDiag_36[33] , 
        \wPDiag_36[32] , \wPDiag_36[31] , \wPDiag_36[30] , \wPDiag_36[29] , 
        \wPDiag_36[28] , \wPDiag_36[27] , \wPDiag_36[26] , \wPDiag_36[25] , 
        \wPDiag_36[24] , \wPDiag_36[23] , \wPDiag_36[22] , \wPDiag_36[21] , 
        \wPDiag_36[20] , \wPDiag_36[19] , \wPDiag_36[18] , \wPDiag_36[17] , 
        \wPDiag_36[16] , \wPDiag_36[15] , \wPDiag_36[14] , \wPDiag_36[13] , 
        \wPDiag_36[12] , \wPDiag_36[11] , \wPDiag_36[10] , \wPDiag_36[9] , 
        \wPDiag_36[8] , \wPDiag_36[7] , \wPDiag_36[6] , \wPDiag_36[5] , 
        \wPDiag_36[4] , \wPDiag_36[3] , \wPDiag_36[2] , \wPDiag_36[1] , 
        \wPDiag_36[0] }), .NDiagIn({\wNDiag_36[63] , \wNDiag_36[62] , 
        \wNDiag_36[61] , \wNDiag_36[60] , \wNDiag_36[59] , \wNDiag_36[58] , 
        \wNDiag_36[57] , \wNDiag_36[56] , \wNDiag_36[55] , \wNDiag_36[54] , 
        \wNDiag_36[53] , \wNDiag_36[52] , \wNDiag_36[51] , \wNDiag_36[50] , 
        \wNDiag_36[49] , \wNDiag_36[48] , \wNDiag_36[47] , \wNDiag_36[46] , 
        \wNDiag_36[45] , \wNDiag_36[44] , \wNDiag_36[43] , \wNDiag_36[42] , 
        \wNDiag_36[41] , \wNDiag_36[40] , \wNDiag_36[39] , \wNDiag_36[38] , 
        \wNDiag_36[37] , \wNDiag_36[36] , \wNDiag_36[35] , \wNDiag_36[34] , 
        \wNDiag_36[33] , \wNDiag_36[32] , \wNDiag_36[31] , \wNDiag_36[30] , 
        \wNDiag_36[29] , \wNDiag_36[28] , \wNDiag_36[27] , \wNDiag_36[26] , 
        \wNDiag_36[25] , \wNDiag_36[24] , \wNDiag_36[23] , \wNDiag_36[22] , 
        \wNDiag_36[21] , \wNDiag_36[20] , \wNDiag_36[19] , \wNDiag_36[18] , 
        \wNDiag_36[17] , \wNDiag_36[16] , \wNDiag_36[15] , \wNDiag_36[14] , 
        \wNDiag_36[13] , \wNDiag_36[12] , \wNDiag_36[11] , \wNDiag_36[10] , 
        \wNDiag_36[9] , \wNDiag_36[8] , \wNDiag_36[7] , \wNDiag_36[6] , 
        \wNDiag_36[5] , \wNDiag_36[4] , \wNDiag_36[3] , \wNDiag_36[2] , 
        \wNDiag_36[1] , \wNDiag_36[0] }), .CallOut(\wCall_37[0] ), .ReturnOut(
        \wReturn_36[0] ), .ColOut({\wColumn_37[63] , \wColumn_37[62] , 
        \wColumn_37[61] , \wColumn_37[60] , \wColumn_37[59] , \wColumn_37[58] , 
        \wColumn_37[57] , \wColumn_37[56] , \wColumn_37[55] , \wColumn_37[54] , 
        \wColumn_37[53] , \wColumn_37[52] , \wColumn_37[51] , \wColumn_37[50] , 
        \wColumn_37[49] , \wColumn_37[48] , \wColumn_37[47] , \wColumn_37[46] , 
        \wColumn_37[45] , \wColumn_37[44] , \wColumn_37[43] , \wColumn_37[42] , 
        \wColumn_37[41] , \wColumn_37[40] , \wColumn_37[39] , \wColumn_37[38] , 
        \wColumn_37[37] , \wColumn_37[36] , \wColumn_37[35] , \wColumn_37[34] , 
        \wColumn_37[33] , \wColumn_37[32] , \wColumn_37[31] , \wColumn_37[30] , 
        \wColumn_37[29] , \wColumn_37[28] , \wColumn_37[27] , \wColumn_37[26] , 
        \wColumn_37[25] , \wColumn_37[24] , \wColumn_37[23] , \wColumn_37[22] , 
        \wColumn_37[21] , \wColumn_37[20] , \wColumn_37[19] , \wColumn_37[18] , 
        \wColumn_37[17] , \wColumn_37[16] , \wColumn_37[15] , \wColumn_37[14] , 
        \wColumn_37[13] , \wColumn_37[12] , \wColumn_37[11] , \wColumn_37[10] , 
        \wColumn_37[9] , \wColumn_37[8] , \wColumn_37[7] , \wColumn_37[6] , 
        \wColumn_37[5] , \wColumn_37[4] , \wColumn_37[3] , \wColumn_37[2] , 
        \wColumn_37[1] , \wColumn_37[0] }), .PDiagOut({\wPDiag_37[63] , 
        \wPDiag_37[62] , \wPDiag_37[61] , \wPDiag_37[60] , \wPDiag_37[59] , 
        \wPDiag_37[58] , \wPDiag_37[57] , \wPDiag_37[56] , \wPDiag_37[55] , 
        \wPDiag_37[54] , \wPDiag_37[53] , \wPDiag_37[52] , \wPDiag_37[51] , 
        \wPDiag_37[50] , \wPDiag_37[49] , \wPDiag_37[48] , \wPDiag_37[47] , 
        \wPDiag_37[46] , \wPDiag_37[45] , \wPDiag_37[44] , \wPDiag_37[43] , 
        \wPDiag_37[42] , \wPDiag_37[41] , \wPDiag_37[40] , \wPDiag_37[39] , 
        \wPDiag_37[38] , \wPDiag_37[37] , \wPDiag_37[36] , \wPDiag_37[35] , 
        \wPDiag_37[34] , \wPDiag_37[33] , \wPDiag_37[32] , \wPDiag_37[31] , 
        \wPDiag_37[30] , \wPDiag_37[29] , \wPDiag_37[28] , \wPDiag_37[27] , 
        \wPDiag_37[26] , \wPDiag_37[25] , \wPDiag_37[24] , \wPDiag_37[23] , 
        \wPDiag_37[22] , \wPDiag_37[21] , \wPDiag_37[20] , \wPDiag_37[19] , 
        \wPDiag_37[18] , \wPDiag_37[17] , \wPDiag_37[16] , \wPDiag_37[15] , 
        \wPDiag_37[14] , \wPDiag_37[13] , \wPDiag_37[12] , \wPDiag_37[11] , 
        \wPDiag_37[10] , \wPDiag_37[9] , \wPDiag_37[8] , \wPDiag_37[7] , 
        \wPDiag_37[6] , \wPDiag_37[5] , \wPDiag_37[4] , \wPDiag_37[3] , 
        \wPDiag_37[2] , \wPDiag_37[1] , \wPDiag_37[0] }), .NDiagOut({
        \wNDiag_37[63] , \wNDiag_37[62] , \wNDiag_37[61] , \wNDiag_37[60] , 
        \wNDiag_37[59] , \wNDiag_37[58] , \wNDiag_37[57] , \wNDiag_37[56] , 
        \wNDiag_37[55] , \wNDiag_37[54] , \wNDiag_37[53] , \wNDiag_37[52] , 
        \wNDiag_37[51] , \wNDiag_37[50] , \wNDiag_37[49] , \wNDiag_37[48] , 
        \wNDiag_37[47] , \wNDiag_37[46] , \wNDiag_37[45] , \wNDiag_37[44] , 
        \wNDiag_37[43] , \wNDiag_37[42] , \wNDiag_37[41] , \wNDiag_37[40] , 
        \wNDiag_37[39] , \wNDiag_37[38] , \wNDiag_37[37] , \wNDiag_37[36] , 
        \wNDiag_37[35] , \wNDiag_37[34] , \wNDiag_37[33] , \wNDiag_37[32] , 
        \wNDiag_37[31] , \wNDiag_37[30] , \wNDiag_37[29] , \wNDiag_37[28] , 
        \wNDiag_37[27] , \wNDiag_37[26] , \wNDiag_37[25] , \wNDiag_37[24] , 
        \wNDiag_37[23] , \wNDiag_37[22] , \wNDiag_37[21] , \wNDiag_37[20] , 
        \wNDiag_37[19] , \wNDiag_37[18] , \wNDiag_37[17] , \wNDiag_37[16] , 
        \wNDiag_37[15] , \wNDiag_37[14] , \wNDiag_37[13] , \wNDiag_37[12] , 
        \wNDiag_37[11] , \wNDiag_37[10] , \wNDiag_37[9] , \wNDiag_37[8] , 
        \wNDiag_37[7] , \wNDiag_37[6] , \wNDiag_37[5] , \wNDiag_37[4] , 
        \wNDiag_37[3] , \wNDiag_37[2] , \wNDiag_37[1] , \wNDiag_37[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_1 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_2[6] , \wScan_2[5] , \wScan_2[4] , 
        \wScan_2[3] , \wScan_2[2] , \wScan_2[1] , \wScan_2[0] }), .ScanOut({
        \wScan_1[6] , \wScan_1[5] , \wScan_1[4] , \wScan_1[3] , \wScan_1[2] , 
        \wScan_1[1] , \wScan_1[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_1[0] ), 
        .ReturnIn(\wReturn_2[0] ), .ColIn({\wColumn_1[63] , \wColumn_1[62] , 
        \wColumn_1[61] , \wColumn_1[60] , \wColumn_1[59] , \wColumn_1[58] , 
        \wColumn_1[57] , \wColumn_1[56] , \wColumn_1[55] , \wColumn_1[54] , 
        \wColumn_1[53] , \wColumn_1[52] , \wColumn_1[51] , \wColumn_1[50] , 
        \wColumn_1[49] , \wColumn_1[48] , \wColumn_1[47] , \wColumn_1[46] , 
        \wColumn_1[45] , \wColumn_1[44] , \wColumn_1[43] , \wColumn_1[42] , 
        \wColumn_1[41] , \wColumn_1[40] , \wColumn_1[39] , \wColumn_1[38] , 
        \wColumn_1[37] , \wColumn_1[36] , \wColumn_1[35] , \wColumn_1[34] , 
        \wColumn_1[33] , \wColumn_1[32] , \wColumn_1[31] , \wColumn_1[30] , 
        \wColumn_1[29] , \wColumn_1[28] , \wColumn_1[27] , \wColumn_1[26] , 
        \wColumn_1[25] , \wColumn_1[24] , \wColumn_1[23] , \wColumn_1[22] , 
        \wColumn_1[21] , \wColumn_1[20] , \wColumn_1[19] , \wColumn_1[18] , 
        \wColumn_1[17] , \wColumn_1[16] , \wColumn_1[15] , \wColumn_1[14] , 
        \wColumn_1[13] , \wColumn_1[12] , \wColumn_1[11] , \wColumn_1[10] , 
        \wColumn_1[9] , \wColumn_1[8] , \wColumn_1[7] , \wColumn_1[6] , 
        \wColumn_1[5] , \wColumn_1[4] , \wColumn_1[3] , \wColumn_1[2] , 
        \wColumn_1[1] , \wColumn_1[0] }), .PDiagIn({\wPDiag_1[63] , 
        \wPDiag_1[62] , \wPDiag_1[61] , \wPDiag_1[60] , \wPDiag_1[59] , 
        \wPDiag_1[58] , \wPDiag_1[57] , \wPDiag_1[56] , \wPDiag_1[55] , 
        \wPDiag_1[54] , \wPDiag_1[53] , \wPDiag_1[52] , \wPDiag_1[51] , 
        \wPDiag_1[50] , \wPDiag_1[49] , \wPDiag_1[48] , \wPDiag_1[47] , 
        \wPDiag_1[46] , \wPDiag_1[45] , \wPDiag_1[44] , \wPDiag_1[43] , 
        \wPDiag_1[42] , \wPDiag_1[41] , \wPDiag_1[40] , \wPDiag_1[39] , 
        \wPDiag_1[38] , \wPDiag_1[37] , \wPDiag_1[36] , \wPDiag_1[35] , 
        \wPDiag_1[34] , \wPDiag_1[33] , \wPDiag_1[32] , \wPDiag_1[31] , 
        \wPDiag_1[30] , \wPDiag_1[29] , \wPDiag_1[28] , \wPDiag_1[27] , 
        \wPDiag_1[26] , \wPDiag_1[25] , \wPDiag_1[24] , \wPDiag_1[23] , 
        \wPDiag_1[22] , \wPDiag_1[21] , \wPDiag_1[20] , \wPDiag_1[19] , 
        \wPDiag_1[18] , \wPDiag_1[17] , \wPDiag_1[16] , \wPDiag_1[15] , 
        \wPDiag_1[14] , \wPDiag_1[13] , \wPDiag_1[12] , \wPDiag_1[11] , 
        \wPDiag_1[10] , \wPDiag_1[9] , \wPDiag_1[8] , \wPDiag_1[7] , 
        \wPDiag_1[6] , \wPDiag_1[5] , \wPDiag_1[4] , \wPDiag_1[3] , 
        \wPDiag_1[2] , \wPDiag_1[1] , \wPDiag_1[0] }), .NDiagIn({
        \wNDiag_1[63] , \wNDiag_1[62] , \wNDiag_1[61] , \wNDiag_1[60] , 
        \wNDiag_1[59] , \wNDiag_1[58] , \wNDiag_1[57] , \wNDiag_1[56] , 
        \wNDiag_1[55] , \wNDiag_1[54] , \wNDiag_1[53] , \wNDiag_1[52] , 
        \wNDiag_1[51] , \wNDiag_1[50] , \wNDiag_1[49] , \wNDiag_1[48] , 
        \wNDiag_1[47] , \wNDiag_1[46] , \wNDiag_1[45] , \wNDiag_1[44] , 
        \wNDiag_1[43] , \wNDiag_1[42] , \wNDiag_1[41] , \wNDiag_1[40] , 
        \wNDiag_1[39] , \wNDiag_1[38] , \wNDiag_1[37] , \wNDiag_1[36] , 
        \wNDiag_1[35] , \wNDiag_1[34] , \wNDiag_1[33] , \wNDiag_1[32] , 
        \wNDiag_1[31] , \wNDiag_1[30] , \wNDiag_1[29] , \wNDiag_1[28] , 
        \wNDiag_1[27] , \wNDiag_1[26] , \wNDiag_1[25] , \wNDiag_1[24] , 
        \wNDiag_1[23] , \wNDiag_1[22] , \wNDiag_1[21] , \wNDiag_1[20] , 
        \wNDiag_1[19] , \wNDiag_1[18] , \wNDiag_1[17] , \wNDiag_1[16] , 
        \wNDiag_1[15] , \wNDiag_1[14] , \wNDiag_1[13] , \wNDiag_1[12] , 
        \wNDiag_1[11] , \wNDiag_1[10] , \wNDiag_1[9] , \wNDiag_1[8] , 
        \wNDiag_1[7] , \wNDiag_1[6] , \wNDiag_1[5] , \wNDiag_1[4] , 
        \wNDiag_1[3] , \wNDiag_1[2] , \wNDiag_1[1] , \wNDiag_1[0] }), 
        .CallOut(\wCall_2[0] ), .ReturnOut(\wReturn_1[0] ), .ColOut({
        \wColumn_2[63] , \wColumn_2[62] , \wColumn_2[61] , \wColumn_2[60] , 
        \wColumn_2[59] , \wColumn_2[58] , \wColumn_2[57] , \wColumn_2[56] , 
        \wColumn_2[55] , \wColumn_2[54] , \wColumn_2[53] , \wColumn_2[52] , 
        \wColumn_2[51] , \wColumn_2[50] , \wColumn_2[49] , \wColumn_2[48] , 
        \wColumn_2[47] , \wColumn_2[46] , \wColumn_2[45] , \wColumn_2[44] , 
        \wColumn_2[43] , \wColumn_2[42] , \wColumn_2[41] , \wColumn_2[40] , 
        \wColumn_2[39] , \wColumn_2[38] , \wColumn_2[37] , \wColumn_2[36] , 
        \wColumn_2[35] , \wColumn_2[34] , \wColumn_2[33] , \wColumn_2[32] , 
        \wColumn_2[31] , \wColumn_2[30] , \wColumn_2[29] , \wColumn_2[28] , 
        \wColumn_2[27] , \wColumn_2[26] , \wColumn_2[25] , \wColumn_2[24] , 
        \wColumn_2[23] , \wColumn_2[22] , \wColumn_2[21] , \wColumn_2[20] , 
        \wColumn_2[19] , \wColumn_2[18] , \wColumn_2[17] , \wColumn_2[16] , 
        \wColumn_2[15] , \wColumn_2[14] , \wColumn_2[13] , \wColumn_2[12] , 
        \wColumn_2[11] , \wColumn_2[10] , \wColumn_2[9] , \wColumn_2[8] , 
        \wColumn_2[7] , \wColumn_2[6] , \wColumn_2[5] , \wColumn_2[4] , 
        \wColumn_2[3] , \wColumn_2[2] , \wColumn_2[1] , \wColumn_2[0] }), 
        .PDiagOut({\wPDiag_2[63] , \wPDiag_2[62] , \wPDiag_2[61] , 
        \wPDiag_2[60] , \wPDiag_2[59] , \wPDiag_2[58] , \wPDiag_2[57] , 
        \wPDiag_2[56] , \wPDiag_2[55] , \wPDiag_2[54] , \wPDiag_2[53] , 
        \wPDiag_2[52] , \wPDiag_2[51] , \wPDiag_2[50] , \wPDiag_2[49] , 
        \wPDiag_2[48] , \wPDiag_2[47] , \wPDiag_2[46] , \wPDiag_2[45] , 
        \wPDiag_2[44] , \wPDiag_2[43] , \wPDiag_2[42] , \wPDiag_2[41] , 
        \wPDiag_2[40] , \wPDiag_2[39] , \wPDiag_2[38] , \wPDiag_2[37] , 
        \wPDiag_2[36] , \wPDiag_2[35] , \wPDiag_2[34] , \wPDiag_2[33] , 
        \wPDiag_2[32] , \wPDiag_2[31] , \wPDiag_2[30] , \wPDiag_2[29] , 
        \wPDiag_2[28] , \wPDiag_2[27] , \wPDiag_2[26] , \wPDiag_2[25] , 
        \wPDiag_2[24] , \wPDiag_2[23] , \wPDiag_2[22] , \wPDiag_2[21] , 
        \wPDiag_2[20] , \wPDiag_2[19] , \wPDiag_2[18] , \wPDiag_2[17] , 
        \wPDiag_2[16] , \wPDiag_2[15] , \wPDiag_2[14] , \wPDiag_2[13] , 
        \wPDiag_2[12] , \wPDiag_2[11] , \wPDiag_2[10] , \wPDiag_2[9] , 
        \wPDiag_2[8] , \wPDiag_2[7] , \wPDiag_2[6] , \wPDiag_2[5] , 
        \wPDiag_2[4] , \wPDiag_2[3] , \wPDiag_2[2] , \wPDiag_2[1] , 
        \wPDiag_2[0] }), .NDiagOut({\wNDiag_2[63] , \wNDiag_2[62] , 
        \wNDiag_2[61] , \wNDiag_2[60] , \wNDiag_2[59] , \wNDiag_2[58] , 
        \wNDiag_2[57] , \wNDiag_2[56] , \wNDiag_2[55] , \wNDiag_2[54] , 
        \wNDiag_2[53] , \wNDiag_2[52] , \wNDiag_2[51] , \wNDiag_2[50] , 
        \wNDiag_2[49] , \wNDiag_2[48] , \wNDiag_2[47] , \wNDiag_2[46] , 
        \wNDiag_2[45] , \wNDiag_2[44] , \wNDiag_2[43] , \wNDiag_2[42] , 
        \wNDiag_2[41] , \wNDiag_2[40] , \wNDiag_2[39] , \wNDiag_2[38] , 
        \wNDiag_2[37] , \wNDiag_2[36] , \wNDiag_2[35] , \wNDiag_2[34] , 
        \wNDiag_2[33] , \wNDiag_2[32] , \wNDiag_2[31] , \wNDiag_2[30] , 
        \wNDiag_2[29] , \wNDiag_2[28] , \wNDiag_2[27] , \wNDiag_2[26] , 
        \wNDiag_2[25] , \wNDiag_2[24] , \wNDiag_2[23] , \wNDiag_2[22] , 
        \wNDiag_2[21] , \wNDiag_2[20] , \wNDiag_2[19] , \wNDiag_2[18] , 
        \wNDiag_2[17] , \wNDiag_2[16] , \wNDiag_2[15] , \wNDiag_2[14] , 
        \wNDiag_2[13] , \wNDiag_2[12] , \wNDiag_2[11] , \wNDiag_2[10] , 
        \wNDiag_2[9] , \wNDiag_2[8] , \wNDiag_2[7] , \wNDiag_2[6] , 
        \wNDiag_2[5] , \wNDiag_2[4] , \wNDiag_2[3] , \wNDiag_2[2] , 
        \wNDiag_2[1] , \wNDiag_2[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_6 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_7[6] , \wScan_7[5] , \wScan_7[4] , 
        \wScan_7[3] , \wScan_7[2] , \wScan_7[1] , \wScan_7[0] }), .ScanOut({
        \wScan_6[6] , \wScan_6[5] , \wScan_6[4] , \wScan_6[3] , \wScan_6[2] , 
        \wScan_6[1] , \wScan_6[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_6[0] ), 
        .ReturnIn(\wReturn_7[0] ), .ColIn({\wColumn_6[63] , \wColumn_6[62] , 
        \wColumn_6[61] , \wColumn_6[60] , \wColumn_6[59] , \wColumn_6[58] , 
        \wColumn_6[57] , \wColumn_6[56] , \wColumn_6[55] , \wColumn_6[54] , 
        \wColumn_6[53] , \wColumn_6[52] , \wColumn_6[51] , \wColumn_6[50] , 
        \wColumn_6[49] , \wColumn_6[48] , \wColumn_6[47] , \wColumn_6[46] , 
        \wColumn_6[45] , \wColumn_6[44] , \wColumn_6[43] , \wColumn_6[42] , 
        \wColumn_6[41] , \wColumn_6[40] , \wColumn_6[39] , \wColumn_6[38] , 
        \wColumn_6[37] , \wColumn_6[36] , \wColumn_6[35] , \wColumn_6[34] , 
        \wColumn_6[33] , \wColumn_6[32] , \wColumn_6[31] , \wColumn_6[30] , 
        \wColumn_6[29] , \wColumn_6[28] , \wColumn_6[27] , \wColumn_6[26] , 
        \wColumn_6[25] , \wColumn_6[24] , \wColumn_6[23] , \wColumn_6[22] , 
        \wColumn_6[21] , \wColumn_6[20] , \wColumn_6[19] , \wColumn_6[18] , 
        \wColumn_6[17] , \wColumn_6[16] , \wColumn_6[15] , \wColumn_6[14] , 
        \wColumn_6[13] , \wColumn_6[12] , \wColumn_6[11] , \wColumn_6[10] , 
        \wColumn_6[9] , \wColumn_6[8] , \wColumn_6[7] , \wColumn_6[6] , 
        \wColumn_6[5] , \wColumn_6[4] , \wColumn_6[3] , \wColumn_6[2] , 
        \wColumn_6[1] , \wColumn_6[0] }), .PDiagIn({\wPDiag_6[63] , 
        \wPDiag_6[62] , \wPDiag_6[61] , \wPDiag_6[60] , \wPDiag_6[59] , 
        \wPDiag_6[58] , \wPDiag_6[57] , \wPDiag_6[56] , \wPDiag_6[55] , 
        \wPDiag_6[54] , \wPDiag_6[53] , \wPDiag_6[52] , \wPDiag_6[51] , 
        \wPDiag_6[50] , \wPDiag_6[49] , \wPDiag_6[48] , \wPDiag_6[47] , 
        \wPDiag_6[46] , \wPDiag_6[45] , \wPDiag_6[44] , \wPDiag_6[43] , 
        \wPDiag_6[42] , \wPDiag_6[41] , \wPDiag_6[40] , \wPDiag_6[39] , 
        \wPDiag_6[38] , \wPDiag_6[37] , \wPDiag_6[36] , \wPDiag_6[35] , 
        \wPDiag_6[34] , \wPDiag_6[33] , \wPDiag_6[32] , \wPDiag_6[31] , 
        \wPDiag_6[30] , \wPDiag_6[29] , \wPDiag_6[28] , \wPDiag_6[27] , 
        \wPDiag_6[26] , \wPDiag_6[25] , \wPDiag_6[24] , \wPDiag_6[23] , 
        \wPDiag_6[22] , \wPDiag_6[21] , \wPDiag_6[20] , \wPDiag_6[19] , 
        \wPDiag_6[18] , \wPDiag_6[17] , \wPDiag_6[16] , \wPDiag_6[15] , 
        \wPDiag_6[14] , \wPDiag_6[13] , \wPDiag_6[12] , \wPDiag_6[11] , 
        \wPDiag_6[10] , \wPDiag_6[9] , \wPDiag_6[8] , \wPDiag_6[7] , 
        \wPDiag_6[6] , \wPDiag_6[5] , \wPDiag_6[4] , \wPDiag_6[3] , 
        \wPDiag_6[2] , \wPDiag_6[1] , \wPDiag_6[0] }), .NDiagIn({
        \wNDiag_6[63] , \wNDiag_6[62] , \wNDiag_6[61] , \wNDiag_6[60] , 
        \wNDiag_6[59] , \wNDiag_6[58] , \wNDiag_6[57] , \wNDiag_6[56] , 
        \wNDiag_6[55] , \wNDiag_6[54] , \wNDiag_6[53] , \wNDiag_6[52] , 
        \wNDiag_6[51] , \wNDiag_6[50] , \wNDiag_6[49] , \wNDiag_6[48] , 
        \wNDiag_6[47] , \wNDiag_6[46] , \wNDiag_6[45] , \wNDiag_6[44] , 
        \wNDiag_6[43] , \wNDiag_6[42] , \wNDiag_6[41] , \wNDiag_6[40] , 
        \wNDiag_6[39] , \wNDiag_6[38] , \wNDiag_6[37] , \wNDiag_6[36] , 
        \wNDiag_6[35] , \wNDiag_6[34] , \wNDiag_6[33] , \wNDiag_6[32] , 
        \wNDiag_6[31] , \wNDiag_6[30] , \wNDiag_6[29] , \wNDiag_6[28] , 
        \wNDiag_6[27] , \wNDiag_6[26] , \wNDiag_6[25] , \wNDiag_6[24] , 
        \wNDiag_6[23] , \wNDiag_6[22] , \wNDiag_6[21] , \wNDiag_6[20] , 
        \wNDiag_6[19] , \wNDiag_6[18] , \wNDiag_6[17] , \wNDiag_6[16] , 
        \wNDiag_6[15] , \wNDiag_6[14] , \wNDiag_6[13] , \wNDiag_6[12] , 
        \wNDiag_6[11] , \wNDiag_6[10] , \wNDiag_6[9] , \wNDiag_6[8] , 
        \wNDiag_6[7] , \wNDiag_6[6] , \wNDiag_6[5] , \wNDiag_6[4] , 
        \wNDiag_6[3] , \wNDiag_6[2] , \wNDiag_6[1] , \wNDiag_6[0] }), 
        .CallOut(\wCall_7[0] ), .ReturnOut(\wReturn_6[0] ), .ColOut({
        \wColumn_7[63] , \wColumn_7[62] , \wColumn_7[61] , \wColumn_7[60] , 
        \wColumn_7[59] , \wColumn_7[58] , \wColumn_7[57] , \wColumn_7[56] , 
        \wColumn_7[55] , \wColumn_7[54] , \wColumn_7[53] , \wColumn_7[52] , 
        \wColumn_7[51] , \wColumn_7[50] , \wColumn_7[49] , \wColumn_7[48] , 
        \wColumn_7[47] , \wColumn_7[46] , \wColumn_7[45] , \wColumn_7[44] , 
        \wColumn_7[43] , \wColumn_7[42] , \wColumn_7[41] , \wColumn_7[40] , 
        \wColumn_7[39] , \wColumn_7[38] , \wColumn_7[37] , \wColumn_7[36] , 
        \wColumn_7[35] , \wColumn_7[34] , \wColumn_7[33] , \wColumn_7[32] , 
        \wColumn_7[31] , \wColumn_7[30] , \wColumn_7[29] , \wColumn_7[28] , 
        \wColumn_7[27] , \wColumn_7[26] , \wColumn_7[25] , \wColumn_7[24] , 
        \wColumn_7[23] , \wColumn_7[22] , \wColumn_7[21] , \wColumn_7[20] , 
        \wColumn_7[19] , \wColumn_7[18] , \wColumn_7[17] , \wColumn_7[16] , 
        \wColumn_7[15] , \wColumn_7[14] , \wColumn_7[13] , \wColumn_7[12] , 
        \wColumn_7[11] , \wColumn_7[10] , \wColumn_7[9] , \wColumn_7[8] , 
        \wColumn_7[7] , \wColumn_7[6] , \wColumn_7[5] , \wColumn_7[4] , 
        \wColumn_7[3] , \wColumn_7[2] , \wColumn_7[1] , \wColumn_7[0] }), 
        .PDiagOut({\wPDiag_7[63] , \wPDiag_7[62] , \wPDiag_7[61] , 
        \wPDiag_7[60] , \wPDiag_7[59] , \wPDiag_7[58] , \wPDiag_7[57] , 
        \wPDiag_7[56] , \wPDiag_7[55] , \wPDiag_7[54] , \wPDiag_7[53] , 
        \wPDiag_7[52] , \wPDiag_7[51] , \wPDiag_7[50] , \wPDiag_7[49] , 
        \wPDiag_7[48] , \wPDiag_7[47] , \wPDiag_7[46] , \wPDiag_7[45] , 
        \wPDiag_7[44] , \wPDiag_7[43] , \wPDiag_7[42] , \wPDiag_7[41] , 
        \wPDiag_7[40] , \wPDiag_7[39] , \wPDiag_7[38] , \wPDiag_7[37] , 
        \wPDiag_7[36] , \wPDiag_7[35] , \wPDiag_7[34] , \wPDiag_7[33] , 
        \wPDiag_7[32] , \wPDiag_7[31] , \wPDiag_7[30] , \wPDiag_7[29] , 
        \wPDiag_7[28] , \wPDiag_7[27] , \wPDiag_7[26] , \wPDiag_7[25] , 
        \wPDiag_7[24] , \wPDiag_7[23] , \wPDiag_7[22] , \wPDiag_7[21] , 
        \wPDiag_7[20] , \wPDiag_7[19] , \wPDiag_7[18] , \wPDiag_7[17] , 
        \wPDiag_7[16] , \wPDiag_7[15] , \wPDiag_7[14] , \wPDiag_7[13] , 
        \wPDiag_7[12] , \wPDiag_7[11] , \wPDiag_7[10] , \wPDiag_7[9] , 
        \wPDiag_7[8] , \wPDiag_7[7] , \wPDiag_7[6] , \wPDiag_7[5] , 
        \wPDiag_7[4] , \wPDiag_7[3] , \wPDiag_7[2] , \wPDiag_7[1] , 
        \wPDiag_7[0] }), .NDiagOut({\wNDiag_7[63] , \wNDiag_7[62] , 
        \wNDiag_7[61] , \wNDiag_7[60] , \wNDiag_7[59] , \wNDiag_7[58] , 
        \wNDiag_7[57] , \wNDiag_7[56] , \wNDiag_7[55] , \wNDiag_7[54] , 
        \wNDiag_7[53] , \wNDiag_7[52] , \wNDiag_7[51] , \wNDiag_7[50] , 
        \wNDiag_7[49] , \wNDiag_7[48] , \wNDiag_7[47] , \wNDiag_7[46] , 
        \wNDiag_7[45] , \wNDiag_7[44] , \wNDiag_7[43] , \wNDiag_7[42] , 
        \wNDiag_7[41] , \wNDiag_7[40] , \wNDiag_7[39] , \wNDiag_7[38] , 
        \wNDiag_7[37] , \wNDiag_7[36] , \wNDiag_7[35] , \wNDiag_7[34] , 
        \wNDiag_7[33] , \wNDiag_7[32] , \wNDiag_7[31] , \wNDiag_7[30] , 
        \wNDiag_7[29] , \wNDiag_7[28] , \wNDiag_7[27] , \wNDiag_7[26] , 
        \wNDiag_7[25] , \wNDiag_7[24] , \wNDiag_7[23] , \wNDiag_7[22] , 
        \wNDiag_7[21] , \wNDiag_7[20] , \wNDiag_7[19] , \wNDiag_7[18] , 
        \wNDiag_7[17] , \wNDiag_7[16] , \wNDiag_7[15] , \wNDiag_7[14] , 
        \wNDiag_7[13] , \wNDiag_7[12] , \wNDiag_7[11] , \wNDiag_7[10] , 
        \wNDiag_7[9] , \wNDiag_7[8] , \wNDiag_7[7] , \wNDiag_7[6] , 
        \wNDiag_7[5] , \wNDiag_7[4] , \wNDiag_7[3] , \wNDiag_7[2] , 
        \wNDiag_7[1] , \wNDiag_7[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_7 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_8[6] , \wScan_8[5] , \wScan_8[4] , 
        \wScan_8[3] , \wScan_8[2] , \wScan_8[1] , \wScan_8[0] }), .ScanOut({
        \wScan_7[6] , \wScan_7[5] , \wScan_7[4] , \wScan_7[3] , \wScan_7[2] , 
        \wScan_7[1] , \wScan_7[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_7[0] ), 
        .ReturnIn(\wReturn_8[0] ), .ColIn({\wColumn_7[63] , \wColumn_7[62] , 
        \wColumn_7[61] , \wColumn_7[60] , \wColumn_7[59] , \wColumn_7[58] , 
        \wColumn_7[57] , \wColumn_7[56] , \wColumn_7[55] , \wColumn_7[54] , 
        \wColumn_7[53] , \wColumn_7[52] , \wColumn_7[51] , \wColumn_7[50] , 
        \wColumn_7[49] , \wColumn_7[48] , \wColumn_7[47] , \wColumn_7[46] , 
        \wColumn_7[45] , \wColumn_7[44] , \wColumn_7[43] , \wColumn_7[42] , 
        \wColumn_7[41] , \wColumn_7[40] , \wColumn_7[39] , \wColumn_7[38] , 
        \wColumn_7[37] , \wColumn_7[36] , \wColumn_7[35] , \wColumn_7[34] , 
        \wColumn_7[33] , \wColumn_7[32] , \wColumn_7[31] , \wColumn_7[30] , 
        \wColumn_7[29] , \wColumn_7[28] , \wColumn_7[27] , \wColumn_7[26] , 
        \wColumn_7[25] , \wColumn_7[24] , \wColumn_7[23] , \wColumn_7[22] , 
        \wColumn_7[21] , \wColumn_7[20] , \wColumn_7[19] , \wColumn_7[18] , 
        \wColumn_7[17] , \wColumn_7[16] , \wColumn_7[15] , \wColumn_7[14] , 
        \wColumn_7[13] , \wColumn_7[12] , \wColumn_7[11] , \wColumn_7[10] , 
        \wColumn_7[9] , \wColumn_7[8] , \wColumn_7[7] , \wColumn_7[6] , 
        \wColumn_7[5] , \wColumn_7[4] , \wColumn_7[3] , \wColumn_7[2] , 
        \wColumn_7[1] , \wColumn_7[0] }), .PDiagIn({\wPDiag_7[63] , 
        \wPDiag_7[62] , \wPDiag_7[61] , \wPDiag_7[60] , \wPDiag_7[59] , 
        \wPDiag_7[58] , \wPDiag_7[57] , \wPDiag_7[56] , \wPDiag_7[55] , 
        \wPDiag_7[54] , \wPDiag_7[53] , \wPDiag_7[52] , \wPDiag_7[51] , 
        \wPDiag_7[50] , \wPDiag_7[49] , \wPDiag_7[48] , \wPDiag_7[47] , 
        \wPDiag_7[46] , \wPDiag_7[45] , \wPDiag_7[44] , \wPDiag_7[43] , 
        \wPDiag_7[42] , \wPDiag_7[41] , \wPDiag_7[40] , \wPDiag_7[39] , 
        \wPDiag_7[38] , \wPDiag_7[37] , \wPDiag_7[36] , \wPDiag_7[35] , 
        \wPDiag_7[34] , \wPDiag_7[33] , \wPDiag_7[32] , \wPDiag_7[31] , 
        \wPDiag_7[30] , \wPDiag_7[29] , \wPDiag_7[28] , \wPDiag_7[27] , 
        \wPDiag_7[26] , \wPDiag_7[25] , \wPDiag_7[24] , \wPDiag_7[23] , 
        \wPDiag_7[22] , \wPDiag_7[21] , \wPDiag_7[20] , \wPDiag_7[19] , 
        \wPDiag_7[18] , \wPDiag_7[17] , \wPDiag_7[16] , \wPDiag_7[15] , 
        \wPDiag_7[14] , \wPDiag_7[13] , \wPDiag_7[12] , \wPDiag_7[11] , 
        \wPDiag_7[10] , \wPDiag_7[9] , \wPDiag_7[8] , \wPDiag_7[7] , 
        \wPDiag_7[6] , \wPDiag_7[5] , \wPDiag_7[4] , \wPDiag_7[3] , 
        \wPDiag_7[2] , \wPDiag_7[1] , \wPDiag_7[0] }), .NDiagIn({
        \wNDiag_7[63] , \wNDiag_7[62] , \wNDiag_7[61] , \wNDiag_7[60] , 
        \wNDiag_7[59] , \wNDiag_7[58] , \wNDiag_7[57] , \wNDiag_7[56] , 
        \wNDiag_7[55] , \wNDiag_7[54] , \wNDiag_7[53] , \wNDiag_7[52] , 
        \wNDiag_7[51] , \wNDiag_7[50] , \wNDiag_7[49] , \wNDiag_7[48] , 
        \wNDiag_7[47] , \wNDiag_7[46] , \wNDiag_7[45] , \wNDiag_7[44] , 
        \wNDiag_7[43] , \wNDiag_7[42] , \wNDiag_7[41] , \wNDiag_7[40] , 
        \wNDiag_7[39] , \wNDiag_7[38] , \wNDiag_7[37] , \wNDiag_7[36] , 
        \wNDiag_7[35] , \wNDiag_7[34] , \wNDiag_7[33] , \wNDiag_7[32] , 
        \wNDiag_7[31] , \wNDiag_7[30] , \wNDiag_7[29] , \wNDiag_7[28] , 
        \wNDiag_7[27] , \wNDiag_7[26] , \wNDiag_7[25] , \wNDiag_7[24] , 
        \wNDiag_7[23] , \wNDiag_7[22] , \wNDiag_7[21] , \wNDiag_7[20] , 
        \wNDiag_7[19] , \wNDiag_7[18] , \wNDiag_7[17] , \wNDiag_7[16] , 
        \wNDiag_7[15] , \wNDiag_7[14] , \wNDiag_7[13] , \wNDiag_7[12] , 
        \wNDiag_7[11] , \wNDiag_7[10] , \wNDiag_7[9] , \wNDiag_7[8] , 
        \wNDiag_7[7] , \wNDiag_7[6] , \wNDiag_7[5] , \wNDiag_7[4] , 
        \wNDiag_7[3] , \wNDiag_7[2] , \wNDiag_7[1] , \wNDiag_7[0] }), 
        .CallOut(\wCall_8[0] ), .ReturnOut(\wReturn_7[0] ), .ColOut({
        \wColumn_8[63] , \wColumn_8[62] , \wColumn_8[61] , \wColumn_8[60] , 
        \wColumn_8[59] , \wColumn_8[58] , \wColumn_8[57] , \wColumn_8[56] , 
        \wColumn_8[55] , \wColumn_8[54] , \wColumn_8[53] , \wColumn_8[52] , 
        \wColumn_8[51] , \wColumn_8[50] , \wColumn_8[49] , \wColumn_8[48] , 
        \wColumn_8[47] , \wColumn_8[46] , \wColumn_8[45] , \wColumn_8[44] , 
        \wColumn_8[43] , \wColumn_8[42] , \wColumn_8[41] , \wColumn_8[40] , 
        \wColumn_8[39] , \wColumn_8[38] , \wColumn_8[37] , \wColumn_8[36] , 
        \wColumn_8[35] , \wColumn_8[34] , \wColumn_8[33] , \wColumn_8[32] , 
        \wColumn_8[31] , \wColumn_8[30] , \wColumn_8[29] , \wColumn_8[28] , 
        \wColumn_8[27] , \wColumn_8[26] , \wColumn_8[25] , \wColumn_8[24] , 
        \wColumn_8[23] , \wColumn_8[22] , \wColumn_8[21] , \wColumn_8[20] , 
        \wColumn_8[19] , \wColumn_8[18] , \wColumn_8[17] , \wColumn_8[16] , 
        \wColumn_8[15] , \wColumn_8[14] , \wColumn_8[13] , \wColumn_8[12] , 
        \wColumn_8[11] , \wColumn_8[10] , \wColumn_8[9] , \wColumn_8[8] , 
        \wColumn_8[7] , \wColumn_8[6] , \wColumn_8[5] , \wColumn_8[4] , 
        \wColumn_8[3] , \wColumn_8[2] , \wColumn_8[1] , \wColumn_8[0] }), 
        .PDiagOut({\wPDiag_8[63] , \wPDiag_8[62] , \wPDiag_8[61] , 
        \wPDiag_8[60] , \wPDiag_8[59] , \wPDiag_8[58] , \wPDiag_8[57] , 
        \wPDiag_8[56] , \wPDiag_8[55] , \wPDiag_8[54] , \wPDiag_8[53] , 
        \wPDiag_8[52] , \wPDiag_8[51] , \wPDiag_8[50] , \wPDiag_8[49] , 
        \wPDiag_8[48] , \wPDiag_8[47] , \wPDiag_8[46] , \wPDiag_8[45] , 
        \wPDiag_8[44] , \wPDiag_8[43] , \wPDiag_8[42] , \wPDiag_8[41] , 
        \wPDiag_8[40] , \wPDiag_8[39] , \wPDiag_8[38] , \wPDiag_8[37] , 
        \wPDiag_8[36] , \wPDiag_8[35] , \wPDiag_8[34] , \wPDiag_8[33] , 
        \wPDiag_8[32] , \wPDiag_8[31] , \wPDiag_8[30] , \wPDiag_8[29] , 
        \wPDiag_8[28] , \wPDiag_8[27] , \wPDiag_8[26] , \wPDiag_8[25] , 
        \wPDiag_8[24] , \wPDiag_8[23] , \wPDiag_8[22] , \wPDiag_8[21] , 
        \wPDiag_8[20] , \wPDiag_8[19] , \wPDiag_8[18] , \wPDiag_8[17] , 
        \wPDiag_8[16] , \wPDiag_8[15] , \wPDiag_8[14] , \wPDiag_8[13] , 
        \wPDiag_8[12] , \wPDiag_8[11] , \wPDiag_8[10] , \wPDiag_8[9] , 
        \wPDiag_8[8] , \wPDiag_8[7] , \wPDiag_8[6] , \wPDiag_8[5] , 
        \wPDiag_8[4] , \wPDiag_8[3] , \wPDiag_8[2] , \wPDiag_8[1] , 
        \wPDiag_8[0] }), .NDiagOut({\wNDiag_8[63] , \wNDiag_8[62] , 
        \wNDiag_8[61] , \wNDiag_8[60] , \wNDiag_8[59] , \wNDiag_8[58] , 
        \wNDiag_8[57] , \wNDiag_8[56] , \wNDiag_8[55] , \wNDiag_8[54] , 
        \wNDiag_8[53] , \wNDiag_8[52] , \wNDiag_8[51] , \wNDiag_8[50] , 
        \wNDiag_8[49] , \wNDiag_8[48] , \wNDiag_8[47] , \wNDiag_8[46] , 
        \wNDiag_8[45] , \wNDiag_8[44] , \wNDiag_8[43] , \wNDiag_8[42] , 
        \wNDiag_8[41] , \wNDiag_8[40] , \wNDiag_8[39] , \wNDiag_8[38] , 
        \wNDiag_8[37] , \wNDiag_8[36] , \wNDiag_8[35] , \wNDiag_8[34] , 
        \wNDiag_8[33] , \wNDiag_8[32] , \wNDiag_8[31] , \wNDiag_8[30] , 
        \wNDiag_8[29] , \wNDiag_8[28] , \wNDiag_8[27] , \wNDiag_8[26] , 
        \wNDiag_8[25] , \wNDiag_8[24] , \wNDiag_8[23] , \wNDiag_8[22] , 
        \wNDiag_8[21] , \wNDiag_8[20] , \wNDiag_8[19] , \wNDiag_8[18] , 
        \wNDiag_8[17] , \wNDiag_8[16] , \wNDiag_8[15] , \wNDiag_8[14] , 
        \wNDiag_8[13] , \wNDiag_8[12] , \wNDiag_8[11] , \wNDiag_8[10] , 
        \wNDiag_8[9] , \wNDiag_8[8] , \wNDiag_8[7] , \wNDiag_8[6] , 
        \wNDiag_8[5] , \wNDiag_8[4] , \wNDiag_8[3] , \wNDiag_8[2] , 
        \wNDiag_8[1] , \wNDiag_8[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_18 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_19[6] , \wScan_19[5] , \wScan_19[4] , 
        \wScan_19[3] , \wScan_19[2] , \wScan_19[1] , \wScan_19[0] }), 
        .ScanOut({\wScan_18[6] , \wScan_18[5] , \wScan_18[4] , \wScan_18[3] , 
        \wScan_18[2] , \wScan_18[1] , \wScan_18[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_18[0] ), .ReturnIn(\wReturn_19[0] ), .ColIn({
        \wColumn_18[63] , \wColumn_18[62] , \wColumn_18[61] , \wColumn_18[60] , 
        \wColumn_18[59] , \wColumn_18[58] , \wColumn_18[57] , \wColumn_18[56] , 
        \wColumn_18[55] , \wColumn_18[54] , \wColumn_18[53] , \wColumn_18[52] , 
        \wColumn_18[51] , \wColumn_18[50] , \wColumn_18[49] , \wColumn_18[48] , 
        \wColumn_18[47] , \wColumn_18[46] , \wColumn_18[45] , \wColumn_18[44] , 
        \wColumn_18[43] , \wColumn_18[42] , \wColumn_18[41] , \wColumn_18[40] , 
        \wColumn_18[39] , \wColumn_18[38] , \wColumn_18[37] , \wColumn_18[36] , 
        \wColumn_18[35] , \wColumn_18[34] , \wColumn_18[33] , \wColumn_18[32] , 
        \wColumn_18[31] , \wColumn_18[30] , \wColumn_18[29] , \wColumn_18[28] , 
        \wColumn_18[27] , \wColumn_18[26] , \wColumn_18[25] , \wColumn_18[24] , 
        \wColumn_18[23] , \wColumn_18[22] , \wColumn_18[21] , \wColumn_18[20] , 
        \wColumn_18[19] , \wColumn_18[18] , \wColumn_18[17] , \wColumn_18[16] , 
        \wColumn_18[15] , \wColumn_18[14] , \wColumn_18[13] , \wColumn_18[12] , 
        \wColumn_18[11] , \wColumn_18[10] , \wColumn_18[9] , \wColumn_18[8] , 
        \wColumn_18[7] , \wColumn_18[6] , \wColumn_18[5] , \wColumn_18[4] , 
        \wColumn_18[3] , \wColumn_18[2] , \wColumn_18[1] , \wColumn_18[0] }), 
        .PDiagIn({\wPDiag_18[63] , \wPDiag_18[62] , \wPDiag_18[61] , 
        \wPDiag_18[60] , \wPDiag_18[59] , \wPDiag_18[58] , \wPDiag_18[57] , 
        \wPDiag_18[56] , \wPDiag_18[55] , \wPDiag_18[54] , \wPDiag_18[53] , 
        \wPDiag_18[52] , \wPDiag_18[51] , \wPDiag_18[50] , \wPDiag_18[49] , 
        \wPDiag_18[48] , \wPDiag_18[47] , \wPDiag_18[46] , \wPDiag_18[45] , 
        \wPDiag_18[44] , \wPDiag_18[43] , \wPDiag_18[42] , \wPDiag_18[41] , 
        \wPDiag_18[40] , \wPDiag_18[39] , \wPDiag_18[38] , \wPDiag_18[37] , 
        \wPDiag_18[36] , \wPDiag_18[35] , \wPDiag_18[34] , \wPDiag_18[33] , 
        \wPDiag_18[32] , \wPDiag_18[31] , \wPDiag_18[30] , \wPDiag_18[29] , 
        \wPDiag_18[28] , \wPDiag_18[27] , \wPDiag_18[26] , \wPDiag_18[25] , 
        \wPDiag_18[24] , \wPDiag_18[23] , \wPDiag_18[22] , \wPDiag_18[21] , 
        \wPDiag_18[20] , \wPDiag_18[19] , \wPDiag_18[18] , \wPDiag_18[17] , 
        \wPDiag_18[16] , \wPDiag_18[15] , \wPDiag_18[14] , \wPDiag_18[13] , 
        \wPDiag_18[12] , \wPDiag_18[11] , \wPDiag_18[10] , \wPDiag_18[9] , 
        \wPDiag_18[8] , \wPDiag_18[7] , \wPDiag_18[6] , \wPDiag_18[5] , 
        \wPDiag_18[4] , \wPDiag_18[3] , \wPDiag_18[2] , \wPDiag_18[1] , 
        \wPDiag_18[0] }), .NDiagIn({\wNDiag_18[63] , \wNDiag_18[62] , 
        \wNDiag_18[61] , \wNDiag_18[60] , \wNDiag_18[59] , \wNDiag_18[58] , 
        \wNDiag_18[57] , \wNDiag_18[56] , \wNDiag_18[55] , \wNDiag_18[54] , 
        \wNDiag_18[53] , \wNDiag_18[52] , \wNDiag_18[51] , \wNDiag_18[50] , 
        \wNDiag_18[49] , \wNDiag_18[48] , \wNDiag_18[47] , \wNDiag_18[46] , 
        \wNDiag_18[45] , \wNDiag_18[44] , \wNDiag_18[43] , \wNDiag_18[42] , 
        \wNDiag_18[41] , \wNDiag_18[40] , \wNDiag_18[39] , \wNDiag_18[38] , 
        \wNDiag_18[37] , \wNDiag_18[36] , \wNDiag_18[35] , \wNDiag_18[34] , 
        \wNDiag_18[33] , \wNDiag_18[32] , \wNDiag_18[31] , \wNDiag_18[30] , 
        \wNDiag_18[29] , \wNDiag_18[28] , \wNDiag_18[27] , \wNDiag_18[26] , 
        \wNDiag_18[25] , \wNDiag_18[24] , \wNDiag_18[23] , \wNDiag_18[22] , 
        \wNDiag_18[21] , \wNDiag_18[20] , \wNDiag_18[19] , \wNDiag_18[18] , 
        \wNDiag_18[17] , \wNDiag_18[16] , \wNDiag_18[15] , \wNDiag_18[14] , 
        \wNDiag_18[13] , \wNDiag_18[12] , \wNDiag_18[11] , \wNDiag_18[10] , 
        \wNDiag_18[9] , \wNDiag_18[8] , \wNDiag_18[7] , \wNDiag_18[6] , 
        \wNDiag_18[5] , \wNDiag_18[4] , \wNDiag_18[3] , \wNDiag_18[2] , 
        \wNDiag_18[1] , \wNDiag_18[0] }), .CallOut(\wCall_19[0] ), .ReturnOut(
        \wReturn_18[0] ), .ColOut({\wColumn_19[63] , \wColumn_19[62] , 
        \wColumn_19[61] , \wColumn_19[60] , \wColumn_19[59] , \wColumn_19[58] , 
        \wColumn_19[57] , \wColumn_19[56] , \wColumn_19[55] , \wColumn_19[54] , 
        \wColumn_19[53] , \wColumn_19[52] , \wColumn_19[51] , \wColumn_19[50] , 
        \wColumn_19[49] , \wColumn_19[48] , \wColumn_19[47] , \wColumn_19[46] , 
        \wColumn_19[45] , \wColumn_19[44] , \wColumn_19[43] , \wColumn_19[42] , 
        \wColumn_19[41] , \wColumn_19[40] , \wColumn_19[39] , \wColumn_19[38] , 
        \wColumn_19[37] , \wColumn_19[36] , \wColumn_19[35] , \wColumn_19[34] , 
        \wColumn_19[33] , \wColumn_19[32] , \wColumn_19[31] , \wColumn_19[30] , 
        \wColumn_19[29] , \wColumn_19[28] , \wColumn_19[27] , \wColumn_19[26] , 
        \wColumn_19[25] , \wColumn_19[24] , \wColumn_19[23] , \wColumn_19[22] , 
        \wColumn_19[21] , \wColumn_19[20] , \wColumn_19[19] , \wColumn_19[18] , 
        \wColumn_19[17] , \wColumn_19[16] , \wColumn_19[15] , \wColumn_19[14] , 
        \wColumn_19[13] , \wColumn_19[12] , \wColumn_19[11] , \wColumn_19[10] , 
        \wColumn_19[9] , \wColumn_19[8] , \wColumn_19[7] , \wColumn_19[6] , 
        \wColumn_19[5] , \wColumn_19[4] , \wColumn_19[3] , \wColumn_19[2] , 
        \wColumn_19[1] , \wColumn_19[0] }), .PDiagOut({\wPDiag_19[63] , 
        \wPDiag_19[62] , \wPDiag_19[61] , \wPDiag_19[60] , \wPDiag_19[59] , 
        \wPDiag_19[58] , \wPDiag_19[57] , \wPDiag_19[56] , \wPDiag_19[55] , 
        \wPDiag_19[54] , \wPDiag_19[53] , \wPDiag_19[52] , \wPDiag_19[51] , 
        \wPDiag_19[50] , \wPDiag_19[49] , \wPDiag_19[48] , \wPDiag_19[47] , 
        \wPDiag_19[46] , \wPDiag_19[45] , \wPDiag_19[44] , \wPDiag_19[43] , 
        \wPDiag_19[42] , \wPDiag_19[41] , \wPDiag_19[40] , \wPDiag_19[39] , 
        \wPDiag_19[38] , \wPDiag_19[37] , \wPDiag_19[36] , \wPDiag_19[35] , 
        \wPDiag_19[34] , \wPDiag_19[33] , \wPDiag_19[32] , \wPDiag_19[31] , 
        \wPDiag_19[30] , \wPDiag_19[29] , \wPDiag_19[28] , \wPDiag_19[27] , 
        \wPDiag_19[26] , \wPDiag_19[25] , \wPDiag_19[24] , \wPDiag_19[23] , 
        \wPDiag_19[22] , \wPDiag_19[21] , \wPDiag_19[20] , \wPDiag_19[19] , 
        \wPDiag_19[18] , \wPDiag_19[17] , \wPDiag_19[16] , \wPDiag_19[15] , 
        \wPDiag_19[14] , \wPDiag_19[13] , \wPDiag_19[12] , \wPDiag_19[11] , 
        \wPDiag_19[10] , \wPDiag_19[9] , \wPDiag_19[8] , \wPDiag_19[7] , 
        \wPDiag_19[6] , \wPDiag_19[5] , \wPDiag_19[4] , \wPDiag_19[3] , 
        \wPDiag_19[2] , \wPDiag_19[1] , \wPDiag_19[0] }), .NDiagOut({
        \wNDiag_19[63] , \wNDiag_19[62] , \wNDiag_19[61] , \wNDiag_19[60] , 
        \wNDiag_19[59] , \wNDiag_19[58] , \wNDiag_19[57] , \wNDiag_19[56] , 
        \wNDiag_19[55] , \wNDiag_19[54] , \wNDiag_19[53] , \wNDiag_19[52] , 
        \wNDiag_19[51] , \wNDiag_19[50] , \wNDiag_19[49] , \wNDiag_19[48] , 
        \wNDiag_19[47] , \wNDiag_19[46] , \wNDiag_19[45] , \wNDiag_19[44] , 
        \wNDiag_19[43] , \wNDiag_19[42] , \wNDiag_19[41] , \wNDiag_19[40] , 
        \wNDiag_19[39] , \wNDiag_19[38] , \wNDiag_19[37] , \wNDiag_19[36] , 
        \wNDiag_19[35] , \wNDiag_19[34] , \wNDiag_19[33] , \wNDiag_19[32] , 
        \wNDiag_19[31] , \wNDiag_19[30] , \wNDiag_19[29] , \wNDiag_19[28] , 
        \wNDiag_19[27] , \wNDiag_19[26] , \wNDiag_19[25] , \wNDiag_19[24] , 
        \wNDiag_19[23] , \wNDiag_19[22] , \wNDiag_19[21] , \wNDiag_19[20] , 
        \wNDiag_19[19] , \wNDiag_19[18] , \wNDiag_19[17] , \wNDiag_19[16] , 
        \wNDiag_19[15] , \wNDiag_19[14] , \wNDiag_19[13] , \wNDiag_19[12] , 
        \wNDiag_19[11] , \wNDiag_19[10] , \wNDiag_19[9] , \wNDiag_19[8] , 
        \wNDiag_19[7] , \wNDiag_19[6] , \wNDiag_19[5] , \wNDiag_19[4] , 
        \wNDiag_19[3] , \wNDiag_19[2] , \wNDiag_19[1] , \wNDiag_19[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_51 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_52[6] , \wScan_52[5] , \wScan_52[4] , 
        \wScan_52[3] , \wScan_52[2] , \wScan_52[1] , \wScan_52[0] }), 
        .ScanOut({\wScan_51[6] , \wScan_51[5] , \wScan_51[4] , \wScan_51[3] , 
        \wScan_51[2] , \wScan_51[1] , \wScan_51[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_51[0] ), .ReturnIn(\wReturn_52[0] ), .ColIn({
        \wColumn_51[63] , \wColumn_51[62] , \wColumn_51[61] , \wColumn_51[60] , 
        \wColumn_51[59] , \wColumn_51[58] , \wColumn_51[57] , \wColumn_51[56] , 
        \wColumn_51[55] , \wColumn_51[54] , \wColumn_51[53] , \wColumn_51[52] , 
        \wColumn_51[51] , \wColumn_51[50] , \wColumn_51[49] , \wColumn_51[48] , 
        \wColumn_51[47] , \wColumn_51[46] , \wColumn_51[45] , \wColumn_51[44] , 
        \wColumn_51[43] , \wColumn_51[42] , \wColumn_51[41] , \wColumn_51[40] , 
        \wColumn_51[39] , \wColumn_51[38] , \wColumn_51[37] , \wColumn_51[36] , 
        \wColumn_51[35] , \wColumn_51[34] , \wColumn_51[33] , \wColumn_51[32] , 
        \wColumn_51[31] , \wColumn_51[30] , \wColumn_51[29] , \wColumn_51[28] , 
        \wColumn_51[27] , \wColumn_51[26] , \wColumn_51[25] , \wColumn_51[24] , 
        \wColumn_51[23] , \wColumn_51[22] , \wColumn_51[21] , \wColumn_51[20] , 
        \wColumn_51[19] , \wColumn_51[18] , \wColumn_51[17] , \wColumn_51[16] , 
        \wColumn_51[15] , \wColumn_51[14] , \wColumn_51[13] , \wColumn_51[12] , 
        \wColumn_51[11] , \wColumn_51[10] , \wColumn_51[9] , \wColumn_51[8] , 
        \wColumn_51[7] , \wColumn_51[6] , \wColumn_51[5] , \wColumn_51[4] , 
        \wColumn_51[3] , \wColumn_51[2] , \wColumn_51[1] , \wColumn_51[0] }), 
        .PDiagIn({\wPDiag_51[63] , \wPDiag_51[62] , \wPDiag_51[61] , 
        \wPDiag_51[60] , \wPDiag_51[59] , \wPDiag_51[58] , \wPDiag_51[57] , 
        \wPDiag_51[56] , \wPDiag_51[55] , \wPDiag_51[54] , \wPDiag_51[53] , 
        \wPDiag_51[52] , \wPDiag_51[51] , \wPDiag_51[50] , \wPDiag_51[49] , 
        \wPDiag_51[48] , \wPDiag_51[47] , \wPDiag_51[46] , \wPDiag_51[45] , 
        \wPDiag_51[44] , \wPDiag_51[43] , \wPDiag_51[42] , \wPDiag_51[41] , 
        \wPDiag_51[40] , \wPDiag_51[39] , \wPDiag_51[38] , \wPDiag_51[37] , 
        \wPDiag_51[36] , \wPDiag_51[35] , \wPDiag_51[34] , \wPDiag_51[33] , 
        \wPDiag_51[32] , \wPDiag_51[31] , \wPDiag_51[30] , \wPDiag_51[29] , 
        \wPDiag_51[28] , \wPDiag_51[27] , \wPDiag_51[26] , \wPDiag_51[25] , 
        \wPDiag_51[24] , \wPDiag_51[23] , \wPDiag_51[22] , \wPDiag_51[21] , 
        \wPDiag_51[20] , \wPDiag_51[19] , \wPDiag_51[18] , \wPDiag_51[17] , 
        \wPDiag_51[16] , \wPDiag_51[15] , \wPDiag_51[14] , \wPDiag_51[13] , 
        \wPDiag_51[12] , \wPDiag_51[11] , \wPDiag_51[10] , \wPDiag_51[9] , 
        \wPDiag_51[8] , \wPDiag_51[7] , \wPDiag_51[6] , \wPDiag_51[5] , 
        \wPDiag_51[4] , \wPDiag_51[3] , \wPDiag_51[2] , \wPDiag_51[1] , 
        \wPDiag_51[0] }), .NDiagIn({\wNDiag_51[63] , \wNDiag_51[62] , 
        \wNDiag_51[61] , \wNDiag_51[60] , \wNDiag_51[59] , \wNDiag_51[58] , 
        \wNDiag_51[57] , \wNDiag_51[56] , \wNDiag_51[55] , \wNDiag_51[54] , 
        \wNDiag_51[53] , \wNDiag_51[52] , \wNDiag_51[51] , \wNDiag_51[50] , 
        \wNDiag_51[49] , \wNDiag_51[48] , \wNDiag_51[47] , \wNDiag_51[46] , 
        \wNDiag_51[45] , \wNDiag_51[44] , \wNDiag_51[43] , \wNDiag_51[42] , 
        \wNDiag_51[41] , \wNDiag_51[40] , \wNDiag_51[39] , \wNDiag_51[38] , 
        \wNDiag_51[37] , \wNDiag_51[36] , \wNDiag_51[35] , \wNDiag_51[34] , 
        \wNDiag_51[33] , \wNDiag_51[32] , \wNDiag_51[31] , \wNDiag_51[30] , 
        \wNDiag_51[29] , \wNDiag_51[28] , \wNDiag_51[27] , \wNDiag_51[26] , 
        \wNDiag_51[25] , \wNDiag_51[24] , \wNDiag_51[23] , \wNDiag_51[22] , 
        \wNDiag_51[21] , \wNDiag_51[20] , \wNDiag_51[19] , \wNDiag_51[18] , 
        \wNDiag_51[17] , \wNDiag_51[16] , \wNDiag_51[15] , \wNDiag_51[14] , 
        \wNDiag_51[13] , \wNDiag_51[12] , \wNDiag_51[11] , \wNDiag_51[10] , 
        \wNDiag_51[9] , \wNDiag_51[8] , \wNDiag_51[7] , \wNDiag_51[6] , 
        \wNDiag_51[5] , \wNDiag_51[4] , \wNDiag_51[3] , \wNDiag_51[2] , 
        \wNDiag_51[1] , \wNDiag_51[0] }), .CallOut(\wCall_52[0] ), .ReturnOut(
        \wReturn_51[0] ), .ColOut({\wColumn_52[63] , \wColumn_52[62] , 
        \wColumn_52[61] , \wColumn_52[60] , \wColumn_52[59] , \wColumn_52[58] , 
        \wColumn_52[57] , \wColumn_52[56] , \wColumn_52[55] , \wColumn_52[54] , 
        \wColumn_52[53] , \wColumn_52[52] , \wColumn_52[51] , \wColumn_52[50] , 
        \wColumn_52[49] , \wColumn_52[48] , \wColumn_52[47] , \wColumn_52[46] , 
        \wColumn_52[45] , \wColumn_52[44] , \wColumn_52[43] , \wColumn_52[42] , 
        \wColumn_52[41] , \wColumn_52[40] , \wColumn_52[39] , \wColumn_52[38] , 
        \wColumn_52[37] , \wColumn_52[36] , \wColumn_52[35] , \wColumn_52[34] , 
        \wColumn_52[33] , \wColumn_52[32] , \wColumn_52[31] , \wColumn_52[30] , 
        \wColumn_52[29] , \wColumn_52[28] , \wColumn_52[27] , \wColumn_52[26] , 
        \wColumn_52[25] , \wColumn_52[24] , \wColumn_52[23] , \wColumn_52[22] , 
        \wColumn_52[21] , \wColumn_52[20] , \wColumn_52[19] , \wColumn_52[18] , 
        \wColumn_52[17] , \wColumn_52[16] , \wColumn_52[15] , \wColumn_52[14] , 
        \wColumn_52[13] , \wColumn_52[12] , \wColumn_52[11] , \wColumn_52[10] , 
        \wColumn_52[9] , \wColumn_52[8] , \wColumn_52[7] , \wColumn_52[6] , 
        \wColumn_52[5] , \wColumn_52[4] , \wColumn_52[3] , \wColumn_52[2] , 
        \wColumn_52[1] , \wColumn_52[0] }), .PDiagOut({\wPDiag_52[63] , 
        \wPDiag_52[62] , \wPDiag_52[61] , \wPDiag_52[60] , \wPDiag_52[59] , 
        \wPDiag_52[58] , \wPDiag_52[57] , \wPDiag_52[56] , \wPDiag_52[55] , 
        \wPDiag_52[54] , \wPDiag_52[53] , \wPDiag_52[52] , \wPDiag_52[51] , 
        \wPDiag_52[50] , \wPDiag_52[49] , \wPDiag_52[48] , \wPDiag_52[47] , 
        \wPDiag_52[46] , \wPDiag_52[45] , \wPDiag_52[44] , \wPDiag_52[43] , 
        \wPDiag_52[42] , \wPDiag_52[41] , \wPDiag_52[40] , \wPDiag_52[39] , 
        \wPDiag_52[38] , \wPDiag_52[37] , \wPDiag_52[36] , \wPDiag_52[35] , 
        \wPDiag_52[34] , \wPDiag_52[33] , \wPDiag_52[32] , \wPDiag_52[31] , 
        \wPDiag_52[30] , \wPDiag_52[29] , \wPDiag_52[28] , \wPDiag_52[27] , 
        \wPDiag_52[26] , \wPDiag_52[25] , \wPDiag_52[24] , \wPDiag_52[23] , 
        \wPDiag_52[22] , \wPDiag_52[21] , \wPDiag_52[20] , \wPDiag_52[19] , 
        \wPDiag_52[18] , \wPDiag_52[17] , \wPDiag_52[16] , \wPDiag_52[15] , 
        \wPDiag_52[14] , \wPDiag_52[13] , \wPDiag_52[12] , \wPDiag_52[11] , 
        \wPDiag_52[10] , \wPDiag_52[9] , \wPDiag_52[8] , \wPDiag_52[7] , 
        \wPDiag_52[6] , \wPDiag_52[5] , \wPDiag_52[4] , \wPDiag_52[3] , 
        \wPDiag_52[2] , \wPDiag_52[1] , \wPDiag_52[0] }), .NDiagOut({
        \wNDiag_52[63] , \wNDiag_52[62] , \wNDiag_52[61] , \wNDiag_52[60] , 
        \wNDiag_52[59] , \wNDiag_52[58] , \wNDiag_52[57] , \wNDiag_52[56] , 
        \wNDiag_52[55] , \wNDiag_52[54] , \wNDiag_52[53] , \wNDiag_52[52] , 
        \wNDiag_52[51] , \wNDiag_52[50] , \wNDiag_52[49] , \wNDiag_52[48] , 
        \wNDiag_52[47] , \wNDiag_52[46] , \wNDiag_52[45] , \wNDiag_52[44] , 
        \wNDiag_52[43] , \wNDiag_52[42] , \wNDiag_52[41] , \wNDiag_52[40] , 
        \wNDiag_52[39] , \wNDiag_52[38] , \wNDiag_52[37] , \wNDiag_52[36] , 
        \wNDiag_52[35] , \wNDiag_52[34] , \wNDiag_52[33] , \wNDiag_52[32] , 
        \wNDiag_52[31] , \wNDiag_52[30] , \wNDiag_52[29] , \wNDiag_52[28] , 
        \wNDiag_52[27] , \wNDiag_52[26] , \wNDiag_52[25] , \wNDiag_52[24] , 
        \wNDiag_52[23] , \wNDiag_52[22] , \wNDiag_52[21] , \wNDiag_52[20] , 
        \wNDiag_52[19] , \wNDiag_52[18] , \wNDiag_52[17] , \wNDiag_52[16] , 
        \wNDiag_52[15] , \wNDiag_52[14] , \wNDiag_52[13] , \wNDiag_52[12] , 
        \wNDiag_52[11] , \wNDiag_52[10] , \wNDiag_52[9] , \wNDiag_52[8] , 
        \wNDiag_52[7] , \wNDiag_52[6] , \wNDiag_52[5] , \wNDiag_52[4] , 
        \wNDiag_52[3] , \wNDiag_52[2] , \wNDiag_52[1] , \wNDiag_52[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_38 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_39[6] , \wScan_39[5] , \wScan_39[4] , 
        \wScan_39[3] , \wScan_39[2] , \wScan_39[1] , \wScan_39[0] }), 
        .ScanOut({\wScan_38[6] , \wScan_38[5] , \wScan_38[4] , \wScan_38[3] , 
        \wScan_38[2] , \wScan_38[1] , \wScan_38[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_38[0] ), .ReturnIn(\wReturn_39[0] ), .ColIn({
        \wColumn_38[63] , \wColumn_38[62] , \wColumn_38[61] , \wColumn_38[60] , 
        \wColumn_38[59] , \wColumn_38[58] , \wColumn_38[57] , \wColumn_38[56] , 
        \wColumn_38[55] , \wColumn_38[54] , \wColumn_38[53] , \wColumn_38[52] , 
        \wColumn_38[51] , \wColumn_38[50] , \wColumn_38[49] , \wColumn_38[48] , 
        \wColumn_38[47] , \wColumn_38[46] , \wColumn_38[45] , \wColumn_38[44] , 
        \wColumn_38[43] , \wColumn_38[42] , \wColumn_38[41] , \wColumn_38[40] , 
        \wColumn_38[39] , \wColumn_38[38] , \wColumn_38[37] , \wColumn_38[36] , 
        \wColumn_38[35] , \wColumn_38[34] , \wColumn_38[33] , \wColumn_38[32] , 
        \wColumn_38[31] , \wColumn_38[30] , \wColumn_38[29] , \wColumn_38[28] , 
        \wColumn_38[27] , \wColumn_38[26] , \wColumn_38[25] , \wColumn_38[24] , 
        \wColumn_38[23] , \wColumn_38[22] , \wColumn_38[21] , \wColumn_38[20] , 
        \wColumn_38[19] , \wColumn_38[18] , \wColumn_38[17] , \wColumn_38[16] , 
        \wColumn_38[15] , \wColumn_38[14] , \wColumn_38[13] , \wColumn_38[12] , 
        \wColumn_38[11] , \wColumn_38[10] , \wColumn_38[9] , \wColumn_38[8] , 
        \wColumn_38[7] , \wColumn_38[6] , \wColumn_38[5] , \wColumn_38[4] , 
        \wColumn_38[3] , \wColumn_38[2] , \wColumn_38[1] , \wColumn_38[0] }), 
        .PDiagIn({\wPDiag_38[63] , \wPDiag_38[62] , \wPDiag_38[61] , 
        \wPDiag_38[60] , \wPDiag_38[59] , \wPDiag_38[58] , \wPDiag_38[57] , 
        \wPDiag_38[56] , \wPDiag_38[55] , \wPDiag_38[54] , \wPDiag_38[53] , 
        \wPDiag_38[52] , \wPDiag_38[51] , \wPDiag_38[50] , \wPDiag_38[49] , 
        \wPDiag_38[48] , \wPDiag_38[47] , \wPDiag_38[46] , \wPDiag_38[45] , 
        \wPDiag_38[44] , \wPDiag_38[43] , \wPDiag_38[42] , \wPDiag_38[41] , 
        \wPDiag_38[40] , \wPDiag_38[39] , \wPDiag_38[38] , \wPDiag_38[37] , 
        \wPDiag_38[36] , \wPDiag_38[35] , \wPDiag_38[34] , \wPDiag_38[33] , 
        \wPDiag_38[32] , \wPDiag_38[31] , \wPDiag_38[30] , \wPDiag_38[29] , 
        \wPDiag_38[28] , \wPDiag_38[27] , \wPDiag_38[26] , \wPDiag_38[25] , 
        \wPDiag_38[24] , \wPDiag_38[23] , \wPDiag_38[22] , \wPDiag_38[21] , 
        \wPDiag_38[20] , \wPDiag_38[19] , \wPDiag_38[18] , \wPDiag_38[17] , 
        \wPDiag_38[16] , \wPDiag_38[15] , \wPDiag_38[14] , \wPDiag_38[13] , 
        \wPDiag_38[12] , \wPDiag_38[11] , \wPDiag_38[10] , \wPDiag_38[9] , 
        \wPDiag_38[8] , \wPDiag_38[7] , \wPDiag_38[6] , \wPDiag_38[5] , 
        \wPDiag_38[4] , \wPDiag_38[3] , \wPDiag_38[2] , \wPDiag_38[1] , 
        \wPDiag_38[0] }), .NDiagIn({\wNDiag_38[63] , \wNDiag_38[62] , 
        \wNDiag_38[61] , \wNDiag_38[60] , \wNDiag_38[59] , \wNDiag_38[58] , 
        \wNDiag_38[57] , \wNDiag_38[56] , \wNDiag_38[55] , \wNDiag_38[54] , 
        \wNDiag_38[53] , \wNDiag_38[52] , \wNDiag_38[51] , \wNDiag_38[50] , 
        \wNDiag_38[49] , \wNDiag_38[48] , \wNDiag_38[47] , \wNDiag_38[46] , 
        \wNDiag_38[45] , \wNDiag_38[44] , \wNDiag_38[43] , \wNDiag_38[42] , 
        \wNDiag_38[41] , \wNDiag_38[40] , \wNDiag_38[39] , \wNDiag_38[38] , 
        \wNDiag_38[37] , \wNDiag_38[36] , \wNDiag_38[35] , \wNDiag_38[34] , 
        \wNDiag_38[33] , \wNDiag_38[32] , \wNDiag_38[31] , \wNDiag_38[30] , 
        \wNDiag_38[29] , \wNDiag_38[28] , \wNDiag_38[27] , \wNDiag_38[26] , 
        \wNDiag_38[25] , \wNDiag_38[24] , \wNDiag_38[23] , \wNDiag_38[22] , 
        \wNDiag_38[21] , \wNDiag_38[20] , \wNDiag_38[19] , \wNDiag_38[18] , 
        \wNDiag_38[17] , \wNDiag_38[16] , \wNDiag_38[15] , \wNDiag_38[14] , 
        \wNDiag_38[13] , \wNDiag_38[12] , \wNDiag_38[11] , \wNDiag_38[10] , 
        \wNDiag_38[9] , \wNDiag_38[8] , \wNDiag_38[7] , \wNDiag_38[6] , 
        \wNDiag_38[5] , \wNDiag_38[4] , \wNDiag_38[3] , \wNDiag_38[2] , 
        \wNDiag_38[1] , \wNDiag_38[0] }), .CallOut(\wCall_39[0] ), .ReturnOut(
        \wReturn_38[0] ), .ColOut({\wColumn_39[63] , \wColumn_39[62] , 
        \wColumn_39[61] , \wColumn_39[60] , \wColumn_39[59] , \wColumn_39[58] , 
        \wColumn_39[57] , \wColumn_39[56] , \wColumn_39[55] , \wColumn_39[54] , 
        \wColumn_39[53] , \wColumn_39[52] , \wColumn_39[51] , \wColumn_39[50] , 
        \wColumn_39[49] , \wColumn_39[48] , \wColumn_39[47] , \wColumn_39[46] , 
        \wColumn_39[45] , \wColumn_39[44] , \wColumn_39[43] , \wColumn_39[42] , 
        \wColumn_39[41] , \wColumn_39[40] , \wColumn_39[39] , \wColumn_39[38] , 
        \wColumn_39[37] , \wColumn_39[36] , \wColumn_39[35] , \wColumn_39[34] , 
        \wColumn_39[33] , \wColumn_39[32] , \wColumn_39[31] , \wColumn_39[30] , 
        \wColumn_39[29] , \wColumn_39[28] , \wColumn_39[27] , \wColumn_39[26] , 
        \wColumn_39[25] , \wColumn_39[24] , \wColumn_39[23] , \wColumn_39[22] , 
        \wColumn_39[21] , \wColumn_39[20] , \wColumn_39[19] , \wColumn_39[18] , 
        \wColumn_39[17] , \wColumn_39[16] , \wColumn_39[15] , \wColumn_39[14] , 
        \wColumn_39[13] , \wColumn_39[12] , \wColumn_39[11] , \wColumn_39[10] , 
        \wColumn_39[9] , \wColumn_39[8] , \wColumn_39[7] , \wColumn_39[6] , 
        \wColumn_39[5] , \wColumn_39[4] , \wColumn_39[3] , \wColumn_39[2] , 
        \wColumn_39[1] , \wColumn_39[0] }), .PDiagOut({\wPDiag_39[63] , 
        \wPDiag_39[62] , \wPDiag_39[61] , \wPDiag_39[60] , \wPDiag_39[59] , 
        \wPDiag_39[58] , \wPDiag_39[57] , \wPDiag_39[56] , \wPDiag_39[55] , 
        \wPDiag_39[54] , \wPDiag_39[53] , \wPDiag_39[52] , \wPDiag_39[51] , 
        \wPDiag_39[50] , \wPDiag_39[49] , \wPDiag_39[48] , \wPDiag_39[47] , 
        \wPDiag_39[46] , \wPDiag_39[45] , \wPDiag_39[44] , \wPDiag_39[43] , 
        \wPDiag_39[42] , \wPDiag_39[41] , \wPDiag_39[40] , \wPDiag_39[39] , 
        \wPDiag_39[38] , \wPDiag_39[37] , \wPDiag_39[36] , \wPDiag_39[35] , 
        \wPDiag_39[34] , \wPDiag_39[33] , \wPDiag_39[32] , \wPDiag_39[31] , 
        \wPDiag_39[30] , \wPDiag_39[29] , \wPDiag_39[28] , \wPDiag_39[27] , 
        \wPDiag_39[26] , \wPDiag_39[25] , \wPDiag_39[24] , \wPDiag_39[23] , 
        \wPDiag_39[22] , \wPDiag_39[21] , \wPDiag_39[20] , \wPDiag_39[19] , 
        \wPDiag_39[18] , \wPDiag_39[17] , \wPDiag_39[16] , \wPDiag_39[15] , 
        \wPDiag_39[14] , \wPDiag_39[13] , \wPDiag_39[12] , \wPDiag_39[11] , 
        \wPDiag_39[10] , \wPDiag_39[9] , \wPDiag_39[8] , \wPDiag_39[7] , 
        \wPDiag_39[6] , \wPDiag_39[5] , \wPDiag_39[4] , \wPDiag_39[3] , 
        \wPDiag_39[2] , \wPDiag_39[1] , \wPDiag_39[0] }), .NDiagOut({
        \wNDiag_39[63] , \wNDiag_39[62] , \wNDiag_39[61] , \wNDiag_39[60] , 
        \wNDiag_39[59] , \wNDiag_39[58] , \wNDiag_39[57] , \wNDiag_39[56] , 
        \wNDiag_39[55] , \wNDiag_39[54] , \wNDiag_39[53] , \wNDiag_39[52] , 
        \wNDiag_39[51] , \wNDiag_39[50] , \wNDiag_39[49] , \wNDiag_39[48] , 
        \wNDiag_39[47] , \wNDiag_39[46] , \wNDiag_39[45] , \wNDiag_39[44] , 
        \wNDiag_39[43] , \wNDiag_39[42] , \wNDiag_39[41] , \wNDiag_39[40] , 
        \wNDiag_39[39] , \wNDiag_39[38] , \wNDiag_39[37] , \wNDiag_39[36] , 
        \wNDiag_39[35] , \wNDiag_39[34] , \wNDiag_39[33] , \wNDiag_39[32] , 
        \wNDiag_39[31] , \wNDiag_39[30] , \wNDiag_39[29] , \wNDiag_39[28] , 
        \wNDiag_39[27] , \wNDiag_39[26] , \wNDiag_39[25] , \wNDiag_39[24] , 
        \wNDiag_39[23] , \wNDiag_39[22] , \wNDiag_39[21] , \wNDiag_39[20] , 
        \wNDiag_39[19] , \wNDiag_39[18] , \wNDiag_39[17] , \wNDiag_39[16] , 
        \wNDiag_39[15] , \wNDiag_39[14] , \wNDiag_39[13] , \wNDiag_39[12] , 
        \wNDiag_39[11] , \wNDiag_39[10] , \wNDiag_39[9] , \wNDiag_39[8] , 
        \wNDiag_39[7] , \wNDiag_39[6] , \wNDiag_39[5] , \wNDiag_39[4] , 
        \wNDiag_39[3] , \wNDiag_39[2] , \wNDiag_39[1] , \wNDiag_39[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_56 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_57[6] , \wScan_57[5] , \wScan_57[4] , 
        \wScan_57[3] , \wScan_57[2] , \wScan_57[1] , \wScan_57[0] }), 
        .ScanOut({\wScan_56[6] , \wScan_56[5] , \wScan_56[4] , \wScan_56[3] , 
        \wScan_56[2] , \wScan_56[1] , \wScan_56[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_56[0] ), .ReturnIn(\wReturn_57[0] ), .ColIn({
        \wColumn_56[63] , \wColumn_56[62] , \wColumn_56[61] , \wColumn_56[60] , 
        \wColumn_56[59] , \wColumn_56[58] , \wColumn_56[57] , \wColumn_56[56] , 
        \wColumn_56[55] , \wColumn_56[54] , \wColumn_56[53] , \wColumn_56[52] , 
        \wColumn_56[51] , \wColumn_56[50] , \wColumn_56[49] , \wColumn_56[48] , 
        \wColumn_56[47] , \wColumn_56[46] , \wColumn_56[45] , \wColumn_56[44] , 
        \wColumn_56[43] , \wColumn_56[42] , \wColumn_56[41] , \wColumn_56[40] , 
        \wColumn_56[39] , \wColumn_56[38] , \wColumn_56[37] , \wColumn_56[36] , 
        \wColumn_56[35] , \wColumn_56[34] , \wColumn_56[33] , \wColumn_56[32] , 
        \wColumn_56[31] , \wColumn_56[30] , \wColumn_56[29] , \wColumn_56[28] , 
        \wColumn_56[27] , \wColumn_56[26] , \wColumn_56[25] , \wColumn_56[24] , 
        \wColumn_56[23] , \wColumn_56[22] , \wColumn_56[21] , \wColumn_56[20] , 
        \wColumn_56[19] , \wColumn_56[18] , \wColumn_56[17] , \wColumn_56[16] , 
        \wColumn_56[15] , \wColumn_56[14] , \wColumn_56[13] , \wColumn_56[12] , 
        \wColumn_56[11] , \wColumn_56[10] , \wColumn_56[9] , \wColumn_56[8] , 
        \wColumn_56[7] , \wColumn_56[6] , \wColumn_56[5] , \wColumn_56[4] , 
        \wColumn_56[3] , \wColumn_56[2] , \wColumn_56[1] , \wColumn_56[0] }), 
        .PDiagIn({\wPDiag_56[63] , \wPDiag_56[62] , \wPDiag_56[61] , 
        \wPDiag_56[60] , \wPDiag_56[59] , \wPDiag_56[58] , \wPDiag_56[57] , 
        \wPDiag_56[56] , \wPDiag_56[55] , \wPDiag_56[54] , \wPDiag_56[53] , 
        \wPDiag_56[52] , \wPDiag_56[51] , \wPDiag_56[50] , \wPDiag_56[49] , 
        \wPDiag_56[48] , \wPDiag_56[47] , \wPDiag_56[46] , \wPDiag_56[45] , 
        \wPDiag_56[44] , \wPDiag_56[43] , \wPDiag_56[42] , \wPDiag_56[41] , 
        \wPDiag_56[40] , \wPDiag_56[39] , \wPDiag_56[38] , \wPDiag_56[37] , 
        \wPDiag_56[36] , \wPDiag_56[35] , \wPDiag_56[34] , \wPDiag_56[33] , 
        \wPDiag_56[32] , \wPDiag_56[31] , \wPDiag_56[30] , \wPDiag_56[29] , 
        \wPDiag_56[28] , \wPDiag_56[27] , \wPDiag_56[26] , \wPDiag_56[25] , 
        \wPDiag_56[24] , \wPDiag_56[23] , \wPDiag_56[22] , \wPDiag_56[21] , 
        \wPDiag_56[20] , \wPDiag_56[19] , \wPDiag_56[18] , \wPDiag_56[17] , 
        \wPDiag_56[16] , \wPDiag_56[15] , \wPDiag_56[14] , \wPDiag_56[13] , 
        \wPDiag_56[12] , \wPDiag_56[11] , \wPDiag_56[10] , \wPDiag_56[9] , 
        \wPDiag_56[8] , \wPDiag_56[7] , \wPDiag_56[6] , \wPDiag_56[5] , 
        \wPDiag_56[4] , \wPDiag_56[3] , \wPDiag_56[2] , \wPDiag_56[1] , 
        \wPDiag_56[0] }), .NDiagIn({\wNDiag_56[63] , \wNDiag_56[62] , 
        \wNDiag_56[61] , \wNDiag_56[60] , \wNDiag_56[59] , \wNDiag_56[58] , 
        \wNDiag_56[57] , \wNDiag_56[56] , \wNDiag_56[55] , \wNDiag_56[54] , 
        \wNDiag_56[53] , \wNDiag_56[52] , \wNDiag_56[51] , \wNDiag_56[50] , 
        \wNDiag_56[49] , \wNDiag_56[48] , \wNDiag_56[47] , \wNDiag_56[46] , 
        \wNDiag_56[45] , \wNDiag_56[44] , \wNDiag_56[43] , \wNDiag_56[42] , 
        \wNDiag_56[41] , \wNDiag_56[40] , \wNDiag_56[39] , \wNDiag_56[38] , 
        \wNDiag_56[37] , \wNDiag_56[36] , \wNDiag_56[35] , \wNDiag_56[34] , 
        \wNDiag_56[33] , \wNDiag_56[32] , \wNDiag_56[31] , \wNDiag_56[30] , 
        \wNDiag_56[29] , \wNDiag_56[28] , \wNDiag_56[27] , \wNDiag_56[26] , 
        \wNDiag_56[25] , \wNDiag_56[24] , \wNDiag_56[23] , \wNDiag_56[22] , 
        \wNDiag_56[21] , \wNDiag_56[20] , \wNDiag_56[19] , \wNDiag_56[18] , 
        \wNDiag_56[17] , \wNDiag_56[16] , \wNDiag_56[15] , \wNDiag_56[14] , 
        \wNDiag_56[13] , \wNDiag_56[12] , \wNDiag_56[11] , \wNDiag_56[10] , 
        \wNDiag_56[9] , \wNDiag_56[8] , \wNDiag_56[7] , \wNDiag_56[6] , 
        \wNDiag_56[5] , \wNDiag_56[4] , \wNDiag_56[3] , \wNDiag_56[2] , 
        \wNDiag_56[1] , \wNDiag_56[0] }), .CallOut(\wCall_57[0] ), .ReturnOut(
        \wReturn_56[0] ), .ColOut({\wColumn_57[63] , \wColumn_57[62] , 
        \wColumn_57[61] , \wColumn_57[60] , \wColumn_57[59] , \wColumn_57[58] , 
        \wColumn_57[57] , \wColumn_57[56] , \wColumn_57[55] , \wColumn_57[54] , 
        \wColumn_57[53] , \wColumn_57[52] , \wColumn_57[51] , \wColumn_57[50] , 
        \wColumn_57[49] , \wColumn_57[48] , \wColumn_57[47] , \wColumn_57[46] , 
        \wColumn_57[45] , \wColumn_57[44] , \wColumn_57[43] , \wColumn_57[42] , 
        \wColumn_57[41] , \wColumn_57[40] , \wColumn_57[39] , \wColumn_57[38] , 
        \wColumn_57[37] , \wColumn_57[36] , \wColumn_57[35] , \wColumn_57[34] , 
        \wColumn_57[33] , \wColumn_57[32] , \wColumn_57[31] , \wColumn_57[30] , 
        \wColumn_57[29] , \wColumn_57[28] , \wColumn_57[27] , \wColumn_57[26] , 
        \wColumn_57[25] , \wColumn_57[24] , \wColumn_57[23] , \wColumn_57[22] , 
        \wColumn_57[21] , \wColumn_57[20] , \wColumn_57[19] , \wColumn_57[18] , 
        \wColumn_57[17] , \wColumn_57[16] , \wColumn_57[15] , \wColumn_57[14] , 
        \wColumn_57[13] , \wColumn_57[12] , \wColumn_57[11] , \wColumn_57[10] , 
        \wColumn_57[9] , \wColumn_57[8] , \wColumn_57[7] , \wColumn_57[6] , 
        \wColumn_57[5] , \wColumn_57[4] , \wColumn_57[3] , \wColumn_57[2] , 
        \wColumn_57[1] , \wColumn_57[0] }), .PDiagOut({\wPDiag_57[63] , 
        \wPDiag_57[62] , \wPDiag_57[61] , \wPDiag_57[60] , \wPDiag_57[59] , 
        \wPDiag_57[58] , \wPDiag_57[57] , \wPDiag_57[56] , \wPDiag_57[55] , 
        \wPDiag_57[54] , \wPDiag_57[53] , \wPDiag_57[52] , \wPDiag_57[51] , 
        \wPDiag_57[50] , \wPDiag_57[49] , \wPDiag_57[48] , \wPDiag_57[47] , 
        \wPDiag_57[46] , \wPDiag_57[45] , \wPDiag_57[44] , \wPDiag_57[43] , 
        \wPDiag_57[42] , \wPDiag_57[41] , \wPDiag_57[40] , \wPDiag_57[39] , 
        \wPDiag_57[38] , \wPDiag_57[37] , \wPDiag_57[36] , \wPDiag_57[35] , 
        \wPDiag_57[34] , \wPDiag_57[33] , \wPDiag_57[32] , \wPDiag_57[31] , 
        \wPDiag_57[30] , \wPDiag_57[29] , \wPDiag_57[28] , \wPDiag_57[27] , 
        \wPDiag_57[26] , \wPDiag_57[25] , \wPDiag_57[24] , \wPDiag_57[23] , 
        \wPDiag_57[22] , \wPDiag_57[21] , \wPDiag_57[20] , \wPDiag_57[19] , 
        \wPDiag_57[18] , \wPDiag_57[17] , \wPDiag_57[16] , \wPDiag_57[15] , 
        \wPDiag_57[14] , \wPDiag_57[13] , \wPDiag_57[12] , \wPDiag_57[11] , 
        \wPDiag_57[10] , \wPDiag_57[9] , \wPDiag_57[8] , \wPDiag_57[7] , 
        \wPDiag_57[6] , \wPDiag_57[5] , \wPDiag_57[4] , \wPDiag_57[3] , 
        \wPDiag_57[2] , \wPDiag_57[1] , \wPDiag_57[0] }), .NDiagOut({
        \wNDiag_57[63] , \wNDiag_57[62] , \wNDiag_57[61] , \wNDiag_57[60] , 
        \wNDiag_57[59] , \wNDiag_57[58] , \wNDiag_57[57] , \wNDiag_57[56] , 
        \wNDiag_57[55] , \wNDiag_57[54] , \wNDiag_57[53] , \wNDiag_57[52] , 
        \wNDiag_57[51] , \wNDiag_57[50] , \wNDiag_57[49] , \wNDiag_57[48] , 
        \wNDiag_57[47] , \wNDiag_57[46] , \wNDiag_57[45] , \wNDiag_57[44] , 
        \wNDiag_57[43] , \wNDiag_57[42] , \wNDiag_57[41] , \wNDiag_57[40] , 
        \wNDiag_57[39] , \wNDiag_57[38] , \wNDiag_57[37] , \wNDiag_57[36] , 
        \wNDiag_57[35] , \wNDiag_57[34] , \wNDiag_57[33] , \wNDiag_57[32] , 
        \wNDiag_57[31] , \wNDiag_57[30] , \wNDiag_57[29] , \wNDiag_57[28] , 
        \wNDiag_57[27] , \wNDiag_57[26] , \wNDiag_57[25] , \wNDiag_57[24] , 
        \wNDiag_57[23] , \wNDiag_57[22] , \wNDiag_57[21] , \wNDiag_57[20] , 
        \wNDiag_57[19] , \wNDiag_57[18] , \wNDiag_57[17] , \wNDiag_57[16] , 
        \wNDiag_57[15] , \wNDiag_57[14] , \wNDiag_57[13] , \wNDiag_57[12] , 
        \wNDiag_57[11] , \wNDiag_57[10] , \wNDiag_57[9] , \wNDiag_57[8] , 
        \wNDiag_57[7] , \wNDiag_57[6] , \wNDiag_57[5] , \wNDiag_57[4] , 
        \wNDiag_57[3] , \wNDiag_57[2] , \wNDiag_57[1] , \wNDiag_57[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_16 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_17[6] , \wScan_17[5] , \wScan_17[4] , 
        \wScan_17[3] , \wScan_17[2] , \wScan_17[1] , \wScan_17[0] }), 
        .ScanOut({\wScan_16[6] , \wScan_16[5] , \wScan_16[4] , \wScan_16[3] , 
        \wScan_16[2] , \wScan_16[1] , \wScan_16[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_16[0] ), .ReturnIn(\wReturn_17[0] ), .ColIn({
        \wColumn_16[63] , \wColumn_16[62] , \wColumn_16[61] , \wColumn_16[60] , 
        \wColumn_16[59] , \wColumn_16[58] , \wColumn_16[57] , \wColumn_16[56] , 
        \wColumn_16[55] , \wColumn_16[54] , \wColumn_16[53] , \wColumn_16[52] , 
        \wColumn_16[51] , \wColumn_16[50] , \wColumn_16[49] , \wColumn_16[48] , 
        \wColumn_16[47] , \wColumn_16[46] , \wColumn_16[45] , \wColumn_16[44] , 
        \wColumn_16[43] , \wColumn_16[42] , \wColumn_16[41] , \wColumn_16[40] , 
        \wColumn_16[39] , \wColumn_16[38] , \wColumn_16[37] , \wColumn_16[36] , 
        \wColumn_16[35] , \wColumn_16[34] , \wColumn_16[33] , \wColumn_16[32] , 
        \wColumn_16[31] , \wColumn_16[30] , \wColumn_16[29] , \wColumn_16[28] , 
        \wColumn_16[27] , \wColumn_16[26] , \wColumn_16[25] , \wColumn_16[24] , 
        \wColumn_16[23] , \wColumn_16[22] , \wColumn_16[21] , \wColumn_16[20] , 
        \wColumn_16[19] , \wColumn_16[18] , \wColumn_16[17] , \wColumn_16[16] , 
        \wColumn_16[15] , \wColumn_16[14] , \wColumn_16[13] , \wColumn_16[12] , 
        \wColumn_16[11] , \wColumn_16[10] , \wColumn_16[9] , \wColumn_16[8] , 
        \wColumn_16[7] , \wColumn_16[6] , \wColumn_16[5] , \wColumn_16[4] , 
        \wColumn_16[3] , \wColumn_16[2] , \wColumn_16[1] , \wColumn_16[0] }), 
        .PDiagIn({\wPDiag_16[63] , \wPDiag_16[62] , \wPDiag_16[61] , 
        \wPDiag_16[60] , \wPDiag_16[59] , \wPDiag_16[58] , \wPDiag_16[57] , 
        \wPDiag_16[56] , \wPDiag_16[55] , \wPDiag_16[54] , \wPDiag_16[53] , 
        \wPDiag_16[52] , \wPDiag_16[51] , \wPDiag_16[50] , \wPDiag_16[49] , 
        \wPDiag_16[48] , \wPDiag_16[47] , \wPDiag_16[46] , \wPDiag_16[45] , 
        \wPDiag_16[44] , \wPDiag_16[43] , \wPDiag_16[42] , \wPDiag_16[41] , 
        \wPDiag_16[40] , \wPDiag_16[39] , \wPDiag_16[38] , \wPDiag_16[37] , 
        \wPDiag_16[36] , \wPDiag_16[35] , \wPDiag_16[34] , \wPDiag_16[33] , 
        \wPDiag_16[32] , \wPDiag_16[31] , \wPDiag_16[30] , \wPDiag_16[29] , 
        \wPDiag_16[28] , \wPDiag_16[27] , \wPDiag_16[26] , \wPDiag_16[25] , 
        \wPDiag_16[24] , \wPDiag_16[23] , \wPDiag_16[22] , \wPDiag_16[21] , 
        \wPDiag_16[20] , \wPDiag_16[19] , \wPDiag_16[18] , \wPDiag_16[17] , 
        \wPDiag_16[16] , \wPDiag_16[15] , \wPDiag_16[14] , \wPDiag_16[13] , 
        \wPDiag_16[12] , \wPDiag_16[11] , \wPDiag_16[10] , \wPDiag_16[9] , 
        \wPDiag_16[8] , \wPDiag_16[7] , \wPDiag_16[6] , \wPDiag_16[5] , 
        \wPDiag_16[4] , \wPDiag_16[3] , \wPDiag_16[2] , \wPDiag_16[1] , 
        \wPDiag_16[0] }), .NDiagIn({\wNDiag_16[63] , \wNDiag_16[62] , 
        \wNDiag_16[61] , \wNDiag_16[60] , \wNDiag_16[59] , \wNDiag_16[58] , 
        \wNDiag_16[57] , \wNDiag_16[56] , \wNDiag_16[55] , \wNDiag_16[54] , 
        \wNDiag_16[53] , \wNDiag_16[52] , \wNDiag_16[51] , \wNDiag_16[50] , 
        \wNDiag_16[49] , \wNDiag_16[48] , \wNDiag_16[47] , \wNDiag_16[46] , 
        \wNDiag_16[45] , \wNDiag_16[44] , \wNDiag_16[43] , \wNDiag_16[42] , 
        \wNDiag_16[41] , \wNDiag_16[40] , \wNDiag_16[39] , \wNDiag_16[38] , 
        \wNDiag_16[37] , \wNDiag_16[36] , \wNDiag_16[35] , \wNDiag_16[34] , 
        \wNDiag_16[33] , \wNDiag_16[32] , \wNDiag_16[31] , \wNDiag_16[30] , 
        \wNDiag_16[29] , \wNDiag_16[28] , \wNDiag_16[27] , \wNDiag_16[26] , 
        \wNDiag_16[25] , \wNDiag_16[24] , \wNDiag_16[23] , \wNDiag_16[22] , 
        \wNDiag_16[21] , \wNDiag_16[20] , \wNDiag_16[19] , \wNDiag_16[18] , 
        \wNDiag_16[17] , \wNDiag_16[16] , \wNDiag_16[15] , \wNDiag_16[14] , 
        \wNDiag_16[13] , \wNDiag_16[12] , \wNDiag_16[11] , \wNDiag_16[10] , 
        \wNDiag_16[9] , \wNDiag_16[8] , \wNDiag_16[7] , \wNDiag_16[6] , 
        \wNDiag_16[5] , \wNDiag_16[4] , \wNDiag_16[3] , \wNDiag_16[2] , 
        \wNDiag_16[1] , \wNDiag_16[0] }), .CallOut(\wCall_17[0] ), .ReturnOut(
        \wReturn_16[0] ), .ColOut({\wColumn_17[63] , \wColumn_17[62] , 
        \wColumn_17[61] , \wColumn_17[60] , \wColumn_17[59] , \wColumn_17[58] , 
        \wColumn_17[57] , \wColumn_17[56] , \wColumn_17[55] , \wColumn_17[54] , 
        \wColumn_17[53] , \wColumn_17[52] , \wColumn_17[51] , \wColumn_17[50] , 
        \wColumn_17[49] , \wColumn_17[48] , \wColumn_17[47] , \wColumn_17[46] , 
        \wColumn_17[45] , \wColumn_17[44] , \wColumn_17[43] , \wColumn_17[42] , 
        \wColumn_17[41] , \wColumn_17[40] , \wColumn_17[39] , \wColumn_17[38] , 
        \wColumn_17[37] , \wColumn_17[36] , \wColumn_17[35] , \wColumn_17[34] , 
        \wColumn_17[33] , \wColumn_17[32] , \wColumn_17[31] , \wColumn_17[30] , 
        \wColumn_17[29] , \wColumn_17[28] , \wColumn_17[27] , \wColumn_17[26] , 
        \wColumn_17[25] , \wColumn_17[24] , \wColumn_17[23] , \wColumn_17[22] , 
        \wColumn_17[21] , \wColumn_17[20] , \wColumn_17[19] , \wColumn_17[18] , 
        \wColumn_17[17] , \wColumn_17[16] , \wColumn_17[15] , \wColumn_17[14] , 
        \wColumn_17[13] , \wColumn_17[12] , \wColumn_17[11] , \wColumn_17[10] , 
        \wColumn_17[9] , \wColumn_17[8] , \wColumn_17[7] , \wColumn_17[6] , 
        \wColumn_17[5] , \wColumn_17[4] , \wColumn_17[3] , \wColumn_17[2] , 
        \wColumn_17[1] , \wColumn_17[0] }), .PDiagOut({\wPDiag_17[63] , 
        \wPDiag_17[62] , \wPDiag_17[61] , \wPDiag_17[60] , \wPDiag_17[59] , 
        \wPDiag_17[58] , \wPDiag_17[57] , \wPDiag_17[56] , \wPDiag_17[55] , 
        \wPDiag_17[54] , \wPDiag_17[53] , \wPDiag_17[52] , \wPDiag_17[51] , 
        \wPDiag_17[50] , \wPDiag_17[49] , \wPDiag_17[48] , \wPDiag_17[47] , 
        \wPDiag_17[46] , \wPDiag_17[45] , \wPDiag_17[44] , \wPDiag_17[43] , 
        \wPDiag_17[42] , \wPDiag_17[41] , \wPDiag_17[40] , \wPDiag_17[39] , 
        \wPDiag_17[38] , \wPDiag_17[37] , \wPDiag_17[36] , \wPDiag_17[35] , 
        \wPDiag_17[34] , \wPDiag_17[33] , \wPDiag_17[32] , \wPDiag_17[31] , 
        \wPDiag_17[30] , \wPDiag_17[29] , \wPDiag_17[28] , \wPDiag_17[27] , 
        \wPDiag_17[26] , \wPDiag_17[25] , \wPDiag_17[24] , \wPDiag_17[23] , 
        \wPDiag_17[22] , \wPDiag_17[21] , \wPDiag_17[20] , \wPDiag_17[19] , 
        \wPDiag_17[18] , \wPDiag_17[17] , \wPDiag_17[16] , \wPDiag_17[15] , 
        \wPDiag_17[14] , \wPDiag_17[13] , \wPDiag_17[12] , \wPDiag_17[11] , 
        \wPDiag_17[10] , \wPDiag_17[9] , \wPDiag_17[8] , \wPDiag_17[7] , 
        \wPDiag_17[6] , \wPDiag_17[5] , \wPDiag_17[4] , \wPDiag_17[3] , 
        \wPDiag_17[2] , \wPDiag_17[1] , \wPDiag_17[0] }), .NDiagOut({
        \wNDiag_17[63] , \wNDiag_17[62] , \wNDiag_17[61] , \wNDiag_17[60] , 
        \wNDiag_17[59] , \wNDiag_17[58] , \wNDiag_17[57] , \wNDiag_17[56] , 
        \wNDiag_17[55] , \wNDiag_17[54] , \wNDiag_17[53] , \wNDiag_17[52] , 
        \wNDiag_17[51] , \wNDiag_17[50] , \wNDiag_17[49] , \wNDiag_17[48] , 
        \wNDiag_17[47] , \wNDiag_17[46] , \wNDiag_17[45] , \wNDiag_17[44] , 
        \wNDiag_17[43] , \wNDiag_17[42] , \wNDiag_17[41] , \wNDiag_17[40] , 
        \wNDiag_17[39] , \wNDiag_17[38] , \wNDiag_17[37] , \wNDiag_17[36] , 
        \wNDiag_17[35] , \wNDiag_17[34] , \wNDiag_17[33] , \wNDiag_17[32] , 
        \wNDiag_17[31] , \wNDiag_17[30] , \wNDiag_17[29] , \wNDiag_17[28] , 
        \wNDiag_17[27] , \wNDiag_17[26] , \wNDiag_17[25] , \wNDiag_17[24] , 
        \wNDiag_17[23] , \wNDiag_17[22] , \wNDiag_17[21] , \wNDiag_17[20] , 
        \wNDiag_17[19] , \wNDiag_17[18] , \wNDiag_17[17] , \wNDiag_17[16] , 
        \wNDiag_17[15] , \wNDiag_17[14] , \wNDiag_17[13] , \wNDiag_17[12] , 
        \wNDiag_17[11] , \wNDiag_17[10] , \wNDiag_17[9] , \wNDiag_17[8] , 
        \wNDiag_17[7] , \wNDiag_17[6] , \wNDiag_17[5] , \wNDiag_17[4] , 
        \wNDiag_17[3] , \wNDiag_17[2] , \wNDiag_17[1] , \wNDiag_17[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_23 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_24[6] , \wScan_24[5] , \wScan_24[4] , 
        \wScan_24[3] , \wScan_24[2] , \wScan_24[1] , \wScan_24[0] }), 
        .ScanOut({\wScan_23[6] , \wScan_23[5] , \wScan_23[4] , \wScan_23[3] , 
        \wScan_23[2] , \wScan_23[1] , \wScan_23[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_23[0] ), .ReturnIn(\wReturn_24[0] ), .ColIn({
        \wColumn_23[63] , \wColumn_23[62] , \wColumn_23[61] , \wColumn_23[60] , 
        \wColumn_23[59] , \wColumn_23[58] , \wColumn_23[57] , \wColumn_23[56] , 
        \wColumn_23[55] , \wColumn_23[54] , \wColumn_23[53] , \wColumn_23[52] , 
        \wColumn_23[51] , \wColumn_23[50] , \wColumn_23[49] , \wColumn_23[48] , 
        \wColumn_23[47] , \wColumn_23[46] , \wColumn_23[45] , \wColumn_23[44] , 
        \wColumn_23[43] , \wColumn_23[42] , \wColumn_23[41] , \wColumn_23[40] , 
        \wColumn_23[39] , \wColumn_23[38] , \wColumn_23[37] , \wColumn_23[36] , 
        \wColumn_23[35] , \wColumn_23[34] , \wColumn_23[33] , \wColumn_23[32] , 
        \wColumn_23[31] , \wColumn_23[30] , \wColumn_23[29] , \wColumn_23[28] , 
        \wColumn_23[27] , \wColumn_23[26] , \wColumn_23[25] , \wColumn_23[24] , 
        \wColumn_23[23] , \wColumn_23[22] , \wColumn_23[21] , \wColumn_23[20] , 
        \wColumn_23[19] , \wColumn_23[18] , \wColumn_23[17] , \wColumn_23[16] , 
        \wColumn_23[15] , \wColumn_23[14] , \wColumn_23[13] , \wColumn_23[12] , 
        \wColumn_23[11] , \wColumn_23[10] , \wColumn_23[9] , \wColumn_23[8] , 
        \wColumn_23[7] , \wColumn_23[6] , \wColumn_23[5] , \wColumn_23[4] , 
        \wColumn_23[3] , \wColumn_23[2] , \wColumn_23[1] , \wColumn_23[0] }), 
        .PDiagIn({\wPDiag_23[63] , \wPDiag_23[62] , \wPDiag_23[61] , 
        \wPDiag_23[60] , \wPDiag_23[59] , \wPDiag_23[58] , \wPDiag_23[57] , 
        \wPDiag_23[56] , \wPDiag_23[55] , \wPDiag_23[54] , \wPDiag_23[53] , 
        \wPDiag_23[52] , \wPDiag_23[51] , \wPDiag_23[50] , \wPDiag_23[49] , 
        \wPDiag_23[48] , \wPDiag_23[47] , \wPDiag_23[46] , \wPDiag_23[45] , 
        \wPDiag_23[44] , \wPDiag_23[43] , \wPDiag_23[42] , \wPDiag_23[41] , 
        \wPDiag_23[40] , \wPDiag_23[39] , \wPDiag_23[38] , \wPDiag_23[37] , 
        \wPDiag_23[36] , \wPDiag_23[35] , \wPDiag_23[34] , \wPDiag_23[33] , 
        \wPDiag_23[32] , \wPDiag_23[31] , \wPDiag_23[30] , \wPDiag_23[29] , 
        \wPDiag_23[28] , \wPDiag_23[27] , \wPDiag_23[26] , \wPDiag_23[25] , 
        \wPDiag_23[24] , \wPDiag_23[23] , \wPDiag_23[22] , \wPDiag_23[21] , 
        \wPDiag_23[20] , \wPDiag_23[19] , \wPDiag_23[18] , \wPDiag_23[17] , 
        \wPDiag_23[16] , \wPDiag_23[15] , \wPDiag_23[14] , \wPDiag_23[13] , 
        \wPDiag_23[12] , \wPDiag_23[11] , \wPDiag_23[10] , \wPDiag_23[9] , 
        \wPDiag_23[8] , \wPDiag_23[7] , \wPDiag_23[6] , \wPDiag_23[5] , 
        \wPDiag_23[4] , \wPDiag_23[3] , \wPDiag_23[2] , \wPDiag_23[1] , 
        \wPDiag_23[0] }), .NDiagIn({\wNDiag_23[63] , \wNDiag_23[62] , 
        \wNDiag_23[61] , \wNDiag_23[60] , \wNDiag_23[59] , \wNDiag_23[58] , 
        \wNDiag_23[57] , \wNDiag_23[56] , \wNDiag_23[55] , \wNDiag_23[54] , 
        \wNDiag_23[53] , \wNDiag_23[52] , \wNDiag_23[51] , \wNDiag_23[50] , 
        \wNDiag_23[49] , \wNDiag_23[48] , \wNDiag_23[47] , \wNDiag_23[46] , 
        \wNDiag_23[45] , \wNDiag_23[44] , \wNDiag_23[43] , \wNDiag_23[42] , 
        \wNDiag_23[41] , \wNDiag_23[40] , \wNDiag_23[39] , \wNDiag_23[38] , 
        \wNDiag_23[37] , \wNDiag_23[36] , \wNDiag_23[35] , \wNDiag_23[34] , 
        \wNDiag_23[33] , \wNDiag_23[32] , \wNDiag_23[31] , \wNDiag_23[30] , 
        \wNDiag_23[29] , \wNDiag_23[28] , \wNDiag_23[27] , \wNDiag_23[26] , 
        \wNDiag_23[25] , \wNDiag_23[24] , \wNDiag_23[23] , \wNDiag_23[22] , 
        \wNDiag_23[21] , \wNDiag_23[20] , \wNDiag_23[19] , \wNDiag_23[18] , 
        \wNDiag_23[17] , \wNDiag_23[16] , \wNDiag_23[15] , \wNDiag_23[14] , 
        \wNDiag_23[13] , \wNDiag_23[12] , \wNDiag_23[11] , \wNDiag_23[10] , 
        \wNDiag_23[9] , \wNDiag_23[8] , \wNDiag_23[7] , \wNDiag_23[6] , 
        \wNDiag_23[5] , \wNDiag_23[4] , \wNDiag_23[3] , \wNDiag_23[2] , 
        \wNDiag_23[1] , \wNDiag_23[0] }), .CallOut(\wCall_24[0] ), .ReturnOut(
        \wReturn_23[0] ), .ColOut({\wColumn_24[63] , \wColumn_24[62] , 
        \wColumn_24[61] , \wColumn_24[60] , \wColumn_24[59] , \wColumn_24[58] , 
        \wColumn_24[57] , \wColumn_24[56] , \wColumn_24[55] , \wColumn_24[54] , 
        \wColumn_24[53] , \wColumn_24[52] , \wColumn_24[51] , \wColumn_24[50] , 
        \wColumn_24[49] , \wColumn_24[48] , \wColumn_24[47] , \wColumn_24[46] , 
        \wColumn_24[45] , \wColumn_24[44] , \wColumn_24[43] , \wColumn_24[42] , 
        \wColumn_24[41] , \wColumn_24[40] , \wColumn_24[39] , \wColumn_24[38] , 
        \wColumn_24[37] , \wColumn_24[36] , \wColumn_24[35] , \wColumn_24[34] , 
        \wColumn_24[33] , \wColumn_24[32] , \wColumn_24[31] , \wColumn_24[30] , 
        \wColumn_24[29] , \wColumn_24[28] , \wColumn_24[27] , \wColumn_24[26] , 
        \wColumn_24[25] , \wColumn_24[24] , \wColumn_24[23] , \wColumn_24[22] , 
        \wColumn_24[21] , \wColumn_24[20] , \wColumn_24[19] , \wColumn_24[18] , 
        \wColumn_24[17] , \wColumn_24[16] , \wColumn_24[15] , \wColumn_24[14] , 
        \wColumn_24[13] , \wColumn_24[12] , \wColumn_24[11] , \wColumn_24[10] , 
        \wColumn_24[9] , \wColumn_24[8] , \wColumn_24[7] , \wColumn_24[6] , 
        \wColumn_24[5] , \wColumn_24[4] , \wColumn_24[3] , \wColumn_24[2] , 
        \wColumn_24[1] , \wColumn_24[0] }), .PDiagOut({\wPDiag_24[63] , 
        \wPDiag_24[62] , \wPDiag_24[61] , \wPDiag_24[60] , \wPDiag_24[59] , 
        \wPDiag_24[58] , \wPDiag_24[57] , \wPDiag_24[56] , \wPDiag_24[55] , 
        \wPDiag_24[54] , \wPDiag_24[53] , \wPDiag_24[52] , \wPDiag_24[51] , 
        \wPDiag_24[50] , \wPDiag_24[49] , \wPDiag_24[48] , \wPDiag_24[47] , 
        \wPDiag_24[46] , \wPDiag_24[45] , \wPDiag_24[44] , \wPDiag_24[43] , 
        \wPDiag_24[42] , \wPDiag_24[41] , \wPDiag_24[40] , \wPDiag_24[39] , 
        \wPDiag_24[38] , \wPDiag_24[37] , \wPDiag_24[36] , \wPDiag_24[35] , 
        \wPDiag_24[34] , \wPDiag_24[33] , \wPDiag_24[32] , \wPDiag_24[31] , 
        \wPDiag_24[30] , \wPDiag_24[29] , \wPDiag_24[28] , \wPDiag_24[27] , 
        \wPDiag_24[26] , \wPDiag_24[25] , \wPDiag_24[24] , \wPDiag_24[23] , 
        \wPDiag_24[22] , \wPDiag_24[21] , \wPDiag_24[20] , \wPDiag_24[19] , 
        \wPDiag_24[18] , \wPDiag_24[17] , \wPDiag_24[16] , \wPDiag_24[15] , 
        \wPDiag_24[14] , \wPDiag_24[13] , \wPDiag_24[12] , \wPDiag_24[11] , 
        \wPDiag_24[10] , \wPDiag_24[9] , \wPDiag_24[8] , \wPDiag_24[7] , 
        \wPDiag_24[6] , \wPDiag_24[5] , \wPDiag_24[4] , \wPDiag_24[3] , 
        \wPDiag_24[2] , \wPDiag_24[1] , \wPDiag_24[0] }), .NDiagOut({
        \wNDiag_24[63] , \wNDiag_24[62] , \wNDiag_24[61] , \wNDiag_24[60] , 
        \wNDiag_24[59] , \wNDiag_24[58] , \wNDiag_24[57] , \wNDiag_24[56] , 
        \wNDiag_24[55] , \wNDiag_24[54] , \wNDiag_24[53] , \wNDiag_24[52] , 
        \wNDiag_24[51] , \wNDiag_24[50] , \wNDiag_24[49] , \wNDiag_24[48] , 
        \wNDiag_24[47] , \wNDiag_24[46] , \wNDiag_24[45] , \wNDiag_24[44] , 
        \wNDiag_24[43] , \wNDiag_24[42] , \wNDiag_24[41] , \wNDiag_24[40] , 
        \wNDiag_24[39] , \wNDiag_24[38] , \wNDiag_24[37] , \wNDiag_24[36] , 
        \wNDiag_24[35] , \wNDiag_24[34] , \wNDiag_24[33] , \wNDiag_24[32] , 
        \wNDiag_24[31] , \wNDiag_24[30] , \wNDiag_24[29] , \wNDiag_24[28] , 
        \wNDiag_24[27] , \wNDiag_24[26] , \wNDiag_24[25] , \wNDiag_24[24] , 
        \wNDiag_24[23] , \wNDiag_24[22] , \wNDiag_24[21] , \wNDiag_24[20] , 
        \wNDiag_24[19] , \wNDiag_24[18] , \wNDiag_24[17] , \wNDiag_24[16] , 
        \wNDiag_24[15] , \wNDiag_24[14] , \wNDiag_24[13] , \wNDiag_24[12] , 
        \wNDiag_24[11] , \wNDiag_24[10] , \wNDiag_24[9] , \wNDiag_24[8] , 
        \wNDiag_24[7] , \wNDiag_24[6] , \wNDiag_24[5] , \wNDiag_24[4] , 
        \wNDiag_24[3] , \wNDiag_24[2] , \wNDiag_24[1] , \wNDiag_24[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_31 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_32[6] , \wScan_32[5] , \wScan_32[4] , 
        \wScan_32[3] , \wScan_32[2] , \wScan_32[1] , \wScan_32[0] }), 
        .ScanOut({\wScan_31[6] , \wScan_31[5] , \wScan_31[4] , \wScan_31[3] , 
        \wScan_31[2] , \wScan_31[1] , \wScan_31[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_31[0] ), .ReturnIn(\wReturn_32[0] ), .ColIn({
        \wColumn_31[63] , \wColumn_31[62] , \wColumn_31[61] , \wColumn_31[60] , 
        \wColumn_31[59] , \wColumn_31[58] , \wColumn_31[57] , \wColumn_31[56] , 
        \wColumn_31[55] , \wColumn_31[54] , \wColumn_31[53] , \wColumn_31[52] , 
        \wColumn_31[51] , \wColumn_31[50] , \wColumn_31[49] , \wColumn_31[48] , 
        \wColumn_31[47] , \wColumn_31[46] , \wColumn_31[45] , \wColumn_31[44] , 
        \wColumn_31[43] , \wColumn_31[42] , \wColumn_31[41] , \wColumn_31[40] , 
        \wColumn_31[39] , \wColumn_31[38] , \wColumn_31[37] , \wColumn_31[36] , 
        \wColumn_31[35] , \wColumn_31[34] , \wColumn_31[33] , \wColumn_31[32] , 
        \wColumn_31[31] , \wColumn_31[30] , \wColumn_31[29] , \wColumn_31[28] , 
        \wColumn_31[27] , \wColumn_31[26] , \wColumn_31[25] , \wColumn_31[24] , 
        \wColumn_31[23] , \wColumn_31[22] , \wColumn_31[21] , \wColumn_31[20] , 
        \wColumn_31[19] , \wColumn_31[18] , \wColumn_31[17] , \wColumn_31[16] , 
        \wColumn_31[15] , \wColumn_31[14] , \wColumn_31[13] , \wColumn_31[12] , 
        \wColumn_31[11] , \wColumn_31[10] , \wColumn_31[9] , \wColumn_31[8] , 
        \wColumn_31[7] , \wColumn_31[6] , \wColumn_31[5] , \wColumn_31[4] , 
        \wColumn_31[3] , \wColumn_31[2] , \wColumn_31[1] , \wColumn_31[0] }), 
        .PDiagIn({\wPDiag_31[63] , \wPDiag_31[62] , \wPDiag_31[61] , 
        \wPDiag_31[60] , \wPDiag_31[59] , \wPDiag_31[58] , \wPDiag_31[57] , 
        \wPDiag_31[56] , \wPDiag_31[55] , \wPDiag_31[54] , \wPDiag_31[53] , 
        \wPDiag_31[52] , \wPDiag_31[51] , \wPDiag_31[50] , \wPDiag_31[49] , 
        \wPDiag_31[48] , \wPDiag_31[47] , \wPDiag_31[46] , \wPDiag_31[45] , 
        \wPDiag_31[44] , \wPDiag_31[43] , \wPDiag_31[42] , \wPDiag_31[41] , 
        \wPDiag_31[40] , \wPDiag_31[39] , \wPDiag_31[38] , \wPDiag_31[37] , 
        \wPDiag_31[36] , \wPDiag_31[35] , \wPDiag_31[34] , \wPDiag_31[33] , 
        \wPDiag_31[32] , \wPDiag_31[31] , \wPDiag_31[30] , \wPDiag_31[29] , 
        \wPDiag_31[28] , \wPDiag_31[27] , \wPDiag_31[26] , \wPDiag_31[25] , 
        \wPDiag_31[24] , \wPDiag_31[23] , \wPDiag_31[22] , \wPDiag_31[21] , 
        \wPDiag_31[20] , \wPDiag_31[19] , \wPDiag_31[18] , \wPDiag_31[17] , 
        \wPDiag_31[16] , \wPDiag_31[15] , \wPDiag_31[14] , \wPDiag_31[13] , 
        \wPDiag_31[12] , \wPDiag_31[11] , \wPDiag_31[10] , \wPDiag_31[9] , 
        \wPDiag_31[8] , \wPDiag_31[7] , \wPDiag_31[6] , \wPDiag_31[5] , 
        \wPDiag_31[4] , \wPDiag_31[3] , \wPDiag_31[2] , \wPDiag_31[1] , 
        \wPDiag_31[0] }), .NDiagIn({\wNDiag_31[63] , \wNDiag_31[62] , 
        \wNDiag_31[61] , \wNDiag_31[60] , \wNDiag_31[59] , \wNDiag_31[58] , 
        \wNDiag_31[57] , \wNDiag_31[56] , \wNDiag_31[55] , \wNDiag_31[54] , 
        \wNDiag_31[53] , \wNDiag_31[52] , \wNDiag_31[51] , \wNDiag_31[50] , 
        \wNDiag_31[49] , \wNDiag_31[48] , \wNDiag_31[47] , \wNDiag_31[46] , 
        \wNDiag_31[45] , \wNDiag_31[44] , \wNDiag_31[43] , \wNDiag_31[42] , 
        \wNDiag_31[41] , \wNDiag_31[40] , \wNDiag_31[39] , \wNDiag_31[38] , 
        \wNDiag_31[37] , \wNDiag_31[36] , \wNDiag_31[35] , \wNDiag_31[34] , 
        \wNDiag_31[33] , \wNDiag_31[32] , \wNDiag_31[31] , \wNDiag_31[30] , 
        \wNDiag_31[29] , \wNDiag_31[28] , \wNDiag_31[27] , \wNDiag_31[26] , 
        \wNDiag_31[25] , \wNDiag_31[24] , \wNDiag_31[23] , \wNDiag_31[22] , 
        \wNDiag_31[21] , \wNDiag_31[20] , \wNDiag_31[19] , \wNDiag_31[18] , 
        \wNDiag_31[17] , \wNDiag_31[16] , \wNDiag_31[15] , \wNDiag_31[14] , 
        \wNDiag_31[13] , \wNDiag_31[12] , \wNDiag_31[11] , \wNDiag_31[10] , 
        \wNDiag_31[9] , \wNDiag_31[8] , \wNDiag_31[7] , \wNDiag_31[6] , 
        \wNDiag_31[5] , \wNDiag_31[4] , \wNDiag_31[3] , \wNDiag_31[2] , 
        \wNDiag_31[1] , \wNDiag_31[0] }), .CallOut(\wCall_32[0] ), .ReturnOut(
        \wReturn_31[0] ), .ColOut({\wColumn_32[63] , \wColumn_32[62] , 
        \wColumn_32[61] , \wColumn_32[60] , \wColumn_32[59] , \wColumn_32[58] , 
        \wColumn_32[57] , \wColumn_32[56] , \wColumn_32[55] , \wColumn_32[54] , 
        \wColumn_32[53] , \wColumn_32[52] , \wColumn_32[51] , \wColumn_32[50] , 
        \wColumn_32[49] , \wColumn_32[48] , \wColumn_32[47] , \wColumn_32[46] , 
        \wColumn_32[45] , \wColumn_32[44] , \wColumn_32[43] , \wColumn_32[42] , 
        \wColumn_32[41] , \wColumn_32[40] , \wColumn_32[39] , \wColumn_32[38] , 
        \wColumn_32[37] , \wColumn_32[36] , \wColumn_32[35] , \wColumn_32[34] , 
        \wColumn_32[33] , \wColumn_32[32] , \wColumn_32[31] , \wColumn_32[30] , 
        \wColumn_32[29] , \wColumn_32[28] , \wColumn_32[27] , \wColumn_32[26] , 
        \wColumn_32[25] , \wColumn_32[24] , \wColumn_32[23] , \wColumn_32[22] , 
        \wColumn_32[21] , \wColumn_32[20] , \wColumn_32[19] , \wColumn_32[18] , 
        \wColumn_32[17] , \wColumn_32[16] , \wColumn_32[15] , \wColumn_32[14] , 
        \wColumn_32[13] , \wColumn_32[12] , \wColumn_32[11] , \wColumn_32[10] , 
        \wColumn_32[9] , \wColumn_32[8] , \wColumn_32[7] , \wColumn_32[6] , 
        \wColumn_32[5] , \wColumn_32[4] , \wColumn_32[3] , \wColumn_32[2] , 
        \wColumn_32[1] , \wColumn_32[0] }), .PDiagOut({\wPDiag_32[63] , 
        \wPDiag_32[62] , \wPDiag_32[61] , \wPDiag_32[60] , \wPDiag_32[59] , 
        \wPDiag_32[58] , \wPDiag_32[57] , \wPDiag_32[56] , \wPDiag_32[55] , 
        \wPDiag_32[54] , \wPDiag_32[53] , \wPDiag_32[52] , \wPDiag_32[51] , 
        \wPDiag_32[50] , \wPDiag_32[49] , \wPDiag_32[48] , \wPDiag_32[47] , 
        \wPDiag_32[46] , \wPDiag_32[45] , \wPDiag_32[44] , \wPDiag_32[43] , 
        \wPDiag_32[42] , \wPDiag_32[41] , \wPDiag_32[40] , \wPDiag_32[39] , 
        \wPDiag_32[38] , \wPDiag_32[37] , \wPDiag_32[36] , \wPDiag_32[35] , 
        \wPDiag_32[34] , \wPDiag_32[33] , \wPDiag_32[32] , \wPDiag_32[31] , 
        \wPDiag_32[30] , \wPDiag_32[29] , \wPDiag_32[28] , \wPDiag_32[27] , 
        \wPDiag_32[26] , \wPDiag_32[25] , \wPDiag_32[24] , \wPDiag_32[23] , 
        \wPDiag_32[22] , \wPDiag_32[21] , \wPDiag_32[20] , \wPDiag_32[19] , 
        \wPDiag_32[18] , \wPDiag_32[17] , \wPDiag_32[16] , \wPDiag_32[15] , 
        \wPDiag_32[14] , \wPDiag_32[13] , \wPDiag_32[12] , \wPDiag_32[11] , 
        \wPDiag_32[10] , \wPDiag_32[9] , \wPDiag_32[8] , \wPDiag_32[7] , 
        \wPDiag_32[6] , \wPDiag_32[5] , \wPDiag_32[4] , \wPDiag_32[3] , 
        \wPDiag_32[2] , \wPDiag_32[1] , \wPDiag_32[0] }), .NDiagOut({
        \wNDiag_32[63] , \wNDiag_32[62] , \wNDiag_32[61] , \wNDiag_32[60] , 
        \wNDiag_32[59] , \wNDiag_32[58] , \wNDiag_32[57] , \wNDiag_32[56] , 
        \wNDiag_32[55] , \wNDiag_32[54] , \wNDiag_32[53] , \wNDiag_32[52] , 
        \wNDiag_32[51] , \wNDiag_32[50] , \wNDiag_32[49] , \wNDiag_32[48] , 
        \wNDiag_32[47] , \wNDiag_32[46] , \wNDiag_32[45] , \wNDiag_32[44] , 
        \wNDiag_32[43] , \wNDiag_32[42] , \wNDiag_32[41] , \wNDiag_32[40] , 
        \wNDiag_32[39] , \wNDiag_32[38] , \wNDiag_32[37] , \wNDiag_32[36] , 
        \wNDiag_32[35] , \wNDiag_32[34] , \wNDiag_32[33] , \wNDiag_32[32] , 
        \wNDiag_32[31] , \wNDiag_32[30] , \wNDiag_32[29] , \wNDiag_32[28] , 
        \wNDiag_32[27] , \wNDiag_32[26] , \wNDiag_32[25] , \wNDiag_32[24] , 
        \wNDiag_32[23] , \wNDiag_32[22] , \wNDiag_32[21] , \wNDiag_32[20] , 
        \wNDiag_32[19] , \wNDiag_32[18] , \wNDiag_32[17] , \wNDiag_32[16] , 
        \wNDiag_32[15] , \wNDiag_32[14] , \wNDiag_32[13] , \wNDiag_32[12] , 
        \wNDiag_32[11] , \wNDiag_32[10] , \wNDiag_32[9] , \wNDiag_32[8] , 
        \wNDiag_32[7] , \wNDiag_32[6] , \wNDiag_32[5] , \wNDiag_32[4] , 
        \wNDiag_32[3] , \wNDiag_32[2] , \wNDiag_32[1] , \wNDiag_32[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_22 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_23[6] , \wScan_23[5] , \wScan_23[4] , 
        \wScan_23[3] , \wScan_23[2] , \wScan_23[1] , \wScan_23[0] }), 
        .ScanOut({\wScan_22[6] , \wScan_22[5] , \wScan_22[4] , \wScan_22[3] , 
        \wScan_22[2] , \wScan_22[1] , \wScan_22[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_22[0] ), .ReturnIn(\wReturn_23[0] ), .ColIn({
        \wColumn_22[63] , \wColumn_22[62] , \wColumn_22[61] , \wColumn_22[60] , 
        \wColumn_22[59] , \wColumn_22[58] , \wColumn_22[57] , \wColumn_22[56] , 
        \wColumn_22[55] , \wColumn_22[54] , \wColumn_22[53] , \wColumn_22[52] , 
        \wColumn_22[51] , \wColumn_22[50] , \wColumn_22[49] , \wColumn_22[48] , 
        \wColumn_22[47] , \wColumn_22[46] , \wColumn_22[45] , \wColumn_22[44] , 
        \wColumn_22[43] , \wColumn_22[42] , \wColumn_22[41] , \wColumn_22[40] , 
        \wColumn_22[39] , \wColumn_22[38] , \wColumn_22[37] , \wColumn_22[36] , 
        \wColumn_22[35] , \wColumn_22[34] , \wColumn_22[33] , \wColumn_22[32] , 
        \wColumn_22[31] , \wColumn_22[30] , \wColumn_22[29] , \wColumn_22[28] , 
        \wColumn_22[27] , \wColumn_22[26] , \wColumn_22[25] , \wColumn_22[24] , 
        \wColumn_22[23] , \wColumn_22[22] , \wColumn_22[21] , \wColumn_22[20] , 
        \wColumn_22[19] , \wColumn_22[18] , \wColumn_22[17] , \wColumn_22[16] , 
        \wColumn_22[15] , \wColumn_22[14] , \wColumn_22[13] , \wColumn_22[12] , 
        \wColumn_22[11] , \wColumn_22[10] , \wColumn_22[9] , \wColumn_22[8] , 
        \wColumn_22[7] , \wColumn_22[6] , \wColumn_22[5] , \wColumn_22[4] , 
        \wColumn_22[3] , \wColumn_22[2] , \wColumn_22[1] , \wColumn_22[0] }), 
        .PDiagIn({\wPDiag_22[63] , \wPDiag_22[62] , \wPDiag_22[61] , 
        \wPDiag_22[60] , \wPDiag_22[59] , \wPDiag_22[58] , \wPDiag_22[57] , 
        \wPDiag_22[56] , \wPDiag_22[55] , \wPDiag_22[54] , \wPDiag_22[53] , 
        \wPDiag_22[52] , \wPDiag_22[51] , \wPDiag_22[50] , \wPDiag_22[49] , 
        \wPDiag_22[48] , \wPDiag_22[47] , \wPDiag_22[46] , \wPDiag_22[45] , 
        \wPDiag_22[44] , \wPDiag_22[43] , \wPDiag_22[42] , \wPDiag_22[41] , 
        \wPDiag_22[40] , \wPDiag_22[39] , \wPDiag_22[38] , \wPDiag_22[37] , 
        \wPDiag_22[36] , \wPDiag_22[35] , \wPDiag_22[34] , \wPDiag_22[33] , 
        \wPDiag_22[32] , \wPDiag_22[31] , \wPDiag_22[30] , \wPDiag_22[29] , 
        \wPDiag_22[28] , \wPDiag_22[27] , \wPDiag_22[26] , \wPDiag_22[25] , 
        \wPDiag_22[24] , \wPDiag_22[23] , \wPDiag_22[22] , \wPDiag_22[21] , 
        \wPDiag_22[20] , \wPDiag_22[19] , \wPDiag_22[18] , \wPDiag_22[17] , 
        \wPDiag_22[16] , \wPDiag_22[15] , \wPDiag_22[14] , \wPDiag_22[13] , 
        \wPDiag_22[12] , \wPDiag_22[11] , \wPDiag_22[10] , \wPDiag_22[9] , 
        \wPDiag_22[8] , \wPDiag_22[7] , \wPDiag_22[6] , \wPDiag_22[5] , 
        \wPDiag_22[4] , \wPDiag_22[3] , \wPDiag_22[2] , \wPDiag_22[1] , 
        \wPDiag_22[0] }), .NDiagIn({\wNDiag_22[63] , \wNDiag_22[62] , 
        \wNDiag_22[61] , \wNDiag_22[60] , \wNDiag_22[59] , \wNDiag_22[58] , 
        \wNDiag_22[57] , \wNDiag_22[56] , \wNDiag_22[55] , \wNDiag_22[54] , 
        \wNDiag_22[53] , \wNDiag_22[52] , \wNDiag_22[51] , \wNDiag_22[50] , 
        \wNDiag_22[49] , \wNDiag_22[48] , \wNDiag_22[47] , \wNDiag_22[46] , 
        \wNDiag_22[45] , \wNDiag_22[44] , \wNDiag_22[43] , \wNDiag_22[42] , 
        \wNDiag_22[41] , \wNDiag_22[40] , \wNDiag_22[39] , \wNDiag_22[38] , 
        \wNDiag_22[37] , \wNDiag_22[36] , \wNDiag_22[35] , \wNDiag_22[34] , 
        \wNDiag_22[33] , \wNDiag_22[32] , \wNDiag_22[31] , \wNDiag_22[30] , 
        \wNDiag_22[29] , \wNDiag_22[28] , \wNDiag_22[27] , \wNDiag_22[26] , 
        \wNDiag_22[25] , \wNDiag_22[24] , \wNDiag_22[23] , \wNDiag_22[22] , 
        \wNDiag_22[21] , \wNDiag_22[20] , \wNDiag_22[19] , \wNDiag_22[18] , 
        \wNDiag_22[17] , \wNDiag_22[16] , \wNDiag_22[15] , \wNDiag_22[14] , 
        \wNDiag_22[13] , \wNDiag_22[12] , \wNDiag_22[11] , \wNDiag_22[10] , 
        \wNDiag_22[9] , \wNDiag_22[8] , \wNDiag_22[7] , \wNDiag_22[6] , 
        \wNDiag_22[5] , \wNDiag_22[4] , \wNDiag_22[3] , \wNDiag_22[2] , 
        \wNDiag_22[1] , \wNDiag_22[0] }), .CallOut(\wCall_23[0] ), .ReturnOut(
        \wReturn_22[0] ), .ColOut({\wColumn_23[63] , \wColumn_23[62] , 
        \wColumn_23[61] , \wColumn_23[60] , \wColumn_23[59] , \wColumn_23[58] , 
        \wColumn_23[57] , \wColumn_23[56] , \wColumn_23[55] , \wColumn_23[54] , 
        \wColumn_23[53] , \wColumn_23[52] , \wColumn_23[51] , \wColumn_23[50] , 
        \wColumn_23[49] , \wColumn_23[48] , \wColumn_23[47] , \wColumn_23[46] , 
        \wColumn_23[45] , \wColumn_23[44] , \wColumn_23[43] , \wColumn_23[42] , 
        \wColumn_23[41] , \wColumn_23[40] , \wColumn_23[39] , \wColumn_23[38] , 
        \wColumn_23[37] , \wColumn_23[36] , \wColumn_23[35] , \wColumn_23[34] , 
        \wColumn_23[33] , \wColumn_23[32] , \wColumn_23[31] , \wColumn_23[30] , 
        \wColumn_23[29] , \wColumn_23[28] , \wColumn_23[27] , \wColumn_23[26] , 
        \wColumn_23[25] , \wColumn_23[24] , \wColumn_23[23] , \wColumn_23[22] , 
        \wColumn_23[21] , \wColumn_23[20] , \wColumn_23[19] , \wColumn_23[18] , 
        \wColumn_23[17] , \wColumn_23[16] , \wColumn_23[15] , \wColumn_23[14] , 
        \wColumn_23[13] , \wColumn_23[12] , \wColumn_23[11] , \wColumn_23[10] , 
        \wColumn_23[9] , \wColumn_23[8] , \wColumn_23[7] , \wColumn_23[6] , 
        \wColumn_23[5] , \wColumn_23[4] , \wColumn_23[3] , \wColumn_23[2] , 
        \wColumn_23[1] , \wColumn_23[0] }), .PDiagOut({\wPDiag_23[63] , 
        \wPDiag_23[62] , \wPDiag_23[61] , \wPDiag_23[60] , \wPDiag_23[59] , 
        \wPDiag_23[58] , \wPDiag_23[57] , \wPDiag_23[56] , \wPDiag_23[55] , 
        \wPDiag_23[54] , \wPDiag_23[53] , \wPDiag_23[52] , \wPDiag_23[51] , 
        \wPDiag_23[50] , \wPDiag_23[49] , \wPDiag_23[48] , \wPDiag_23[47] , 
        \wPDiag_23[46] , \wPDiag_23[45] , \wPDiag_23[44] , \wPDiag_23[43] , 
        \wPDiag_23[42] , \wPDiag_23[41] , \wPDiag_23[40] , \wPDiag_23[39] , 
        \wPDiag_23[38] , \wPDiag_23[37] , \wPDiag_23[36] , \wPDiag_23[35] , 
        \wPDiag_23[34] , \wPDiag_23[33] , \wPDiag_23[32] , \wPDiag_23[31] , 
        \wPDiag_23[30] , \wPDiag_23[29] , \wPDiag_23[28] , \wPDiag_23[27] , 
        \wPDiag_23[26] , \wPDiag_23[25] , \wPDiag_23[24] , \wPDiag_23[23] , 
        \wPDiag_23[22] , \wPDiag_23[21] , \wPDiag_23[20] , \wPDiag_23[19] , 
        \wPDiag_23[18] , \wPDiag_23[17] , \wPDiag_23[16] , \wPDiag_23[15] , 
        \wPDiag_23[14] , \wPDiag_23[13] , \wPDiag_23[12] , \wPDiag_23[11] , 
        \wPDiag_23[10] , \wPDiag_23[9] , \wPDiag_23[8] , \wPDiag_23[7] , 
        \wPDiag_23[6] , \wPDiag_23[5] , \wPDiag_23[4] , \wPDiag_23[3] , 
        \wPDiag_23[2] , \wPDiag_23[1] , \wPDiag_23[0] }), .NDiagOut({
        \wNDiag_23[63] , \wNDiag_23[62] , \wNDiag_23[61] , \wNDiag_23[60] , 
        \wNDiag_23[59] , \wNDiag_23[58] , \wNDiag_23[57] , \wNDiag_23[56] , 
        \wNDiag_23[55] , \wNDiag_23[54] , \wNDiag_23[53] , \wNDiag_23[52] , 
        \wNDiag_23[51] , \wNDiag_23[50] , \wNDiag_23[49] , \wNDiag_23[48] , 
        \wNDiag_23[47] , \wNDiag_23[46] , \wNDiag_23[45] , \wNDiag_23[44] , 
        \wNDiag_23[43] , \wNDiag_23[42] , \wNDiag_23[41] , \wNDiag_23[40] , 
        \wNDiag_23[39] , \wNDiag_23[38] , \wNDiag_23[37] , \wNDiag_23[36] , 
        \wNDiag_23[35] , \wNDiag_23[34] , \wNDiag_23[33] , \wNDiag_23[32] , 
        \wNDiag_23[31] , \wNDiag_23[30] , \wNDiag_23[29] , \wNDiag_23[28] , 
        \wNDiag_23[27] , \wNDiag_23[26] , \wNDiag_23[25] , \wNDiag_23[24] , 
        \wNDiag_23[23] , \wNDiag_23[22] , \wNDiag_23[21] , \wNDiag_23[20] , 
        \wNDiag_23[19] , \wNDiag_23[18] , \wNDiag_23[17] , \wNDiag_23[16] , 
        \wNDiag_23[15] , \wNDiag_23[14] , \wNDiag_23[13] , \wNDiag_23[12] , 
        \wNDiag_23[11] , \wNDiag_23[10] , \wNDiag_23[9] , \wNDiag_23[8] , 
        \wNDiag_23[7] , \wNDiag_23[6] , \wNDiag_23[5] , \wNDiag_23[4] , 
        \wNDiag_23[3] , \wNDiag_23[2] , \wNDiag_23[1] , \wNDiag_23[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_44 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_45[6] , \wScan_45[5] , \wScan_45[4] , 
        \wScan_45[3] , \wScan_45[2] , \wScan_45[1] , \wScan_45[0] }), 
        .ScanOut({\wScan_44[6] , \wScan_44[5] , \wScan_44[4] , \wScan_44[3] , 
        \wScan_44[2] , \wScan_44[1] , \wScan_44[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_44[0] ), .ReturnIn(\wReturn_45[0] ), .ColIn({
        \wColumn_44[63] , \wColumn_44[62] , \wColumn_44[61] , \wColumn_44[60] , 
        \wColumn_44[59] , \wColumn_44[58] , \wColumn_44[57] , \wColumn_44[56] , 
        \wColumn_44[55] , \wColumn_44[54] , \wColumn_44[53] , \wColumn_44[52] , 
        \wColumn_44[51] , \wColumn_44[50] , \wColumn_44[49] , \wColumn_44[48] , 
        \wColumn_44[47] , \wColumn_44[46] , \wColumn_44[45] , \wColumn_44[44] , 
        \wColumn_44[43] , \wColumn_44[42] , \wColumn_44[41] , \wColumn_44[40] , 
        \wColumn_44[39] , \wColumn_44[38] , \wColumn_44[37] , \wColumn_44[36] , 
        \wColumn_44[35] , \wColumn_44[34] , \wColumn_44[33] , \wColumn_44[32] , 
        \wColumn_44[31] , \wColumn_44[30] , \wColumn_44[29] , \wColumn_44[28] , 
        \wColumn_44[27] , \wColumn_44[26] , \wColumn_44[25] , \wColumn_44[24] , 
        \wColumn_44[23] , \wColumn_44[22] , \wColumn_44[21] , \wColumn_44[20] , 
        \wColumn_44[19] , \wColumn_44[18] , \wColumn_44[17] , \wColumn_44[16] , 
        \wColumn_44[15] , \wColumn_44[14] , \wColumn_44[13] , \wColumn_44[12] , 
        \wColumn_44[11] , \wColumn_44[10] , \wColumn_44[9] , \wColumn_44[8] , 
        \wColumn_44[7] , \wColumn_44[6] , \wColumn_44[5] , \wColumn_44[4] , 
        \wColumn_44[3] , \wColumn_44[2] , \wColumn_44[1] , \wColumn_44[0] }), 
        .PDiagIn({\wPDiag_44[63] , \wPDiag_44[62] , \wPDiag_44[61] , 
        \wPDiag_44[60] , \wPDiag_44[59] , \wPDiag_44[58] , \wPDiag_44[57] , 
        \wPDiag_44[56] , \wPDiag_44[55] , \wPDiag_44[54] , \wPDiag_44[53] , 
        \wPDiag_44[52] , \wPDiag_44[51] , \wPDiag_44[50] , \wPDiag_44[49] , 
        \wPDiag_44[48] , \wPDiag_44[47] , \wPDiag_44[46] , \wPDiag_44[45] , 
        \wPDiag_44[44] , \wPDiag_44[43] , \wPDiag_44[42] , \wPDiag_44[41] , 
        \wPDiag_44[40] , \wPDiag_44[39] , \wPDiag_44[38] , \wPDiag_44[37] , 
        \wPDiag_44[36] , \wPDiag_44[35] , \wPDiag_44[34] , \wPDiag_44[33] , 
        \wPDiag_44[32] , \wPDiag_44[31] , \wPDiag_44[30] , \wPDiag_44[29] , 
        \wPDiag_44[28] , \wPDiag_44[27] , \wPDiag_44[26] , \wPDiag_44[25] , 
        \wPDiag_44[24] , \wPDiag_44[23] , \wPDiag_44[22] , \wPDiag_44[21] , 
        \wPDiag_44[20] , \wPDiag_44[19] , \wPDiag_44[18] , \wPDiag_44[17] , 
        \wPDiag_44[16] , \wPDiag_44[15] , \wPDiag_44[14] , \wPDiag_44[13] , 
        \wPDiag_44[12] , \wPDiag_44[11] , \wPDiag_44[10] , \wPDiag_44[9] , 
        \wPDiag_44[8] , \wPDiag_44[7] , \wPDiag_44[6] , \wPDiag_44[5] , 
        \wPDiag_44[4] , \wPDiag_44[3] , \wPDiag_44[2] , \wPDiag_44[1] , 
        \wPDiag_44[0] }), .NDiagIn({\wNDiag_44[63] , \wNDiag_44[62] , 
        \wNDiag_44[61] , \wNDiag_44[60] , \wNDiag_44[59] , \wNDiag_44[58] , 
        \wNDiag_44[57] , \wNDiag_44[56] , \wNDiag_44[55] , \wNDiag_44[54] , 
        \wNDiag_44[53] , \wNDiag_44[52] , \wNDiag_44[51] , \wNDiag_44[50] , 
        \wNDiag_44[49] , \wNDiag_44[48] , \wNDiag_44[47] , \wNDiag_44[46] , 
        \wNDiag_44[45] , \wNDiag_44[44] , \wNDiag_44[43] , \wNDiag_44[42] , 
        \wNDiag_44[41] , \wNDiag_44[40] , \wNDiag_44[39] , \wNDiag_44[38] , 
        \wNDiag_44[37] , \wNDiag_44[36] , \wNDiag_44[35] , \wNDiag_44[34] , 
        \wNDiag_44[33] , \wNDiag_44[32] , \wNDiag_44[31] , \wNDiag_44[30] , 
        \wNDiag_44[29] , \wNDiag_44[28] , \wNDiag_44[27] , \wNDiag_44[26] , 
        \wNDiag_44[25] , \wNDiag_44[24] , \wNDiag_44[23] , \wNDiag_44[22] , 
        \wNDiag_44[21] , \wNDiag_44[20] , \wNDiag_44[19] , \wNDiag_44[18] , 
        \wNDiag_44[17] , \wNDiag_44[16] , \wNDiag_44[15] , \wNDiag_44[14] , 
        \wNDiag_44[13] , \wNDiag_44[12] , \wNDiag_44[11] , \wNDiag_44[10] , 
        \wNDiag_44[9] , \wNDiag_44[8] , \wNDiag_44[7] , \wNDiag_44[6] , 
        \wNDiag_44[5] , \wNDiag_44[4] , \wNDiag_44[3] , \wNDiag_44[2] , 
        \wNDiag_44[1] , \wNDiag_44[0] }), .CallOut(\wCall_45[0] ), .ReturnOut(
        \wReturn_44[0] ), .ColOut({\wColumn_45[63] , \wColumn_45[62] , 
        \wColumn_45[61] , \wColumn_45[60] , \wColumn_45[59] , \wColumn_45[58] , 
        \wColumn_45[57] , \wColumn_45[56] , \wColumn_45[55] , \wColumn_45[54] , 
        \wColumn_45[53] , \wColumn_45[52] , \wColumn_45[51] , \wColumn_45[50] , 
        \wColumn_45[49] , \wColumn_45[48] , \wColumn_45[47] , \wColumn_45[46] , 
        \wColumn_45[45] , \wColumn_45[44] , \wColumn_45[43] , \wColumn_45[42] , 
        \wColumn_45[41] , \wColumn_45[40] , \wColumn_45[39] , \wColumn_45[38] , 
        \wColumn_45[37] , \wColumn_45[36] , \wColumn_45[35] , \wColumn_45[34] , 
        \wColumn_45[33] , \wColumn_45[32] , \wColumn_45[31] , \wColumn_45[30] , 
        \wColumn_45[29] , \wColumn_45[28] , \wColumn_45[27] , \wColumn_45[26] , 
        \wColumn_45[25] , \wColumn_45[24] , \wColumn_45[23] , \wColumn_45[22] , 
        \wColumn_45[21] , \wColumn_45[20] , \wColumn_45[19] , \wColumn_45[18] , 
        \wColumn_45[17] , \wColumn_45[16] , \wColumn_45[15] , \wColumn_45[14] , 
        \wColumn_45[13] , \wColumn_45[12] , \wColumn_45[11] , \wColumn_45[10] , 
        \wColumn_45[9] , \wColumn_45[8] , \wColumn_45[7] , \wColumn_45[6] , 
        \wColumn_45[5] , \wColumn_45[4] , \wColumn_45[3] , \wColumn_45[2] , 
        \wColumn_45[1] , \wColumn_45[0] }), .PDiagOut({\wPDiag_45[63] , 
        \wPDiag_45[62] , \wPDiag_45[61] , \wPDiag_45[60] , \wPDiag_45[59] , 
        \wPDiag_45[58] , \wPDiag_45[57] , \wPDiag_45[56] , \wPDiag_45[55] , 
        \wPDiag_45[54] , \wPDiag_45[53] , \wPDiag_45[52] , \wPDiag_45[51] , 
        \wPDiag_45[50] , \wPDiag_45[49] , \wPDiag_45[48] , \wPDiag_45[47] , 
        \wPDiag_45[46] , \wPDiag_45[45] , \wPDiag_45[44] , \wPDiag_45[43] , 
        \wPDiag_45[42] , \wPDiag_45[41] , \wPDiag_45[40] , \wPDiag_45[39] , 
        \wPDiag_45[38] , \wPDiag_45[37] , \wPDiag_45[36] , \wPDiag_45[35] , 
        \wPDiag_45[34] , \wPDiag_45[33] , \wPDiag_45[32] , \wPDiag_45[31] , 
        \wPDiag_45[30] , \wPDiag_45[29] , \wPDiag_45[28] , \wPDiag_45[27] , 
        \wPDiag_45[26] , \wPDiag_45[25] , \wPDiag_45[24] , \wPDiag_45[23] , 
        \wPDiag_45[22] , \wPDiag_45[21] , \wPDiag_45[20] , \wPDiag_45[19] , 
        \wPDiag_45[18] , \wPDiag_45[17] , \wPDiag_45[16] , \wPDiag_45[15] , 
        \wPDiag_45[14] , \wPDiag_45[13] , \wPDiag_45[12] , \wPDiag_45[11] , 
        \wPDiag_45[10] , \wPDiag_45[9] , \wPDiag_45[8] , \wPDiag_45[7] , 
        \wPDiag_45[6] , \wPDiag_45[5] , \wPDiag_45[4] , \wPDiag_45[3] , 
        \wPDiag_45[2] , \wPDiag_45[1] , \wPDiag_45[0] }), .NDiagOut({
        \wNDiag_45[63] , \wNDiag_45[62] , \wNDiag_45[61] , \wNDiag_45[60] , 
        \wNDiag_45[59] , \wNDiag_45[58] , \wNDiag_45[57] , \wNDiag_45[56] , 
        \wNDiag_45[55] , \wNDiag_45[54] , \wNDiag_45[53] , \wNDiag_45[52] , 
        \wNDiag_45[51] , \wNDiag_45[50] , \wNDiag_45[49] , \wNDiag_45[48] , 
        \wNDiag_45[47] , \wNDiag_45[46] , \wNDiag_45[45] , \wNDiag_45[44] , 
        \wNDiag_45[43] , \wNDiag_45[42] , \wNDiag_45[41] , \wNDiag_45[40] , 
        \wNDiag_45[39] , \wNDiag_45[38] , \wNDiag_45[37] , \wNDiag_45[36] , 
        \wNDiag_45[35] , \wNDiag_45[34] , \wNDiag_45[33] , \wNDiag_45[32] , 
        \wNDiag_45[31] , \wNDiag_45[30] , \wNDiag_45[29] , \wNDiag_45[28] , 
        \wNDiag_45[27] , \wNDiag_45[26] , \wNDiag_45[25] , \wNDiag_45[24] , 
        \wNDiag_45[23] , \wNDiag_45[22] , \wNDiag_45[21] , \wNDiag_45[20] , 
        \wNDiag_45[19] , \wNDiag_45[18] , \wNDiag_45[17] , \wNDiag_45[16] , 
        \wNDiag_45[15] , \wNDiag_45[14] , \wNDiag_45[13] , \wNDiag_45[12] , 
        \wNDiag_45[11] , \wNDiag_45[10] , \wNDiag_45[9] , \wNDiag_45[8] , 
        \wNDiag_45[7] , \wNDiag_45[6] , \wNDiag_45[5] , \wNDiag_45[4] , 
        \wNDiag_45[3] , \wNDiag_45[2] , \wNDiag_45[1] , \wNDiag_45[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_63 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_64[6] , \wScan_64[5] , \wScan_64[4] , 
        \wScan_64[3] , \wScan_64[2] , \wScan_64[1] , \wScan_64[0] }), 
        .ScanOut({\wScan_63[6] , \wScan_63[5] , \wScan_63[4] , \wScan_63[3] , 
        \wScan_63[2] , \wScan_63[1] , \wScan_63[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_63[0] ), .ReturnIn(1'b0), .ColIn({\wColumn_63[63] , 
        \wColumn_63[62] , \wColumn_63[61] , \wColumn_63[60] , \wColumn_63[59] , 
        \wColumn_63[58] , \wColumn_63[57] , \wColumn_63[56] , \wColumn_63[55] , 
        \wColumn_63[54] , \wColumn_63[53] , \wColumn_63[52] , \wColumn_63[51] , 
        \wColumn_63[50] , \wColumn_63[49] , \wColumn_63[48] , \wColumn_63[47] , 
        \wColumn_63[46] , \wColumn_63[45] , \wColumn_63[44] , \wColumn_63[43] , 
        \wColumn_63[42] , \wColumn_63[41] , \wColumn_63[40] , \wColumn_63[39] , 
        \wColumn_63[38] , \wColumn_63[37] , \wColumn_63[36] , \wColumn_63[35] , 
        \wColumn_63[34] , \wColumn_63[33] , \wColumn_63[32] , \wColumn_63[31] , 
        \wColumn_63[30] , \wColumn_63[29] , \wColumn_63[28] , \wColumn_63[27] , 
        \wColumn_63[26] , \wColumn_63[25] , \wColumn_63[24] , \wColumn_63[23] , 
        \wColumn_63[22] , \wColumn_63[21] , \wColumn_63[20] , \wColumn_63[19] , 
        \wColumn_63[18] , \wColumn_63[17] , \wColumn_63[16] , \wColumn_63[15] , 
        \wColumn_63[14] , \wColumn_63[13] , \wColumn_63[12] , \wColumn_63[11] , 
        \wColumn_63[10] , \wColumn_63[9] , \wColumn_63[8] , \wColumn_63[7] , 
        \wColumn_63[6] , \wColumn_63[5] , \wColumn_63[4] , \wColumn_63[3] , 
        \wColumn_63[2] , \wColumn_63[1] , \wColumn_63[0] }), .PDiagIn({
        \wPDiag_63[63] , \wPDiag_63[62] , \wPDiag_63[61] , \wPDiag_63[60] , 
        \wPDiag_63[59] , \wPDiag_63[58] , \wPDiag_63[57] , \wPDiag_63[56] , 
        \wPDiag_63[55] , \wPDiag_63[54] , \wPDiag_63[53] , \wPDiag_63[52] , 
        \wPDiag_63[51] , \wPDiag_63[50] , \wPDiag_63[49] , \wPDiag_63[48] , 
        \wPDiag_63[47] , \wPDiag_63[46] , \wPDiag_63[45] , \wPDiag_63[44] , 
        \wPDiag_63[43] , \wPDiag_63[42] , \wPDiag_63[41] , \wPDiag_63[40] , 
        \wPDiag_63[39] , \wPDiag_63[38] , \wPDiag_63[37] , \wPDiag_63[36] , 
        \wPDiag_63[35] , \wPDiag_63[34] , \wPDiag_63[33] , \wPDiag_63[32] , 
        \wPDiag_63[31] , \wPDiag_63[30] , \wPDiag_63[29] , \wPDiag_63[28] , 
        \wPDiag_63[27] , \wPDiag_63[26] , \wPDiag_63[25] , \wPDiag_63[24] , 
        \wPDiag_63[23] , \wPDiag_63[22] , \wPDiag_63[21] , \wPDiag_63[20] , 
        \wPDiag_63[19] , \wPDiag_63[18] , \wPDiag_63[17] , \wPDiag_63[16] , 
        \wPDiag_63[15] , \wPDiag_63[14] , \wPDiag_63[13] , \wPDiag_63[12] , 
        \wPDiag_63[11] , \wPDiag_63[10] , \wPDiag_63[9] , \wPDiag_63[8] , 
        \wPDiag_63[7] , \wPDiag_63[6] , \wPDiag_63[5] , \wPDiag_63[4] , 
        \wPDiag_63[3] , \wPDiag_63[2] , \wPDiag_63[1] , \wPDiag_63[0] }), 
        .NDiagIn({\wNDiag_63[63] , \wNDiag_63[62] , \wNDiag_63[61] , 
        \wNDiag_63[60] , \wNDiag_63[59] , \wNDiag_63[58] , \wNDiag_63[57] , 
        \wNDiag_63[56] , \wNDiag_63[55] , \wNDiag_63[54] , \wNDiag_63[53] , 
        \wNDiag_63[52] , \wNDiag_63[51] , \wNDiag_63[50] , \wNDiag_63[49] , 
        \wNDiag_63[48] , \wNDiag_63[47] , \wNDiag_63[46] , \wNDiag_63[45] , 
        \wNDiag_63[44] , \wNDiag_63[43] , \wNDiag_63[42] , \wNDiag_63[41] , 
        \wNDiag_63[40] , \wNDiag_63[39] , \wNDiag_63[38] , \wNDiag_63[37] , 
        \wNDiag_63[36] , \wNDiag_63[35] , \wNDiag_63[34] , \wNDiag_63[33] , 
        \wNDiag_63[32] , \wNDiag_63[31] , \wNDiag_63[30] , \wNDiag_63[29] , 
        \wNDiag_63[28] , \wNDiag_63[27] , \wNDiag_63[26] , \wNDiag_63[25] , 
        \wNDiag_63[24] , \wNDiag_63[23] , \wNDiag_63[22] , \wNDiag_63[21] , 
        \wNDiag_63[20] , \wNDiag_63[19] , \wNDiag_63[18] , \wNDiag_63[17] , 
        \wNDiag_63[16] , \wNDiag_63[15] , \wNDiag_63[14] , \wNDiag_63[13] , 
        \wNDiag_63[12] , \wNDiag_63[11] , \wNDiag_63[10] , \wNDiag_63[9] , 
        \wNDiag_63[8] , \wNDiag_63[7] , \wNDiag_63[6] , \wNDiag_63[5] , 
        \wNDiag_63[4] , \wNDiag_63[3] , \wNDiag_63[2] , \wNDiag_63[1] , 
        \wNDiag_63[0] }), .CallOut(\wCall_64[0] ), .ReturnOut(\wReturn_63[0] )
         );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_57 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_58[6] , \wScan_58[5] , \wScan_58[4] , 
        \wScan_58[3] , \wScan_58[2] , \wScan_58[1] , \wScan_58[0] }), 
        .ScanOut({\wScan_57[6] , \wScan_57[5] , \wScan_57[4] , \wScan_57[3] , 
        \wScan_57[2] , \wScan_57[1] , \wScan_57[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_57[0] ), .ReturnIn(\wReturn_58[0] ), .ColIn({
        \wColumn_57[63] , \wColumn_57[62] , \wColumn_57[61] , \wColumn_57[60] , 
        \wColumn_57[59] , \wColumn_57[58] , \wColumn_57[57] , \wColumn_57[56] , 
        \wColumn_57[55] , \wColumn_57[54] , \wColumn_57[53] , \wColumn_57[52] , 
        \wColumn_57[51] , \wColumn_57[50] , \wColumn_57[49] , \wColumn_57[48] , 
        \wColumn_57[47] , \wColumn_57[46] , \wColumn_57[45] , \wColumn_57[44] , 
        \wColumn_57[43] , \wColumn_57[42] , \wColumn_57[41] , \wColumn_57[40] , 
        \wColumn_57[39] , \wColumn_57[38] , \wColumn_57[37] , \wColumn_57[36] , 
        \wColumn_57[35] , \wColumn_57[34] , \wColumn_57[33] , \wColumn_57[32] , 
        \wColumn_57[31] , \wColumn_57[30] , \wColumn_57[29] , \wColumn_57[28] , 
        \wColumn_57[27] , \wColumn_57[26] , \wColumn_57[25] , \wColumn_57[24] , 
        \wColumn_57[23] , \wColumn_57[22] , \wColumn_57[21] , \wColumn_57[20] , 
        \wColumn_57[19] , \wColumn_57[18] , \wColumn_57[17] , \wColumn_57[16] , 
        \wColumn_57[15] , \wColumn_57[14] , \wColumn_57[13] , \wColumn_57[12] , 
        \wColumn_57[11] , \wColumn_57[10] , \wColumn_57[9] , \wColumn_57[8] , 
        \wColumn_57[7] , \wColumn_57[6] , \wColumn_57[5] , \wColumn_57[4] , 
        \wColumn_57[3] , \wColumn_57[2] , \wColumn_57[1] , \wColumn_57[0] }), 
        .PDiagIn({\wPDiag_57[63] , \wPDiag_57[62] , \wPDiag_57[61] , 
        \wPDiag_57[60] , \wPDiag_57[59] , \wPDiag_57[58] , \wPDiag_57[57] , 
        \wPDiag_57[56] , \wPDiag_57[55] , \wPDiag_57[54] , \wPDiag_57[53] , 
        \wPDiag_57[52] , \wPDiag_57[51] , \wPDiag_57[50] , \wPDiag_57[49] , 
        \wPDiag_57[48] , \wPDiag_57[47] , \wPDiag_57[46] , \wPDiag_57[45] , 
        \wPDiag_57[44] , \wPDiag_57[43] , \wPDiag_57[42] , \wPDiag_57[41] , 
        \wPDiag_57[40] , \wPDiag_57[39] , \wPDiag_57[38] , \wPDiag_57[37] , 
        \wPDiag_57[36] , \wPDiag_57[35] , \wPDiag_57[34] , \wPDiag_57[33] , 
        \wPDiag_57[32] , \wPDiag_57[31] , \wPDiag_57[30] , \wPDiag_57[29] , 
        \wPDiag_57[28] , \wPDiag_57[27] , \wPDiag_57[26] , \wPDiag_57[25] , 
        \wPDiag_57[24] , \wPDiag_57[23] , \wPDiag_57[22] , \wPDiag_57[21] , 
        \wPDiag_57[20] , \wPDiag_57[19] , \wPDiag_57[18] , \wPDiag_57[17] , 
        \wPDiag_57[16] , \wPDiag_57[15] , \wPDiag_57[14] , \wPDiag_57[13] , 
        \wPDiag_57[12] , \wPDiag_57[11] , \wPDiag_57[10] , \wPDiag_57[9] , 
        \wPDiag_57[8] , \wPDiag_57[7] , \wPDiag_57[6] , \wPDiag_57[5] , 
        \wPDiag_57[4] , \wPDiag_57[3] , \wPDiag_57[2] , \wPDiag_57[1] , 
        \wPDiag_57[0] }), .NDiagIn({\wNDiag_57[63] , \wNDiag_57[62] , 
        \wNDiag_57[61] , \wNDiag_57[60] , \wNDiag_57[59] , \wNDiag_57[58] , 
        \wNDiag_57[57] , \wNDiag_57[56] , \wNDiag_57[55] , \wNDiag_57[54] , 
        \wNDiag_57[53] , \wNDiag_57[52] , \wNDiag_57[51] , \wNDiag_57[50] , 
        \wNDiag_57[49] , \wNDiag_57[48] , \wNDiag_57[47] , \wNDiag_57[46] , 
        \wNDiag_57[45] , \wNDiag_57[44] , \wNDiag_57[43] , \wNDiag_57[42] , 
        \wNDiag_57[41] , \wNDiag_57[40] , \wNDiag_57[39] , \wNDiag_57[38] , 
        \wNDiag_57[37] , \wNDiag_57[36] , \wNDiag_57[35] , \wNDiag_57[34] , 
        \wNDiag_57[33] , \wNDiag_57[32] , \wNDiag_57[31] , \wNDiag_57[30] , 
        \wNDiag_57[29] , \wNDiag_57[28] , \wNDiag_57[27] , \wNDiag_57[26] , 
        \wNDiag_57[25] , \wNDiag_57[24] , \wNDiag_57[23] , \wNDiag_57[22] , 
        \wNDiag_57[21] , \wNDiag_57[20] , \wNDiag_57[19] , \wNDiag_57[18] , 
        \wNDiag_57[17] , \wNDiag_57[16] , \wNDiag_57[15] , \wNDiag_57[14] , 
        \wNDiag_57[13] , \wNDiag_57[12] , \wNDiag_57[11] , \wNDiag_57[10] , 
        \wNDiag_57[9] , \wNDiag_57[8] , \wNDiag_57[7] , \wNDiag_57[6] , 
        \wNDiag_57[5] , \wNDiag_57[4] , \wNDiag_57[3] , \wNDiag_57[2] , 
        \wNDiag_57[1] , \wNDiag_57[0] }), .CallOut(\wCall_58[0] ), .ReturnOut(
        \wReturn_57[0] ), .ColOut({\wColumn_58[63] , \wColumn_58[62] , 
        \wColumn_58[61] , \wColumn_58[60] , \wColumn_58[59] , \wColumn_58[58] , 
        \wColumn_58[57] , \wColumn_58[56] , \wColumn_58[55] , \wColumn_58[54] , 
        \wColumn_58[53] , \wColumn_58[52] , \wColumn_58[51] , \wColumn_58[50] , 
        \wColumn_58[49] , \wColumn_58[48] , \wColumn_58[47] , \wColumn_58[46] , 
        \wColumn_58[45] , \wColumn_58[44] , \wColumn_58[43] , \wColumn_58[42] , 
        \wColumn_58[41] , \wColumn_58[40] , \wColumn_58[39] , \wColumn_58[38] , 
        \wColumn_58[37] , \wColumn_58[36] , \wColumn_58[35] , \wColumn_58[34] , 
        \wColumn_58[33] , \wColumn_58[32] , \wColumn_58[31] , \wColumn_58[30] , 
        \wColumn_58[29] , \wColumn_58[28] , \wColumn_58[27] , \wColumn_58[26] , 
        \wColumn_58[25] , \wColumn_58[24] , \wColumn_58[23] , \wColumn_58[22] , 
        \wColumn_58[21] , \wColumn_58[20] , \wColumn_58[19] , \wColumn_58[18] , 
        \wColumn_58[17] , \wColumn_58[16] , \wColumn_58[15] , \wColumn_58[14] , 
        \wColumn_58[13] , \wColumn_58[12] , \wColumn_58[11] , \wColumn_58[10] , 
        \wColumn_58[9] , \wColumn_58[8] , \wColumn_58[7] , \wColumn_58[6] , 
        \wColumn_58[5] , \wColumn_58[4] , \wColumn_58[3] , \wColumn_58[2] , 
        \wColumn_58[1] , \wColumn_58[0] }), .PDiagOut({\wPDiag_58[63] , 
        \wPDiag_58[62] , \wPDiag_58[61] , \wPDiag_58[60] , \wPDiag_58[59] , 
        \wPDiag_58[58] , \wPDiag_58[57] , \wPDiag_58[56] , \wPDiag_58[55] , 
        \wPDiag_58[54] , \wPDiag_58[53] , \wPDiag_58[52] , \wPDiag_58[51] , 
        \wPDiag_58[50] , \wPDiag_58[49] , \wPDiag_58[48] , \wPDiag_58[47] , 
        \wPDiag_58[46] , \wPDiag_58[45] , \wPDiag_58[44] , \wPDiag_58[43] , 
        \wPDiag_58[42] , \wPDiag_58[41] , \wPDiag_58[40] , \wPDiag_58[39] , 
        \wPDiag_58[38] , \wPDiag_58[37] , \wPDiag_58[36] , \wPDiag_58[35] , 
        \wPDiag_58[34] , \wPDiag_58[33] , \wPDiag_58[32] , \wPDiag_58[31] , 
        \wPDiag_58[30] , \wPDiag_58[29] , \wPDiag_58[28] , \wPDiag_58[27] , 
        \wPDiag_58[26] , \wPDiag_58[25] , \wPDiag_58[24] , \wPDiag_58[23] , 
        \wPDiag_58[22] , \wPDiag_58[21] , \wPDiag_58[20] , \wPDiag_58[19] , 
        \wPDiag_58[18] , \wPDiag_58[17] , \wPDiag_58[16] , \wPDiag_58[15] , 
        \wPDiag_58[14] , \wPDiag_58[13] , \wPDiag_58[12] , \wPDiag_58[11] , 
        \wPDiag_58[10] , \wPDiag_58[9] , \wPDiag_58[8] , \wPDiag_58[7] , 
        \wPDiag_58[6] , \wPDiag_58[5] , \wPDiag_58[4] , \wPDiag_58[3] , 
        \wPDiag_58[2] , \wPDiag_58[1] , \wPDiag_58[0] }), .NDiagOut({
        \wNDiag_58[63] , \wNDiag_58[62] , \wNDiag_58[61] , \wNDiag_58[60] , 
        \wNDiag_58[59] , \wNDiag_58[58] , \wNDiag_58[57] , \wNDiag_58[56] , 
        \wNDiag_58[55] , \wNDiag_58[54] , \wNDiag_58[53] , \wNDiag_58[52] , 
        \wNDiag_58[51] , \wNDiag_58[50] , \wNDiag_58[49] , \wNDiag_58[48] , 
        \wNDiag_58[47] , \wNDiag_58[46] , \wNDiag_58[45] , \wNDiag_58[44] , 
        \wNDiag_58[43] , \wNDiag_58[42] , \wNDiag_58[41] , \wNDiag_58[40] , 
        \wNDiag_58[39] , \wNDiag_58[38] , \wNDiag_58[37] , \wNDiag_58[36] , 
        \wNDiag_58[35] , \wNDiag_58[34] , \wNDiag_58[33] , \wNDiag_58[32] , 
        \wNDiag_58[31] , \wNDiag_58[30] , \wNDiag_58[29] , \wNDiag_58[28] , 
        \wNDiag_58[27] , \wNDiag_58[26] , \wNDiag_58[25] , \wNDiag_58[24] , 
        \wNDiag_58[23] , \wNDiag_58[22] , \wNDiag_58[21] , \wNDiag_58[20] , 
        \wNDiag_58[19] , \wNDiag_58[18] , \wNDiag_58[17] , \wNDiag_58[16] , 
        \wNDiag_58[15] , \wNDiag_58[14] , \wNDiag_58[13] , \wNDiag_58[12] , 
        \wNDiag_58[11] , \wNDiag_58[10] , \wNDiag_58[9] , \wNDiag_58[8] , 
        \wNDiag_58[7] , \wNDiag_58[6] , \wNDiag_58[5] , \wNDiag_58[4] , 
        \wNDiag_58[3] , \wNDiag_58[2] , \wNDiag_58[1] , \wNDiag_58[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_8 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_9[6] , \wScan_9[5] , \wScan_9[4] , 
        \wScan_9[3] , \wScan_9[2] , \wScan_9[1] , \wScan_9[0] }), .ScanOut({
        \wScan_8[6] , \wScan_8[5] , \wScan_8[4] , \wScan_8[3] , \wScan_8[2] , 
        \wScan_8[1] , \wScan_8[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_8[0] ), 
        .ReturnIn(\wReturn_9[0] ), .ColIn({\wColumn_8[63] , \wColumn_8[62] , 
        \wColumn_8[61] , \wColumn_8[60] , \wColumn_8[59] , \wColumn_8[58] , 
        \wColumn_8[57] , \wColumn_8[56] , \wColumn_8[55] , \wColumn_8[54] , 
        \wColumn_8[53] , \wColumn_8[52] , \wColumn_8[51] , \wColumn_8[50] , 
        \wColumn_8[49] , \wColumn_8[48] , \wColumn_8[47] , \wColumn_8[46] , 
        \wColumn_8[45] , \wColumn_8[44] , \wColumn_8[43] , \wColumn_8[42] , 
        \wColumn_8[41] , \wColumn_8[40] , \wColumn_8[39] , \wColumn_8[38] , 
        \wColumn_8[37] , \wColumn_8[36] , \wColumn_8[35] , \wColumn_8[34] , 
        \wColumn_8[33] , \wColumn_8[32] , \wColumn_8[31] , \wColumn_8[30] , 
        \wColumn_8[29] , \wColumn_8[28] , \wColumn_8[27] , \wColumn_8[26] , 
        \wColumn_8[25] , \wColumn_8[24] , \wColumn_8[23] , \wColumn_8[22] , 
        \wColumn_8[21] , \wColumn_8[20] , \wColumn_8[19] , \wColumn_8[18] , 
        \wColumn_8[17] , \wColumn_8[16] , \wColumn_8[15] , \wColumn_8[14] , 
        \wColumn_8[13] , \wColumn_8[12] , \wColumn_8[11] , \wColumn_8[10] , 
        \wColumn_8[9] , \wColumn_8[8] , \wColumn_8[7] , \wColumn_8[6] , 
        \wColumn_8[5] , \wColumn_8[4] , \wColumn_8[3] , \wColumn_8[2] , 
        \wColumn_8[1] , \wColumn_8[0] }), .PDiagIn({\wPDiag_8[63] , 
        \wPDiag_8[62] , \wPDiag_8[61] , \wPDiag_8[60] , \wPDiag_8[59] , 
        \wPDiag_8[58] , \wPDiag_8[57] , \wPDiag_8[56] , \wPDiag_8[55] , 
        \wPDiag_8[54] , \wPDiag_8[53] , \wPDiag_8[52] , \wPDiag_8[51] , 
        \wPDiag_8[50] , \wPDiag_8[49] , \wPDiag_8[48] , \wPDiag_8[47] , 
        \wPDiag_8[46] , \wPDiag_8[45] , \wPDiag_8[44] , \wPDiag_8[43] , 
        \wPDiag_8[42] , \wPDiag_8[41] , \wPDiag_8[40] , \wPDiag_8[39] , 
        \wPDiag_8[38] , \wPDiag_8[37] , \wPDiag_8[36] , \wPDiag_8[35] , 
        \wPDiag_8[34] , \wPDiag_8[33] , \wPDiag_8[32] , \wPDiag_8[31] , 
        \wPDiag_8[30] , \wPDiag_8[29] , \wPDiag_8[28] , \wPDiag_8[27] , 
        \wPDiag_8[26] , \wPDiag_8[25] , \wPDiag_8[24] , \wPDiag_8[23] , 
        \wPDiag_8[22] , \wPDiag_8[21] , \wPDiag_8[20] , \wPDiag_8[19] , 
        \wPDiag_8[18] , \wPDiag_8[17] , \wPDiag_8[16] , \wPDiag_8[15] , 
        \wPDiag_8[14] , \wPDiag_8[13] , \wPDiag_8[12] , \wPDiag_8[11] , 
        \wPDiag_8[10] , \wPDiag_8[9] , \wPDiag_8[8] , \wPDiag_8[7] , 
        \wPDiag_8[6] , \wPDiag_8[5] , \wPDiag_8[4] , \wPDiag_8[3] , 
        \wPDiag_8[2] , \wPDiag_8[1] , \wPDiag_8[0] }), .NDiagIn({
        \wNDiag_8[63] , \wNDiag_8[62] , \wNDiag_8[61] , \wNDiag_8[60] , 
        \wNDiag_8[59] , \wNDiag_8[58] , \wNDiag_8[57] , \wNDiag_8[56] , 
        \wNDiag_8[55] , \wNDiag_8[54] , \wNDiag_8[53] , \wNDiag_8[52] , 
        \wNDiag_8[51] , \wNDiag_8[50] , \wNDiag_8[49] , \wNDiag_8[48] , 
        \wNDiag_8[47] , \wNDiag_8[46] , \wNDiag_8[45] , \wNDiag_8[44] , 
        \wNDiag_8[43] , \wNDiag_8[42] , \wNDiag_8[41] , \wNDiag_8[40] , 
        \wNDiag_8[39] , \wNDiag_8[38] , \wNDiag_8[37] , \wNDiag_8[36] , 
        \wNDiag_8[35] , \wNDiag_8[34] , \wNDiag_8[33] , \wNDiag_8[32] , 
        \wNDiag_8[31] , \wNDiag_8[30] , \wNDiag_8[29] , \wNDiag_8[28] , 
        \wNDiag_8[27] , \wNDiag_8[26] , \wNDiag_8[25] , \wNDiag_8[24] , 
        \wNDiag_8[23] , \wNDiag_8[22] , \wNDiag_8[21] , \wNDiag_8[20] , 
        \wNDiag_8[19] , \wNDiag_8[18] , \wNDiag_8[17] , \wNDiag_8[16] , 
        \wNDiag_8[15] , \wNDiag_8[14] , \wNDiag_8[13] , \wNDiag_8[12] , 
        \wNDiag_8[11] , \wNDiag_8[10] , \wNDiag_8[9] , \wNDiag_8[8] , 
        \wNDiag_8[7] , \wNDiag_8[6] , \wNDiag_8[5] , \wNDiag_8[4] , 
        \wNDiag_8[3] , \wNDiag_8[2] , \wNDiag_8[1] , \wNDiag_8[0] }), 
        .CallOut(\wCall_9[0] ), .ReturnOut(\wReturn_8[0] ), .ColOut({
        \wColumn_9[63] , \wColumn_9[62] , \wColumn_9[61] , \wColumn_9[60] , 
        \wColumn_9[59] , \wColumn_9[58] , \wColumn_9[57] , \wColumn_9[56] , 
        \wColumn_9[55] , \wColumn_9[54] , \wColumn_9[53] , \wColumn_9[52] , 
        \wColumn_9[51] , \wColumn_9[50] , \wColumn_9[49] , \wColumn_9[48] , 
        \wColumn_9[47] , \wColumn_9[46] , \wColumn_9[45] , \wColumn_9[44] , 
        \wColumn_9[43] , \wColumn_9[42] , \wColumn_9[41] , \wColumn_9[40] , 
        \wColumn_9[39] , \wColumn_9[38] , \wColumn_9[37] , \wColumn_9[36] , 
        \wColumn_9[35] , \wColumn_9[34] , \wColumn_9[33] , \wColumn_9[32] , 
        \wColumn_9[31] , \wColumn_9[30] , \wColumn_9[29] , \wColumn_9[28] , 
        \wColumn_9[27] , \wColumn_9[26] , \wColumn_9[25] , \wColumn_9[24] , 
        \wColumn_9[23] , \wColumn_9[22] , \wColumn_9[21] , \wColumn_9[20] , 
        \wColumn_9[19] , \wColumn_9[18] , \wColumn_9[17] , \wColumn_9[16] , 
        \wColumn_9[15] , \wColumn_9[14] , \wColumn_9[13] , \wColumn_9[12] , 
        \wColumn_9[11] , \wColumn_9[10] , \wColumn_9[9] , \wColumn_9[8] , 
        \wColumn_9[7] , \wColumn_9[6] , \wColumn_9[5] , \wColumn_9[4] , 
        \wColumn_9[3] , \wColumn_9[2] , \wColumn_9[1] , \wColumn_9[0] }), 
        .PDiagOut({\wPDiag_9[63] , \wPDiag_9[62] , \wPDiag_9[61] , 
        \wPDiag_9[60] , \wPDiag_9[59] , \wPDiag_9[58] , \wPDiag_9[57] , 
        \wPDiag_9[56] , \wPDiag_9[55] , \wPDiag_9[54] , \wPDiag_9[53] , 
        \wPDiag_9[52] , \wPDiag_9[51] , \wPDiag_9[50] , \wPDiag_9[49] , 
        \wPDiag_9[48] , \wPDiag_9[47] , \wPDiag_9[46] , \wPDiag_9[45] , 
        \wPDiag_9[44] , \wPDiag_9[43] , \wPDiag_9[42] , \wPDiag_9[41] , 
        \wPDiag_9[40] , \wPDiag_9[39] , \wPDiag_9[38] , \wPDiag_9[37] , 
        \wPDiag_9[36] , \wPDiag_9[35] , \wPDiag_9[34] , \wPDiag_9[33] , 
        \wPDiag_9[32] , \wPDiag_9[31] , \wPDiag_9[30] , \wPDiag_9[29] , 
        \wPDiag_9[28] , \wPDiag_9[27] , \wPDiag_9[26] , \wPDiag_9[25] , 
        \wPDiag_9[24] , \wPDiag_9[23] , \wPDiag_9[22] , \wPDiag_9[21] , 
        \wPDiag_9[20] , \wPDiag_9[19] , \wPDiag_9[18] , \wPDiag_9[17] , 
        \wPDiag_9[16] , \wPDiag_9[15] , \wPDiag_9[14] , \wPDiag_9[13] , 
        \wPDiag_9[12] , \wPDiag_9[11] , \wPDiag_9[10] , \wPDiag_9[9] , 
        \wPDiag_9[8] , \wPDiag_9[7] , \wPDiag_9[6] , \wPDiag_9[5] , 
        \wPDiag_9[4] , \wPDiag_9[3] , \wPDiag_9[2] , \wPDiag_9[1] , 
        \wPDiag_9[0] }), .NDiagOut({\wNDiag_9[63] , \wNDiag_9[62] , 
        \wNDiag_9[61] , \wNDiag_9[60] , \wNDiag_9[59] , \wNDiag_9[58] , 
        \wNDiag_9[57] , \wNDiag_9[56] , \wNDiag_9[55] , \wNDiag_9[54] , 
        \wNDiag_9[53] , \wNDiag_9[52] , \wNDiag_9[51] , \wNDiag_9[50] , 
        \wNDiag_9[49] , \wNDiag_9[48] , \wNDiag_9[47] , \wNDiag_9[46] , 
        \wNDiag_9[45] , \wNDiag_9[44] , \wNDiag_9[43] , \wNDiag_9[42] , 
        \wNDiag_9[41] , \wNDiag_9[40] , \wNDiag_9[39] , \wNDiag_9[38] , 
        \wNDiag_9[37] , \wNDiag_9[36] , \wNDiag_9[35] , \wNDiag_9[34] , 
        \wNDiag_9[33] , \wNDiag_9[32] , \wNDiag_9[31] , \wNDiag_9[30] , 
        \wNDiag_9[29] , \wNDiag_9[28] , \wNDiag_9[27] , \wNDiag_9[26] , 
        \wNDiag_9[25] , \wNDiag_9[24] , \wNDiag_9[23] , \wNDiag_9[22] , 
        \wNDiag_9[21] , \wNDiag_9[20] , \wNDiag_9[19] , \wNDiag_9[18] , 
        \wNDiag_9[17] , \wNDiag_9[16] , \wNDiag_9[15] , \wNDiag_9[14] , 
        \wNDiag_9[13] , \wNDiag_9[12] , \wNDiag_9[11] , \wNDiag_9[10] , 
        \wNDiag_9[9] , \wNDiag_9[8] , \wNDiag_9[7] , \wNDiag_9[6] , 
        \wNDiag_9[5] , \wNDiag_9[4] , \wNDiag_9[3] , \wNDiag_9[2] , 
        \wNDiag_9[1] , \wNDiag_9[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_10 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_11[6] , \wScan_11[5] , \wScan_11[4] , 
        \wScan_11[3] , \wScan_11[2] , \wScan_11[1] , \wScan_11[0] }), 
        .ScanOut({\wScan_10[6] , \wScan_10[5] , \wScan_10[4] , \wScan_10[3] , 
        \wScan_10[2] , \wScan_10[1] , \wScan_10[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_10[0] ), .ReturnIn(\wReturn_11[0] ), .ColIn({
        \wColumn_10[63] , \wColumn_10[62] , \wColumn_10[61] , \wColumn_10[60] , 
        \wColumn_10[59] , \wColumn_10[58] , \wColumn_10[57] , \wColumn_10[56] , 
        \wColumn_10[55] , \wColumn_10[54] , \wColumn_10[53] , \wColumn_10[52] , 
        \wColumn_10[51] , \wColumn_10[50] , \wColumn_10[49] , \wColumn_10[48] , 
        \wColumn_10[47] , \wColumn_10[46] , \wColumn_10[45] , \wColumn_10[44] , 
        \wColumn_10[43] , \wColumn_10[42] , \wColumn_10[41] , \wColumn_10[40] , 
        \wColumn_10[39] , \wColumn_10[38] , \wColumn_10[37] , \wColumn_10[36] , 
        \wColumn_10[35] , \wColumn_10[34] , \wColumn_10[33] , \wColumn_10[32] , 
        \wColumn_10[31] , \wColumn_10[30] , \wColumn_10[29] , \wColumn_10[28] , 
        \wColumn_10[27] , \wColumn_10[26] , \wColumn_10[25] , \wColumn_10[24] , 
        \wColumn_10[23] , \wColumn_10[22] , \wColumn_10[21] , \wColumn_10[20] , 
        \wColumn_10[19] , \wColumn_10[18] , \wColumn_10[17] , \wColumn_10[16] , 
        \wColumn_10[15] , \wColumn_10[14] , \wColumn_10[13] , \wColumn_10[12] , 
        \wColumn_10[11] , \wColumn_10[10] , \wColumn_10[9] , \wColumn_10[8] , 
        \wColumn_10[7] , \wColumn_10[6] , \wColumn_10[5] , \wColumn_10[4] , 
        \wColumn_10[3] , \wColumn_10[2] , \wColumn_10[1] , \wColumn_10[0] }), 
        .PDiagIn({\wPDiag_10[63] , \wPDiag_10[62] , \wPDiag_10[61] , 
        \wPDiag_10[60] , \wPDiag_10[59] , \wPDiag_10[58] , \wPDiag_10[57] , 
        \wPDiag_10[56] , \wPDiag_10[55] , \wPDiag_10[54] , \wPDiag_10[53] , 
        \wPDiag_10[52] , \wPDiag_10[51] , \wPDiag_10[50] , \wPDiag_10[49] , 
        \wPDiag_10[48] , \wPDiag_10[47] , \wPDiag_10[46] , \wPDiag_10[45] , 
        \wPDiag_10[44] , \wPDiag_10[43] , \wPDiag_10[42] , \wPDiag_10[41] , 
        \wPDiag_10[40] , \wPDiag_10[39] , \wPDiag_10[38] , \wPDiag_10[37] , 
        \wPDiag_10[36] , \wPDiag_10[35] , \wPDiag_10[34] , \wPDiag_10[33] , 
        \wPDiag_10[32] , \wPDiag_10[31] , \wPDiag_10[30] , \wPDiag_10[29] , 
        \wPDiag_10[28] , \wPDiag_10[27] , \wPDiag_10[26] , \wPDiag_10[25] , 
        \wPDiag_10[24] , \wPDiag_10[23] , \wPDiag_10[22] , \wPDiag_10[21] , 
        \wPDiag_10[20] , \wPDiag_10[19] , \wPDiag_10[18] , \wPDiag_10[17] , 
        \wPDiag_10[16] , \wPDiag_10[15] , \wPDiag_10[14] , \wPDiag_10[13] , 
        \wPDiag_10[12] , \wPDiag_10[11] , \wPDiag_10[10] , \wPDiag_10[9] , 
        \wPDiag_10[8] , \wPDiag_10[7] , \wPDiag_10[6] , \wPDiag_10[5] , 
        \wPDiag_10[4] , \wPDiag_10[3] , \wPDiag_10[2] , \wPDiag_10[1] , 
        \wPDiag_10[0] }), .NDiagIn({\wNDiag_10[63] , \wNDiag_10[62] , 
        \wNDiag_10[61] , \wNDiag_10[60] , \wNDiag_10[59] , \wNDiag_10[58] , 
        \wNDiag_10[57] , \wNDiag_10[56] , \wNDiag_10[55] , \wNDiag_10[54] , 
        \wNDiag_10[53] , \wNDiag_10[52] , \wNDiag_10[51] , \wNDiag_10[50] , 
        \wNDiag_10[49] , \wNDiag_10[48] , \wNDiag_10[47] , \wNDiag_10[46] , 
        \wNDiag_10[45] , \wNDiag_10[44] , \wNDiag_10[43] , \wNDiag_10[42] , 
        \wNDiag_10[41] , \wNDiag_10[40] , \wNDiag_10[39] , \wNDiag_10[38] , 
        \wNDiag_10[37] , \wNDiag_10[36] , \wNDiag_10[35] , \wNDiag_10[34] , 
        \wNDiag_10[33] , \wNDiag_10[32] , \wNDiag_10[31] , \wNDiag_10[30] , 
        \wNDiag_10[29] , \wNDiag_10[28] , \wNDiag_10[27] , \wNDiag_10[26] , 
        \wNDiag_10[25] , \wNDiag_10[24] , \wNDiag_10[23] , \wNDiag_10[22] , 
        \wNDiag_10[21] , \wNDiag_10[20] , \wNDiag_10[19] , \wNDiag_10[18] , 
        \wNDiag_10[17] , \wNDiag_10[16] , \wNDiag_10[15] , \wNDiag_10[14] , 
        \wNDiag_10[13] , \wNDiag_10[12] , \wNDiag_10[11] , \wNDiag_10[10] , 
        \wNDiag_10[9] , \wNDiag_10[8] , \wNDiag_10[7] , \wNDiag_10[6] , 
        \wNDiag_10[5] , \wNDiag_10[4] , \wNDiag_10[3] , \wNDiag_10[2] , 
        \wNDiag_10[1] , \wNDiag_10[0] }), .CallOut(\wCall_11[0] ), .ReturnOut(
        \wReturn_10[0] ), .ColOut({\wColumn_11[63] , \wColumn_11[62] , 
        \wColumn_11[61] , \wColumn_11[60] , \wColumn_11[59] , \wColumn_11[58] , 
        \wColumn_11[57] , \wColumn_11[56] , \wColumn_11[55] , \wColumn_11[54] , 
        \wColumn_11[53] , \wColumn_11[52] , \wColumn_11[51] , \wColumn_11[50] , 
        \wColumn_11[49] , \wColumn_11[48] , \wColumn_11[47] , \wColumn_11[46] , 
        \wColumn_11[45] , \wColumn_11[44] , \wColumn_11[43] , \wColumn_11[42] , 
        \wColumn_11[41] , \wColumn_11[40] , \wColumn_11[39] , \wColumn_11[38] , 
        \wColumn_11[37] , \wColumn_11[36] , \wColumn_11[35] , \wColumn_11[34] , 
        \wColumn_11[33] , \wColumn_11[32] , \wColumn_11[31] , \wColumn_11[30] , 
        \wColumn_11[29] , \wColumn_11[28] , \wColumn_11[27] , \wColumn_11[26] , 
        \wColumn_11[25] , \wColumn_11[24] , \wColumn_11[23] , \wColumn_11[22] , 
        \wColumn_11[21] , \wColumn_11[20] , \wColumn_11[19] , \wColumn_11[18] , 
        \wColumn_11[17] , \wColumn_11[16] , \wColumn_11[15] , \wColumn_11[14] , 
        \wColumn_11[13] , \wColumn_11[12] , \wColumn_11[11] , \wColumn_11[10] , 
        \wColumn_11[9] , \wColumn_11[8] , \wColumn_11[7] , \wColumn_11[6] , 
        \wColumn_11[5] , \wColumn_11[4] , \wColumn_11[3] , \wColumn_11[2] , 
        \wColumn_11[1] , \wColumn_11[0] }), .PDiagOut({\wPDiag_11[63] , 
        \wPDiag_11[62] , \wPDiag_11[61] , \wPDiag_11[60] , \wPDiag_11[59] , 
        \wPDiag_11[58] , \wPDiag_11[57] , \wPDiag_11[56] , \wPDiag_11[55] , 
        \wPDiag_11[54] , \wPDiag_11[53] , \wPDiag_11[52] , \wPDiag_11[51] , 
        \wPDiag_11[50] , \wPDiag_11[49] , \wPDiag_11[48] , \wPDiag_11[47] , 
        \wPDiag_11[46] , \wPDiag_11[45] , \wPDiag_11[44] , \wPDiag_11[43] , 
        \wPDiag_11[42] , \wPDiag_11[41] , \wPDiag_11[40] , \wPDiag_11[39] , 
        \wPDiag_11[38] , \wPDiag_11[37] , \wPDiag_11[36] , \wPDiag_11[35] , 
        \wPDiag_11[34] , \wPDiag_11[33] , \wPDiag_11[32] , \wPDiag_11[31] , 
        \wPDiag_11[30] , \wPDiag_11[29] , \wPDiag_11[28] , \wPDiag_11[27] , 
        \wPDiag_11[26] , \wPDiag_11[25] , \wPDiag_11[24] , \wPDiag_11[23] , 
        \wPDiag_11[22] , \wPDiag_11[21] , \wPDiag_11[20] , \wPDiag_11[19] , 
        \wPDiag_11[18] , \wPDiag_11[17] , \wPDiag_11[16] , \wPDiag_11[15] , 
        \wPDiag_11[14] , \wPDiag_11[13] , \wPDiag_11[12] , \wPDiag_11[11] , 
        \wPDiag_11[10] , \wPDiag_11[9] , \wPDiag_11[8] , \wPDiag_11[7] , 
        \wPDiag_11[6] , \wPDiag_11[5] , \wPDiag_11[4] , \wPDiag_11[3] , 
        \wPDiag_11[2] , \wPDiag_11[1] , \wPDiag_11[0] }), .NDiagOut({
        \wNDiag_11[63] , \wNDiag_11[62] , \wNDiag_11[61] , \wNDiag_11[60] , 
        \wNDiag_11[59] , \wNDiag_11[58] , \wNDiag_11[57] , \wNDiag_11[56] , 
        \wNDiag_11[55] , \wNDiag_11[54] , \wNDiag_11[53] , \wNDiag_11[52] , 
        \wNDiag_11[51] , \wNDiag_11[50] , \wNDiag_11[49] , \wNDiag_11[48] , 
        \wNDiag_11[47] , \wNDiag_11[46] , \wNDiag_11[45] , \wNDiag_11[44] , 
        \wNDiag_11[43] , \wNDiag_11[42] , \wNDiag_11[41] , \wNDiag_11[40] , 
        \wNDiag_11[39] , \wNDiag_11[38] , \wNDiag_11[37] , \wNDiag_11[36] , 
        \wNDiag_11[35] , \wNDiag_11[34] , \wNDiag_11[33] , \wNDiag_11[32] , 
        \wNDiag_11[31] , \wNDiag_11[30] , \wNDiag_11[29] , \wNDiag_11[28] , 
        \wNDiag_11[27] , \wNDiag_11[26] , \wNDiag_11[25] , \wNDiag_11[24] , 
        \wNDiag_11[23] , \wNDiag_11[22] , \wNDiag_11[21] , \wNDiag_11[20] , 
        \wNDiag_11[19] , \wNDiag_11[18] , \wNDiag_11[17] , \wNDiag_11[16] , 
        \wNDiag_11[15] , \wNDiag_11[14] , \wNDiag_11[13] , \wNDiag_11[12] , 
        \wNDiag_11[11] , \wNDiag_11[10] , \wNDiag_11[9] , \wNDiag_11[8] , 
        \wNDiag_11[7] , \wNDiag_11[6] , \wNDiag_11[5] , \wNDiag_11[4] , 
        \wNDiag_11[3] , \wNDiag_11[2] , \wNDiag_11[1] , \wNDiag_11[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_17 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_18[6] , \wScan_18[5] , \wScan_18[4] , 
        \wScan_18[3] , \wScan_18[2] , \wScan_18[1] , \wScan_18[0] }), 
        .ScanOut({\wScan_17[6] , \wScan_17[5] , \wScan_17[4] , \wScan_17[3] , 
        \wScan_17[2] , \wScan_17[1] , \wScan_17[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_17[0] ), .ReturnIn(\wReturn_18[0] ), .ColIn({
        \wColumn_17[63] , \wColumn_17[62] , \wColumn_17[61] , \wColumn_17[60] , 
        \wColumn_17[59] , \wColumn_17[58] , \wColumn_17[57] , \wColumn_17[56] , 
        \wColumn_17[55] , \wColumn_17[54] , \wColumn_17[53] , \wColumn_17[52] , 
        \wColumn_17[51] , \wColumn_17[50] , \wColumn_17[49] , \wColumn_17[48] , 
        \wColumn_17[47] , \wColumn_17[46] , \wColumn_17[45] , \wColumn_17[44] , 
        \wColumn_17[43] , \wColumn_17[42] , \wColumn_17[41] , \wColumn_17[40] , 
        \wColumn_17[39] , \wColumn_17[38] , \wColumn_17[37] , \wColumn_17[36] , 
        \wColumn_17[35] , \wColumn_17[34] , \wColumn_17[33] , \wColumn_17[32] , 
        \wColumn_17[31] , \wColumn_17[30] , \wColumn_17[29] , \wColumn_17[28] , 
        \wColumn_17[27] , \wColumn_17[26] , \wColumn_17[25] , \wColumn_17[24] , 
        \wColumn_17[23] , \wColumn_17[22] , \wColumn_17[21] , \wColumn_17[20] , 
        \wColumn_17[19] , \wColumn_17[18] , \wColumn_17[17] , \wColumn_17[16] , 
        \wColumn_17[15] , \wColumn_17[14] , \wColumn_17[13] , \wColumn_17[12] , 
        \wColumn_17[11] , \wColumn_17[10] , \wColumn_17[9] , \wColumn_17[8] , 
        \wColumn_17[7] , \wColumn_17[6] , \wColumn_17[5] , \wColumn_17[4] , 
        \wColumn_17[3] , \wColumn_17[2] , \wColumn_17[1] , \wColumn_17[0] }), 
        .PDiagIn({\wPDiag_17[63] , \wPDiag_17[62] , \wPDiag_17[61] , 
        \wPDiag_17[60] , \wPDiag_17[59] , \wPDiag_17[58] , \wPDiag_17[57] , 
        \wPDiag_17[56] , \wPDiag_17[55] , \wPDiag_17[54] , \wPDiag_17[53] , 
        \wPDiag_17[52] , \wPDiag_17[51] , \wPDiag_17[50] , \wPDiag_17[49] , 
        \wPDiag_17[48] , \wPDiag_17[47] , \wPDiag_17[46] , \wPDiag_17[45] , 
        \wPDiag_17[44] , \wPDiag_17[43] , \wPDiag_17[42] , \wPDiag_17[41] , 
        \wPDiag_17[40] , \wPDiag_17[39] , \wPDiag_17[38] , \wPDiag_17[37] , 
        \wPDiag_17[36] , \wPDiag_17[35] , \wPDiag_17[34] , \wPDiag_17[33] , 
        \wPDiag_17[32] , \wPDiag_17[31] , \wPDiag_17[30] , \wPDiag_17[29] , 
        \wPDiag_17[28] , \wPDiag_17[27] , \wPDiag_17[26] , \wPDiag_17[25] , 
        \wPDiag_17[24] , \wPDiag_17[23] , \wPDiag_17[22] , \wPDiag_17[21] , 
        \wPDiag_17[20] , \wPDiag_17[19] , \wPDiag_17[18] , \wPDiag_17[17] , 
        \wPDiag_17[16] , \wPDiag_17[15] , \wPDiag_17[14] , \wPDiag_17[13] , 
        \wPDiag_17[12] , \wPDiag_17[11] , \wPDiag_17[10] , \wPDiag_17[9] , 
        \wPDiag_17[8] , \wPDiag_17[7] , \wPDiag_17[6] , \wPDiag_17[5] , 
        \wPDiag_17[4] , \wPDiag_17[3] , \wPDiag_17[2] , \wPDiag_17[1] , 
        \wPDiag_17[0] }), .NDiagIn({\wNDiag_17[63] , \wNDiag_17[62] , 
        \wNDiag_17[61] , \wNDiag_17[60] , \wNDiag_17[59] , \wNDiag_17[58] , 
        \wNDiag_17[57] , \wNDiag_17[56] , \wNDiag_17[55] , \wNDiag_17[54] , 
        \wNDiag_17[53] , \wNDiag_17[52] , \wNDiag_17[51] , \wNDiag_17[50] , 
        \wNDiag_17[49] , \wNDiag_17[48] , \wNDiag_17[47] , \wNDiag_17[46] , 
        \wNDiag_17[45] , \wNDiag_17[44] , \wNDiag_17[43] , \wNDiag_17[42] , 
        \wNDiag_17[41] , \wNDiag_17[40] , \wNDiag_17[39] , \wNDiag_17[38] , 
        \wNDiag_17[37] , \wNDiag_17[36] , \wNDiag_17[35] , \wNDiag_17[34] , 
        \wNDiag_17[33] , \wNDiag_17[32] , \wNDiag_17[31] , \wNDiag_17[30] , 
        \wNDiag_17[29] , \wNDiag_17[28] , \wNDiag_17[27] , \wNDiag_17[26] , 
        \wNDiag_17[25] , \wNDiag_17[24] , \wNDiag_17[23] , \wNDiag_17[22] , 
        \wNDiag_17[21] , \wNDiag_17[20] , \wNDiag_17[19] , \wNDiag_17[18] , 
        \wNDiag_17[17] , \wNDiag_17[16] , \wNDiag_17[15] , \wNDiag_17[14] , 
        \wNDiag_17[13] , \wNDiag_17[12] , \wNDiag_17[11] , \wNDiag_17[10] , 
        \wNDiag_17[9] , \wNDiag_17[8] , \wNDiag_17[7] , \wNDiag_17[6] , 
        \wNDiag_17[5] , \wNDiag_17[4] , \wNDiag_17[3] , \wNDiag_17[2] , 
        \wNDiag_17[1] , \wNDiag_17[0] }), .CallOut(\wCall_18[0] ), .ReturnOut(
        \wReturn_17[0] ), .ColOut({\wColumn_18[63] , \wColumn_18[62] , 
        \wColumn_18[61] , \wColumn_18[60] , \wColumn_18[59] , \wColumn_18[58] , 
        \wColumn_18[57] , \wColumn_18[56] , \wColumn_18[55] , \wColumn_18[54] , 
        \wColumn_18[53] , \wColumn_18[52] , \wColumn_18[51] , \wColumn_18[50] , 
        \wColumn_18[49] , \wColumn_18[48] , \wColumn_18[47] , \wColumn_18[46] , 
        \wColumn_18[45] , \wColumn_18[44] , \wColumn_18[43] , \wColumn_18[42] , 
        \wColumn_18[41] , \wColumn_18[40] , \wColumn_18[39] , \wColumn_18[38] , 
        \wColumn_18[37] , \wColumn_18[36] , \wColumn_18[35] , \wColumn_18[34] , 
        \wColumn_18[33] , \wColumn_18[32] , \wColumn_18[31] , \wColumn_18[30] , 
        \wColumn_18[29] , \wColumn_18[28] , \wColumn_18[27] , \wColumn_18[26] , 
        \wColumn_18[25] , \wColumn_18[24] , \wColumn_18[23] , \wColumn_18[22] , 
        \wColumn_18[21] , \wColumn_18[20] , \wColumn_18[19] , \wColumn_18[18] , 
        \wColumn_18[17] , \wColumn_18[16] , \wColumn_18[15] , \wColumn_18[14] , 
        \wColumn_18[13] , \wColumn_18[12] , \wColumn_18[11] , \wColumn_18[10] , 
        \wColumn_18[9] , \wColumn_18[8] , \wColumn_18[7] , \wColumn_18[6] , 
        \wColumn_18[5] , \wColumn_18[4] , \wColumn_18[3] , \wColumn_18[2] , 
        \wColumn_18[1] , \wColumn_18[0] }), .PDiagOut({\wPDiag_18[63] , 
        \wPDiag_18[62] , \wPDiag_18[61] , \wPDiag_18[60] , \wPDiag_18[59] , 
        \wPDiag_18[58] , \wPDiag_18[57] , \wPDiag_18[56] , \wPDiag_18[55] , 
        \wPDiag_18[54] , \wPDiag_18[53] , \wPDiag_18[52] , \wPDiag_18[51] , 
        \wPDiag_18[50] , \wPDiag_18[49] , \wPDiag_18[48] , \wPDiag_18[47] , 
        \wPDiag_18[46] , \wPDiag_18[45] , \wPDiag_18[44] , \wPDiag_18[43] , 
        \wPDiag_18[42] , \wPDiag_18[41] , \wPDiag_18[40] , \wPDiag_18[39] , 
        \wPDiag_18[38] , \wPDiag_18[37] , \wPDiag_18[36] , \wPDiag_18[35] , 
        \wPDiag_18[34] , \wPDiag_18[33] , \wPDiag_18[32] , \wPDiag_18[31] , 
        \wPDiag_18[30] , \wPDiag_18[29] , \wPDiag_18[28] , \wPDiag_18[27] , 
        \wPDiag_18[26] , \wPDiag_18[25] , \wPDiag_18[24] , \wPDiag_18[23] , 
        \wPDiag_18[22] , \wPDiag_18[21] , \wPDiag_18[20] , \wPDiag_18[19] , 
        \wPDiag_18[18] , \wPDiag_18[17] , \wPDiag_18[16] , \wPDiag_18[15] , 
        \wPDiag_18[14] , \wPDiag_18[13] , \wPDiag_18[12] , \wPDiag_18[11] , 
        \wPDiag_18[10] , \wPDiag_18[9] , \wPDiag_18[8] , \wPDiag_18[7] , 
        \wPDiag_18[6] , \wPDiag_18[5] , \wPDiag_18[4] , \wPDiag_18[3] , 
        \wPDiag_18[2] , \wPDiag_18[1] , \wPDiag_18[0] }), .NDiagOut({
        \wNDiag_18[63] , \wNDiag_18[62] , \wNDiag_18[61] , \wNDiag_18[60] , 
        \wNDiag_18[59] , \wNDiag_18[58] , \wNDiag_18[57] , \wNDiag_18[56] , 
        \wNDiag_18[55] , \wNDiag_18[54] , \wNDiag_18[53] , \wNDiag_18[52] , 
        \wNDiag_18[51] , \wNDiag_18[50] , \wNDiag_18[49] , \wNDiag_18[48] , 
        \wNDiag_18[47] , \wNDiag_18[46] , \wNDiag_18[45] , \wNDiag_18[44] , 
        \wNDiag_18[43] , \wNDiag_18[42] , \wNDiag_18[41] , \wNDiag_18[40] , 
        \wNDiag_18[39] , \wNDiag_18[38] , \wNDiag_18[37] , \wNDiag_18[36] , 
        \wNDiag_18[35] , \wNDiag_18[34] , \wNDiag_18[33] , \wNDiag_18[32] , 
        \wNDiag_18[31] , \wNDiag_18[30] , \wNDiag_18[29] , \wNDiag_18[28] , 
        \wNDiag_18[27] , \wNDiag_18[26] , \wNDiag_18[25] , \wNDiag_18[24] , 
        \wNDiag_18[23] , \wNDiag_18[22] , \wNDiag_18[21] , \wNDiag_18[20] , 
        \wNDiag_18[19] , \wNDiag_18[18] , \wNDiag_18[17] , \wNDiag_18[16] , 
        \wNDiag_18[15] , \wNDiag_18[14] , \wNDiag_18[13] , \wNDiag_18[12] , 
        \wNDiag_18[11] , \wNDiag_18[10] , \wNDiag_18[9] , \wNDiag_18[8] , 
        \wNDiag_18[7] , \wNDiag_18[6] , \wNDiag_18[5] , \wNDiag_18[4] , 
        \wNDiag_18[3] , \wNDiag_18[2] , \wNDiag_18[1] , \wNDiag_18[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_30 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_31[6] , \wScan_31[5] , \wScan_31[4] , 
        \wScan_31[3] , \wScan_31[2] , \wScan_31[1] , \wScan_31[0] }), 
        .ScanOut({\wScan_30[6] , \wScan_30[5] , \wScan_30[4] , \wScan_30[3] , 
        \wScan_30[2] , \wScan_30[1] , \wScan_30[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_30[0] ), .ReturnIn(\wReturn_31[0] ), .ColIn({
        \wColumn_30[63] , \wColumn_30[62] , \wColumn_30[61] , \wColumn_30[60] , 
        \wColumn_30[59] , \wColumn_30[58] , \wColumn_30[57] , \wColumn_30[56] , 
        \wColumn_30[55] , \wColumn_30[54] , \wColumn_30[53] , \wColumn_30[52] , 
        \wColumn_30[51] , \wColumn_30[50] , \wColumn_30[49] , \wColumn_30[48] , 
        \wColumn_30[47] , \wColumn_30[46] , \wColumn_30[45] , \wColumn_30[44] , 
        \wColumn_30[43] , \wColumn_30[42] , \wColumn_30[41] , \wColumn_30[40] , 
        \wColumn_30[39] , \wColumn_30[38] , \wColumn_30[37] , \wColumn_30[36] , 
        \wColumn_30[35] , \wColumn_30[34] , \wColumn_30[33] , \wColumn_30[32] , 
        \wColumn_30[31] , \wColumn_30[30] , \wColumn_30[29] , \wColumn_30[28] , 
        \wColumn_30[27] , \wColumn_30[26] , \wColumn_30[25] , \wColumn_30[24] , 
        \wColumn_30[23] , \wColumn_30[22] , \wColumn_30[21] , \wColumn_30[20] , 
        \wColumn_30[19] , \wColumn_30[18] , \wColumn_30[17] , \wColumn_30[16] , 
        \wColumn_30[15] , \wColumn_30[14] , \wColumn_30[13] , \wColumn_30[12] , 
        \wColumn_30[11] , \wColumn_30[10] , \wColumn_30[9] , \wColumn_30[8] , 
        \wColumn_30[7] , \wColumn_30[6] , \wColumn_30[5] , \wColumn_30[4] , 
        \wColumn_30[3] , \wColumn_30[2] , \wColumn_30[1] , \wColumn_30[0] }), 
        .PDiagIn({\wPDiag_30[63] , \wPDiag_30[62] , \wPDiag_30[61] , 
        \wPDiag_30[60] , \wPDiag_30[59] , \wPDiag_30[58] , \wPDiag_30[57] , 
        \wPDiag_30[56] , \wPDiag_30[55] , \wPDiag_30[54] , \wPDiag_30[53] , 
        \wPDiag_30[52] , \wPDiag_30[51] , \wPDiag_30[50] , \wPDiag_30[49] , 
        \wPDiag_30[48] , \wPDiag_30[47] , \wPDiag_30[46] , \wPDiag_30[45] , 
        \wPDiag_30[44] , \wPDiag_30[43] , \wPDiag_30[42] , \wPDiag_30[41] , 
        \wPDiag_30[40] , \wPDiag_30[39] , \wPDiag_30[38] , \wPDiag_30[37] , 
        \wPDiag_30[36] , \wPDiag_30[35] , \wPDiag_30[34] , \wPDiag_30[33] , 
        \wPDiag_30[32] , \wPDiag_30[31] , \wPDiag_30[30] , \wPDiag_30[29] , 
        \wPDiag_30[28] , \wPDiag_30[27] , \wPDiag_30[26] , \wPDiag_30[25] , 
        \wPDiag_30[24] , \wPDiag_30[23] , \wPDiag_30[22] , \wPDiag_30[21] , 
        \wPDiag_30[20] , \wPDiag_30[19] , \wPDiag_30[18] , \wPDiag_30[17] , 
        \wPDiag_30[16] , \wPDiag_30[15] , \wPDiag_30[14] , \wPDiag_30[13] , 
        \wPDiag_30[12] , \wPDiag_30[11] , \wPDiag_30[10] , \wPDiag_30[9] , 
        \wPDiag_30[8] , \wPDiag_30[7] , \wPDiag_30[6] , \wPDiag_30[5] , 
        \wPDiag_30[4] , \wPDiag_30[3] , \wPDiag_30[2] , \wPDiag_30[1] , 
        \wPDiag_30[0] }), .NDiagIn({\wNDiag_30[63] , \wNDiag_30[62] , 
        \wNDiag_30[61] , \wNDiag_30[60] , \wNDiag_30[59] , \wNDiag_30[58] , 
        \wNDiag_30[57] , \wNDiag_30[56] , \wNDiag_30[55] , \wNDiag_30[54] , 
        \wNDiag_30[53] , \wNDiag_30[52] , \wNDiag_30[51] , \wNDiag_30[50] , 
        \wNDiag_30[49] , \wNDiag_30[48] , \wNDiag_30[47] , \wNDiag_30[46] , 
        \wNDiag_30[45] , \wNDiag_30[44] , \wNDiag_30[43] , \wNDiag_30[42] , 
        \wNDiag_30[41] , \wNDiag_30[40] , \wNDiag_30[39] , \wNDiag_30[38] , 
        \wNDiag_30[37] , \wNDiag_30[36] , \wNDiag_30[35] , \wNDiag_30[34] , 
        \wNDiag_30[33] , \wNDiag_30[32] , \wNDiag_30[31] , \wNDiag_30[30] , 
        \wNDiag_30[29] , \wNDiag_30[28] , \wNDiag_30[27] , \wNDiag_30[26] , 
        \wNDiag_30[25] , \wNDiag_30[24] , \wNDiag_30[23] , \wNDiag_30[22] , 
        \wNDiag_30[21] , \wNDiag_30[20] , \wNDiag_30[19] , \wNDiag_30[18] , 
        \wNDiag_30[17] , \wNDiag_30[16] , \wNDiag_30[15] , \wNDiag_30[14] , 
        \wNDiag_30[13] , \wNDiag_30[12] , \wNDiag_30[11] , \wNDiag_30[10] , 
        \wNDiag_30[9] , \wNDiag_30[8] , \wNDiag_30[7] , \wNDiag_30[6] , 
        \wNDiag_30[5] , \wNDiag_30[4] , \wNDiag_30[3] , \wNDiag_30[2] , 
        \wNDiag_30[1] , \wNDiag_30[0] }), .CallOut(\wCall_31[0] ), .ReturnOut(
        \wReturn_30[0] ), .ColOut({\wColumn_31[63] , \wColumn_31[62] , 
        \wColumn_31[61] , \wColumn_31[60] , \wColumn_31[59] , \wColumn_31[58] , 
        \wColumn_31[57] , \wColumn_31[56] , \wColumn_31[55] , \wColumn_31[54] , 
        \wColumn_31[53] , \wColumn_31[52] , \wColumn_31[51] , \wColumn_31[50] , 
        \wColumn_31[49] , \wColumn_31[48] , \wColumn_31[47] , \wColumn_31[46] , 
        \wColumn_31[45] , \wColumn_31[44] , \wColumn_31[43] , \wColumn_31[42] , 
        \wColumn_31[41] , \wColumn_31[40] , \wColumn_31[39] , \wColumn_31[38] , 
        \wColumn_31[37] , \wColumn_31[36] , \wColumn_31[35] , \wColumn_31[34] , 
        \wColumn_31[33] , \wColumn_31[32] , \wColumn_31[31] , \wColumn_31[30] , 
        \wColumn_31[29] , \wColumn_31[28] , \wColumn_31[27] , \wColumn_31[26] , 
        \wColumn_31[25] , \wColumn_31[24] , \wColumn_31[23] , \wColumn_31[22] , 
        \wColumn_31[21] , \wColumn_31[20] , \wColumn_31[19] , \wColumn_31[18] , 
        \wColumn_31[17] , \wColumn_31[16] , \wColumn_31[15] , \wColumn_31[14] , 
        \wColumn_31[13] , \wColumn_31[12] , \wColumn_31[11] , \wColumn_31[10] , 
        \wColumn_31[9] , \wColumn_31[8] , \wColumn_31[7] , \wColumn_31[6] , 
        \wColumn_31[5] , \wColumn_31[4] , \wColumn_31[3] , \wColumn_31[2] , 
        \wColumn_31[1] , \wColumn_31[0] }), .PDiagOut({\wPDiag_31[63] , 
        \wPDiag_31[62] , \wPDiag_31[61] , \wPDiag_31[60] , \wPDiag_31[59] , 
        \wPDiag_31[58] , \wPDiag_31[57] , \wPDiag_31[56] , \wPDiag_31[55] , 
        \wPDiag_31[54] , \wPDiag_31[53] , \wPDiag_31[52] , \wPDiag_31[51] , 
        \wPDiag_31[50] , \wPDiag_31[49] , \wPDiag_31[48] , \wPDiag_31[47] , 
        \wPDiag_31[46] , \wPDiag_31[45] , \wPDiag_31[44] , \wPDiag_31[43] , 
        \wPDiag_31[42] , \wPDiag_31[41] , \wPDiag_31[40] , \wPDiag_31[39] , 
        \wPDiag_31[38] , \wPDiag_31[37] , \wPDiag_31[36] , \wPDiag_31[35] , 
        \wPDiag_31[34] , \wPDiag_31[33] , \wPDiag_31[32] , \wPDiag_31[31] , 
        \wPDiag_31[30] , \wPDiag_31[29] , \wPDiag_31[28] , \wPDiag_31[27] , 
        \wPDiag_31[26] , \wPDiag_31[25] , \wPDiag_31[24] , \wPDiag_31[23] , 
        \wPDiag_31[22] , \wPDiag_31[21] , \wPDiag_31[20] , \wPDiag_31[19] , 
        \wPDiag_31[18] , \wPDiag_31[17] , \wPDiag_31[16] , \wPDiag_31[15] , 
        \wPDiag_31[14] , \wPDiag_31[13] , \wPDiag_31[12] , \wPDiag_31[11] , 
        \wPDiag_31[10] , \wPDiag_31[9] , \wPDiag_31[8] , \wPDiag_31[7] , 
        \wPDiag_31[6] , \wPDiag_31[5] , \wPDiag_31[4] , \wPDiag_31[3] , 
        \wPDiag_31[2] , \wPDiag_31[1] , \wPDiag_31[0] }), .NDiagOut({
        \wNDiag_31[63] , \wNDiag_31[62] , \wNDiag_31[61] , \wNDiag_31[60] , 
        \wNDiag_31[59] , \wNDiag_31[58] , \wNDiag_31[57] , \wNDiag_31[56] , 
        \wNDiag_31[55] , \wNDiag_31[54] , \wNDiag_31[53] , \wNDiag_31[52] , 
        \wNDiag_31[51] , \wNDiag_31[50] , \wNDiag_31[49] , \wNDiag_31[48] , 
        \wNDiag_31[47] , \wNDiag_31[46] , \wNDiag_31[45] , \wNDiag_31[44] , 
        \wNDiag_31[43] , \wNDiag_31[42] , \wNDiag_31[41] , \wNDiag_31[40] , 
        \wNDiag_31[39] , \wNDiag_31[38] , \wNDiag_31[37] , \wNDiag_31[36] , 
        \wNDiag_31[35] , \wNDiag_31[34] , \wNDiag_31[33] , \wNDiag_31[32] , 
        \wNDiag_31[31] , \wNDiag_31[30] , \wNDiag_31[29] , \wNDiag_31[28] , 
        \wNDiag_31[27] , \wNDiag_31[26] , \wNDiag_31[25] , \wNDiag_31[24] , 
        \wNDiag_31[23] , \wNDiag_31[22] , \wNDiag_31[21] , \wNDiag_31[20] , 
        \wNDiag_31[19] , \wNDiag_31[18] , \wNDiag_31[17] , \wNDiag_31[16] , 
        \wNDiag_31[15] , \wNDiag_31[14] , \wNDiag_31[13] , \wNDiag_31[12] , 
        \wNDiag_31[11] , \wNDiag_31[10] , \wNDiag_31[9] , \wNDiag_31[8] , 
        \wNDiag_31[7] , \wNDiag_31[6] , \wNDiag_31[5] , \wNDiag_31[4] , 
        \wNDiag_31[3] , \wNDiag_31[2] , \wNDiag_31[1] , \wNDiag_31[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_39 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_40[6] , \wScan_40[5] , \wScan_40[4] , 
        \wScan_40[3] , \wScan_40[2] , \wScan_40[1] , \wScan_40[0] }), 
        .ScanOut({\wScan_39[6] , \wScan_39[5] , \wScan_39[4] , \wScan_39[3] , 
        \wScan_39[2] , \wScan_39[1] , \wScan_39[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_39[0] ), .ReturnIn(\wReturn_40[0] ), .ColIn({
        \wColumn_39[63] , \wColumn_39[62] , \wColumn_39[61] , \wColumn_39[60] , 
        \wColumn_39[59] , \wColumn_39[58] , \wColumn_39[57] , \wColumn_39[56] , 
        \wColumn_39[55] , \wColumn_39[54] , \wColumn_39[53] , \wColumn_39[52] , 
        \wColumn_39[51] , \wColumn_39[50] , \wColumn_39[49] , \wColumn_39[48] , 
        \wColumn_39[47] , \wColumn_39[46] , \wColumn_39[45] , \wColumn_39[44] , 
        \wColumn_39[43] , \wColumn_39[42] , \wColumn_39[41] , \wColumn_39[40] , 
        \wColumn_39[39] , \wColumn_39[38] , \wColumn_39[37] , \wColumn_39[36] , 
        \wColumn_39[35] , \wColumn_39[34] , \wColumn_39[33] , \wColumn_39[32] , 
        \wColumn_39[31] , \wColumn_39[30] , \wColumn_39[29] , \wColumn_39[28] , 
        \wColumn_39[27] , \wColumn_39[26] , \wColumn_39[25] , \wColumn_39[24] , 
        \wColumn_39[23] , \wColumn_39[22] , \wColumn_39[21] , \wColumn_39[20] , 
        \wColumn_39[19] , \wColumn_39[18] , \wColumn_39[17] , \wColumn_39[16] , 
        \wColumn_39[15] , \wColumn_39[14] , \wColumn_39[13] , \wColumn_39[12] , 
        \wColumn_39[11] , \wColumn_39[10] , \wColumn_39[9] , \wColumn_39[8] , 
        \wColumn_39[7] , \wColumn_39[6] , \wColumn_39[5] , \wColumn_39[4] , 
        \wColumn_39[3] , \wColumn_39[2] , \wColumn_39[1] , \wColumn_39[0] }), 
        .PDiagIn({\wPDiag_39[63] , \wPDiag_39[62] , \wPDiag_39[61] , 
        \wPDiag_39[60] , \wPDiag_39[59] , \wPDiag_39[58] , \wPDiag_39[57] , 
        \wPDiag_39[56] , \wPDiag_39[55] , \wPDiag_39[54] , \wPDiag_39[53] , 
        \wPDiag_39[52] , \wPDiag_39[51] , \wPDiag_39[50] , \wPDiag_39[49] , 
        \wPDiag_39[48] , \wPDiag_39[47] , \wPDiag_39[46] , \wPDiag_39[45] , 
        \wPDiag_39[44] , \wPDiag_39[43] , \wPDiag_39[42] , \wPDiag_39[41] , 
        \wPDiag_39[40] , \wPDiag_39[39] , \wPDiag_39[38] , \wPDiag_39[37] , 
        \wPDiag_39[36] , \wPDiag_39[35] , \wPDiag_39[34] , \wPDiag_39[33] , 
        \wPDiag_39[32] , \wPDiag_39[31] , \wPDiag_39[30] , \wPDiag_39[29] , 
        \wPDiag_39[28] , \wPDiag_39[27] , \wPDiag_39[26] , \wPDiag_39[25] , 
        \wPDiag_39[24] , \wPDiag_39[23] , \wPDiag_39[22] , \wPDiag_39[21] , 
        \wPDiag_39[20] , \wPDiag_39[19] , \wPDiag_39[18] , \wPDiag_39[17] , 
        \wPDiag_39[16] , \wPDiag_39[15] , \wPDiag_39[14] , \wPDiag_39[13] , 
        \wPDiag_39[12] , \wPDiag_39[11] , \wPDiag_39[10] , \wPDiag_39[9] , 
        \wPDiag_39[8] , \wPDiag_39[7] , \wPDiag_39[6] , \wPDiag_39[5] , 
        \wPDiag_39[4] , \wPDiag_39[3] , \wPDiag_39[2] , \wPDiag_39[1] , 
        \wPDiag_39[0] }), .NDiagIn({\wNDiag_39[63] , \wNDiag_39[62] , 
        \wNDiag_39[61] , \wNDiag_39[60] , \wNDiag_39[59] , \wNDiag_39[58] , 
        \wNDiag_39[57] , \wNDiag_39[56] , \wNDiag_39[55] , \wNDiag_39[54] , 
        \wNDiag_39[53] , \wNDiag_39[52] , \wNDiag_39[51] , \wNDiag_39[50] , 
        \wNDiag_39[49] , \wNDiag_39[48] , \wNDiag_39[47] , \wNDiag_39[46] , 
        \wNDiag_39[45] , \wNDiag_39[44] , \wNDiag_39[43] , \wNDiag_39[42] , 
        \wNDiag_39[41] , \wNDiag_39[40] , \wNDiag_39[39] , \wNDiag_39[38] , 
        \wNDiag_39[37] , \wNDiag_39[36] , \wNDiag_39[35] , \wNDiag_39[34] , 
        \wNDiag_39[33] , \wNDiag_39[32] , \wNDiag_39[31] , \wNDiag_39[30] , 
        \wNDiag_39[29] , \wNDiag_39[28] , \wNDiag_39[27] , \wNDiag_39[26] , 
        \wNDiag_39[25] , \wNDiag_39[24] , \wNDiag_39[23] , \wNDiag_39[22] , 
        \wNDiag_39[21] , \wNDiag_39[20] , \wNDiag_39[19] , \wNDiag_39[18] , 
        \wNDiag_39[17] , \wNDiag_39[16] , \wNDiag_39[15] , \wNDiag_39[14] , 
        \wNDiag_39[13] , \wNDiag_39[12] , \wNDiag_39[11] , \wNDiag_39[10] , 
        \wNDiag_39[9] , \wNDiag_39[8] , \wNDiag_39[7] , \wNDiag_39[6] , 
        \wNDiag_39[5] , \wNDiag_39[4] , \wNDiag_39[3] , \wNDiag_39[2] , 
        \wNDiag_39[1] , \wNDiag_39[0] }), .CallOut(\wCall_40[0] ), .ReturnOut(
        \wReturn_39[0] ), .ColOut({\wColumn_40[63] , \wColumn_40[62] , 
        \wColumn_40[61] , \wColumn_40[60] , \wColumn_40[59] , \wColumn_40[58] , 
        \wColumn_40[57] , \wColumn_40[56] , \wColumn_40[55] , \wColumn_40[54] , 
        \wColumn_40[53] , \wColumn_40[52] , \wColumn_40[51] , \wColumn_40[50] , 
        \wColumn_40[49] , \wColumn_40[48] , \wColumn_40[47] , \wColumn_40[46] , 
        \wColumn_40[45] , \wColumn_40[44] , \wColumn_40[43] , \wColumn_40[42] , 
        \wColumn_40[41] , \wColumn_40[40] , \wColumn_40[39] , \wColumn_40[38] , 
        \wColumn_40[37] , \wColumn_40[36] , \wColumn_40[35] , \wColumn_40[34] , 
        \wColumn_40[33] , \wColumn_40[32] , \wColumn_40[31] , \wColumn_40[30] , 
        \wColumn_40[29] , \wColumn_40[28] , \wColumn_40[27] , \wColumn_40[26] , 
        \wColumn_40[25] , \wColumn_40[24] , \wColumn_40[23] , \wColumn_40[22] , 
        \wColumn_40[21] , \wColumn_40[20] , \wColumn_40[19] , \wColumn_40[18] , 
        \wColumn_40[17] , \wColumn_40[16] , \wColumn_40[15] , \wColumn_40[14] , 
        \wColumn_40[13] , \wColumn_40[12] , \wColumn_40[11] , \wColumn_40[10] , 
        \wColumn_40[9] , \wColumn_40[8] , \wColumn_40[7] , \wColumn_40[6] , 
        \wColumn_40[5] , \wColumn_40[4] , \wColumn_40[3] , \wColumn_40[2] , 
        \wColumn_40[1] , \wColumn_40[0] }), .PDiagOut({\wPDiag_40[63] , 
        \wPDiag_40[62] , \wPDiag_40[61] , \wPDiag_40[60] , \wPDiag_40[59] , 
        \wPDiag_40[58] , \wPDiag_40[57] , \wPDiag_40[56] , \wPDiag_40[55] , 
        \wPDiag_40[54] , \wPDiag_40[53] , \wPDiag_40[52] , \wPDiag_40[51] , 
        \wPDiag_40[50] , \wPDiag_40[49] , \wPDiag_40[48] , \wPDiag_40[47] , 
        \wPDiag_40[46] , \wPDiag_40[45] , \wPDiag_40[44] , \wPDiag_40[43] , 
        \wPDiag_40[42] , \wPDiag_40[41] , \wPDiag_40[40] , \wPDiag_40[39] , 
        \wPDiag_40[38] , \wPDiag_40[37] , \wPDiag_40[36] , \wPDiag_40[35] , 
        \wPDiag_40[34] , \wPDiag_40[33] , \wPDiag_40[32] , \wPDiag_40[31] , 
        \wPDiag_40[30] , \wPDiag_40[29] , \wPDiag_40[28] , \wPDiag_40[27] , 
        \wPDiag_40[26] , \wPDiag_40[25] , \wPDiag_40[24] , \wPDiag_40[23] , 
        \wPDiag_40[22] , \wPDiag_40[21] , \wPDiag_40[20] , \wPDiag_40[19] , 
        \wPDiag_40[18] , \wPDiag_40[17] , \wPDiag_40[16] , \wPDiag_40[15] , 
        \wPDiag_40[14] , \wPDiag_40[13] , \wPDiag_40[12] , \wPDiag_40[11] , 
        \wPDiag_40[10] , \wPDiag_40[9] , \wPDiag_40[8] , \wPDiag_40[7] , 
        \wPDiag_40[6] , \wPDiag_40[5] , \wPDiag_40[4] , \wPDiag_40[3] , 
        \wPDiag_40[2] , \wPDiag_40[1] , \wPDiag_40[0] }), .NDiagOut({
        \wNDiag_40[63] , \wNDiag_40[62] , \wNDiag_40[61] , \wNDiag_40[60] , 
        \wNDiag_40[59] , \wNDiag_40[58] , \wNDiag_40[57] , \wNDiag_40[56] , 
        \wNDiag_40[55] , \wNDiag_40[54] , \wNDiag_40[53] , \wNDiag_40[52] , 
        \wNDiag_40[51] , \wNDiag_40[50] , \wNDiag_40[49] , \wNDiag_40[48] , 
        \wNDiag_40[47] , \wNDiag_40[46] , \wNDiag_40[45] , \wNDiag_40[44] , 
        \wNDiag_40[43] , \wNDiag_40[42] , \wNDiag_40[41] , \wNDiag_40[40] , 
        \wNDiag_40[39] , \wNDiag_40[38] , \wNDiag_40[37] , \wNDiag_40[36] , 
        \wNDiag_40[35] , \wNDiag_40[34] , \wNDiag_40[33] , \wNDiag_40[32] , 
        \wNDiag_40[31] , \wNDiag_40[30] , \wNDiag_40[29] , \wNDiag_40[28] , 
        \wNDiag_40[27] , \wNDiag_40[26] , \wNDiag_40[25] , \wNDiag_40[24] , 
        \wNDiag_40[23] , \wNDiag_40[22] , \wNDiag_40[21] , \wNDiag_40[20] , 
        \wNDiag_40[19] , \wNDiag_40[18] , \wNDiag_40[17] , \wNDiag_40[16] , 
        \wNDiag_40[15] , \wNDiag_40[14] , \wNDiag_40[13] , \wNDiag_40[12] , 
        \wNDiag_40[11] , \wNDiag_40[10] , \wNDiag_40[9] , \wNDiag_40[8] , 
        \wNDiag_40[7] , \wNDiag_40[6] , \wNDiag_40[5] , \wNDiag_40[4] , 
        \wNDiag_40[3] , \wNDiag_40[2] , \wNDiag_40[1] , \wNDiag_40[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_45 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_46[6] , \wScan_46[5] , \wScan_46[4] , 
        \wScan_46[3] , \wScan_46[2] , \wScan_46[1] , \wScan_46[0] }), 
        .ScanOut({\wScan_45[6] , \wScan_45[5] , \wScan_45[4] , \wScan_45[3] , 
        \wScan_45[2] , \wScan_45[1] , \wScan_45[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_45[0] ), .ReturnIn(\wReturn_46[0] ), .ColIn({
        \wColumn_45[63] , \wColumn_45[62] , \wColumn_45[61] , \wColumn_45[60] , 
        \wColumn_45[59] , \wColumn_45[58] , \wColumn_45[57] , \wColumn_45[56] , 
        \wColumn_45[55] , \wColumn_45[54] , \wColumn_45[53] , \wColumn_45[52] , 
        \wColumn_45[51] , \wColumn_45[50] , \wColumn_45[49] , \wColumn_45[48] , 
        \wColumn_45[47] , \wColumn_45[46] , \wColumn_45[45] , \wColumn_45[44] , 
        \wColumn_45[43] , \wColumn_45[42] , \wColumn_45[41] , \wColumn_45[40] , 
        \wColumn_45[39] , \wColumn_45[38] , \wColumn_45[37] , \wColumn_45[36] , 
        \wColumn_45[35] , \wColumn_45[34] , \wColumn_45[33] , \wColumn_45[32] , 
        \wColumn_45[31] , \wColumn_45[30] , \wColumn_45[29] , \wColumn_45[28] , 
        \wColumn_45[27] , \wColumn_45[26] , \wColumn_45[25] , \wColumn_45[24] , 
        \wColumn_45[23] , \wColumn_45[22] , \wColumn_45[21] , \wColumn_45[20] , 
        \wColumn_45[19] , \wColumn_45[18] , \wColumn_45[17] , \wColumn_45[16] , 
        \wColumn_45[15] , \wColumn_45[14] , \wColumn_45[13] , \wColumn_45[12] , 
        \wColumn_45[11] , \wColumn_45[10] , \wColumn_45[9] , \wColumn_45[8] , 
        \wColumn_45[7] , \wColumn_45[6] , \wColumn_45[5] , \wColumn_45[4] , 
        \wColumn_45[3] , \wColumn_45[2] , \wColumn_45[1] , \wColumn_45[0] }), 
        .PDiagIn({\wPDiag_45[63] , \wPDiag_45[62] , \wPDiag_45[61] , 
        \wPDiag_45[60] , \wPDiag_45[59] , \wPDiag_45[58] , \wPDiag_45[57] , 
        \wPDiag_45[56] , \wPDiag_45[55] , \wPDiag_45[54] , \wPDiag_45[53] , 
        \wPDiag_45[52] , \wPDiag_45[51] , \wPDiag_45[50] , \wPDiag_45[49] , 
        \wPDiag_45[48] , \wPDiag_45[47] , \wPDiag_45[46] , \wPDiag_45[45] , 
        \wPDiag_45[44] , \wPDiag_45[43] , \wPDiag_45[42] , \wPDiag_45[41] , 
        \wPDiag_45[40] , \wPDiag_45[39] , \wPDiag_45[38] , \wPDiag_45[37] , 
        \wPDiag_45[36] , \wPDiag_45[35] , \wPDiag_45[34] , \wPDiag_45[33] , 
        \wPDiag_45[32] , \wPDiag_45[31] , \wPDiag_45[30] , \wPDiag_45[29] , 
        \wPDiag_45[28] , \wPDiag_45[27] , \wPDiag_45[26] , \wPDiag_45[25] , 
        \wPDiag_45[24] , \wPDiag_45[23] , \wPDiag_45[22] , \wPDiag_45[21] , 
        \wPDiag_45[20] , \wPDiag_45[19] , \wPDiag_45[18] , \wPDiag_45[17] , 
        \wPDiag_45[16] , \wPDiag_45[15] , \wPDiag_45[14] , \wPDiag_45[13] , 
        \wPDiag_45[12] , \wPDiag_45[11] , \wPDiag_45[10] , \wPDiag_45[9] , 
        \wPDiag_45[8] , \wPDiag_45[7] , \wPDiag_45[6] , \wPDiag_45[5] , 
        \wPDiag_45[4] , \wPDiag_45[3] , \wPDiag_45[2] , \wPDiag_45[1] , 
        \wPDiag_45[0] }), .NDiagIn({\wNDiag_45[63] , \wNDiag_45[62] , 
        \wNDiag_45[61] , \wNDiag_45[60] , \wNDiag_45[59] , \wNDiag_45[58] , 
        \wNDiag_45[57] , \wNDiag_45[56] , \wNDiag_45[55] , \wNDiag_45[54] , 
        \wNDiag_45[53] , \wNDiag_45[52] , \wNDiag_45[51] , \wNDiag_45[50] , 
        \wNDiag_45[49] , \wNDiag_45[48] , \wNDiag_45[47] , \wNDiag_45[46] , 
        \wNDiag_45[45] , \wNDiag_45[44] , \wNDiag_45[43] , \wNDiag_45[42] , 
        \wNDiag_45[41] , \wNDiag_45[40] , \wNDiag_45[39] , \wNDiag_45[38] , 
        \wNDiag_45[37] , \wNDiag_45[36] , \wNDiag_45[35] , \wNDiag_45[34] , 
        \wNDiag_45[33] , \wNDiag_45[32] , \wNDiag_45[31] , \wNDiag_45[30] , 
        \wNDiag_45[29] , \wNDiag_45[28] , \wNDiag_45[27] , \wNDiag_45[26] , 
        \wNDiag_45[25] , \wNDiag_45[24] , \wNDiag_45[23] , \wNDiag_45[22] , 
        \wNDiag_45[21] , \wNDiag_45[20] , \wNDiag_45[19] , \wNDiag_45[18] , 
        \wNDiag_45[17] , \wNDiag_45[16] , \wNDiag_45[15] , \wNDiag_45[14] , 
        \wNDiag_45[13] , \wNDiag_45[12] , \wNDiag_45[11] , \wNDiag_45[10] , 
        \wNDiag_45[9] , \wNDiag_45[8] , \wNDiag_45[7] , \wNDiag_45[6] , 
        \wNDiag_45[5] , \wNDiag_45[4] , \wNDiag_45[3] , \wNDiag_45[2] , 
        \wNDiag_45[1] , \wNDiag_45[0] }), .CallOut(\wCall_46[0] ), .ReturnOut(
        \wReturn_45[0] ), .ColOut({\wColumn_46[63] , \wColumn_46[62] , 
        \wColumn_46[61] , \wColumn_46[60] , \wColumn_46[59] , \wColumn_46[58] , 
        \wColumn_46[57] , \wColumn_46[56] , \wColumn_46[55] , \wColumn_46[54] , 
        \wColumn_46[53] , \wColumn_46[52] , \wColumn_46[51] , \wColumn_46[50] , 
        \wColumn_46[49] , \wColumn_46[48] , \wColumn_46[47] , \wColumn_46[46] , 
        \wColumn_46[45] , \wColumn_46[44] , \wColumn_46[43] , \wColumn_46[42] , 
        \wColumn_46[41] , \wColumn_46[40] , \wColumn_46[39] , \wColumn_46[38] , 
        \wColumn_46[37] , \wColumn_46[36] , \wColumn_46[35] , \wColumn_46[34] , 
        \wColumn_46[33] , \wColumn_46[32] , \wColumn_46[31] , \wColumn_46[30] , 
        \wColumn_46[29] , \wColumn_46[28] , \wColumn_46[27] , \wColumn_46[26] , 
        \wColumn_46[25] , \wColumn_46[24] , \wColumn_46[23] , \wColumn_46[22] , 
        \wColumn_46[21] , \wColumn_46[20] , \wColumn_46[19] , \wColumn_46[18] , 
        \wColumn_46[17] , \wColumn_46[16] , \wColumn_46[15] , \wColumn_46[14] , 
        \wColumn_46[13] , \wColumn_46[12] , \wColumn_46[11] , \wColumn_46[10] , 
        \wColumn_46[9] , \wColumn_46[8] , \wColumn_46[7] , \wColumn_46[6] , 
        \wColumn_46[5] , \wColumn_46[4] , \wColumn_46[3] , \wColumn_46[2] , 
        \wColumn_46[1] , \wColumn_46[0] }), .PDiagOut({\wPDiag_46[63] , 
        \wPDiag_46[62] , \wPDiag_46[61] , \wPDiag_46[60] , \wPDiag_46[59] , 
        \wPDiag_46[58] , \wPDiag_46[57] , \wPDiag_46[56] , \wPDiag_46[55] , 
        \wPDiag_46[54] , \wPDiag_46[53] , \wPDiag_46[52] , \wPDiag_46[51] , 
        \wPDiag_46[50] , \wPDiag_46[49] , \wPDiag_46[48] , \wPDiag_46[47] , 
        \wPDiag_46[46] , \wPDiag_46[45] , \wPDiag_46[44] , \wPDiag_46[43] , 
        \wPDiag_46[42] , \wPDiag_46[41] , \wPDiag_46[40] , \wPDiag_46[39] , 
        \wPDiag_46[38] , \wPDiag_46[37] , \wPDiag_46[36] , \wPDiag_46[35] , 
        \wPDiag_46[34] , \wPDiag_46[33] , \wPDiag_46[32] , \wPDiag_46[31] , 
        \wPDiag_46[30] , \wPDiag_46[29] , \wPDiag_46[28] , \wPDiag_46[27] , 
        \wPDiag_46[26] , \wPDiag_46[25] , \wPDiag_46[24] , \wPDiag_46[23] , 
        \wPDiag_46[22] , \wPDiag_46[21] , \wPDiag_46[20] , \wPDiag_46[19] , 
        \wPDiag_46[18] , \wPDiag_46[17] , \wPDiag_46[16] , \wPDiag_46[15] , 
        \wPDiag_46[14] , \wPDiag_46[13] , \wPDiag_46[12] , \wPDiag_46[11] , 
        \wPDiag_46[10] , \wPDiag_46[9] , \wPDiag_46[8] , \wPDiag_46[7] , 
        \wPDiag_46[6] , \wPDiag_46[5] , \wPDiag_46[4] , \wPDiag_46[3] , 
        \wPDiag_46[2] , \wPDiag_46[1] , \wPDiag_46[0] }), .NDiagOut({
        \wNDiag_46[63] , \wNDiag_46[62] , \wNDiag_46[61] , \wNDiag_46[60] , 
        \wNDiag_46[59] , \wNDiag_46[58] , \wNDiag_46[57] , \wNDiag_46[56] , 
        \wNDiag_46[55] , \wNDiag_46[54] , \wNDiag_46[53] , \wNDiag_46[52] , 
        \wNDiag_46[51] , \wNDiag_46[50] , \wNDiag_46[49] , \wNDiag_46[48] , 
        \wNDiag_46[47] , \wNDiag_46[46] , \wNDiag_46[45] , \wNDiag_46[44] , 
        \wNDiag_46[43] , \wNDiag_46[42] , \wNDiag_46[41] , \wNDiag_46[40] , 
        \wNDiag_46[39] , \wNDiag_46[38] , \wNDiag_46[37] , \wNDiag_46[36] , 
        \wNDiag_46[35] , \wNDiag_46[34] , \wNDiag_46[33] , \wNDiag_46[32] , 
        \wNDiag_46[31] , \wNDiag_46[30] , \wNDiag_46[29] , \wNDiag_46[28] , 
        \wNDiag_46[27] , \wNDiag_46[26] , \wNDiag_46[25] , \wNDiag_46[24] , 
        \wNDiag_46[23] , \wNDiag_46[22] , \wNDiag_46[21] , \wNDiag_46[20] , 
        \wNDiag_46[19] , \wNDiag_46[18] , \wNDiag_46[17] , \wNDiag_46[16] , 
        \wNDiag_46[15] , \wNDiag_46[14] , \wNDiag_46[13] , \wNDiag_46[12] , 
        \wNDiag_46[11] , \wNDiag_46[10] , \wNDiag_46[9] , \wNDiag_46[8] , 
        \wNDiag_46[7] , \wNDiag_46[6] , \wNDiag_46[5] , \wNDiag_46[4] , 
        \wNDiag_46[3] , \wNDiag_46[2] , \wNDiag_46[1] , \wNDiag_46[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_62 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_63[6] , \wScan_63[5] , \wScan_63[4] , 
        \wScan_63[3] , \wScan_63[2] , \wScan_63[1] , \wScan_63[0] }), 
        .ScanOut({\wScan_62[6] , \wScan_62[5] , \wScan_62[4] , \wScan_62[3] , 
        \wScan_62[2] , \wScan_62[1] , \wScan_62[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_62[0] ), .ReturnIn(\wReturn_63[0] ), .ColIn({
        \wColumn_62[63] , \wColumn_62[62] , \wColumn_62[61] , \wColumn_62[60] , 
        \wColumn_62[59] , \wColumn_62[58] , \wColumn_62[57] , \wColumn_62[56] , 
        \wColumn_62[55] , \wColumn_62[54] , \wColumn_62[53] , \wColumn_62[52] , 
        \wColumn_62[51] , \wColumn_62[50] , \wColumn_62[49] , \wColumn_62[48] , 
        \wColumn_62[47] , \wColumn_62[46] , \wColumn_62[45] , \wColumn_62[44] , 
        \wColumn_62[43] , \wColumn_62[42] , \wColumn_62[41] , \wColumn_62[40] , 
        \wColumn_62[39] , \wColumn_62[38] , \wColumn_62[37] , \wColumn_62[36] , 
        \wColumn_62[35] , \wColumn_62[34] , \wColumn_62[33] , \wColumn_62[32] , 
        \wColumn_62[31] , \wColumn_62[30] , \wColumn_62[29] , \wColumn_62[28] , 
        \wColumn_62[27] , \wColumn_62[26] , \wColumn_62[25] , \wColumn_62[24] , 
        \wColumn_62[23] , \wColumn_62[22] , \wColumn_62[21] , \wColumn_62[20] , 
        \wColumn_62[19] , \wColumn_62[18] , \wColumn_62[17] , \wColumn_62[16] , 
        \wColumn_62[15] , \wColumn_62[14] , \wColumn_62[13] , \wColumn_62[12] , 
        \wColumn_62[11] , \wColumn_62[10] , \wColumn_62[9] , \wColumn_62[8] , 
        \wColumn_62[7] , \wColumn_62[6] , \wColumn_62[5] , \wColumn_62[4] , 
        \wColumn_62[3] , \wColumn_62[2] , \wColumn_62[1] , \wColumn_62[0] }), 
        .PDiagIn({\wPDiag_62[63] , \wPDiag_62[62] , \wPDiag_62[61] , 
        \wPDiag_62[60] , \wPDiag_62[59] , \wPDiag_62[58] , \wPDiag_62[57] , 
        \wPDiag_62[56] , \wPDiag_62[55] , \wPDiag_62[54] , \wPDiag_62[53] , 
        \wPDiag_62[52] , \wPDiag_62[51] , \wPDiag_62[50] , \wPDiag_62[49] , 
        \wPDiag_62[48] , \wPDiag_62[47] , \wPDiag_62[46] , \wPDiag_62[45] , 
        \wPDiag_62[44] , \wPDiag_62[43] , \wPDiag_62[42] , \wPDiag_62[41] , 
        \wPDiag_62[40] , \wPDiag_62[39] , \wPDiag_62[38] , \wPDiag_62[37] , 
        \wPDiag_62[36] , \wPDiag_62[35] , \wPDiag_62[34] , \wPDiag_62[33] , 
        \wPDiag_62[32] , \wPDiag_62[31] , \wPDiag_62[30] , \wPDiag_62[29] , 
        \wPDiag_62[28] , \wPDiag_62[27] , \wPDiag_62[26] , \wPDiag_62[25] , 
        \wPDiag_62[24] , \wPDiag_62[23] , \wPDiag_62[22] , \wPDiag_62[21] , 
        \wPDiag_62[20] , \wPDiag_62[19] , \wPDiag_62[18] , \wPDiag_62[17] , 
        \wPDiag_62[16] , \wPDiag_62[15] , \wPDiag_62[14] , \wPDiag_62[13] , 
        \wPDiag_62[12] , \wPDiag_62[11] , \wPDiag_62[10] , \wPDiag_62[9] , 
        \wPDiag_62[8] , \wPDiag_62[7] , \wPDiag_62[6] , \wPDiag_62[5] , 
        \wPDiag_62[4] , \wPDiag_62[3] , \wPDiag_62[2] , \wPDiag_62[1] , 
        \wPDiag_62[0] }), .NDiagIn({\wNDiag_62[63] , \wNDiag_62[62] , 
        \wNDiag_62[61] , \wNDiag_62[60] , \wNDiag_62[59] , \wNDiag_62[58] , 
        \wNDiag_62[57] , \wNDiag_62[56] , \wNDiag_62[55] , \wNDiag_62[54] , 
        \wNDiag_62[53] , \wNDiag_62[52] , \wNDiag_62[51] , \wNDiag_62[50] , 
        \wNDiag_62[49] , \wNDiag_62[48] , \wNDiag_62[47] , \wNDiag_62[46] , 
        \wNDiag_62[45] , \wNDiag_62[44] , \wNDiag_62[43] , \wNDiag_62[42] , 
        \wNDiag_62[41] , \wNDiag_62[40] , \wNDiag_62[39] , \wNDiag_62[38] , 
        \wNDiag_62[37] , \wNDiag_62[36] , \wNDiag_62[35] , \wNDiag_62[34] , 
        \wNDiag_62[33] , \wNDiag_62[32] , \wNDiag_62[31] , \wNDiag_62[30] , 
        \wNDiag_62[29] , \wNDiag_62[28] , \wNDiag_62[27] , \wNDiag_62[26] , 
        \wNDiag_62[25] , \wNDiag_62[24] , \wNDiag_62[23] , \wNDiag_62[22] , 
        \wNDiag_62[21] , \wNDiag_62[20] , \wNDiag_62[19] , \wNDiag_62[18] , 
        \wNDiag_62[17] , \wNDiag_62[16] , \wNDiag_62[15] , \wNDiag_62[14] , 
        \wNDiag_62[13] , \wNDiag_62[12] , \wNDiag_62[11] , \wNDiag_62[10] , 
        \wNDiag_62[9] , \wNDiag_62[8] , \wNDiag_62[7] , \wNDiag_62[6] , 
        \wNDiag_62[5] , \wNDiag_62[4] , \wNDiag_62[3] , \wNDiag_62[2] , 
        \wNDiag_62[1] , \wNDiag_62[0] }), .CallOut(\wCall_63[0] ), .ReturnOut(
        \wReturn_62[0] ), .ColOut({\wColumn_63[63] , \wColumn_63[62] , 
        \wColumn_63[61] , \wColumn_63[60] , \wColumn_63[59] , \wColumn_63[58] , 
        \wColumn_63[57] , \wColumn_63[56] , \wColumn_63[55] , \wColumn_63[54] , 
        \wColumn_63[53] , \wColumn_63[52] , \wColumn_63[51] , \wColumn_63[50] , 
        \wColumn_63[49] , \wColumn_63[48] , \wColumn_63[47] , \wColumn_63[46] , 
        \wColumn_63[45] , \wColumn_63[44] , \wColumn_63[43] , \wColumn_63[42] , 
        \wColumn_63[41] , \wColumn_63[40] , \wColumn_63[39] , \wColumn_63[38] , 
        \wColumn_63[37] , \wColumn_63[36] , \wColumn_63[35] , \wColumn_63[34] , 
        \wColumn_63[33] , \wColumn_63[32] , \wColumn_63[31] , \wColumn_63[30] , 
        \wColumn_63[29] , \wColumn_63[28] , \wColumn_63[27] , \wColumn_63[26] , 
        \wColumn_63[25] , \wColumn_63[24] , \wColumn_63[23] , \wColumn_63[22] , 
        \wColumn_63[21] , \wColumn_63[20] , \wColumn_63[19] , \wColumn_63[18] , 
        \wColumn_63[17] , \wColumn_63[16] , \wColumn_63[15] , \wColumn_63[14] , 
        \wColumn_63[13] , \wColumn_63[12] , \wColumn_63[11] , \wColumn_63[10] , 
        \wColumn_63[9] , \wColumn_63[8] , \wColumn_63[7] , \wColumn_63[6] , 
        \wColumn_63[5] , \wColumn_63[4] , \wColumn_63[3] , \wColumn_63[2] , 
        \wColumn_63[1] , \wColumn_63[0] }), .PDiagOut({\wPDiag_63[63] , 
        \wPDiag_63[62] , \wPDiag_63[61] , \wPDiag_63[60] , \wPDiag_63[59] , 
        \wPDiag_63[58] , \wPDiag_63[57] , \wPDiag_63[56] , \wPDiag_63[55] , 
        \wPDiag_63[54] , \wPDiag_63[53] , \wPDiag_63[52] , \wPDiag_63[51] , 
        \wPDiag_63[50] , \wPDiag_63[49] , \wPDiag_63[48] , \wPDiag_63[47] , 
        \wPDiag_63[46] , \wPDiag_63[45] , \wPDiag_63[44] , \wPDiag_63[43] , 
        \wPDiag_63[42] , \wPDiag_63[41] , \wPDiag_63[40] , \wPDiag_63[39] , 
        \wPDiag_63[38] , \wPDiag_63[37] , \wPDiag_63[36] , \wPDiag_63[35] , 
        \wPDiag_63[34] , \wPDiag_63[33] , \wPDiag_63[32] , \wPDiag_63[31] , 
        \wPDiag_63[30] , \wPDiag_63[29] , \wPDiag_63[28] , \wPDiag_63[27] , 
        \wPDiag_63[26] , \wPDiag_63[25] , \wPDiag_63[24] , \wPDiag_63[23] , 
        \wPDiag_63[22] , \wPDiag_63[21] , \wPDiag_63[20] , \wPDiag_63[19] , 
        \wPDiag_63[18] , \wPDiag_63[17] , \wPDiag_63[16] , \wPDiag_63[15] , 
        \wPDiag_63[14] , \wPDiag_63[13] , \wPDiag_63[12] , \wPDiag_63[11] , 
        \wPDiag_63[10] , \wPDiag_63[9] , \wPDiag_63[8] , \wPDiag_63[7] , 
        \wPDiag_63[6] , \wPDiag_63[5] , \wPDiag_63[4] , \wPDiag_63[3] , 
        \wPDiag_63[2] , \wPDiag_63[1] , \wPDiag_63[0] }), .NDiagOut({
        \wNDiag_63[63] , \wNDiag_63[62] , \wNDiag_63[61] , \wNDiag_63[60] , 
        \wNDiag_63[59] , \wNDiag_63[58] , \wNDiag_63[57] , \wNDiag_63[56] , 
        \wNDiag_63[55] , \wNDiag_63[54] , \wNDiag_63[53] , \wNDiag_63[52] , 
        \wNDiag_63[51] , \wNDiag_63[50] , \wNDiag_63[49] , \wNDiag_63[48] , 
        \wNDiag_63[47] , \wNDiag_63[46] , \wNDiag_63[45] , \wNDiag_63[44] , 
        \wNDiag_63[43] , \wNDiag_63[42] , \wNDiag_63[41] , \wNDiag_63[40] , 
        \wNDiag_63[39] , \wNDiag_63[38] , \wNDiag_63[37] , \wNDiag_63[36] , 
        \wNDiag_63[35] , \wNDiag_63[34] , \wNDiag_63[33] , \wNDiag_63[32] , 
        \wNDiag_63[31] , \wNDiag_63[30] , \wNDiag_63[29] , \wNDiag_63[28] , 
        \wNDiag_63[27] , \wNDiag_63[26] , \wNDiag_63[25] , \wNDiag_63[24] , 
        \wNDiag_63[23] , \wNDiag_63[22] , \wNDiag_63[21] , \wNDiag_63[20] , 
        \wNDiag_63[19] , \wNDiag_63[18] , \wNDiag_63[17] , \wNDiag_63[16] , 
        \wNDiag_63[15] , \wNDiag_63[14] , \wNDiag_63[13] , \wNDiag_63[12] , 
        \wNDiag_63[11] , \wNDiag_63[10] , \wNDiag_63[9] , \wNDiag_63[8] , 
        \wNDiag_63[7] , \wNDiag_63[6] , \wNDiag_63[5] , \wNDiag_63[4] , 
        \wNDiag_63[3] , \wNDiag_63[2] , \wNDiag_63[1] , \wNDiag_63[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_37 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_38[6] , \wScan_38[5] , \wScan_38[4] , 
        \wScan_38[3] , \wScan_38[2] , \wScan_38[1] , \wScan_38[0] }), 
        .ScanOut({\wScan_37[6] , \wScan_37[5] , \wScan_37[4] , \wScan_37[3] , 
        \wScan_37[2] , \wScan_37[1] , \wScan_37[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_37[0] ), .ReturnIn(\wReturn_38[0] ), .ColIn({
        \wColumn_37[63] , \wColumn_37[62] , \wColumn_37[61] , \wColumn_37[60] , 
        \wColumn_37[59] , \wColumn_37[58] , \wColumn_37[57] , \wColumn_37[56] , 
        \wColumn_37[55] , \wColumn_37[54] , \wColumn_37[53] , \wColumn_37[52] , 
        \wColumn_37[51] , \wColumn_37[50] , \wColumn_37[49] , \wColumn_37[48] , 
        \wColumn_37[47] , \wColumn_37[46] , \wColumn_37[45] , \wColumn_37[44] , 
        \wColumn_37[43] , \wColumn_37[42] , \wColumn_37[41] , \wColumn_37[40] , 
        \wColumn_37[39] , \wColumn_37[38] , \wColumn_37[37] , \wColumn_37[36] , 
        \wColumn_37[35] , \wColumn_37[34] , \wColumn_37[33] , \wColumn_37[32] , 
        \wColumn_37[31] , \wColumn_37[30] , \wColumn_37[29] , \wColumn_37[28] , 
        \wColumn_37[27] , \wColumn_37[26] , \wColumn_37[25] , \wColumn_37[24] , 
        \wColumn_37[23] , \wColumn_37[22] , \wColumn_37[21] , \wColumn_37[20] , 
        \wColumn_37[19] , \wColumn_37[18] , \wColumn_37[17] , \wColumn_37[16] , 
        \wColumn_37[15] , \wColumn_37[14] , \wColumn_37[13] , \wColumn_37[12] , 
        \wColumn_37[11] , \wColumn_37[10] , \wColumn_37[9] , \wColumn_37[8] , 
        \wColumn_37[7] , \wColumn_37[6] , \wColumn_37[5] , \wColumn_37[4] , 
        \wColumn_37[3] , \wColumn_37[2] , \wColumn_37[1] , \wColumn_37[0] }), 
        .PDiagIn({\wPDiag_37[63] , \wPDiag_37[62] , \wPDiag_37[61] , 
        \wPDiag_37[60] , \wPDiag_37[59] , \wPDiag_37[58] , \wPDiag_37[57] , 
        \wPDiag_37[56] , \wPDiag_37[55] , \wPDiag_37[54] , \wPDiag_37[53] , 
        \wPDiag_37[52] , \wPDiag_37[51] , \wPDiag_37[50] , \wPDiag_37[49] , 
        \wPDiag_37[48] , \wPDiag_37[47] , \wPDiag_37[46] , \wPDiag_37[45] , 
        \wPDiag_37[44] , \wPDiag_37[43] , \wPDiag_37[42] , \wPDiag_37[41] , 
        \wPDiag_37[40] , \wPDiag_37[39] , \wPDiag_37[38] , \wPDiag_37[37] , 
        \wPDiag_37[36] , \wPDiag_37[35] , \wPDiag_37[34] , \wPDiag_37[33] , 
        \wPDiag_37[32] , \wPDiag_37[31] , \wPDiag_37[30] , \wPDiag_37[29] , 
        \wPDiag_37[28] , \wPDiag_37[27] , \wPDiag_37[26] , \wPDiag_37[25] , 
        \wPDiag_37[24] , \wPDiag_37[23] , \wPDiag_37[22] , \wPDiag_37[21] , 
        \wPDiag_37[20] , \wPDiag_37[19] , \wPDiag_37[18] , \wPDiag_37[17] , 
        \wPDiag_37[16] , \wPDiag_37[15] , \wPDiag_37[14] , \wPDiag_37[13] , 
        \wPDiag_37[12] , \wPDiag_37[11] , \wPDiag_37[10] , \wPDiag_37[9] , 
        \wPDiag_37[8] , \wPDiag_37[7] , \wPDiag_37[6] , \wPDiag_37[5] , 
        \wPDiag_37[4] , \wPDiag_37[3] , \wPDiag_37[2] , \wPDiag_37[1] , 
        \wPDiag_37[0] }), .NDiagIn({\wNDiag_37[63] , \wNDiag_37[62] , 
        \wNDiag_37[61] , \wNDiag_37[60] , \wNDiag_37[59] , \wNDiag_37[58] , 
        \wNDiag_37[57] , \wNDiag_37[56] , \wNDiag_37[55] , \wNDiag_37[54] , 
        \wNDiag_37[53] , \wNDiag_37[52] , \wNDiag_37[51] , \wNDiag_37[50] , 
        \wNDiag_37[49] , \wNDiag_37[48] , \wNDiag_37[47] , \wNDiag_37[46] , 
        \wNDiag_37[45] , \wNDiag_37[44] , \wNDiag_37[43] , \wNDiag_37[42] , 
        \wNDiag_37[41] , \wNDiag_37[40] , \wNDiag_37[39] , \wNDiag_37[38] , 
        \wNDiag_37[37] , \wNDiag_37[36] , \wNDiag_37[35] , \wNDiag_37[34] , 
        \wNDiag_37[33] , \wNDiag_37[32] , \wNDiag_37[31] , \wNDiag_37[30] , 
        \wNDiag_37[29] , \wNDiag_37[28] , \wNDiag_37[27] , \wNDiag_37[26] , 
        \wNDiag_37[25] , \wNDiag_37[24] , \wNDiag_37[23] , \wNDiag_37[22] , 
        \wNDiag_37[21] , \wNDiag_37[20] , \wNDiag_37[19] , \wNDiag_37[18] , 
        \wNDiag_37[17] , \wNDiag_37[16] , \wNDiag_37[15] , \wNDiag_37[14] , 
        \wNDiag_37[13] , \wNDiag_37[12] , \wNDiag_37[11] , \wNDiag_37[10] , 
        \wNDiag_37[9] , \wNDiag_37[8] , \wNDiag_37[7] , \wNDiag_37[6] , 
        \wNDiag_37[5] , \wNDiag_37[4] , \wNDiag_37[3] , \wNDiag_37[2] , 
        \wNDiag_37[1] , \wNDiag_37[0] }), .CallOut(\wCall_38[0] ), .ReturnOut(
        \wReturn_37[0] ), .ColOut({\wColumn_38[63] , \wColumn_38[62] , 
        \wColumn_38[61] , \wColumn_38[60] , \wColumn_38[59] , \wColumn_38[58] , 
        \wColumn_38[57] , \wColumn_38[56] , \wColumn_38[55] , \wColumn_38[54] , 
        \wColumn_38[53] , \wColumn_38[52] , \wColumn_38[51] , \wColumn_38[50] , 
        \wColumn_38[49] , \wColumn_38[48] , \wColumn_38[47] , \wColumn_38[46] , 
        \wColumn_38[45] , \wColumn_38[44] , \wColumn_38[43] , \wColumn_38[42] , 
        \wColumn_38[41] , \wColumn_38[40] , \wColumn_38[39] , \wColumn_38[38] , 
        \wColumn_38[37] , \wColumn_38[36] , \wColumn_38[35] , \wColumn_38[34] , 
        \wColumn_38[33] , \wColumn_38[32] , \wColumn_38[31] , \wColumn_38[30] , 
        \wColumn_38[29] , \wColumn_38[28] , \wColumn_38[27] , \wColumn_38[26] , 
        \wColumn_38[25] , \wColumn_38[24] , \wColumn_38[23] , \wColumn_38[22] , 
        \wColumn_38[21] , \wColumn_38[20] , \wColumn_38[19] , \wColumn_38[18] , 
        \wColumn_38[17] , \wColumn_38[16] , \wColumn_38[15] , \wColumn_38[14] , 
        \wColumn_38[13] , \wColumn_38[12] , \wColumn_38[11] , \wColumn_38[10] , 
        \wColumn_38[9] , \wColumn_38[8] , \wColumn_38[7] , \wColumn_38[6] , 
        \wColumn_38[5] , \wColumn_38[4] , \wColumn_38[3] , \wColumn_38[2] , 
        \wColumn_38[1] , \wColumn_38[0] }), .PDiagOut({\wPDiag_38[63] , 
        \wPDiag_38[62] , \wPDiag_38[61] , \wPDiag_38[60] , \wPDiag_38[59] , 
        \wPDiag_38[58] , \wPDiag_38[57] , \wPDiag_38[56] , \wPDiag_38[55] , 
        \wPDiag_38[54] , \wPDiag_38[53] , \wPDiag_38[52] , \wPDiag_38[51] , 
        \wPDiag_38[50] , \wPDiag_38[49] , \wPDiag_38[48] , \wPDiag_38[47] , 
        \wPDiag_38[46] , \wPDiag_38[45] , \wPDiag_38[44] , \wPDiag_38[43] , 
        \wPDiag_38[42] , \wPDiag_38[41] , \wPDiag_38[40] , \wPDiag_38[39] , 
        \wPDiag_38[38] , \wPDiag_38[37] , \wPDiag_38[36] , \wPDiag_38[35] , 
        \wPDiag_38[34] , \wPDiag_38[33] , \wPDiag_38[32] , \wPDiag_38[31] , 
        \wPDiag_38[30] , \wPDiag_38[29] , \wPDiag_38[28] , \wPDiag_38[27] , 
        \wPDiag_38[26] , \wPDiag_38[25] , \wPDiag_38[24] , \wPDiag_38[23] , 
        \wPDiag_38[22] , \wPDiag_38[21] , \wPDiag_38[20] , \wPDiag_38[19] , 
        \wPDiag_38[18] , \wPDiag_38[17] , \wPDiag_38[16] , \wPDiag_38[15] , 
        \wPDiag_38[14] , \wPDiag_38[13] , \wPDiag_38[12] , \wPDiag_38[11] , 
        \wPDiag_38[10] , \wPDiag_38[9] , \wPDiag_38[8] , \wPDiag_38[7] , 
        \wPDiag_38[6] , \wPDiag_38[5] , \wPDiag_38[4] , \wPDiag_38[3] , 
        \wPDiag_38[2] , \wPDiag_38[1] , \wPDiag_38[0] }), .NDiagOut({
        \wNDiag_38[63] , \wNDiag_38[62] , \wNDiag_38[61] , \wNDiag_38[60] , 
        \wNDiag_38[59] , \wNDiag_38[58] , \wNDiag_38[57] , \wNDiag_38[56] , 
        \wNDiag_38[55] , \wNDiag_38[54] , \wNDiag_38[53] , \wNDiag_38[52] , 
        \wNDiag_38[51] , \wNDiag_38[50] , \wNDiag_38[49] , \wNDiag_38[48] , 
        \wNDiag_38[47] , \wNDiag_38[46] , \wNDiag_38[45] , \wNDiag_38[44] , 
        \wNDiag_38[43] , \wNDiag_38[42] , \wNDiag_38[41] , \wNDiag_38[40] , 
        \wNDiag_38[39] , \wNDiag_38[38] , \wNDiag_38[37] , \wNDiag_38[36] , 
        \wNDiag_38[35] , \wNDiag_38[34] , \wNDiag_38[33] , \wNDiag_38[32] , 
        \wNDiag_38[31] , \wNDiag_38[30] , \wNDiag_38[29] , \wNDiag_38[28] , 
        \wNDiag_38[27] , \wNDiag_38[26] , \wNDiag_38[25] , \wNDiag_38[24] , 
        \wNDiag_38[23] , \wNDiag_38[22] , \wNDiag_38[21] , \wNDiag_38[20] , 
        \wNDiag_38[19] , \wNDiag_38[18] , \wNDiag_38[17] , \wNDiag_38[16] , 
        \wNDiag_38[15] , \wNDiag_38[14] , \wNDiag_38[13] , \wNDiag_38[12] , 
        \wNDiag_38[11] , \wNDiag_38[10] , \wNDiag_38[9] , \wNDiag_38[8] , 
        \wNDiag_38[7] , \wNDiag_38[6] , \wNDiag_38[5] , \wNDiag_38[4] , 
        \wNDiag_38[3] , \wNDiag_38[2] , \wNDiag_38[1] , \wNDiag_38[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_59 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_60[6] , \wScan_60[5] , \wScan_60[4] , 
        \wScan_60[3] , \wScan_60[2] , \wScan_60[1] , \wScan_60[0] }), 
        .ScanOut({\wScan_59[6] , \wScan_59[5] , \wScan_59[4] , \wScan_59[3] , 
        \wScan_59[2] , \wScan_59[1] , \wScan_59[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_59[0] ), .ReturnIn(\wReturn_60[0] ), .ColIn({
        \wColumn_59[63] , \wColumn_59[62] , \wColumn_59[61] , \wColumn_59[60] , 
        \wColumn_59[59] , \wColumn_59[58] , \wColumn_59[57] , \wColumn_59[56] , 
        \wColumn_59[55] , \wColumn_59[54] , \wColumn_59[53] , \wColumn_59[52] , 
        \wColumn_59[51] , \wColumn_59[50] , \wColumn_59[49] , \wColumn_59[48] , 
        \wColumn_59[47] , \wColumn_59[46] , \wColumn_59[45] , \wColumn_59[44] , 
        \wColumn_59[43] , \wColumn_59[42] , \wColumn_59[41] , \wColumn_59[40] , 
        \wColumn_59[39] , \wColumn_59[38] , \wColumn_59[37] , \wColumn_59[36] , 
        \wColumn_59[35] , \wColumn_59[34] , \wColumn_59[33] , \wColumn_59[32] , 
        \wColumn_59[31] , \wColumn_59[30] , \wColumn_59[29] , \wColumn_59[28] , 
        \wColumn_59[27] , \wColumn_59[26] , \wColumn_59[25] , \wColumn_59[24] , 
        \wColumn_59[23] , \wColumn_59[22] , \wColumn_59[21] , \wColumn_59[20] , 
        \wColumn_59[19] , \wColumn_59[18] , \wColumn_59[17] , \wColumn_59[16] , 
        \wColumn_59[15] , \wColumn_59[14] , \wColumn_59[13] , \wColumn_59[12] , 
        \wColumn_59[11] , \wColumn_59[10] , \wColumn_59[9] , \wColumn_59[8] , 
        \wColumn_59[7] , \wColumn_59[6] , \wColumn_59[5] , \wColumn_59[4] , 
        \wColumn_59[3] , \wColumn_59[2] , \wColumn_59[1] , \wColumn_59[0] }), 
        .PDiagIn({\wPDiag_59[63] , \wPDiag_59[62] , \wPDiag_59[61] , 
        \wPDiag_59[60] , \wPDiag_59[59] , \wPDiag_59[58] , \wPDiag_59[57] , 
        \wPDiag_59[56] , \wPDiag_59[55] , \wPDiag_59[54] , \wPDiag_59[53] , 
        \wPDiag_59[52] , \wPDiag_59[51] , \wPDiag_59[50] , \wPDiag_59[49] , 
        \wPDiag_59[48] , \wPDiag_59[47] , \wPDiag_59[46] , \wPDiag_59[45] , 
        \wPDiag_59[44] , \wPDiag_59[43] , \wPDiag_59[42] , \wPDiag_59[41] , 
        \wPDiag_59[40] , \wPDiag_59[39] , \wPDiag_59[38] , \wPDiag_59[37] , 
        \wPDiag_59[36] , \wPDiag_59[35] , \wPDiag_59[34] , \wPDiag_59[33] , 
        \wPDiag_59[32] , \wPDiag_59[31] , \wPDiag_59[30] , \wPDiag_59[29] , 
        \wPDiag_59[28] , \wPDiag_59[27] , \wPDiag_59[26] , \wPDiag_59[25] , 
        \wPDiag_59[24] , \wPDiag_59[23] , \wPDiag_59[22] , \wPDiag_59[21] , 
        \wPDiag_59[20] , \wPDiag_59[19] , \wPDiag_59[18] , \wPDiag_59[17] , 
        \wPDiag_59[16] , \wPDiag_59[15] , \wPDiag_59[14] , \wPDiag_59[13] , 
        \wPDiag_59[12] , \wPDiag_59[11] , \wPDiag_59[10] , \wPDiag_59[9] , 
        \wPDiag_59[8] , \wPDiag_59[7] , \wPDiag_59[6] , \wPDiag_59[5] , 
        \wPDiag_59[4] , \wPDiag_59[3] , \wPDiag_59[2] , \wPDiag_59[1] , 
        \wPDiag_59[0] }), .NDiagIn({\wNDiag_59[63] , \wNDiag_59[62] , 
        \wNDiag_59[61] , \wNDiag_59[60] , \wNDiag_59[59] , \wNDiag_59[58] , 
        \wNDiag_59[57] , \wNDiag_59[56] , \wNDiag_59[55] , \wNDiag_59[54] , 
        \wNDiag_59[53] , \wNDiag_59[52] , \wNDiag_59[51] , \wNDiag_59[50] , 
        \wNDiag_59[49] , \wNDiag_59[48] , \wNDiag_59[47] , \wNDiag_59[46] , 
        \wNDiag_59[45] , \wNDiag_59[44] , \wNDiag_59[43] , \wNDiag_59[42] , 
        \wNDiag_59[41] , \wNDiag_59[40] , \wNDiag_59[39] , \wNDiag_59[38] , 
        \wNDiag_59[37] , \wNDiag_59[36] , \wNDiag_59[35] , \wNDiag_59[34] , 
        \wNDiag_59[33] , \wNDiag_59[32] , \wNDiag_59[31] , \wNDiag_59[30] , 
        \wNDiag_59[29] , \wNDiag_59[28] , \wNDiag_59[27] , \wNDiag_59[26] , 
        \wNDiag_59[25] , \wNDiag_59[24] , \wNDiag_59[23] , \wNDiag_59[22] , 
        \wNDiag_59[21] , \wNDiag_59[20] , \wNDiag_59[19] , \wNDiag_59[18] , 
        \wNDiag_59[17] , \wNDiag_59[16] , \wNDiag_59[15] , \wNDiag_59[14] , 
        \wNDiag_59[13] , \wNDiag_59[12] , \wNDiag_59[11] , \wNDiag_59[10] , 
        \wNDiag_59[9] , \wNDiag_59[8] , \wNDiag_59[7] , \wNDiag_59[6] , 
        \wNDiag_59[5] , \wNDiag_59[4] , \wNDiag_59[3] , \wNDiag_59[2] , 
        \wNDiag_59[1] , \wNDiag_59[0] }), .CallOut(\wCall_60[0] ), .ReturnOut(
        \wReturn_59[0] ), .ColOut({\wColumn_60[63] , \wColumn_60[62] , 
        \wColumn_60[61] , \wColumn_60[60] , \wColumn_60[59] , \wColumn_60[58] , 
        \wColumn_60[57] , \wColumn_60[56] , \wColumn_60[55] , \wColumn_60[54] , 
        \wColumn_60[53] , \wColumn_60[52] , \wColumn_60[51] , \wColumn_60[50] , 
        \wColumn_60[49] , \wColumn_60[48] , \wColumn_60[47] , \wColumn_60[46] , 
        \wColumn_60[45] , \wColumn_60[44] , \wColumn_60[43] , \wColumn_60[42] , 
        \wColumn_60[41] , \wColumn_60[40] , \wColumn_60[39] , \wColumn_60[38] , 
        \wColumn_60[37] , \wColumn_60[36] , \wColumn_60[35] , \wColumn_60[34] , 
        \wColumn_60[33] , \wColumn_60[32] , \wColumn_60[31] , \wColumn_60[30] , 
        \wColumn_60[29] , \wColumn_60[28] , \wColumn_60[27] , \wColumn_60[26] , 
        \wColumn_60[25] , \wColumn_60[24] , \wColumn_60[23] , \wColumn_60[22] , 
        \wColumn_60[21] , \wColumn_60[20] , \wColumn_60[19] , \wColumn_60[18] , 
        \wColumn_60[17] , \wColumn_60[16] , \wColumn_60[15] , \wColumn_60[14] , 
        \wColumn_60[13] , \wColumn_60[12] , \wColumn_60[11] , \wColumn_60[10] , 
        \wColumn_60[9] , \wColumn_60[8] , \wColumn_60[7] , \wColumn_60[6] , 
        \wColumn_60[5] , \wColumn_60[4] , \wColumn_60[3] , \wColumn_60[2] , 
        \wColumn_60[1] , \wColumn_60[0] }), .PDiagOut({\wPDiag_60[63] , 
        \wPDiag_60[62] , \wPDiag_60[61] , \wPDiag_60[60] , \wPDiag_60[59] , 
        \wPDiag_60[58] , \wPDiag_60[57] , \wPDiag_60[56] , \wPDiag_60[55] , 
        \wPDiag_60[54] , \wPDiag_60[53] , \wPDiag_60[52] , \wPDiag_60[51] , 
        \wPDiag_60[50] , \wPDiag_60[49] , \wPDiag_60[48] , \wPDiag_60[47] , 
        \wPDiag_60[46] , \wPDiag_60[45] , \wPDiag_60[44] , \wPDiag_60[43] , 
        \wPDiag_60[42] , \wPDiag_60[41] , \wPDiag_60[40] , \wPDiag_60[39] , 
        \wPDiag_60[38] , \wPDiag_60[37] , \wPDiag_60[36] , \wPDiag_60[35] , 
        \wPDiag_60[34] , \wPDiag_60[33] , \wPDiag_60[32] , \wPDiag_60[31] , 
        \wPDiag_60[30] , \wPDiag_60[29] , \wPDiag_60[28] , \wPDiag_60[27] , 
        \wPDiag_60[26] , \wPDiag_60[25] , \wPDiag_60[24] , \wPDiag_60[23] , 
        \wPDiag_60[22] , \wPDiag_60[21] , \wPDiag_60[20] , \wPDiag_60[19] , 
        \wPDiag_60[18] , \wPDiag_60[17] , \wPDiag_60[16] , \wPDiag_60[15] , 
        \wPDiag_60[14] , \wPDiag_60[13] , \wPDiag_60[12] , \wPDiag_60[11] , 
        \wPDiag_60[10] , \wPDiag_60[9] , \wPDiag_60[8] , \wPDiag_60[7] , 
        \wPDiag_60[6] , \wPDiag_60[5] , \wPDiag_60[4] , \wPDiag_60[3] , 
        \wPDiag_60[2] , \wPDiag_60[1] , \wPDiag_60[0] }), .NDiagOut({
        \wNDiag_60[63] , \wNDiag_60[62] , \wNDiag_60[61] , \wNDiag_60[60] , 
        \wNDiag_60[59] , \wNDiag_60[58] , \wNDiag_60[57] , \wNDiag_60[56] , 
        \wNDiag_60[55] , \wNDiag_60[54] , \wNDiag_60[53] , \wNDiag_60[52] , 
        \wNDiag_60[51] , \wNDiag_60[50] , \wNDiag_60[49] , \wNDiag_60[48] , 
        \wNDiag_60[47] , \wNDiag_60[46] , \wNDiag_60[45] , \wNDiag_60[44] , 
        \wNDiag_60[43] , \wNDiag_60[42] , \wNDiag_60[41] , \wNDiag_60[40] , 
        \wNDiag_60[39] , \wNDiag_60[38] , \wNDiag_60[37] , \wNDiag_60[36] , 
        \wNDiag_60[35] , \wNDiag_60[34] , \wNDiag_60[33] , \wNDiag_60[32] , 
        \wNDiag_60[31] , \wNDiag_60[30] , \wNDiag_60[29] , \wNDiag_60[28] , 
        \wNDiag_60[27] , \wNDiag_60[26] , \wNDiag_60[25] , \wNDiag_60[24] , 
        \wNDiag_60[23] , \wNDiag_60[22] , \wNDiag_60[21] , \wNDiag_60[20] , 
        \wNDiag_60[19] , \wNDiag_60[18] , \wNDiag_60[17] , \wNDiag_60[16] , 
        \wNDiag_60[15] , \wNDiag_60[14] , \wNDiag_60[13] , \wNDiag_60[12] , 
        \wNDiag_60[11] , \wNDiag_60[10] , \wNDiag_60[9] , \wNDiag_60[8] , 
        \wNDiag_60[7] , \wNDiag_60[6] , \wNDiag_60[5] , \wNDiag_60[4] , 
        \wNDiag_60[3] , \wNDiag_60[2] , \wNDiag_60[1] , \wNDiag_60[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_19 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_20[6] , \wScan_20[5] , \wScan_20[4] , 
        \wScan_20[3] , \wScan_20[2] , \wScan_20[1] , \wScan_20[0] }), 
        .ScanOut({\wScan_19[6] , \wScan_19[5] , \wScan_19[4] , \wScan_19[3] , 
        \wScan_19[2] , \wScan_19[1] , \wScan_19[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_19[0] ), .ReturnIn(\wReturn_20[0] ), .ColIn({
        \wColumn_19[63] , \wColumn_19[62] , \wColumn_19[61] , \wColumn_19[60] , 
        \wColumn_19[59] , \wColumn_19[58] , \wColumn_19[57] , \wColumn_19[56] , 
        \wColumn_19[55] , \wColumn_19[54] , \wColumn_19[53] , \wColumn_19[52] , 
        \wColumn_19[51] , \wColumn_19[50] , \wColumn_19[49] , \wColumn_19[48] , 
        \wColumn_19[47] , \wColumn_19[46] , \wColumn_19[45] , \wColumn_19[44] , 
        \wColumn_19[43] , \wColumn_19[42] , \wColumn_19[41] , \wColumn_19[40] , 
        \wColumn_19[39] , \wColumn_19[38] , \wColumn_19[37] , \wColumn_19[36] , 
        \wColumn_19[35] , \wColumn_19[34] , \wColumn_19[33] , \wColumn_19[32] , 
        \wColumn_19[31] , \wColumn_19[30] , \wColumn_19[29] , \wColumn_19[28] , 
        \wColumn_19[27] , \wColumn_19[26] , \wColumn_19[25] , \wColumn_19[24] , 
        \wColumn_19[23] , \wColumn_19[22] , \wColumn_19[21] , \wColumn_19[20] , 
        \wColumn_19[19] , \wColumn_19[18] , \wColumn_19[17] , \wColumn_19[16] , 
        \wColumn_19[15] , \wColumn_19[14] , \wColumn_19[13] , \wColumn_19[12] , 
        \wColumn_19[11] , \wColumn_19[10] , \wColumn_19[9] , \wColumn_19[8] , 
        \wColumn_19[7] , \wColumn_19[6] , \wColumn_19[5] , \wColumn_19[4] , 
        \wColumn_19[3] , \wColumn_19[2] , \wColumn_19[1] , \wColumn_19[0] }), 
        .PDiagIn({\wPDiag_19[63] , \wPDiag_19[62] , \wPDiag_19[61] , 
        \wPDiag_19[60] , \wPDiag_19[59] , \wPDiag_19[58] , \wPDiag_19[57] , 
        \wPDiag_19[56] , \wPDiag_19[55] , \wPDiag_19[54] , \wPDiag_19[53] , 
        \wPDiag_19[52] , \wPDiag_19[51] , \wPDiag_19[50] , \wPDiag_19[49] , 
        \wPDiag_19[48] , \wPDiag_19[47] , \wPDiag_19[46] , \wPDiag_19[45] , 
        \wPDiag_19[44] , \wPDiag_19[43] , \wPDiag_19[42] , \wPDiag_19[41] , 
        \wPDiag_19[40] , \wPDiag_19[39] , \wPDiag_19[38] , \wPDiag_19[37] , 
        \wPDiag_19[36] , \wPDiag_19[35] , \wPDiag_19[34] , \wPDiag_19[33] , 
        \wPDiag_19[32] , \wPDiag_19[31] , \wPDiag_19[30] , \wPDiag_19[29] , 
        \wPDiag_19[28] , \wPDiag_19[27] , \wPDiag_19[26] , \wPDiag_19[25] , 
        \wPDiag_19[24] , \wPDiag_19[23] , \wPDiag_19[22] , \wPDiag_19[21] , 
        \wPDiag_19[20] , \wPDiag_19[19] , \wPDiag_19[18] , \wPDiag_19[17] , 
        \wPDiag_19[16] , \wPDiag_19[15] , \wPDiag_19[14] , \wPDiag_19[13] , 
        \wPDiag_19[12] , \wPDiag_19[11] , \wPDiag_19[10] , \wPDiag_19[9] , 
        \wPDiag_19[8] , \wPDiag_19[7] , \wPDiag_19[6] , \wPDiag_19[5] , 
        \wPDiag_19[4] , \wPDiag_19[3] , \wPDiag_19[2] , \wPDiag_19[1] , 
        \wPDiag_19[0] }), .NDiagIn({\wNDiag_19[63] , \wNDiag_19[62] , 
        \wNDiag_19[61] , \wNDiag_19[60] , \wNDiag_19[59] , \wNDiag_19[58] , 
        \wNDiag_19[57] , \wNDiag_19[56] , \wNDiag_19[55] , \wNDiag_19[54] , 
        \wNDiag_19[53] , \wNDiag_19[52] , \wNDiag_19[51] , \wNDiag_19[50] , 
        \wNDiag_19[49] , \wNDiag_19[48] , \wNDiag_19[47] , \wNDiag_19[46] , 
        \wNDiag_19[45] , \wNDiag_19[44] , \wNDiag_19[43] , \wNDiag_19[42] , 
        \wNDiag_19[41] , \wNDiag_19[40] , \wNDiag_19[39] , \wNDiag_19[38] , 
        \wNDiag_19[37] , \wNDiag_19[36] , \wNDiag_19[35] , \wNDiag_19[34] , 
        \wNDiag_19[33] , \wNDiag_19[32] , \wNDiag_19[31] , \wNDiag_19[30] , 
        \wNDiag_19[29] , \wNDiag_19[28] , \wNDiag_19[27] , \wNDiag_19[26] , 
        \wNDiag_19[25] , \wNDiag_19[24] , \wNDiag_19[23] , \wNDiag_19[22] , 
        \wNDiag_19[21] , \wNDiag_19[20] , \wNDiag_19[19] , \wNDiag_19[18] , 
        \wNDiag_19[17] , \wNDiag_19[16] , \wNDiag_19[15] , \wNDiag_19[14] , 
        \wNDiag_19[13] , \wNDiag_19[12] , \wNDiag_19[11] , \wNDiag_19[10] , 
        \wNDiag_19[9] , \wNDiag_19[8] , \wNDiag_19[7] , \wNDiag_19[6] , 
        \wNDiag_19[5] , \wNDiag_19[4] , \wNDiag_19[3] , \wNDiag_19[2] , 
        \wNDiag_19[1] , \wNDiag_19[0] }), .CallOut(\wCall_20[0] ), .ReturnOut(
        \wReturn_19[0] ), .ColOut({\wColumn_20[63] , \wColumn_20[62] , 
        \wColumn_20[61] , \wColumn_20[60] , \wColumn_20[59] , \wColumn_20[58] , 
        \wColumn_20[57] , \wColumn_20[56] , \wColumn_20[55] , \wColumn_20[54] , 
        \wColumn_20[53] , \wColumn_20[52] , \wColumn_20[51] , \wColumn_20[50] , 
        \wColumn_20[49] , \wColumn_20[48] , \wColumn_20[47] , \wColumn_20[46] , 
        \wColumn_20[45] , \wColumn_20[44] , \wColumn_20[43] , \wColumn_20[42] , 
        \wColumn_20[41] , \wColumn_20[40] , \wColumn_20[39] , \wColumn_20[38] , 
        \wColumn_20[37] , \wColumn_20[36] , \wColumn_20[35] , \wColumn_20[34] , 
        \wColumn_20[33] , \wColumn_20[32] , \wColumn_20[31] , \wColumn_20[30] , 
        \wColumn_20[29] , \wColumn_20[28] , \wColumn_20[27] , \wColumn_20[26] , 
        \wColumn_20[25] , \wColumn_20[24] , \wColumn_20[23] , \wColumn_20[22] , 
        \wColumn_20[21] , \wColumn_20[20] , \wColumn_20[19] , \wColumn_20[18] , 
        \wColumn_20[17] , \wColumn_20[16] , \wColumn_20[15] , \wColumn_20[14] , 
        \wColumn_20[13] , \wColumn_20[12] , \wColumn_20[11] , \wColumn_20[10] , 
        \wColumn_20[9] , \wColumn_20[8] , \wColumn_20[7] , \wColumn_20[6] , 
        \wColumn_20[5] , \wColumn_20[4] , \wColumn_20[3] , \wColumn_20[2] , 
        \wColumn_20[1] , \wColumn_20[0] }), .PDiagOut({\wPDiag_20[63] , 
        \wPDiag_20[62] , \wPDiag_20[61] , \wPDiag_20[60] , \wPDiag_20[59] , 
        \wPDiag_20[58] , \wPDiag_20[57] , \wPDiag_20[56] , \wPDiag_20[55] , 
        \wPDiag_20[54] , \wPDiag_20[53] , \wPDiag_20[52] , \wPDiag_20[51] , 
        \wPDiag_20[50] , \wPDiag_20[49] , \wPDiag_20[48] , \wPDiag_20[47] , 
        \wPDiag_20[46] , \wPDiag_20[45] , \wPDiag_20[44] , \wPDiag_20[43] , 
        \wPDiag_20[42] , \wPDiag_20[41] , \wPDiag_20[40] , \wPDiag_20[39] , 
        \wPDiag_20[38] , \wPDiag_20[37] , \wPDiag_20[36] , \wPDiag_20[35] , 
        \wPDiag_20[34] , \wPDiag_20[33] , \wPDiag_20[32] , \wPDiag_20[31] , 
        \wPDiag_20[30] , \wPDiag_20[29] , \wPDiag_20[28] , \wPDiag_20[27] , 
        \wPDiag_20[26] , \wPDiag_20[25] , \wPDiag_20[24] , \wPDiag_20[23] , 
        \wPDiag_20[22] , \wPDiag_20[21] , \wPDiag_20[20] , \wPDiag_20[19] , 
        \wPDiag_20[18] , \wPDiag_20[17] , \wPDiag_20[16] , \wPDiag_20[15] , 
        \wPDiag_20[14] , \wPDiag_20[13] , \wPDiag_20[12] , \wPDiag_20[11] , 
        \wPDiag_20[10] , \wPDiag_20[9] , \wPDiag_20[8] , \wPDiag_20[7] , 
        \wPDiag_20[6] , \wPDiag_20[5] , \wPDiag_20[4] , \wPDiag_20[3] , 
        \wPDiag_20[2] , \wPDiag_20[1] , \wPDiag_20[0] }), .NDiagOut({
        \wNDiag_20[63] , \wNDiag_20[62] , \wNDiag_20[61] , \wNDiag_20[60] , 
        \wNDiag_20[59] , \wNDiag_20[58] , \wNDiag_20[57] , \wNDiag_20[56] , 
        \wNDiag_20[55] , \wNDiag_20[54] , \wNDiag_20[53] , \wNDiag_20[52] , 
        \wNDiag_20[51] , \wNDiag_20[50] , \wNDiag_20[49] , \wNDiag_20[48] , 
        \wNDiag_20[47] , \wNDiag_20[46] , \wNDiag_20[45] , \wNDiag_20[44] , 
        \wNDiag_20[43] , \wNDiag_20[42] , \wNDiag_20[41] , \wNDiag_20[40] , 
        \wNDiag_20[39] , \wNDiag_20[38] , \wNDiag_20[37] , \wNDiag_20[36] , 
        \wNDiag_20[35] , \wNDiag_20[34] , \wNDiag_20[33] , \wNDiag_20[32] , 
        \wNDiag_20[31] , \wNDiag_20[30] , \wNDiag_20[29] , \wNDiag_20[28] , 
        \wNDiag_20[27] , \wNDiag_20[26] , \wNDiag_20[25] , \wNDiag_20[24] , 
        \wNDiag_20[23] , \wNDiag_20[22] , \wNDiag_20[21] , \wNDiag_20[20] , 
        \wNDiag_20[19] , \wNDiag_20[18] , \wNDiag_20[17] , \wNDiag_20[16] , 
        \wNDiag_20[15] , \wNDiag_20[14] , \wNDiag_20[13] , \wNDiag_20[12] , 
        \wNDiag_20[11] , \wNDiag_20[10] , \wNDiag_20[9] , \wNDiag_20[8] , 
        \wNDiag_20[7] , \wNDiag_20[6] , \wNDiag_20[5] , \wNDiag_20[4] , 
        \wNDiag_20[3] , \wNDiag_20[2] , \wNDiag_20[1] , \wNDiag_20[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_42 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_43[6] , \wScan_43[5] , \wScan_43[4] , 
        \wScan_43[3] , \wScan_43[2] , \wScan_43[1] , \wScan_43[0] }), 
        .ScanOut({\wScan_42[6] , \wScan_42[5] , \wScan_42[4] , \wScan_42[3] , 
        \wScan_42[2] , \wScan_42[1] , \wScan_42[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_42[0] ), .ReturnIn(\wReturn_43[0] ), .ColIn({
        \wColumn_42[63] , \wColumn_42[62] , \wColumn_42[61] , \wColumn_42[60] , 
        \wColumn_42[59] , \wColumn_42[58] , \wColumn_42[57] , \wColumn_42[56] , 
        \wColumn_42[55] , \wColumn_42[54] , \wColumn_42[53] , \wColumn_42[52] , 
        \wColumn_42[51] , \wColumn_42[50] , \wColumn_42[49] , \wColumn_42[48] , 
        \wColumn_42[47] , \wColumn_42[46] , \wColumn_42[45] , \wColumn_42[44] , 
        \wColumn_42[43] , \wColumn_42[42] , \wColumn_42[41] , \wColumn_42[40] , 
        \wColumn_42[39] , \wColumn_42[38] , \wColumn_42[37] , \wColumn_42[36] , 
        \wColumn_42[35] , \wColumn_42[34] , \wColumn_42[33] , \wColumn_42[32] , 
        \wColumn_42[31] , \wColumn_42[30] , \wColumn_42[29] , \wColumn_42[28] , 
        \wColumn_42[27] , \wColumn_42[26] , \wColumn_42[25] , \wColumn_42[24] , 
        \wColumn_42[23] , \wColumn_42[22] , \wColumn_42[21] , \wColumn_42[20] , 
        \wColumn_42[19] , \wColumn_42[18] , \wColumn_42[17] , \wColumn_42[16] , 
        \wColumn_42[15] , \wColumn_42[14] , \wColumn_42[13] , \wColumn_42[12] , 
        \wColumn_42[11] , \wColumn_42[10] , \wColumn_42[9] , \wColumn_42[8] , 
        \wColumn_42[7] , \wColumn_42[6] , \wColumn_42[5] , \wColumn_42[4] , 
        \wColumn_42[3] , \wColumn_42[2] , \wColumn_42[1] , \wColumn_42[0] }), 
        .PDiagIn({\wPDiag_42[63] , \wPDiag_42[62] , \wPDiag_42[61] , 
        \wPDiag_42[60] , \wPDiag_42[59] , \wPDiag_42[58] , \wPDiag_42[57] , 
        \wPDiag_42[56] , \wPDiag_42[55] , \wPDiag_42[54] , \wPDiag_42[53] , 
        \wPDiag_42[52] , \wPDiag_42[51] , \wPDiag_42[50] , \wPDiag_42[49] , 
        \wPDiag_42[48] , \wPDiag_42[47] , \wPDiag_42[46] , \wPDiag_42[45] , 
        \wPDiag_42[44] , \wPDiag_42[43] , \wPDiag_42[42] , \wPDiag_42[41] , 
        \wPDiag_42[40] , \wPDiag_42[39] , \wPDiag_42[38] , \wPDiag_42[37] , 
        \wPDiag_42[36] , \wPDiag_42[35] , \wPDiag_42[34] , \wPDiag_42[33] , 
        \wPDiag_42[32] , \wPDiag_42[31] , \wPDiag_42[30] , \wPDiag_42[29] , 
        \wPDiag_42[28] , \wPDiag_42[27] , \wPDiag_42[26] , \wPDiag_42[25] , 
        \wPDiag_42[24] , \wPDiag_42[23] , \wPDiag_42[22] , \wPDiag_42[21] , 
        \wPDiag_42[20] , \wPDiag_42[19] , \wPDiag_42[18] , \wPDiag_42[17] , 
        \wPDiag_42[16] , \wPDiag_42[15] , \wPDiag_42[14] , \wPDiag_42[13] , 
        \wPDiag_42[12] , \wPDiag_42[11] , \wPDiag_42[10] , \wPDiag_42[9] , 
        \wPDiag_42[8] , \wPDiag_42[7] , \wPDiag_42[6] , \wPDiag_42[5] , 
        \wPDiag_42[4] , \wPDiag_42[3] , \wPDiag_42[2] , \wPDiag_42[1] , 
        \wPDiag_42[0] }), .NDiagIn({\wNDiag_42[63] , \wNDiag_42[62] , 
        \wNDiag_42[61] , \wNDiag_42[60] , \wNDiag_42[59] , \wNDiag_42[58] , 
        \wNDiag_42[57] , \wNDiag_42[56] , \wNDiag_42[55] , \wNDiag_42[54] , 
        \wNDiag_42[53] , \wNDiag_42[52] , \wNDiag_42[51] , \wNDiag_42[50] , 
        \wNDiag_42[49] , \wNDiag_42[48] , \wNDiag_42[47] , \wNDiag_42[46] , 
        \wNDiag_42[45] , \wNDiag_42[44] , \wNDiag_42[43] , \wNDiag_42[42] , 
        \wNDiag_42[41] , \wNDiag_42[40] , \wNDiag_42[39] , \wNDiag_42[38] , 
        \wNDiag_42[37] , \wNDiag_42[36] , \wNDiag_42[35] , \wNDiag_42[34] , 
        \wNDiag_42[33] , \wNDiag_42[32] , \wNDiag_42[31] , \wNDiag_42[30] , 
        \wNDiag_42[29] , \wNDiag_42[28] , \wNDiag_42[27] , \wNDiag_42[26] , 
        \wNDiag_42[25] , \wNDiag_42[24] , \wNDiag_42[23] , \wNDiag_42[22] , 
        \wNDiag_42[21] , \wNDiag_42[20] , \wNDiag_42[19] , \wNDiag_42[18] , 
        \wNDiag_42[17] , \wNDiag_42[16] , \wNDiag_42[15] , \wNDiag_42[14] , 
        \wNDiag_42[13] , \wNDiag_42[12] , \wNDiag_42[11] , \wNDiag_42[10] , 
        \wNDiag_42[9] , \wNDiag_42[8] , \wNDiag_42[7] , \wNDiag_42[6] , 
        \wNDiag_42[5] , \wNDiag_42[4] , \wNDiag_42[3] , \wNDiag_42[2] , 
        \wNDiag_42[1] , \wNDiag_42[0] }), .CallOut(\wCall_43[0] ), .ReturnOut(
        \wReturn_42[0] ), .ColOut({\wColumn_43[63] , \wColumn_43[62] , 
        \wColumn_43[61] , \wColumn_43[60] , \wColumn_43[59] , \wColumn_43[58] , 
        \wColumn_43[57] , \wColumn_43[56] , \wColumn_43[55] , \wColumn_43[54] , 
        \wColumn_43[53] , \wColumn_43[52] , \wColumn_43[51] , \wColumn_43[50] , 
        \wColumn_43[49] , \wColumn_43[48] , \wColumn_43[47] , \wColumn_43[46] , 
        \wColumn_43[45] , \wColumn_43[44] , \wColumn_43[43] , \wColumn_43[42] , 
        \wColumn_43[41] , \wColumn_43[40] , \wColumn_43[39] , \wColumn_43[38] , 
        \wColumn_43[37] , \wColumn_43[36] , \wColumn_43[35] , \wColumn_43[34] , 
        \wColumn_43[33] , \wColumn_43[32] , \wColumn_43[31] , \wColumn_43[30] , 
        \wColumn_43[29] , \wColumn_43[28] , \wColumn_43[27] , \wColumn_43[26] , 
        \wColumn_43[25] , \wColumn_43[24] , \wColumn_43[23] , \wColumn_43[22] , 
        \wColumn_43[21] , \wColumn_43[20] , \wColumn_43[19] , \wColumn_43[18] , 
        \wColumn_43[17] , \wColumn_43[16] , \wColumn_43[15] , \wColumn_43[14] , 
        \wColumn_43[13] , \wColumn_43[12] , \wColumn_43[11] , \wColumn_43[10] , 
        \wColumn_43[9] , \wColumn_43[8] , \wColumn_43[7] , \wColumn_43[6] , 
        \wColumn_43[5] , \wColumn_43[4] , \wColumn_43[3] , \wColumn_43[2] , 
        \wColumn_43[1] , \wColumn_43[0] }), .PDiagOut({\wPDiag_43[63] , 
        \wPDiag_43[62] , \wPDiag_43[61] , \wPDiag_43[60] , \wPDiag_43[59] , 
        \wPDiag_43[58] , \wPDiag_43[57] , \wPDiag_43[56] , \wPDiag_43[55] , 
        \wPDiag_43[54] , \wPDiag_43[53] , \wPDiag_43[52] , \wPDiag_43[51] , 
        \wPDiag_43[50] , \wPDiag_43[49] , \wPDiag_43[48] , \wPDiag_43[47] , 
        \wPDiag_43[46] , \wPDiag_43[45] , \wPDiag_43[44] , \wPDiag_43[43] , 
        \wPDiag_43[42] , \wPDiag_43[41] , \wPDiag_43[40] , \wPDiag_43[39] , 
        \wPDiag_43[38] , \wPDiag_43[37] , \wPDiag_43[36] , \wPDiag_43[35] , 
        \wPDiag_43[34] , \wPDiag_43[33] , \wPDiag_43[32] , \wPDiag_43[31] , 
        \wPDiag_43[30] , \wPDiag_43[29] , \wPDiag_43[28] , \wPDiag_43[27] , 
        \wPDiag_43[26] , \wPDiag_43[25] , \wPDiag_43[24] , \wPDiag_43[23] , 
        \wPDiag_43[22] , \wPDiag_43[21] , \wPDiag_43[20] , \wPDiag_43[19] , 
        \wPDiag_43[18] , \wPDiag_43[17] , \wPDiag_43[16] , \wPDiag_43[15] , 
        \wPDiag_43[14] , \wPDiag_43[13] , \wPDiag_43[12] , \wPDiag_43[11] , 
        \wPDiag_43[10] , \wPDiag_43[9] , \wPDiag_43[8] , \wPDiag_43[7] , 
        \wPDiag_43[6] , \wPDiag_43[5] , \wPDiag_43[4] , \wPDiag_43[3] , 
        \wPDiag_43[2] , \wPDiag_43[1] , \wPDiag_43[0] }), .NDiagOut({
        \wNDiag_43[63] , \wNDiag_43[62] , \wNDiag_43[61] , \wNDiag_43[60] , 
        \wNDiag_43[59] , \wNDiag_43[58] , \wNDiag_43[57] , \wNDiag_43[56] , 
        \wNDiag_43[55] , \wNDiag_43[54] , \wNDiag_43[53] , \wNDiag_43[52] , 
        \wNDiag_43[51] , \wNDiag_43[50] , \wNDiag_43[49] , \wNDiag_43[48] , 
        \wNDiag_43[47] , \wNDiag_43[46] , \wNDiag_43[45] , \wNDiag_43[44] , 
        \wNDiag_43[43] , \wNDiag_43[42] , \wNDiag_43[41] , \wNDiag_43[40] , 
        \wNDiag_43[39] , \wNDiag_43[38] , \wNDiag_43[37] , \wNDiag_43[36] , 
        \wNDiag_43[35] , \wNDiag_43[34] , \wNDiag_43[33] , \wNDiag_43[32] , 
        \wNDiag_43[31] , \wNDiag_43[30] , \wNDiag_43[29] , \wNDiag_43[28] , 
        \wNDiag_43[27] , \wNDiag_43[26] , \wNDiag_43[25] , \wNDiag_43[24] , 
        \wNDiag_43[23] , \wNDiag_43[22] , \wNDiag_43[21] , \wNDiag_43[20] , 
        \wNDiag_43[19] , \wNDiag_43[18] , \wNDiag_43[17] , \wNDiag_43[16] , 
        \wNDiag_43[15] , \wNDiag_43[14] , \wNDiag_43[13] , \wNDiag_43[12] , 
        \wNDiag_43[11] , \wNDiag_43[10] , \wNDiag_43[9] , \wNDiag_43[8] , 
        \wNDiag_43[7] , \wNDiag_43[6] , \wNDiag_43[5] , \wNDiag_43[4] , 
        \wNDiag_43[3] , \wNDiag_43[2] , \wNDiag_43[1] , \wNDiag_43[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_25 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_26[6] , \wScan_26[5] , \wScan_26[4] , 
        \wScan_26[3] , \wScan_26[2] , \wScan_26[1] , \wScan_26[0] }), 
        .ScanOut({\wScan_25[6] , \wScan_25[5] , \wScan_25[4] , \wScan_25[3] , 
        \wScan_25[2] , \wScan_25[1] , \wScan_25[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_25[0] ), .ReturnIn(\wReturn_26[0] ), .ColIn({
        \wColumn_25[63] , \wColumn_25[62] , \wColumn_25[61] , \wColumn_25[60] , 
        \wColumn_25[59] , \wColumn_25[58] , \wColumn_25[57] , \wColumn_25[56] , 
        \wColumn_25[55] , \wColumn_25[54] , \wColumn_25[53] , \wColumn_25[52] , 
        \wColumn_25[51] , \wColumn_25[50] , \wColumn_25[49] , \wColumn_25[48] , 
        \wColumn_25[47] , \wColumn_25[46] , \wColumn_25[45] , \wColumn_25[44] , 
        \wColumn_25[43] , \wColumn_25[42] , \wColumn_25[41] , \wColumn_25[40] , 
        \wColumn_25[39] , \wColumn_25[38] , \wColumn_25[37] , \wColumn_25[36] , 
        \wColumn_25[35] , \wColumn_25[34] , \wColumn_25[33] , \wColumn_25[32] , 
        \wColumn_25[31] , \wColumn_25[30] , \wColumn_25[29] , \wColumn_25[28] , 
        \wColumn_25[27] , \wColumn_25[26] , \wColumn_25[25] , \wColumn_25[24] , 
        \wColumn_25[23] , \wColumn_25[22] , \wColumn_25[21] , \wColumn_25[20] , 
        \wColumn_25[19] , \wColumn_25[18] , \wColumn_25[17] , \wColumn_25[16] , 
        \wColumn_25[15] , \wColumn_25[14] , \wColumn_25[13] , \wColumn_25[12] , 
        \wColumn_25[11] , \wColumn_25[10] , \wColumn_25[9] , \wColumn_25[8] , 
        \wColumn_25[7] , \wColumn_25[6] , \wColumn_25[5] , \wColumn_25[4] , 
        \wColumn_25[3] , \wColumn_25[2] , \wColumn_25[1] , \wColumn_25[0] }), 
        .PDiagIn({\wPDiag_25[63] , \wPDiag_25[62] , \wPDiag_25[61] , 
        \wPDiag_25[60] , \wPDiag_25[59] , \wPDiag_25[58] , \wPDiag_25[57] , 
        \wPDiag_25[56] , \wPDiag_25[55] , \wPDiag_25[54] , \wPDiag_25[53] , 
        \wPDiag_25[52] , \wPDiag_25[51] , \wPDiag_25[50] , \wPDiag_25[49] , 
        \wPDiag_25[48] , \wPDiag_25[47] , \wPDiag_25[46] , \wPDiag_25[45] , 
        \wPDiag_25[44] , \wPDiag_25[43] , \wPDiag_25[42] , \wPDiag_25[41] , 
        \wPDiag_25[40] , \wPDiag_25[39] , \wPDiag_25[38] , \wPDiag_25[37] , 
        \wPDiag_25[36] , \wPDiag_25[35] , \wPDiag_25[34] , \wPDiag_25[33] , 
        \wPDiag_25[32] , \wPDiag_25[31] , \wPDiag_25[30] , \wPDiag_25[29] , 
        \wPDiag_25[28] , \wPDiag_25[27] , \wPDiag_25[26] , \wPDiag_25[25] , 
        \wPDiag_25[24] , \wPDiag_25[23] , \wPDiag_25[22] , \wPDiag_25[21] , 
        \wPDiag_25[20] , \wPDiag_25[19] , \wPDiag_25[18] , \wPDiag_25[17] , 
        \wPDiag_25[16] , \wPDiag_25[15] , \wPDiag_25[14] , \wPDiag_25[13] , 
        \wPDiag_25[12] , \wPDiag_25[11] , \wPDiag_25[10] , \wPDiag_25[9] , 
        \wPDiag_25[8] , \wPDiag_25[7] , \wPDiag_25[6] , \wPDiag_25[5] , 
        \wPDiag_25[4] , \wPDiag_25[3] , \wPDiag_25[2] , \wPDiag_25[1] , 
        \wPDiag_25[0] }), .NDiagIn({\wNDiag_25[63] , \wNDiag_25[62] , 
        \wNDiag_25[61] , \wNDiag_25[60] , \wNDiag_25[59] , \wNDiag_25[58] , 
        \wNDiag_25[57] , \wNDiag_25[56] , \wNDiag_25[55] , \wNDiag_25[54] , 
        \wNDiag_25[53] , \wNDiag_25[52] , \wNDiag_25[51] , \wNDiag_25[50] , 
        \wNDiag_25[49] , \wNDiag_25[48] , \wNDiag_25[47] , \wNDiag_25[46] , 
        \wNDiag_25[45] , \wNDiag_25[44] , \wNDiag_25[43] , \wNDiag_25[42] , 
        \wNDiag_25[41] , \wNDiag_25[40] , \wNDiag_25[39] , \wNDiag_25[38] , 
        \wNDiag_25[37] , \wNDiag_25[36] , \wNDiag_25[35] , \wNDiag_25[34] , 
        \wNDiag_25[33] , \wNDiag_25[32] , \wNDiag_25[31] , \wNDiag_25[30] , 
        \wNDiag_25[29] , \wNDiag_25[28] , \wNDiag_25[27] , \wNDiag_25[26] , 
        \wNDiag_25[25] , \wNDiag_25[24] , \wNDiag_25[23] , \wNDiag_25[22] , 
        \wNDiag_25[21] , \wNDiag_25[20] , \wNDiag_25[19] , \wNDiag_25[18] , 
        \wNDiag_25[17] , \wNDiag_25[16] , \wNDiag_25[15] , \wNDiag_25[14] , 
        \wNDiag_25[13] , \wNDiag_25[12] , \wNDiag_25[11] , \wNDiag_25[10] , 
        \wNDiag_25[9] , \wNDiag_25[8] , \wNDiag_25[7] , \wNDiag_25[6] , 
        \wNDiag_25[5] , \wNDiag_25[4] , \wNDiag_25[3] , \wNDiag_25[2] , 
        \wNDiag_25[1] , \wNDiag_25[0] }), .CallOut(\wCall_26[0] ), .ReturnOut(
        \wReturn_25[0] ), .ColOut({\wColumn_26[63] , \wColumn_26[62] , 
        \wColumn_26[61] , \wColumn_26[60] , \wColumn_26[59] , \wColumn_26[58] , 
        \wColumn_26[57] , \wColumn_26[56] , \wColumn_26[55] , \wColumn_26[54] , 
        \wColumn_26[53] , \wColumn_26[52] , \wColumn_26[51] , \wColumn_26[50] , 
        \wColumn_26[49] , \wColumn_26[48] , \wColumn_26[47] , \wColumn_26[46] , 
        \wColumn_26[45] , \wColumn_26[44] , \wColumn_26[43] , \wColumn_26[42] , 
        \wColumn_26[41] , \wColumn_26[40] , \wColumn_26[39] , \wColumn_26[38] , 
        \wColumn_26[37] , \wColumn_26[36] , \wColumn_26[35] , \wColumn_26[34] , 
        \wColumn_26[33] , \wColumn_26[32] , \wColumn_26[31] , \wColumn_26[30] , 
        \wColumn_26[29] , \wColumn_26[28] , \wColumn_26[27] , \wColumn_26[26] , 
        \wColumn_26[25] , \wColumn_26[24] , \wColumn_26[23] , \wColumn_26[22] , 
        \wColumn_26[21] , \wColumn_26[20] , \wColumn_26[19] , \wColumn_26[18] , 
        \wColumn_26[17] , \wColumn_26[16] , \wColumn_26[15] , \wColumn_26[14] , 
        \wColumn_26[13] , \wColumn_26[12] , \wColumn_26[11] , \wColumn_26[10] , 
        \wColumn_26[9] , \wColumn_26[8] , \wColumn_26[7] , \wColumn_26[6] , 
        \wColumn_26[5] , \wColumn_26[4] , \wColumn_26[3] , \wColumn_26[2] , 
        \wColumn_26[1] , \wColumn_26[0] }), .PDiagOut({\wPDiag_26[63] , 
        \wPDiag_26[62] , \wPDiag_26[61] , \wPDiag_26[60] , \wPDiag_26[59] , 
        \wPDiag_26[58] , \wPDiag_26[57] , \wPDiag_26[56] , \wPDiag_26[55] , 
        \wPDiag_26[54] , \wPDiag_26[53] , \wPDiag_26[52] , \wPDiag_26[51] , 
        \wPDiag_26[50] , \wPDiag_26[49] , \wPDiag_26[48] , \wPDiag_26[47] , 
        \wPDiag_26[46] , \wPDiag_26[45] , \wPDiag_26[44] , \wPDiag_26[43] , 
        \wPDiag_26[42] , \wPDiag_26[41] , \wPDiag_26[40] , \wPDiag_26[39] , 
        \wPDiag_26[38] , \wPDiag_26[37] , \wPDiag_26[36] , \wPDiag_26[35] , 
        \wPDiag_26[34] , \wPDiag_26[33] , \wPDiag_26[32] , \wPDiag_26[31] , 
        \wPDiag_26[30] , \wPDiag_26[29] , \wPDiag_26[28] , \wPDiag_26[27] , 
        \wPDiag_26[26] , \wPDiag_26[25] , \wPDiag_26[24] , \wPDiag_26[23] , 
        \wPDiag_26[22] , \wPDiag_26[21] , \wPDiag_26[20] , \wPDiag_26[19] , 
        \wPDiag_26[18] , \wPDiag_26[17] , \wPDiag_26[16] , \wPDiag_26[15] , 
        \wPDiag_26[14] , \wPDiag_26[13] , \wPDiag_26[12] , \wPDiag_26[11] , 
        \wPDiag_26[10] , \wPDiag_26[9] , \wPDiag_26[8] , \wPDiag_26[7] , 
        \wPDiag_26[6] , \wPDiag_26[5] , \wPDiag_26[4] , \wPDiag_26[3] , 
        \wPDiag_26[2] , \wPDiag_26[1] , \wPDiag_26[0] }), .NDiagOut({
        \wNDiag_26[63] , \wNDiag_26[62] , \wNDiag_26[61] , \wNDiag_26[60] , 
        \wNDiag_26[59] , \wNDiag_26[58] , \wNDiag_26[57] , \wNDiag_26[56] , 
        \wNDiag_26[55] , \wNDiag_26[54] , \wNDiag_26[53] , \wNDiag_26[52] , 
        \wNDiag_26[51] , \wNDiag_26[50] , \wNDiag_26[49] , \wNDiag_26[48] , 
        \wNDiag_26[47] , \wNDiag_26[46] , \wNDiag_26[45] , \wNDiag_26[44] , 
        \wNDiag_26[43] , \wNDiag_26[42] , \wNDiag_26[41] , \wNDiag_26[40] , 
        \wNDiag_26[39] , \wNDiag_26[38] , \wNDiag_26[37] , \wNDiag_26[36] , 
        \wNDiag_26[35] , \wNDiag_26[34] , \wNDiag_26[33] , \wNDiag_26[32] , 
        \wNDiag_26[31] , \wNDiag_26[30] , \wNDiag_26[29] , \wNDiag_26[28] , 
        \wNDiag_26[27] , \wNDiag_26[26] , \wNDiag_26[25] , \wNDiag_26[24] , 
        \wNDiag_26[23] , \wNDiag_26[22] , \wNDiag_26[21] , \wNDiag_26[20] , 
        \wNDiag_26[19] , \wNDiag_26[18] , \wNDiag_26[17] , \wNDiag_26[16] , 
        \wNDiag_26[15] , \wNDiag_26[14] , \wNDiag_26[13] , \wNDiag_26[12] , 
        \wNDiag_26[11] , \wNDiag_26[10] , \wNDiag_26[9] , \wNDiag_26[8] , 
        \wNDiag_26[7] , \wNDiag_26[6] , \wNDiag_26[5] , \wNDiag_26[4] , 
        \wNDiag_26[3] , \wNDiag_26[2] , \wNDiag_26[1] , \wNDiag_26[0] }) );
    NQueens_Node_WIDTH64_IDWIDTH7_SCAN1 U_NQueens_Node_50 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_51[6] , \wScan_51[5] , \wScan_51[4] , 
        \wScan_51[3] , \wScan_51[2] , \wScan_51[1] , \wScan_51[0] }), 
        .ScanOut({\wScan_50[6] , \wScan_50[5] , \wScan_50[4] , \wScan_50[3] , 
        \wScan_50[2] , \wScan_50[1] , \wScan_50[0] }), .ScanEnable(
        \wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CallIn(\wCall_50[0] ), .ReturnIn(\wReturn_51[0] ), .ColIn({
        \wColumn_50[63] , \wColumn_50[62] , \wColumn_50[61] , \wColumn_50[60] , 
        \wColumn_50[59] , \wColumn_50[58] , \wColumn_50[57] , \wColumn_50[56] , 
        \wColumn_50[55] , \wColumn_50[54] , \wColumn_50[53] , \wColumn_50[52] , 
        \wColumn_50[51] , \wColumn_50[50] , \wColumn_50[49] , \wColumn_50[48] , 
        \wColumn_50[47] , \wColumn_50[46] , \wColumn_50[45] , \wColumn_50[44] , 
        \wColumn_50[43] , \wColumn_50[42] , \wColumn_50[41] , \wColumn_50[40] , 
        \wColumn_50[39] , \wColumn_50[38] , \wColumn_50[37] , \wColumn_50[36] , 
        \wColumn_50[35] , \wColumn_50[34] , \wColumn_50[33] , \wColumn_50[32] , 
        \wColumn_50[31] , \wColumn_50[30] , \wColumn_50[29] , \wColumn_50[28] , 
        \wColumn_50[27] , \wColumn_50[26] , \wColumn_50[25] , \wColumn_50[24] , 
        \wColumn_50[23] , \wColumn_50[22] , \wColumn_50[21] , \wColumn_50[20] , 
        \wColumn_50[19] , \wColumn_50[18] , \wColumn_50[17] , \wColumn_50[16] , 
        \wColumn_50[15] , \wColumn_50[14] , \wColumn_50[13] , \wColumn_50[12] , 
        \wColumn_50[11] , \wColumn_50[10] , \wColumn_50[9] , \wColumn_50[8] , 
        \wColumn_50[7] , \wColumn_50[6] , \wColumn_50[5] , \wColumn_50[4] , 
        \wColumn_50[3] , \wColumn_50[2] , \wColumn_50[1] , \wColumn_50[0] }), 
        .PDiagIn({\wPDiag_50[63] , \wPDiag_50[62] , \wPDiag_50[61] , 
        \wPDiag_50[60] , \wPDiag_50[59] , \wPDiag_50[58] , \wPDiag_50[57] , 
        \wPDiag_50[56] , \wPDiag_50[55] , \wPDiag_50[54] , \wPDiag_50[53] , 
        \wPDiag_50[52] , \wPDiag_50[51] , \wPDiag_50[50] , \wPDiag_50[49] , 
        \wPDiag_50[48] , \wPDiag_50[47] , \wPDiag_50[46] , \wPDiag_50[45] , 
        \wPDiag_50[44] , \wPDiag_50[43] , \wPDiag_50[42] , \wPDiag_50[41] , 
        \wPDiag_50[40] , \wPDiag_50[39] , \wPDiag_50[38] , \wPDiag_50[37] , 
        \wPDiag_50[36] , \wPDiag_50[35] , \wPDiag_50[34] , \wPDiag_50[33] , 
        \wPDiag_50[32] , \wPDiag_50[31] , \wPDiag_50[30] , \wPDiag_50[29] , 
        \wPDiag_50[28] , \wPDiag_50[27] , \wPDiag_50[26] , \wPDiag_50[25] , 
        \wPDiag_50[24] , \wPDiag_50[23] , \wPDiag_50[22] , \wPDiag_50[21] , 
        \wPDiag_50[20] , \wPDiag_50[19] , \wPDiag_50[18] , \wPDiag_50[17] , 
        \wPDiag_50[16] , \wPDiag_50[15] , \wPDiag_50[14] , \wPDiag_50[13] , 
        \wPDiag_50[12] , \wPDiag_50[11] , \wPDiag_50[10] , \wPDiag_50[9] , 
        \wPDiag_50[8] , \wPDiag_50[7] , \wPDiag_50[6] , \wPDiag_50[5] , 
        \wPDiag_50[4] , \wPDiag_50[3] , \wPDiag_50[2] , \wPDiag_50[1] , 
        \wPDiag_50[0] }), .NDiagIn({\wNDiag_50[63] , \wNDiag_50[62] , 
        \wNDiag_50[61] , \wNDiag_50[60] , \wNDiag_50[59] , \wNDiag_50[58] , 
        \wNDiag_50[57] , \wNDiag_50[56] , \wNDiag_50[55] , \wNDiag_50[54] , 
        \wNDiag_50[53] , \wNDiag_50[52] , \wNDiag_50[51] , \wNDiag_50[50] , 
        \wNDiag_50[49] , \wNDiag_50[48] , \wNDiag_50[47] , \wNDiag_50[46] , 
        \wNDiag_50[45] , \wNDiag_50[44] , \wNDiag_50[43] , \wNDiag_50[42] , 
        \wNDiag_50[41] , \wNDiag_50[40] , \wNDiag_50[39] , \wNDiag_50[38] , 
        \wNDiag_50[37] , \wNDiag_50[36] , \wNDiag_50[35] , \wNDiag_50[34] , 
        \wNDiag_50[33] , \wNDiag_50[32] , \wNDiag_50[31] , \wNDiag_50[30] , 
        \wNDiag_50[29] , \wNDiag_50[28] , \wNDiag_50[27] , \wNDiag_50[26] , 
        \wNDiag_50[25] , \wNDiag_50[24] , \wNDiag_50[23] , \wNDiag_50[22] , 
        \wNDiag_50[21] , \wNDiag_50[20] , \wNDiag_50[19] , \wNDiag_50[18] , 
        \wNDiag_50[17] , \wNDiag_50[16] , \wNDiag_50[15] , \wNDiag_50[14] , 
        \wNDiag_50[13] , \wNDiag_50[12] , \wNDiag_50[11] , \wNDiag_50[10] , 
        \wNDiag_50[9] , \wNDiag_50[8] , \wNDiag_50[7] , \wNDiag_50[6] , 
        \wNDiag_50[5] , \wNDiag_50[4] , \wNDiag_50[3] , \wNDiag_50[2] , 
        \wNDiag_50[1] , \wNDiag_50[0] }), .CallOut(\wCall_51[0] ), .ReturnOut(
        \wReturn_50[0] ), .ColOut({\wColumn_51[63] , \wColumn_51[62] , 
        \wColumn_51[61] , \wColumn_51[60] , \wColumn_51[59] , \wColumn_51[58] , 
        \wColumn_51[57] , \wColumn_51[56] , \wColumn_51[55] , \wColumn_51[54] , 
        \wColumn_51[53] , \wColumn_51[52] , \wColumn_51[51] , \wColumn_51[50] , 
        \wColumn_51[49] , \wColumn_51[48] , \wColumn_51[47] , \wColumn_51[46] , 
        \wColumn_51[45] , \wColumn_51[44] , \wColumn_51[43] , \wColumn_51[42] , 
        \wColumn_51[41] , \wColumn_51[40] , \wColumn_51[39] , \wColumn_51[38] , 
        \wColumn_51[37] , \wColumn_51[36] , \wColumn_51[35] , \wColumn_51[34] , 
        \wColumn_51[33] , \wColumn_51[32] , \wColumn_51[31] , \wColumn_51[30] , 
        \wColumn_51[29] , \wColumn_51[28] , \wColumn_51[27] , \wColumn_51[26] , 
        \wColumn_51[25] , \wColumn_51[24] , \wColumn_51[23] , \wColumn_51[22] , 
        \wColumn_51[21] , \wColumn_51[20] , \wColumn_51[19] , \wColumn_51[18] , 
        \wColumn_51[17] , \wColumn_51[16] , \wColumn_51[15] , \wColumn_51[14] , 
        \wColumn_51[13] , \wColumn_51[12] , \wColumn_51[11] , \wColumn_51[10] , 
        \wColumn_51[9] , \wColumn_51[8] , \wColumn_51[7] , \wColumn_51[6] , 
        \wColumn_51[5] , \wColumn_51[4] , \wColumn_51[3] , \wColumn_51[2] , 
        \wColumn_51[1] , \wColumn_51[0] }), .PDiagOut({\wPDiag_51[63] , 
        \wPDiag_51[62] , \wPDiag_51[61] , \wPDiag_51[60] , \wPDiag_51[59] , 
        \wPDiag_51[58] , \wPDiag_51[57] , \wPDiag_51[56] , \wPDiag_51[55] , 
        \wPDiag_51[54] , \wPDiag_51[53] , \wPDiag_51[52] , \wPDiag_51[51] , 
        \wPDiag_51[50] , \wPDiag_51[49] , \wPDiag_51[48] , \wPDiag_51[47] , 
        \wPDiag_51[46] , \wPDiag_51[45] , \wPDiag_51[44] , \wPDiag_51[43] , 
        \wPDiag_51[42] , \wPDiag_51[41] , \wPDiag_51[40] , \wPDiag_51[39] , 
        \wPDiag_51[38] , \wPDiag_51[37] , \wPDiag_51[36] , \wPDiag_51[35] , 
        \wPDiag_51[34] , \wPDiag_51[33] , \wPDiag_51[32] , \wPDiag_51[31] , 
        \wPDiag_51[30] , \wPDiag_51[29] , \wPDiag_51[28] , \wPDiag_51[27] , 
        \wPDiag_51[26] , \wPDiag_51[25] , \wPDiag_51[24] , \wPDiag_51[23] , 
        \wPDiag_51[22] , \wPDiag_51[21] , \wPDiag_51[20] , \wPDiag_51[19] , 
        \wPDiag_51[18] , \wPDiag_51[17] , \wPDiag_51[16] , \wPDiag_51[15] , 
        \wPDiag_51[14] , \wPDiag_51[13] , \wPDiag_51[12] , \wPDiag_51[11] , 
        \wPDiag_51[10] , \wPDiag_51[9] , \wPDiag_51[8] , \wPDiag_51[7] , 
        \wPDiag_51[6] , \wPDiag_51[5] , \wPDiag_51[4] , \wPDiag_51[3] , 
        \wPDiag_51[2] , \wPDiag_51[1] , \wPDiag_51[0] }), .NDiagOut({
        \wNDiag_51[63] , \wNDiag_51[62] , \wNDiag_51[61] , \wNDiag_51[60] , 
        \wNDiag_51[59] , \wNDiag_51[58] , \wNDiag_51[57] , \wNDiag_51[56] , 
        \wNDiag_51[55] , \wNDiag_51[54] , \wNDiag_51[53] , \wNDiag_51[52] , 
        \wNDiag_51[51] , \wNDiag_51[50] , \wNDiag_51[49] , \wNDiag_51[48] , 
        \wNDiag_51[47] , \wNDiag_51[46] , \wNDiag_51[45] , \wNDiag_51[44] , 
        \wNDiag_51[43] , \wNDiag_51[42] , \wNDiag_51[41] , \wNDiag_51[40] , 
        \wNDiag_51[39] , \wNDiag_51[38] , \wNDiag_51[37] , \wNDiag_51[36] , 
        \wNDiag_51[35] , \wNDiag_51[34] , \wNDiag_51[33] , \wNDiag_51[32] , 
        \wNDiag_51[31] , \wNDiag_51[30] , \wNDiag_51[29] , \wNDiag_51[28] , 
        \wNDiag_51[27] , \wNDiag_51[26] , \wNDiag_51[25] , \wNDiag_51[24] , 
        \wNDiag_51[23] , \wNDiag_51[22] , \wNDiag_51[21] , \wNDiag_51[20] , 
        \wNDiag_51[19] , \wNDiag_51[18] , \wNDiag_51[17] , \wNDiag_51[16] , 
        \wNDiag_51[15] , \wNDiag_51[14] , \wNDiag_51[13] , \wNDiag_51[12] , 
        \wNDiag_51[11] , \wNDiag_51[10] , \wNDiag_51[9] , \wNDiag_51[8] , 
        \wNDiag_51[7] , \wNDiag_51[6] , \wNDiag_51[5] , \wNDiag_51[4] , 
        \wNDiag_51[3] , \wNDiag_51[2] , \wNDiag_51[1] , \wNDiag_51[0] }) );
    NQueens_Control_IDWIDTH7_SCAN1 U_NQueens_Control ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\wScan_0[6] , \wScan_0[5] , \wScan_0[4] , \wScan_0[3] , 
        \wScan_0[2] , \wScan_0[1] , \wScan_0[0] }), .ScanOut({\wScan_64[6] , 
        \wScan_64[5] , \wScan_64[4] , \wScan_64[3] , \wScan_64[2] , 
        \wScan_64[1] , \wScan_64[0] }), .ScanEnable(\wScanEnable[0] ), .Id({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .ScanId({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(\wCall_64[0] ), .ReturnIn(
        \wReturn_0[0] ), .CallOut(\wCall_0[0] ) );
endmodule

