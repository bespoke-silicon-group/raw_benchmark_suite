
module IntMatMul_Control_pVectorSize16_pWordSize8_pScan1_DW01_cmp2_15_0 ( A, B, 
    LEQ, TC, LT_LE, GE_GT );
input  [14:0] A;
input  [14:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17;
    VMW_NOR4 U3 ( .A(n15), .B(n16), .C(A[5]), .D(A[4]), .Z(LT_LE) );
    VMW_OR4 U5 ( .A(A[11]), .B(A[10]), .C(A[9]), .D(n17), .Z(n15) );
    VMW_OR3 U6 ( .A(A[8]), .B(A[7]), .C(A[6]), .Z(n16) );
    VMW_OR3 U4 ( .A(A[14]), .B(A[13]), .C(A[12]), .Z(n17) );
endmodule


module IntMatMul_Control_pVectorSize16_pWordSize8_pScan1 ( Clk, Reset, RD, WR, 
    Addr, DataIn, DataOut, vectorInput, matrixInput, cOutput );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [127:0] vectorInput;
input  [127:0] cOutput;
output [2047:0] matrixInput;
input  Clk, Reset, RD, WR;
    wire n26979, n25091, n27349, n25949, n27079, n27145, n27275, n25680, 
        n25710, n25101, n26131, n26720, n25231, n25420, n25852, n26862, n26391, 
        n26410, n26580, n26201, n25597, n27252, n25216, n25386, n25407, n26845, 
        n25875, n26437, n26226, n27162, n25737, n25126, n26707, n26086, n26116, 
        n26697, n25278, n25469, n26248, n26459, n25759, n25148, n26769, n26178, 
        n25074, n27327, n26930, n26353, n26542, n25363, n25572, n25890, n26672, 
        n25900, n26063, n27187, n27017, n25642, n26655, n26044, n27030, n25665, 
        n26374, n26887, n26917, n26565, n25344, n25555, n25927, n27290, n27300, 
        n25191, n27390, n25659, n26559, n26669, n25378, n26078, n25569, n26348, 
        n26817, n26987, n26465, n26274, n25244, n25455, n27200, n26755, n25827, 
        n26144, n27130, n25174, n25765, n26772, n26163, n27117, n27087, n25742, 
        n25153, n26830, n26442, n26253, n25263, n25472, n27227, n25800, n25990, 
        n27249, n27179, n26879, n25849, n27062, n25637, n26607, n26797, n26016, 
        n26186, n25286, n25507, n25316, n25497, n25975, n27375, n27352, n26945, 
        n26326, n26537, n25331, n25520, n25952, n26962, n26291, n26510, n26301, 
        n26480, \holder[0] , n27045, n25780, n26620, n25610, n26031, n25625, 
        n27340, n26615, n27070, n26194, n26785, n26004, n25967, n25304, n25485, 
        n25294, n25515, n26525, n26334, n26957, n27382, n27367, n25940, n25323, 
        n25532, n26283, n26313, n26492, n26502, n26970, n25602, n25183, n25792, 
        n27057, n26632, n26023, n26398, n26419, n26589, n26208, n25238, n25429, 
        n26729, n26138, n25689, n25108, n25719, n25098, n26266, n26477, n26995, 
        n26805, n25835, n27212, n25447, n25256, n26156, n26747, n25777, n27299, 
        n25166, n27122, n26760, n26171, n25141, n25750, n27095, n27105, n26450, 
        n26241, n26822, n27235, n25812, n25982, n25271, n25460, n27309, n27039, 
        n25899, n25909, Logic11, n26341, n26939, n26550, n25066, n27335, 
        n26922, n25912, n25882, n25371, n25560, n26660, n26071, n27195, n27005, 
        n25650, \holder[4] , n26647, n26056, n27312, n27282, n25677, n27022, 
        n26366, n26577, n26895, n26905, n25935, n25356, n25547, n25809, n25999, 
        n26839, n25198, n25204, n25083, n27209, n27139, n25692, n25113, n27267, 
        n25702, n27157, n26732, n26123, n25840, n26383, n26402, n25223, n25432, 
        n26592, n26213, n26870, n25394, n25415, n27240, n25867, n25585, n26425, 
        n26234, n26857, n25725, n25134, n27170, n26104, n26629, n26685, n26715, 
        n26094, n26038, n25203, n25619, n25789, n26489, n26298, n26308, n26519, 
        n25338, n25529, n26682, n26712, n26093, n26103, n27177, n26850, n25722, 
        n25133, n26422, n26233, n25061, n25084, n27260, n25393, n25582, n25412, 
        n25860, n27247, n26877, n26214, n26384, n26595, n26405, n25224, n25435, 
        n25847, n26735, n26124, n25705, n27150, n27285, n27315, n25695, n25114, 
        n25639, n26328, n26609, n26799, n26018, n25288, n26188, n25318, n25509, 
        n25499, n26539, n25351, n25540, n25932, n26892, n26902, n26361, n26570, 
        n27025, \holder[6] , n25670, n26640, n26051, n27192, n27002, n25657, 
        n27332, n26667, n26076, n25376, n25567, n25885, n25915, n26925, n26557, 
        n26346, n26819, n26989, n25829, n27385, n27229, n27089, n27119, n25467, 
        n27232, n25276, n25815, n25985, n26825, n26246, n26457, n27092, n27102, 
        n25757, n25146, n26176, n26767, n27125, n25161, n26740, n25770, n26151, 
        n25251, n25440, n25832, n27329, n27215, n26802, n26992, n26261, n26470, 
        n27189, n27019, n26889, n26919, n25929, n26635, n26024, n27050, n25795, 
        n26284, n26977, n25605, n25184, n26505, n26314, n26495, n25324, n25535, 
        n27347, n27360, n25947, n26950, n26333, n26522, n25293, n25303, n25512, 
        n25482, n26612, n26782, n25960, n26003, n26193, n27077, n25622, n26439, 
        n25218, n25388, n25599, n25409, n25739, n26228, n25128, n26699, n26709, 
        n26088, n26118, n27269, n27159, n25869, n26859, n25196, n26036, n26627, 
        n25617, n25068, n25787, n27372, n27042, n26306, n26296, n26487, n26517, 
        n26965, n27355, n25955, n25527, n26321, n26530, n25336, n26942, n25972, 
        n25281, n25311, n25490, n25500, n26600, n26790, n26181, n26011, n27065, 
        n25630, \holder[2] , n26649, n26058, n25073, n25679, n26368, n26579, 
        n25358, n25549, n25997, n25807, n27220, n25264, n25475, n26445, n26254, 
        n26837, n27080, n25745, n25154, n27110, n27297, n26775, n25762, n26164, 
        n25173, n27137, n26752, n26143, n27207, n25820, n26273, n25243, n25452, 
        n26462, n26810, n26980, n26268, n26479, n25258, n25449, n26749, n26158, 
        n25779, n25168, n25920, n27307, n25343, n25552, n26373, n26562, n26910, 
        n26880, n25662, n27037, n26652, n25645, n26043, n27320, n27180, n27010, 
        n26064, n26675, n25907, n25897, n25575, n25364, n26354, n26545, n26937, 
        n25969, n26959, n27369, n27059, n27272, n26690, n26700, n26111, n26081, 
        n25730, n25121, n27165, n26430, n26221, n26842, n27255, n25872, n26396, 
        n25211, n25381, n25400, n25590, n26417, n26587, n26206, n26865, n25855, 
        n25236, n25427, n25185, n26727, n26136, n25687, n25106, n25096, n25717, 
        n27051, n27142, n27346, n27361, n25604, n25794, n26025, n26634, n25534, 
        n25325, n25946, n26976, n26315, n26494, n26504, n26285, n25292, n25302, 
        n25483, n25513, n25961, n26951, n26332, n26523, n27076, n26613, n25623, 
        n26192, n26002, n26783, n26438, n26229, n26698, n25219, n25389, n25408, 
        n25598, n26119, n26708, n26089, n25738, n25129, n27328, n27384, n26824, 
        n26456, n26247, n25277, n25466, n27233, n25814, n25984, n26766, n26177, 
        n27093, n27103, n25147, n25756, n26741, n26150, n27124, n26993, n25771, 
        n25160, n26803, n26260, n26471, n25250, n25441, n25833, n27214, n27188, 
        n27018, n25928, n26888, n26918, n26893, n26903, n26360, n26571, n25060, 
        n27314, n27284, n25350, n25541, n26641, n25933, n26050, n27024, n27333, 
        n25671, n26666, n26077, n27193, n27003, n25656, n26924, n26347, n26556, 
        n25377, n25566, n25884, n25914, n25828, n26818, n26988, n27088, n27118, 
        n27228, n25202, n27176, n25723, n26102, n25132, n26683, n26713, n26092, 
        n25392, n25413, n25583, n25085, n27261, n25861, n27246, n26851, n26423, 
        n26232, n25225, n25434, n25846, n26876, n26385, n26404, n26594, n26215, 
        n25694, n27151, n25115, n25704, n26734, n26125, n26608, n26189, n26798, 
        n26019, n25638, n26329, n26538, n27368, n25289, n25319, n25498, n25508, 
        n26958, n25968, n27058, n27273, n25731, n25120, n27164, n26691, n26701, 
        n26080, n26110, n27254, n26431, n25210, n25591, n25873, n25380, n25401, 
        n26220, n26843, n25854, n25237, n25426, n26416, n26586, n26207, n26397, 
        n26864, n25097, n25686, n25716, n25107, n27143, n26726, n26137, n26269, 
        n26478, n25259, n25448, n25778, n25169, n26748, n26159, n25055, n25072, 
        n27296, n27306, n26372, n26563, n26881, n26911, n25921, n25342, n25553, 
        n26042, n26653, n25663, n27036, n26674, n26065, n25644, n27181, n27011, 
        n27321, n26544, n26355, n26936, n25896, n25906, n25365, n25574, n25069, 
        n25678, n26648, n26059, n25359, n25548, n26369, n26578, n26255, n26444, 
        n26836, n25806, n25996, n27221, n25265, n25474, n26774, n26165, n25744, 
        n27111, n25155, n27081, n26753, n26142, n25763, n25172, n27136, n26272, 
        n26463, n26811, n26981, n27206, n25821, n25242, n25453, n27158, n25197, 
        n27268, n26858, n25868, n25786, n27354, n27373, n25616, n27043, n26626, 
        n26037, n25954, n25337, n25526, n26297, n26516, n26307, n26486, n26964, 
        n25973, n26320, n25280, n25501, n25310, n25491, n26531, n26943, n27064, 
        n25631, n27178, n26601, n26791, n26010, n26180, n27248, n25848, n26878, 
        n26606, n26796, n26187, n27063, n26017, n26944, n25636, n25190, n27353, 
        n26536, n26327, n25287, n25317, n25496, n25506, n25974, n27374, n26290, 
        n26300, n26963, n26481, n26511, n25330, n25521, n25953, n26621, n26030, 
        n27044, n25611, n27391, n25781, n26668, n26079, n25658, n26349, n26558, 
        n25379, n25568, n25454, n27201, n25245, n25075, n25826, n26986, n26816, 
        n26275, n26464, n27131, n25764, n25175, n26145, n26754, n27086, n27116, 
        n25743, n25152, n26773, n26162, n25262, n25473, n27226, n25801, n25991, 
        n26831, n26443, n26252, n26458, n26768, n25279, n26249, n25468, n26179, 
        n25758, n25149, n27326, n25362, n25573, n25901, n25891, n26931, n26352, 
        n26543, n27186, n27016, n25643, n26062, n26673, n27031, n25090, n27291, 
        n25664, n26654, n26045, n25345, n25554, n25926, n27301, n27348, n26916, 
        n26886, n26375, n26564, n25948, n26978, n26721, n27078, n26130, n27144, 
        n25681, n25711, n25100, n27274, n26863, n26390, n26411, n26581, n26200, 
        n25230, n25421, n25853, n25199, n25205, n25082, n26844, n26227, n26436, 
        n25387, n25406, n26696, n27253, n25217, n25596, n25874, n26117, n26706, 
        n26087, n27163, n25736, n25127, n26122, n26733, n25703, n27266, n25693, 
        n25112, n27156, n26382, n26593, n26212, n26403, n26871, n25841, n26424, 
        n25222, n25433, n26235, n26856, n27241, n25866, n25395, n25584, n25414, 
        n26684, n26714, n26095, n26105, n25135, n25724, n27171, n25618, n25788, 
        n25067, n26628, n25339, n26039, n25528, n27334, n26299, n26309, n26518, 
        n26488, n25883, n25913, n26340, n26551, n25370, n25561, n26923, n27194, 
        n25651, n27004, n26661, n25676, n26070, n27313, n27023, n26057, n26646, 
        n27283, n25934, n25546, n25357, n26367, n26576, n26894, n26904, n26838, 
        n25808, n25998, n27138, n27383, n27208, n25834, n27213, n25257, n25446, 
        n26476, n26267, n26804, n26994, n25167, n25776, n27123, n26746, n25751, 
        n26157, n25140, n27094, n27104, n26761, n26170, n27234, n25813, n26451, 
        n25270, n25461, n25983, n26240, n26823, n27298, n27308, n27038, n26938, 
        n25898, n25908, n26614, n26784, n26005, n26195, n25624, n27341, n27071, 
        n26335, n26524, n26956, n25966, n25295, n26282, n25305, n25514, n25484, 
        n26312, n26503, n26493, n26971, n25941, n25189, n27366, n25322, n25533, 
        n26633, n26022, n25793, n25603, n25182, n27056, n26399, n26588, n25239, 
        n25428, n26209, n26418, n25688, n25718, n25099, n25109, n25092, n27251, 
        n26728, n26139, n25876, n25385, n25404, n25215, n25594, n26225, n26434, 
        n26846, n25734, n25125, n27161, n26694, n26115, n26704, n26085, n25683, 
        n25102, n25713, n27276, n27146, n26723, n26132, n25851, n25232, n25423, 
        n26392, n26413, n26583, n26202, n26861, n26638, n26029, n25608, n27388, 
        n25077, n26289, n26319, n25798, n26498, n26508, n25329, n25538, n26656, 
        n26047, n27293, n26566, n27033, n25666, n26377, n26884, n26914, n25924, 
        n27303, n27324, n25347, n25556, n26350, n26541, n26933, n25903, n25360, 
        n25571, n25893, n26671, n26060, n25641, n27184, n27014, n27128, n27218, 
        n27393, n25818, n25988, n26828, n26771, n27084, n25741, n26160, n25150, 
        n27114, n26441, n26833, n26250, n27224, n25803, n25993, n25260, n25471, 
        n26277, n26466, n27203, n26814, n26984, n25824, n25456, n25247, n26147, 
        n26756, n25766, n25177, n27133, n27288, n26928, n25888, n25918, n27318, 
        n25192, n27376, n27028, n25951, n25332, n25523, n26292, n26302, n26483, 
        n26513, n26961, n25613, n25783, n27046, n26623, n26032, n25634, n27061, 
        n27351, n26604, n26794, n26185, n26015, n25976, n25285, n25315, n25494, 
        n25504, n26325, n26534, n26946, n26389, n26408, n26598, n26219, n26738, 
        n25229, n25438, n26129, n25089, n25698, n25708, n25119, n26868, n25858, 
        n27168, n25059, n27343, n27364, n27258, n25320, n25531, n25943, n26973, 
        n26280, n26310, n26501, n26491, n27054, n26631, n25601, n25791, n25180, 
        n26020, n27073, n25626, n26786, n26007, n26616, n26197, n25297, n25516, 
        n25307, n25486, n26954, n25964, n26337, n26526, n25648, n26678, n26069, 
        n26359, n26548, n25369, n25578, n26763, n26172, n27096, n27106, n25753, 
        n25142, n26821, n26453, n26242, n25272, n25463, n27236, n25811, n26806, 
        n25981, n26474, n26996, n26265, n25255, n25444, n27381, n25836, n27211, 
        n26744, n26155, n27121, n25165, n25774, n25207, n25065, n26259, n25269, 
        n25478, n26448, n25748, n25159, n26644, n26778, n26169, n26055, n27021, 
        n25674, n164, n27311, n26896, n26906, n26365, n26574, n25355, n25544, 
        n27336, n27281, n25936, n26921, n26342, n26553, n25372, n25563, n25881, 
        n25911, n26663, n26072, n27196, n27006, n27358, n25653, n27068, n26968, 
        n25958, n25080, n25397, n25586, n25416, n26426, n26854, n27243, n25864, 
        n26237, n27173, n25137, n25726, n26716, n26686, n26097, n26107, n25701, 
        n27154, n27378, n27264, n26731, n25691, n26120, n25110, n25220, n25431, 
        n25843, n26380, n26591, n26873, n26210, n26401, n27263, n27048, n25978, 
        n26948, n26387, n26406, n26596, n26874, n26217, n25844, n25227, n25436, 
        n25200, n25087, n26736, n26127, n25696, n25117, n25706, n27153, n27174, 
        n26681, n26100, n26711, n26090, n25721, n25130, n26421, n26230, n26853, 
        n25863, n25390, n25411, n27244, n25581, n25062, n26279, n26468, n26758, 
        n25249, n25458, n26149, n25768, n25179, n27001, n25654, n27191, n26075, 
        n26664, n25916, n27286, n27331, n25886, n25564, n25375, n26345, n26554, 
        n26926, n27316, n25931, n25352, n25543, n26362, n26573, n26891, n26901, 
        n27386, n25079, n25673, n27026, n26643, n26658, n26052, n26049, n26379, 
        n26568, n25668, n25349, n25558, n25773, n25162, n27126, n26152, n26743, 
        n25831, n27216, n25252, n25443, n26262, n26473, n26991, n26801, n27231, 
        n25986, n25816, n25275, n25464, n26454, n26245, n26826, n25754, n25145, 
        n27091, n27101, n26764, n26175, n25878, n26848, n27278, n27148, n27344, 
        n26330, n26521, n26953, n25290, n25300, n25481, n25963, n25511, n26611, 
        n26190, n26781, n26000, n25621, n27074, n25187, n26636, n26027, n25195, 
        n27356, n27363, n26317, n26496, n27053, n25606, n25796, n26506, n26287, 
        n26974, n25944, n25327, n25536, n26941, n26322, n26533, n25282, n25503, 
        n25312, n25493, n25971, n26603, n26793, n26012, n26182, n27066, n25633, 
        n26624, n26035, n27041, n25784, n25057, n27371, n25614, n26966, n26514, 
        n26295, n26305, n26484, n25335, n25524, n25956, n26428, n25209, n25588, 
        n25399, n25418, n25728, n26239, n25139, n27338, n26688, n26718, n26099, 
        n26109, n26751, n25761, n27134, n25170, n26140, n27204, n25240, n25451, 
        n25823, n26813, n26983, n26270, n26461, n25267, n25476, n26834, n27223, 
        n25804, n25994, n26257, n26446, n27083, n27113, n25746, n25157, n26776, 
        n26167, n26898, n26908, n25938, n27198, n27008, n27183, n27013, n25070, 
        n27294, n27304, n27323, n25646, n26676, n26067, n25367, n25576, n26934, 
        n25894, n25904, n26546, n26357, n25340, n25551, n25923, n26883, n26913, 
        n26370, n26561, n27034, n25661, n26651, n26040, n27098, n27108, n25186, 
        n26808, n27238, n26998, n25838, n26866, n26584, n26205, n26395, n26414, 
        n25424, n25235, n25856, n27271, n26135, n26724, n27141, n25095, n25714, 
        n26703, n25684, n25105, n26082, n26693, n26112, n27166, n25122, n25733, 
        n26841, n26433, n26222, n25212, n25593, n25382, n25403, n27256, n25871, 
        n25628, n26618, n26788, n26009, n26199, n27345, n27279, n26339, n25299, 
        n25518, n25309, n25488, n26528, n26849, n25879, n27149, n25962, n25291, 
        n25301, n25510, n25480, n26331, n26520, n26952, n25620, n27075, 
        \holder[3] , n26780, n26001, n26610, n26191, n25797, n25607, n25078, 
        n27052, n26637, n26026, n27362, n25945, n25326, n25537, n26286, n26507, 
        n26316, n26497, n26975, n25669, n26378, n26659, n26048, n25348, n25559, 
        n26569, n27387, n26742, n26153, n25772, n25163, n27127, n26263, n26472, 
        n26800, n26990, n25830, n27217, n25253, n25442, n26244, n26455, n26827, 
        n27230, n25817, n25987, n25274, n25465, n26765, n26174, n25755, n25144, 
        n27090, n27100, n25063, n26469, n25248, n25459, n26278, n25769, n25178, 
        n26759, n26148, n26665, n26074, n27190, n25655, n27000, n26555, n26344, 
        n26927, n25887, n27287, n27317, n27330, n25917, n25374, n25565, n26363, 
        n26572, n26890, n26900, n25930, n25353, n25542, n26642, n26053, n25672, 
        n27379, n27027, n27049, n25201, n25086, n27262, n26949, n25979, n25845, 
        n25437, n25226, n26216, n26386, n26597, n26407, n26875, n25707, n25697, 
        n25116, n27152, n26126, n26737, n25720, n25131, n27175, n26680, n26710, 
        n26091, n26101, n25862, n27245, n25056, n25094, n25391, n25580, n25410, 
        n26420, n26231, n26852, n25234, n25425, n25857, n27270, n26394, n26867, 
        n26415, n26204, n26585, n27140, n25685, n25715, n25104, n27257, n26725, 
        n26134, n27167, n25732, n25123, n26692, n26702, n26113, n26083, n25213, 
        n25383, n25402, n25592, n25870, n26432, n26840, n26223, n26619, n26789, 
        n26198, n26008, n25629, n26338, n26529, n25298, n25308, n25489, n25519, 
        n26066, n26677, n27012, n27182, n25647, n25071, n27322, n26935, n26356, 
        n26547, n25577, n25366, n27295, n25905, n26912, n25895, n26882, n26371, 
        n26560, n25341, n25550, n25922, n27305, n26650, n26041, n27035, 
        \holder[7] , n25660, n27239, n27099, n27109, n25839, n26809, n26999, 
        n26141, n26750, n25760, n27135, n25171, n26812, n26982, n26271, n26460, 
        n27205, n25241, n25450, n25822, n26835, n26447, n26256, n25266, n25477, 
        n27222, n25805, n25995, n26777, n26166, n27082, n27112, n25156, n25747, 
        n26909, n25939, n25193, n25194, n27339, n26899, n27357, n27199, n27009, 
        n25283, n25313, n25492, n25502, n25970, n26940, n26323, n26532, n27067, 
        n26602, n25632, n26792, n26183, n26013, n27040, n25615, n25208, n27370, 
        n25785, n26034, n26625, n25525, n25334, n26967, n25957, n26294, n26304, 
        n26485, n26515, n26429, n26238, n25398, n25419, n27377, n25589, n26689, 
        n26719, n26108, n26098, n25729, n25138, n26293, n26512, n26303, n26482, 
        n26960, n25950, n25333, n25522, n26622, n25782, n26033, n27392, n25088, 
        n25612, n27047, n26605, n26795, n26014, n26184, n25635, n27060, n26324, 
        n26535, n26947, n25977, n27350, n25284, n25505, n25314, n25495, n26599, 
        n25228, n25439, n26218, n26388, n26409, n25699, n25709, n25118, n26739, 
        n26128, n25740, n27085, n27115, n25151, n26161, n26770, n27225, n25802, 
        n25992, n25261, n25470, n26440, n26251, n26832, n27202, n25825, n25246, 
        n25457, n26276, n26467, n26815, n26985, n25767, n25176, n27132, n26757, 
        n26146, n26929, Logic01, n25076, n27289, n27319, n25889, n25919, 
        n27029, n25667, n27292, n27302, n27032, n26046, n26657, n25925, n27325, 
        n25557, n25346, n26376, n26567, n26885, n26915, n25892, n25902, n25361, 
        n25570, n26351, n26540, n26932, n27389, n25640, \holder[5] , n27185, 
        n27015, n26670, n27129, n26061, n27219, n26829, n25188, n25093, n25819, 
        n25989, n26435, n27250, n26847, n26224, n25877, n25595, n26705, n25214, 
        n25384, n25405, n26084, n26114, n26695, n25124, n25735, n27160, n26722, 
        n26133, n27277, n25682, n25712, n25103, n27147, n26393, n26412, n26582, 
        n26203, n26860, n25850, n25233, n25422, n25799, n27359, n25609, n26288, 
        n26509, n26639, n25328, n26028, n25539, n26499, n26318, n27069, n25959, 
        n26969, n26855, n25206, n26427, n26236, n25396, n25417, n25587, n25058, 
        n25064, n25081, n25865, n27242, n26687, n26106, n26717, n26096, n27172, 
        n25727, n25136, n26730, n26121, n25690, n27155, n25111, n27265, n25700, 
        n26872, n26381, n26400, n26590, n26211, n25221, n25430, n25842, n26449, 
        n26258, n25268, n25479, n26779, n26168, n25749, n25158, n27020, n27310, 
        n27280, n25675, n26645, n26054, n25354, n25545, n25937, n27337, n26897, 
        n26907, n26575, n26364, n25373, n25562, n25910, n25880, n26920, n26343, 
        n26552, n27007, n27197, n26662, n25652, n26073, n26679, n26068, n25649, 
        n26358, n26549, n25368, n25579, n27097, n25752, n27107, n25143, n26762, 
        n26173, n25273, n25462, n27237, n25810, n25980, n26820, n26452, n25445, 
        n26243, n25254, n27380, n27210, n25837, n26807, n26997, n26264, n26475, 
        n27120, n25775, n25164, n26154, n26745, n25859, n26869, n27169, n27365, 
        n27259, n26972, n26281, n26311, n26490, n26500, n25321, n25530, n25942, 
        n26021, n26630, n27055, n25600, n25181, \holder[1] , n26617, n25790, 
        n26196, n26006, n26787, n27072, n25627, n27342, n26955, n26336, n26527, 
        n25487, n25296, n25306, n25517, n25965;
    tri \DataOut[31] , \DataOut[27]1 , \DataOut[14]1 , \DataOut[26]1 , 
        \DataOut[15]1 , \DataOut[18]1 , \DataOut[0]1 , \DataOut[19]1 , 
        \DataOut[1]1 , \DataOut[23]1 , \DataOut[22]1 , \DataOut[11]1 , 
        \DataOut[10]1 , \DataOut[9]1 , \DataOut[8]1 , \DataOut[5]1 , 
        \DataOut[4]1 , \DataOut[21]1 , \DataOut[20]1 , \DataOut[13]1 , 
        \DataOut[12]1 , \DataOut[7]1 , \DataOut[6]1 , \DataOut[25]1 , 
        \DataOut[16]1 , \DataOut[24]1 , \DataOut[17]1 , \DataOut[29]1 , 
        \DataOut[30]1 , \DataOut[2]1 , \DataOut[28]1 , \DataOut[3]1 ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 ;
    assign DataOut[31] = \DataOut[31] ;
    assign DataOut[30] = \DataOut[30]1 ;
    assign DataOut[29] = \DataOut[29]1 ;
    assign DataOut[28] = \DataOut[28]1 ;
    assign DataOut[27] = \DataOut[27]1 ;
    assign DataOut[26] = \DataOut[26]1 ;
    assign DataOut[25] = \DataOut[25]1 ;
    assign DataOut[24] = \DataOut[24]1 ;
    assign DataOut[23] = \DataOut[23]1 ;
    assign DataOut[22] = \DataOut[22]1 ;
    assign DataOut[21] = \DataOut[21]1 ;
    assign DataOut[20] = \DataOut[20]1 ;
    assign DataOut[19] = \DataOut[19]1 ;
    assign DataOut[18] = \DataOut[18]1 ;
    assign DataOut[17] = \DataOut[17]1 ;
    assign DataOut[16] = \DataOut[16]1 ;
    assign DataOut[15] = \DataOut[15]1 ;
    assign DataOut[14] = \DataOut[14]1 ;
    assign DataOut[13] = \DataOut[13]1 ;
    assign DataOut[12] = \DataOut[12]1 ;
    assign DataOut[11] = \DataOut[11]1 ;
    assign DataOut[10] = \DataOut[10]1 ;
    assign DataOut[9] = \DataOut[9]1 ;
    assign DataOut[8] = \DataOut[8]1 ;
    assign DataOut[7] = \DataOut[7]1 ;
    assign DataOut[6] = \DataOut[6]1 ;
    assign DataOut[5] = \DataOut[5]1 ;
    assign DataOut[4] = \DataOut[4]1 ;
    assign DataOut[3] = \DataOut[3]1 ;
    assign DataOut[2] = \DataOut[2]1 ;
    assign DataOut[1] = \DataOut[1]1 ;
    assign DataOut[0] = \DataOut[0]1 ;
    VMW_PULLDOWN U271 ( .Z(n25189) );
    VMW_AO22 U338 ( .A(vectorInput[85]), .B(n25095), .C(vectorInput[77]), .D(
        n25080), .Z(n27307) );
    VMW_AO22 U394 ( .A(vectorInput[34]), .B(n25095), .C(vectorInput[26]), .D(
        n25080), .Z(n27358) );
    VMW_AO22 U415 ( .A(DataIn[2]), .B(n25095), .C(vectorInput[122]), .D(n25080
        ), .Z(n27262) );
    VMW_AO22 U432 ( .A(vectorInput[115]), .B(n25095), .C(vectorInput[107]), 
        .D(n25080), .Z(n27277) );
    VMW_FD \matrixInput_reg[1939]  ( .D(n25317), .CP(Clk), .Q(matrixInput
        [1939]) );
    VMW_FD \matrixInput_reg[1920]  ( .D(n25336), .CP(Clk), .Q(matrixInput
        [1920]) );
    VMW_FD \matrixInput_reg[3]  ( .D(n27253), .CP(Clk), .Q(matrixInput[3]) );
    VMW_AO22 U692 ( .A(matrixInput[782]), .B(n25096), .C(matrixInput[774]), 
        .D(n25081), .Z(n26482) );
    VMW_AO22 U840 ( .A(matrixInput[648]), .B(n25096), .C(matrixInput[640]), 
        .D(n25081), .Z(n26616) );
    VMW_FD \matrixInput_reg[883]  ( .D(n26373), .CP(Clk), .Q(matrixInput[883])
         );
    VMW_AO22 U702 ( .A(matrixInput[773]), .B(n25096), .C(matrixInput[765]), 
        .D(n25081), .Z(n26491) );
    VMW_AO22 U725 ( .A(matrixInput[752]), .B(n25096), .C(matrixInput[744]), 
        .D(n25081), .Z(n26512) );
    VMW_AO22 U1828 ( .A(matrixInput[1603]), .B(n25096), .C(matrixInput[1595]), 
        .D(n25081), .Z(n25661) );
    VMW_FD \matrixInput_reg[1913]  ( .D(n25343), .CP(Clk), .Q(matrixInput
        [1913]) );
    VMW_FD \vectorInput_reg[59]  ( .D(n27325), .CP(Clk), .Q(vectorInput[59])
         );
    VMW_FD \vectorInput_reg[40]  ( .D(n27344), .CP(Clk), .Q(vectorInput[40])
         );
    VMW_FD \matrixInput_reg[939]  ( .D(n26317), .CP(Clk), .Q(matrixInput[939])
         );
    VMW_FD \matrixInput_reg[920]  ( .D(n26336), .CP(Clk), .Q(matrixInput[920])
         );
    VMW_FD \matrixInput_reg[1883]  ( .D(n25373), .CP(Clk), .Q(matrixInput
        [1883]) );
    VMW_FD \vectorInput_reg[73]  ( .D(n27311), .CP(Clk), .Q(vectorInput[73])
         );
    VMW_AO22 U529 ( .A(matrixInput[928]), .B(n25096), .C(matrixInput[920]), 
        .D(n25081), .Z(n26336) );
    VMW_AO22 U585 ( .A(matrixInput[878]), .B(n25096), .C(matrixInput[870]), 
        .D(n25081), .Z(n26386) );
    VMW_AO22 U867 ( .A(matrixInput[624]), .B(n25096), .C(matrixInput[616]), 
        .D(n25081), .Z(n26640) );
    VMW_FD \matrixInput_reg[1370]  ( .D(n25886), .CP(Clk), .Q(matrixInput
        [1370]) );
    VMW_FD \matrixInput_reg[1369]  ( .D(n25887), .CP(Clk), .Q(matrixInput
        [1369]) );
    VMW_FD \matrixInput_reg[913]  ( .D(n26343), .CP(Clk), .Q(matrixInput[913])
         );
    VMW_AO22 U2077 ( .A(matrixInput[1378]), .B(n25096), .C(matrixInput[1370]), 
        .D(n25081), .Z(n25886) );
    VMW_FD \matrixInput_reg[567]  ( .D(n26689), .CP(Clk), .Q(matrixInput[567])
         );
    VMW_AO22 U356 ( .A(vectorInput[68]), .B(n25095), .C(vectorInput[60]), .D(
        n25080), .Z(n27324) );
    VMW_AO22 U371 ( .A(vectorInput[55]), .B(n25095), .C(vectorInput[47]), .D(
        n25080), .Z(n27337) );
    VMW_AO22 U560 ( .A(matrixInput[901]), .B(n25096), .C(matrixInput[893]), 
        .D(n25081), .Z(n26363) );
    VMW_AO22 U619 ( .A(matrixInput[91]), .B(n25096), .C(matrixInput[83]), .D(
        n25081), .Z(n27173) );
    VMW_AO22 U1047 ( .A(matrixInput[462]), .B(n25096), .C(matrixInput[454]), 
        .D(n25081), .Z(n26802) );
    VMW_FD \matrixInput_reg[1073]  ( .D(n26183), .CP(Clk), .Q(matrixInput
        [1073]) );
    VMW_FD \matrixInput_reg[664]  ( .D(n26592), .CP(Clk), .Q(matrixInput[664])
         );
    VMW_AO22 U1656 ( .A(matrixInput[182]), .B(n25096), .C(matrixInput[174]), 
        .D(n25081), .Z(n27082) );
    VMW_AO22 U2556 ( .A(cOutput[80]), .B(n25087), .C(cOutput[64]), .D(n25084), 
        .Z(n25178) );
    VMW_AO22 U650 ( .A(matrixInput[819]), .B(n25096), .C(matrixInput[811]), 
        .D(n25081), .Z(n26445) );
    VMW_AO22 U789 ( .A(matrixInput[695]), .B(n25096), .C(matrixInput[687]), 
        .D(n25081), .Z(n26569) );
    VMW_AO22 U2347 ( .A(matrixInput[1135]), .B(n25096), .C(matrixInput[1127]), 
        .D(n25081), .Z(n26129) );
    VMW_FD \matrixInput_reg[554]  ( .D(n26702), .CP(Clk), .Q(matrixInput[554])
         );
    VMW_AO22 U1060 ( .A(matrixInput[450]), .B(n25096), .C(matrixInput[442]), 
        .D(n25081), .Z(n26814) );
    VMW_AO22 U1350 ( .A(matrixInput[2032]), .B(n25096), .C(matrixInput[2024]), 
        .D(n25081), .Z(n25232) );
    VMW_AO22 U1377 ( .A(matrixInput[9]), .B(n25096), .C(matrixInput[1]), .D(
        n25081), .Z(n27255) );
    VMW_AO22 U1884 ( .A(matrixInput[1552]), .B(n25096), .C(matrixInput[1544]), 
        .D(n25081), .Z(n25712) );
    VMW_FD \matrixInput_reg[1343]  ( .D(n25913), .CP(Clk), .Q(matrixInput
        [1343]) );
    VMW_AO22 U1914 ( .A(matrixInput[1525]), .B(n25096), .C(matrixInput[1517]), 
        .D(n25081), .Z(n25739) );
    VMW_AO22 U1541 ( .A(matrixInput[1861]), .B(n25096), .C(matrixInput[1853]), 
        .D(n25081), .Z(n25403) );
    VMW_AO22 U1566 ( .A(matrixInput[1838]), .B(n25096), .C(matrixInput[1830]), 
        .D(n25081), .Z(n25426) );
    VMW_FD \matrixInput_reg[657]  ( .D(n26599), .CP(Clk), .Q(matrixInput[657])
         );
    VMW_AO22 U1933 ( .A(matrixInput[22]), .B(n25096), .C(matrixInput[14]), .D(
        n25081), .Z(n27242) );
    VMW_AO22 U2360 ( .A(matrixInput[1123]), .B(n25096), .C(matrixInput[1115]), 
        .D(n25081), .Z(n26141) );
    VMW_FD \matrixInput_reg[2003]  ( .D(n25253), .CP(Clk), .Q(matrixInput
        [2003]) );
    VMW_FD \matrixInput_reg[1059]  ( .D(n26197), .CP(Clk), .Q(matrixInput
        [1059]) );
    VMW_FD \matrixInput_reg[1040]  ( .D(n26216), .CP(Clk), .Q(matrixInput
        [1040]) );
    VMW_OAI21 U2571 ( .A(n25119), .B(n25120), .C(n25090), .Z(n25128) );
    VMW_FD \matrixInput_reg[1664]  ( .D(n25592), .CP(Clk), .Q(matrixInput
        [1664]) );
    VMW_FD \matrixInput_reg[1567]  ( .D(n25689), .CP(Clk), .Q(matrixInput
        [1567]) );
    VMW_FD \matrixInput_reg[370]  ( .D(n26886), .CP(Clk), .Q(matrixInput[370])
         );
    VMW_FD \matrixInput_reg[369]  ( .D(n26887), .CP(Clk), .Q(matrixInput[369])
         );
    VMW_AO22 U1671 ( .A(matrixInput[1744]), .B(n25096), .C(matrixInput[1736]), 
        .D(n25081), .Z(n25520) );
    VMW_AO22 U2050 ( .A(matrixInput[1403]), .B(n25096), .C(matrixInput[1395]), 
        .D(n25081), .Z(n25861) );
    VMW_FD \matrixInput_reg[1554]  ( .D(n25702), .CP(Clk), .Q(matrixInput
        [1554]) );
    VMW_FD \matrixInput_reg[343]  ( .D(n26913), .CP(Clk), .Q(matrixInput[343])
         );
    VMW_FD \matrixInput_reg[2030]  ( .D(n25226), .CP(Clk), .Q(matrixInput
        [2030]) );
    VMW_FD \matrixInput_reg[2029]  ( .D(n25227), .CP(Clk), .Q(matrixInput
        [2029]) );
    VMW_FD \matrixInput_reg[1657]  ( .D(n25599), .CP(Clk), .Q(matrixInput
        [1657]) );
    VMW_FD \matrixInput_reg[11]  ( .D(n27245), .CP(Clk), .Q(matrixInput[11])
         );
    VMW_FD \matrixInput_reg[851]  ( .D(n26405), .CP(Clk), .Q(matrixInput[851])
         );
    VMW_FD \matrixInput_reg[848]  ( .D(n26408), .CP(Clk), .Q(matrixInput[848])
         );
    VMW_AO22 U882 ( .A(matrixInput[610]), .B(n25096), .C(matrixInput[602]), 
        .D(n25081), .Z(n26654) );
    VMW_AO22 U912 ( .A(matrixInput[584]), .B(n25096), .C(matrixInput[576]), 
        .D(n25081), .Z(n26680) );
    VMW_AO22 U2019 ( .A(matrixInput[1430]), .B(n25096), .C(matrixInput[1422]), 
        .D(n25081), .Z(n25834) );
    VMW_FD \matrixInput_reg[862]  ( .D(n26394), .CP(Clk), .Q(matrixInput[862])
         );
    VMW_FD \matrixInput_reg[22]  ( .D(n27234), .CP(Clk), .Q(matrixInput[22])
         );
    VMW_FD \vectorInput_reg[111]  ( .D(n27273), .CP(Clk), .Q(vectorInput[111])
         );
    VMW_AO22 U447 ( .A(matrixInput[1003]), .B(n25096), .C(matrixInput[995]), 
        .D(n25081), .Z(n26261) );
    VMW_AO22 U547 ( .A(matrixInput[912]), .B(n25096), .C(matrixInput[904]), 
        .D(n25081), .Z(n26352) );
    VMW_BUFIZ U2608 ( .A(n25185), .E(RD), .Z(\DataOut[27]1 ) );
    VMW_FD \vectorInput_reg[108]  ( .D(n27276), .CP(Clk), .Q(vectorInput[108])
         );
    VMW_AO22 U677 ( .A(matrixInput[796]), .B(n25096), .C(matrixInput[788]), 
        .D(n25081), .Z(n26468) );
    VMW_AO22 U935 ( .A(matrixInput[563]), .B(n25096), .C(matrixInput[555]), 
        .D(n25081), .Z(n26701) );
    VMW_AO22 U2189 ( .A(matrixInput[134]), .B(n25096), .C(matrixInput[126]), 
        .D(n25081), .Z(n27130) );
    VMW_AO22 U1029 ( .A(matrixInput[478]), .B(n25096), .C(matrixInput[470]), 
        .D(n25081), .Z(n26786) );
    VMW_AO22 U1638 ( .A(matrixInput[1774]), .B(n25096), .C(matrixInput[1766]), 
        .D(n25081), .Z(n25490) );
    VMW_FD \matrixInput_reg[1851]  ( .D(n25405), .CP(Clk), .Q(matrixInput
        [1851]) );
    VMW_FD \matrixInput_reg[1848]  ( .D(n25408), .CP(Clk), .Q(matrixInput
        [1848]) );
    VMW_AO22 U2329 ( .A(matrixInput[1151]), .B(n25096), .C(matrixInput[1143]), 
        .D(n25081), .Z(n26113) );
    VMW_AO22 U2538 ( .A(cOutput[82]), .B(n25087), .C(cOutput[66]), .D(n25084), 
        .Z(n25156) );
    VMW_FD \vectorInput_reg[122]  ( .D(n27262), .CP(Clk), .Q(vectorInput[122])
         );
    VMW_AO22 U777 ( .A(matrixInput[706]), .B(n25096), .C(matrixInput[698]), 
        .D(n25081), .Z(n26558) );
    VMW_AO22 U809 ( .A(matrixInput[677]), .B(n25096), .C(matrixInput[669]), 
        .D(n25081), .Z(n26587) );
    VMW_AO22 U999 ( .A(matrixInput[506]), .B(n25096), .C(matrixInput[498]), 
        .D(n25081), .Z(n26758) );
    VMW_AO22 U1085 ( .A(matrixInput[49]), .B(n25096), .C(matrixInput[41]), .D(
        n25081), .Z(n27215) );
    VMW_AO22 U1225 ( .A(matrixInput[302]), .B(n25096), .C(matrixInput[294]), 
        .D(n25081), .Z(n26962) );
    VMW_AO22 U1289 ( .A(matrixInput[244]), .B(n25096), .C(matrixInput[236]), 
        .D(n25081), .Z(n27020) );
    VMW_AO22 U1319 ( .A(matrixInput[217]), .B(n25096), .C(matrixInput[209]), 
        .D(n25081), .Z(n27047) );
    VMW_AO22 U1508 ( .A(matrixInput[1891]), .B(n25096), .C(matrixInput[1883]), 
        .D(n25081), .Z(n25373) );
    VMW_AO22 U1434 ( .A(matrixInput[202]), .B(n25096), .C(matrixInput[194]), 
        .D(n25081), .Z(n27062) );
    VMW_AO22 U1498 ( .A(matrixInput[1900]), .B(n25096), .C(matrixInput[1892]), 
        .D(n25081), .Z(n25364) );
    VMW_AO22 U1846 ( .A(matrixInput[1587]), .B(n25096), .C(matrixInput[1579]), 
        .D(n25081), .Z(n25677) );
    VMW_FD \matrixInput_reg[1862]  ( .D(n25394), .CP(Clk), .Q(matrixInput
        [1862]) );
    VMW_FD \vectorInput_reg[92]  ( .D(n27292), .CP(Clk), .Q(vectorInput[92])
         );
    VMW_FD \matrixInput_reg[1092]  ( .D(n26164), .CP(Clk), .Q(matrixInput
        [1092]) );
    VMW_FD \matrixInput_reg[685]  ( .D(n26571), .CP(Clk), .Q(matrixInput[685])
         );
    VMW_FD \matrixInput_reg[218]  ( .D(n27038), .CP(Clk), .Q(matrixInput[218])
         );
    VMW_FD \matrixInput_reg[201]  ( .D(n27055), .CP(Clk), .Q(matrixInput[201])
         );
    VMW_FD \matrixInput_reg[1416]  ( .D(n25840), .CP(Clk), .Q(matrixInput
        [1416]) );
    VMW_AO22 U1704 ( .A(matrixInput[1714]), .B(n25096), .C(matrixInput[1706]), 
        .D(n25081), .Z(n25550) );
    VMW_AO22 U2215 ( .A(matrixInput[1254]), .B(n25096), .C(matrixInput[1246]), 
        .D(n25081), .Z(n26010) );
    VMW_FD \matrixInput_reg[102]  ( .D(n27154), .CP(Clk), .Q(matrixInput[102])
         );
    VMW_AO22 U2385 ( .A(matrixInput[1101]), .B(n25096), .C(matrixInput[1093]), 
        .D(n25081), .Z(n26163) );
    VMW_OAI21 U2594 ( .A(n25180), .B(n25181), .C(n25094), .Z(n25057) );
    VMW_AO22 U2404 ( .A(matrixInput[1084]), .B(n25096), .C(matrixInput[1076]), 
        .D(n25081), .Z(n26180) );
    VMW_FD \matrixInput_reg[1715]  ( .D(n25541), .CP(Clk), .Q(matrixInput
        [1715]) );
    VMW_FD \matrixInput_reg[1391]  ( .D(n25865), .CP(Clk), .Q(matrixInput
        [1391]) );
    VMW_FD \matrixInput_reg[1388]  ( .D(n25868), .CP(Clk), .Q(matrixInput
        [1388]) );
    VMW_FD \matrixInput_reg[586]  ( .D(n26670), .CP(Clk), .Q(matrixInput[586])
         );
    VMW_FD \matrixInput_reg[1425]  ( .D(n25831), .CP(Clk), .Q(matrixInput
        [1425]) );
    VMW_AO22 U1115 ( .A(matrixInput[401]), .B(n25096), .C(matrixInput[393]), 
        .D(n25081), .Z(n26863) );
    VMW_AO22 U1694 ( .A(matrixInput[1723]), .B(n25096), .C(matrixInput[1715]), 
        .D(n25081), .Z(n25541) );
    VMW_FD \matrixInput_reg[232]  ( .D(n27024), .CP(Clk), .Q(matrixInput[232])
         );
    VMW_AO22 U1132 ( .A(matrixInput[386]), .B(n25096), .C(matrixInput[378]), 
        .D(n25081), .Z(n26878) );
    VMW_AO22 U2125 ( .A(matrixInput[1335]), .B(n25096), .C(matrixInput[1327]), 
        .D(n25081), .Z(n25929) );
    VMW_FD \matrixInput_reg[1726]  ( .D(n25530), .CP(Clk), .Q(matrixInput
        [1726]) );
    VMW_FD \matrixInput_reg[1685]  ( .D(n25571), .CP(Clk), .Q(matrixInput
        [1685]) );
    VMW_FD \matrixInput_reg[131]  ( .D(n27125), .CP(Clk), .Q(matrixInput[131])
         );
    VMW_FD \matrixInput_reg[128]  ( .D(n27128), .CP(Clk), .Q(matrixInput[128])
         );
    VMW_AO22 U1202 ( .A(matrixInput[322]), .B(n25096), .C(matrixInput[314]), 
        .D(n25081), .Z(n26942) );
    VMW_AO22 U1723 ( .A(matrixInput[176]), .B(n25096), .C(matrixInput[168]), 
        .D(n25081), .Z(n27088) );
    VMW_AO22 U1861 ( .A(matrixInput[1573]), .B(n25096), .C(matrixInput[1565]), 
        .D(n25081), .Z(n25691) );
    VMW_AO22 U2092 ( .A(matrixInput[1365]), .B(n25096), .C(matrixInput[1357]), 
        .D(n25081), .Z(n25899) );
    VMW_FD \matrixInput_reg[1586]  ( .D(n25670), .CP(Clk), .Q(matrixInput
        [1586]) );
    VMW_FD \matrixInput_reg[1218]  ( .D(n26038), .CP(Clk), .Q(matrixInput
        [1218]) );
    VMW_FD \matrixInput_reg[1201]  ( .D(n26055), .CP(Clk), .Q(matrixInput
        [1201]) );
    VMW_FD \matrixInput_reg[416]  ( .D(n26840), .CP(Clk), .Q(matrixInput[416])
         );
    VMW_FD \matrixInput_reg[1102]  ( .D(n26154), .CP(Clk), .Q(matrixInput
        [1102]) );
    VMW_FD \matrixInput_reg[715]  ( .D(n26541), .CP(Clk), .Q(matrixInput[715])
         );
    VMW_FD \matrixInput_reg[391]  ( .D(n26865), .CP(Clk), .Q(matrixInput[391])
         );
    VMW_AO22 U2102 ( .A(matrixInput[1356]), .B(n25096), .C(matrixInput[1348]), 
        .D(n25081), .Z(n25908) );
    VMW_FD \matrixInput_reg[388]  ( .D(n26868), .CP(Clk), .Q(matrixInput[388])
         );
    VMW_FD \matrixInput_reg[1232]  ( .D(n26024), .CP(Clk), .Q(matrixInput
        [1232]) );
    VMW_FD \matrixInput_reg[425]  ( .D(n26831), .CP(Clk), .Q(matrixInput[425])
         );
    VMW_AO22 U1392 ( .A(matrixInput[1996]), .B(n25096), .C(matrixInput[1988]), 
        .D(n25081), .Z(n25268) );
    VMW_AO22 U1583 ( .A(matrixInput[1823]), .B(n25096), .C(matrixInput[1815]), 
        .D(n25081), .Z(n25441) );
    VMW_AO22 U1413 ( .A(matrixInput[1977]), .B(n25096), .C(matrixInput[1969]), 
        .D(n25081), .Z(n25287) );
    VMW_AO22 U2232 ( .A(matrixInput[1238]), .B(n25096), .C(matrixInput[1230]), 
        .D(n25081), .Z(n26026) );
    VMW_AO22 U2423 ( .A(matrixInput[1067]), .B(n25096), .C(matrixInput[1059]), 
        .D(n25081), .Z(n26197) );
    VMW_AO22 U2438 ( .A(matrixInput[1053]), .B(n25096), .C(matrixInput[1045]), 
        .D(n25081), .Z(n26211) );
    VMW_FD \matrixInput_reg[1131]  ( .D(n26125), .CP(Clk), .Q(matrixInput
        [1131]) );
    VMW_FD \matrixInput_reg[1128]  ( .D(n26128), .CP(Clk), .Q(matrixInput
        [1128]) );
    VMW_FD \matrixInput_reg[726]  ( .D(n26530), .CP(Clk), .Q(matrixInput[726])
         );
    VMW_FD \vectorInput_reg[5]  ( .D(n27379), .CP(Clk), .Q(vectorInput[5]) );
    VMW_AO22 U1219 ( .A(matrixInput[37]), .B(n25096), .C(matrixInput[29]), .D(
        n25081), .Z(n27227) );
    VMW_AO22 U2229 ( .A(matrixInput[1241]), .B(n25096), .C(matrixInput[1233]), 
        .D(n25081), .Z(n26023) );
    VMW_FD \vectorInput_reg[82]  ( .D(n27302), .CP(Clk), .Q(vectorInput[82])
         );
    VMW_AO22 U1389 ( .A(matrixInput[1998]), .B(n25096), .C(matrixInput[1990]), 
        .D(n25081), .Z(n25266) );
    VMW_AO22 U1598 ( .A(matrixInput[1809]), .B(n25096), .C(matrixInput[1801]), 
        .D(n25081), .Z(n25455) );
    VMW_AO22 U1408 ( .A(matrixInput[1981]), .B(n25096), .C(matrixInput[1973]), 
        .D(n25081), .Z(n25283) );
    VMW_FD \matrixInput_reg[1872]  ( .D(n25384), .CP(Clk), .Q(matrixInput
        [1872]) );
    VMW_FD \vectorInput_reg[118]  ( .D(n27266), .CP(Clk), .Q(vectorInput[118])
         );
    VMW_AO22 U835 ( .A(matrixInput[653]), .B(n25096), .C(matrixInput[645]), 
        .D(n25081), .Z(n26611) );
    VMW_AO22 U2089 ( .A(matrixInput[143]), .B(n25096), .C(matrixInput[135]), 
        .D(n25081), .Z(n27121) );
    VMW_AO22 U2119 ( .A(matrixInput[1340]), .B(n25096), .C(matrixInput[1332]), 
        .D(n25081), .Z(n25924) );
    VMW_FD \vectorInput_reg[101]  ( .D(n27283), .CP(Clk), .Q(vectorInput[101])
         );
    VMW_AO22 U1129 ( .A(matrixInput[388]), .B(n25096), .C(matrixInput[380]), 
        .D(n25081), .Z(n26876) );
    VMW_FD \matrixInput_reg[1858]  ( .D(n25398), .CP(Clk), .Q(matrixInput
        [1858]) );
    VMW_FD \matrixInput_reg[1841]  ( .D(n25415), .CP(Clk), .Q(matrixInput
        [1841]) );
    VMW_AO22 U1738 ( .A(matrixInput[1684]), .B(n25096), .C(matrixInput[1676]), 
        .D(n25081), .Z(n25580) );
    VMW_OAI211 U294 ( .A(n25055), .B(n25056), .C(n25057), .D(n25058), .Z(
        n27392) );
    VMW_AND2 U304 ( .A(n25082), .B(n25085), .Z(n25084) );
    VMW_AO22 U460 ( .A(matrixInput[991]), .B(n25096), .C(matrixInput[983]), 
        .D(n25081), .Z(n26273) );
    VMW_AO22 U485 ( .A(matrixInput[968]), .B(n25096), .C(matrixInput[960]), 
        .D(n25081), .Z(n26296) );
    VMW_AO22 U750 ( .A(matrixInput[729]), .B(n25096), .C(matrixInput[721]), 
        .D(n25081), .Z(n26535) );
    VMW_AO22 U812 ( .A(matrixInput[674]), .B(n25096), .C(matrixInput[666]), 
        .D(n25081), .Z(n26590) );
    VMW_AO22 U982 ( .A(matrixInput[520]), .B(n25096), .C(matrixInput[512]), 
        .D(n25081), .Z(n26744) );
    VMW_FD \matrixInput_reg[32]  ( .D(n27224), .CP(Clk), .Q(matrixInput[32])
         );
    VMW_FD \matrixInput_reg[872]  ( .D(n26384), .CP(Clk), .Q(matrixInput[872])
         );
    VMW_FD \matrixInput_reg[18]  ( .D(n27238), .CP(Clk), .Q(matrixInput[18])
         );
    VMW_AO22 U899 ( .A(matrixInput[596]), .B(n25096), .C(matrixInput[588]), 
        .D(n25081), .Z(n26668) );
    VMW_AO22 U909 ( .A(matrixInput[587]), .B(n25096), .C(matrixInput[579]), 
        .D(n25081), .Z(n26677) );
    VMW_AO22 U1015 ( .A(matrixInput[491]), .B(n25096), .C(matrixInput[483]), 
        .D(n25081), .Z(n26773) );
    VMW_AO22 U1032 ( .A(matrixInput[476]), .B(n25096), .C(matrixInput[468]), 
        .D(n25081), .Z(n26788) );
    VMW_AO22 U1292 ( .A(matrixInput[241]), .B(n25096), .C(matrixInput[233]), 
        .D(n25081), .Z(n27023) );
    VMW_AO22 U1961 ( .A(matrixInput[1483]), .B(n25096), .C(matrixInput[1475]), 
        .D(n25081), .Z(n25781) );
    VMW_FD \matrixInput_reg[858]  ( .D(n26398), .CP(Clk), .Q(matrixInput[858])
         );
    VMW_FD \matrixInput_reg[841]  ( .D(n26415), .CP(Clk), .Q(matrixInput[841])
         );
    VMW_FD \matrixInput_reg[435]  ( .D(n26821), .CP(Clk), .Q(matrixInput[435])
         );
    VMW_FD \matrixInput_reg[1222]  ( .D(n26034), .CP(Clk), .Q(matrixInput
        [1222]) );
    VMW_AO22 U1302 ( .A(matrixInput[232]), .B(n25096), .C(matrixInput[224]), 
        .D(n25081), .Z(n27032) );
    VMW_AO22 U1513 ( .A(matrixInput[1887]), .B(n25096), .C(matrixInput[1879]), 
        .D(n25081), .Z(n25377) );
    VMW_AO22 U1483 ( .A(matrixInput[1913]), .B(n25096), .C(matrixInput[1905]), 
        .D(n25081), .Z(n25351) );
    VMW_AO22 U1623 ( .A(matrixInput[185]), .B(n25096), .C(matrixInput[177]), 
        .D(n25081), .Z(n27079) );
    VMW_AO22 U2332 ( .A(matrixInput[1148]), .B(n25096), .C(matrixInput[1140]), 
        .D(n25081), .Z(n26116) );
    VMW_AO22 U2523 ( .A(cOutput[124]), .B(n25089), .C(cOutput[108]), .D(n25088
        ), .Z(n25137) );
    VMW_FD \matrixInput_reg[1138]  ( .D(n26118), .CP(Clk), .Q(matrixInput
        [1138]) );
    VMW_FD \matrixInput_reg[1121]  ( .D(n26135), .CP(Clk), .Q(matrixInput
        [1121]) );
    VMW_FD \matrixInput_reg[736]  ( .D(n26520), .CP(Clk), .Q(matrixInput[736])
         );
    VMW_AO22 U1794 ( .A(matrixInput[1633]), .B(n25096), .C(matrixInput[1625]), 
        .D(n25081), .Z(n25631) );
    VMW_AO22 U2002 ( .A(matrixInput[1446]), .B(n25096), .C(matrixInput[1438]), 
        .D(n25081), .Z(n25818) );
    VMW_FD \matrixInput_reg[1695]  ( .D(n25561), .CP(Clk), .Q(matrixInput
        [1695]) );
    VMW_FD \matrixInput_reg[1211]  ( .D(n26045), .CP(Clk), .Q(matrixInput
        [1211]) );
    VMW_FD \matrixInput_reg[1208]  ( .D(n26048), .CP(Clk), .Q(matrixInput
        [1208]) );
    VMW_FD \matrixInput_reg[1112]  ( .D(n26144), .CP(Clk), .Q(matrixInput
        [1112]) );
    VMW_FD \matrixInput_reg[406]  ( .D(n26850), .CP(Clk), .Q(matrixInput[406])
         );
    VMW_FD \matrixInput_reg[705]  ( .D(n26551), .CP(Clk), .Q(matrixInput[705])
         );
    VMW_AO22 U2192 ( .A(matrixInput[1275]), .B(n25096), .C(matrixInput[1267]), 
        .D(n25081), .Z(n25989) );
    VMW_BUFIZ U2613 ( .A(n25189), .E(RD), .Z(\DataOut[14]1 ) );
    VMW_FD \matrixInput_reg[398]  ( .D(n26858), .CP(Clk), .Q(matrixInput[398])
         );
    VMW_FD \matrixInput_reg[1596]  ( .D(n25660), .CP(Clk), .Q(matrixInput
        [1596]) );
    VMW_FD \matrixInput_reg[381]  ( .D(n26875), .CP(Clk), .Q(matrixInput[381])
         );
    VMW_FD \matrixInput_reg[222]  ( .D(n27034), .CP(Clk), .Q(matrixInput[222])
         );
    VMW_AO22 U1185 ( .A(matrixInput[40]), .B(n25096), .C(matrixInput[32]), .D(
        n25081), .Z(n27224) );
    VMW_AO22 U1604 ( .A(matrixInput[1805]), .B(n25096), .C(matrixInput[1797]), 
        .D(n25081), .Z(n25459) );
    VMW_FD \matrixInput_reg[1435]  ( .D(n25821), .CP(Clk), .Q(matrixInput
        [1435]) );
    VMW_AO22 U1325 ( .A(DataIn[7]), .B(n25096), .C(matrixInput[2047]), .D(
        n25081), .Z(n25209) );
    VMW_AO22 U1946 ( .A(matrixInput[1497]), .B(n25096), .C(matrixInput[1489]), 
        .D(n25081), .Z(n25767) );
    VMW_AO22 U2025 ( .A(matrixInput[1425]), .B(n25096), .C(matrixInput[1417]), 
        .D(n25081), .Z(n25839) );
    VMW_BUFIZ U2634 ( .A(\holder[5] ), .E(RD), .Z(\DataOut[5]1 ) );
    VMW_FD \matrixInput_reg[1736]  ( .D(n25520), .CP(Clk), .Q(matrixInput
        [1736]) );
    VMW_FD \matrixInput_reg[138]  ( .D(n27118), .CP(Clk), .Q(matrixInput[138])
         );
    VMW_FD \matrixInput_reg[121]  ( .D(n27135), .CP(Clk), .Q(matrixInput[121])
         );
    VMW_FD \matrixInput_reg[695]  ( .D(n26561), .CP(Clk), .Q(matrixInput[695])
         );
    VMW_FD \matrixInput_reg[1082]  ( .D(n26174), .CP(Clk), .Q(matrixInput
        [1082]) );
    VMW_AO22 U1534 ( .A(matrixInput[193]), .B(n25096), .C(matrixInput[185]), 
        .D(n25081), .Z(n27071) );
    VMW_AO22 U2285 ( .A(matrixInput[1191]), .B(n25096), .C(matrixInput[1183]), 
        .D(n25081), .Z(n26073) );
    VMW_FD \matrixInput_reg[1406]  ( .D(n25850), .CP(Clk), .Q(matrixInput
        [1406]) );
    VMW_FD \matrixInput_reg[211]  ( .D(n27045), .CP(Clk), .Q(matrixInput[211])
         );
    VMW_FD \matrixInput_reg[208]  ( .D(n27048), .CP(Clk), .Q(matrixInput[208])
         );
    VMW_AO22 U2315 ( .A(matrixInput[1164]), .B(n25096), .C(matrixInput[1156]), 
        .D(n25081), .Z(n26100) );
    VMW_AO22 U2504 ( .A(cOutput[118]), .B(n25087), .C(cOutput[102]), .D(n25084
        ), .Z(n25114) );
    VMW_FD \matrixInput_reg[1705]  ( .D(n25551), .CP(Clk), .Q(matrixInput
        [1705]) );
    VMW_AO22 U2494 ( .A(cOutput[95]), .B(n25089), .C(cOutput[79]), .D(n25088), 
        .Z(n25102) );
    VMW_FD \matrixInput_reg[1893]  ( .D(n25363), .CP(Clk), .Q(matrixInput
        [1893]) );
    VMW_FD \matrixInput_reg[1398]  ( .D(n25858), .CP(Clk), .Q(matrixInput
        [1398]) );
    VMW_FD \matrixInput_reg[596]  ( .D(n26660), .CP(Clk), .Q(matrixInput[596])
         );
    VMW_FD \matrixInput_reg[112]  ( .D(n27144), .CP(Clk), .Q(matrixInput[112])
         );
    VMW_FD \matrixInput_reg[1381]  ( .D(n25875), .CP(Clk), .Q(matrixInput
        [1381]) );
    VMW_FD \vectorInput_reg[63]  ( .D(n27321), .CP(Clk), .Q(vectorInput[63])
         );
    VMW_AO22 U515 ( .A(matrixInput[941]), .B(n25096), .C(matrixInput[933]), 
        .D(n25081), .Z(n26323) );
    VMW_AO22 U323 ( .A(vectorInput[98]), .B(n25095), .C(vectorInput[90]), .D(
        n25080), .Z(n27294) );
    VMW_AO22 U532 ( .A(matrixInput[926]), .B(n25096), .C(matrixInput[918]), 
        .D(n25081), .Z(n26338) );
    VMW_AO22 U602 ( .A(matrixInput[863]), .B(n25096), .C(matrixInput[855]), 
        .D(n25081), .Z(n26401) );
    VMW_AO22 U625 ( .A(matrixInput[842]), .B(n25096), .C(matrixInput[834]), 
        .D(n25081), .Z(n26422) );
    VMW_AO22 U967 ( .A(matrixInput[534]), .B(n25096), .C(matrixInput[526]), 
        .D(n25081), .Z(n26730) );
    VMW_FD \matrixInput_reg[903]  ( .D(n26353), .CP(Clk), .Q(matrixInput[903])
         );
    VMW_AO22 U1928 ( .A(matrixInput[1512]), .B(n25096), .C(matrixInput[1504]), 
        .D(n25081), .Z(n25752) );
    VMW_FD \matrixInput_reg[930]  ( .D(n26326), .CP(Clk), .Q(matrixInput[930])
         );
    VMW_FD \vectorInput_reg[50]  ( .D(n27334), .CP(Clk), .Q(vectorInput[50])
         );
    VMW_FD \vectorInput_reg[49]  ( .D(n27335), .CP(Clk), .Q(vectorInput[49])
         );
    VMW_FD \matrixInput_reg[929]  ( .D(n26327), .CP(Clk), .Q(matrixInput[929])
         );
    VMW_FD \matrixInput_reg[1903]  ( .D(n25353), .CP(Clk), .Q(matrixInput
        [1903]) );
    VMW_FD \matrixInput_reg[893]  ( .D(n26363), .CP(Clk), .Q(matrixInput[893])
         );
    VMW_AO22 U792 ( .A(matrixInput[692]), .B(n25096), .C(matrixInput[684]), 
        .D(n25081), .Z(n26572) );
    VMW_AO22 U429 ( .A(vectorInput[18]), .B(n25095), .C(vectorInput[10]), .D(
        n25080), .Z(n27374) );
    VMW_AO22 U689 ( .A(matrixInput[785]), .B(n25096), .C(matrixInput[777]), 
        .D(n25081), .Z(n26479) );
    VMW_AO22 U940 ( .A(matrixInput[558]), .B(n25096), .C(matrixInput[550]), 
        .D(n25081), .Z(n26706) );
    VMW_FD \matrixInput_reg[1930]  ( .D(n25326), .CP(Clk), .Q(matrixInput
        [1930]) );
    VMW_FD \matrixInput_reg[1929]  ( .D(n25327), .CP(Clk), .Q(matrixInput
        [1929]) );
    VMW_AO22 U1160 ( .A(matrixInput[360]), .B(n25096), .C(matrixInput[352]), 
        .D(n25081), .Z(n26904) );
    VMW_AO22 U2150 ( .A(matrixInput[1312]), .B(n25096), .C(matrixInput[1304]), 
        .D(n25081), .Z(n25952) );
    VMW_FD \matrixInput_reg[2039]  ( .D(n25217), .CP(Clk), .Q(matrixInput
        [2039]) );
    VMW_FD \matrixInput_reg[2020]  ( .D(n25236), .CP(Clk), .Q(matrixInput
        [2020]) );
    VMW_FD \matrixInput_reg[1544]  ( .D(n25712), .CP(Clk), .Q(matrixInput
        [1544]) );
    VMW_FD \matrixInput_reg[353]  ( .D(n26903), .CP(Clk), .Q(matrixInput[353])
         );
    VMW_AO22 U1250 ( .A(matrixInput[279]), .B(n25096), .C(matrixInput[271]), 
        .D(n25081), .Z(n26985) );
    VMW_AO22 U1771 ( .A(matrixInput[1654]), .B(n25096), .C(matrixInput[1646]), 
        .D(n25081), .Z(n25610) );
    VMW_AO22 U1833 ( .A(matrixInput[1598]), .B(n25096), .C(matrixInput[1590]), 
        .D(n25081), .Z(n25666) );
    VMW_AO22 U2260 ( .A(matrixInput[1213]), .B(n25096), .C(matrixInput[1205]), 
        .D(n25081), .Z(n26051) );
    VMW_AO22 U2471 ( .A(matrixInput[1023]), .B(n25096), .C(matrixInput[1015]), 
        .D(n25081), .Z(n26241) );
    VMW_FD \matrixInput_reg[1647]  ( .D(n25609), .CP(Clk), .Q(matrixInput
        [1647]) );
    VMW_FD \matrixInput_reg[2013]  ( .D(n25243), .CP(Clk), .Q(matrixInput
        [2013]) );
    VMW_FD \matrixInput_reg[1577]  ( .D(n25679), .CP(Clk), .Q(matrixInput
        [1577]) );
    VMW_FD \matrixInput_reg[379]  ( .D(n26877), .CP(Clk), .Q(matrixInput[379])
         );
    VMW_FD \matrixInput_reg[360]  ( .D(n26896), .CP(Clk), .Q(matrixInput[360])
         );
    VMW_FD \matrixInput_reg[1674]  ( .D(n25582), .CP(Clk), .Q(matrixInput
        [1674]) );
    VMW_AO22 U1441 ( .A(matrixInput[1951]), .B(n25096), .C(matrixInput[1943]), 
        .D(n25081), .Z(n25313) );
    VMW_AO22 U2247 ( .A(matrixInput[1225]), .B(n25096), .C(matrixInput[1217]), 
        .D(n25081), .Z(n26039) );
    VMW_FD \matrixInput_reg[1353]  ( .D(n25903), .CP(Clk), .Q(matrixInput
        [1353]) );
    VMW_AO22 U719 ( .A(matrixInput[82]), .B(n25096), .C(matrixInput[74]), .D(
        n25081), .Z(n27182) );
    VMW_AO22 U2456 ( .A(matrixInput[1037]), .B(n25096), .C(matrixInput[1029]), 
        .D(n25081), .Z(n26227) );
    VMW_FD \matrixInput_reg[544]  ( .D(n26712), .CP(Clk), .Q(matrixInput[544])
         );
    VMW_AO22 U1277 ( .A(matrixInput[255]), .B(n25096), .C(matrixInput[247]), 
        .D(n25081), .Z(n27009) );
    VMW_AO22 U1466 ( .A(matrixInput[1928]), .B(n25096), .C(matrixInput[1920]), 
        .D(n25081), .Z(n25336) );
    VMW_AO22 U1814 ( .A(matrixInput[1615]), .B(n25096), .C(matrixInput[1607]), 
        .D(n25081), .Z(n25649) );
    VMW_AO22 U1984 ( .A(matrixInput[1462]), .B(n25096), .C(matrixInput[1454]), 
        .D(n25081), .Z(n25802) );
    VMW_FD \matrixInput_reg[1050]  ( .D(n26206), .CP(Clk), .Q(matrixInput
        [1050]) );
    VMW_FD \matrixInput_reg[1049]  ( .D(n26207), .CP(Clk), .Q(matrixInput
        [1049]) );
    VMW_AO22 U2177 ( .A(matrixInput[1288]), .B(n25096), .C(matrixInput[1280]), 
        .D(n25081), .Z(n25976) );
    VMW_FD \matrixInput_reg[647]  ( .D(n26609), .CP(Clk), .Q(matrixInput[647])
         );
    VMW_FD \matrixInput_reg[577]  ( .D(n26679), .CP(Clk), .Q(matrixInput[577])
         );
    VMW_AO22 U1147 ( .A(matrixInput[372]), .B(n25096), .C(matrixInput[364]), 
        .D(n25081), .Z(n26892) );
    VMW_AO22 U1756 ( .A(matrixInput[173]), .B(n25096), .C(matrixInput[165]), 
        .D(n25081), .Z(n27091) );
    VMW_FD \matrixInput_reg[1379]  ( .D(n25877), .CP(Clk), .Q(matrixInput
        [1379]) );
    VMW_FD \matrixInput_reg[1360]  ( .D(n25896), .CP(Clk), .Q(matrixInput
        [1360]) );
    VMW_FD \matrixInput_reg[674]  ( .D(n26582), .CP(Clk), .Q(matrixInput[674])
         );
    VMW_AO22 U1172 ( .A(matrixInput[349]), .B(n25096), .C(matrixInput[341]), 
        .D(n25081), .Z(n26915) );
    VMW_AO22 U1763 ( .A(matrixInput[1661]), .B(n25096), .C(matrixInput[1653]), 
        .D(n25081), .Z(n25603) );
    VMW_AO22 U2142 ( .A(matrixInput[1319]), .B(n25096), .C(matrixInput[1311]), 
        .D(n25081), .Z(n25945) );
    VMW_FD \matrixInput_reg[1063]  ( .D(n26193), .CP(Clk), .Q(matrixInput
        [1063]) );
    VMW_FD \matrixInput_reg[1582]  ( .D(n25674), .CP(Clk), .Q(matrixInput
        [1582]) );
    VMW_FD \matrixInput_reg[395]  ( .D(n26861), .CP(Clk), .Q(matrixInput[395])
         );
    VMW_FD \matrixInput_reg[1205]  ( .D(n26051), .CP(Clk), .Q(matrixInput
        [1205]) );
    VMW_FD \matrixInput_reg[1106]  ( .D(n26150), .CP(Clk), .Q(matrixInput
        [1106]) );
    VMW_FD \matrixInput_reg[711]  ( .D(n26545), .CP(Clk), .Q(matrixInput[711])
         );
    VMW_FD \matrixInput_reg[708]  ( .D(n26548), .CP(Clk), .Q(matrixInput[708])
         );
    VMW_FD \matrixInput_reg[412]  ( .D(n26844), .CP(Clk), .Q(matrixInput[412])
         );
    VMW_AO22 U1242 ( .A(matrixInput[287]), .B(n25096), .C(matrixInput[279]), 
        .D(n25081), .Z(n26977) );
    VMW_AO22 U1453 ( .A(matrixInput[1940]), .B(n25096), .C(matrixInput[1932]), 
        .D(n25081), .Z(n25324) );
    VMW_AO22 U2272 ( .A(matrixInput[1203]), .B(n25096), .C(matrixInput[1195]), 
        .D(n25081), .Z(n26061) );
    VMW_FD \matrixInput_reg[1698]  ( .D(n25558), .CP(Clk), .Q(matrixInput
        [1698]) );
    VMW_FD \matrixInput_reg[1681]  ( .D(n25575), .CP(Clk), .Q(matrixInput
        [1681]) );
    VMW_FD \matrixInput_reg[1135]  ( .D(n26121), .CP(Clk), .Q(matrixInput
        [1135]) );
    VMW_FD \matrixInput_reg[722]  ( .D(n26534), .CP(Clk), .Q(matrixInput[722])
         );
    VMW_FD \vectorInput_reg[1]  ( .D(n27383), .CP(Clk), .Q(vectorInput[1]) );
    VMW_AO22 U2463 ( .A(matrixInput[1030]), .B(n25096), .C(matrixInput[1022]), 
        .D(n25081), .Z(n26234) );
    VMW_AO22 U1821 ( .A(matrixInput[1608]), .B(n25096), .C(matrixInput[1600]), 
        .D(n25081), .Z(n25656) );
    VMW_FD \matrixInput_reg[438]  ( .D(n26818), .CP(Clk), .Q(matrixInput[438])
         );
    VMW_FD \matrixInput_reg[421]  ( .D(n26835), .CP(Clk), .Q(matrixInput[421])
         );
    VMW_FD \matrixInput_reg[1236]  ( .D(n26020), .CP(Clk), .Q(matrixInput
        [1236]) );
    VMW_PULLDOWN U276 ( .Z(n25194) );
    VMW_PULLDOWN U278 ( .Z(n25196) );
    VMW_PULLDOWN U286 ( .Z(n25204) );
    VMW_AO22 U507 ( .A(matrixInput[948]), .B(n25096), .C(matrixInput[940]), 
        .D(n25081), .Z(n26316) );
    VMW_AO22 U849 ( .A(matrixInput[640]), .B(n25096), .C(matrixInput[632]), 
        .D(n25081), .Z(n26624) );
    VMW_AO22 U1265 ( .A(matrixInput[266]), .B(n25096), .C(matrixInput[258]), 
        .D(n25081), .Z(n26998) );
    VMW_AO22 U2255 ( .A(matrixInput[128]), .B(n25096), .C(matrixInput[120]), 
        .D(n25081), .Z(n27136) );
    VMW_AO22 U2444 ( .A(matrixInput[111]), .B(n25096), .C(matrixInput[103]), 
        .D(n25081), .Z(n27153) );
    VMW_FD \matrixInput_reg[1711]  ( .D(n25545), .CP(Clk), .Q(matrixInput
        [1711]) );
    VMW_FD \matrixInput_reg[1395]  ( .D(n25861), .CP(Clk), .Q(matrixInput
        [1395]) );
    VMW_FD \matrixInput_reg[582]  ( .D(n26674), .CP(Clk), .Q(matrixInput[582])
         );
    VMW_FD \matrixInput_reg[1708]  ( .D(n25548), .CP(Clk), .Q(matrixInput
        [1708]) );
    VMW_FD \matrixInput_reg[106]  ( .D(n27150), .CP(Clk), .Q(matrixInput[106])
         );
    VMW_AO22 U1474 ( .A(matrixInput[1921]), .B(n25096), .C(matrixInput[1913]), 
        .D(n25081), .Z(n25343) );
    VMW_AO22 U1806 ( .A(matrixInput[1622]), .B(n25096), .C(matrixInput[1614]), 
        .D(n25081), .Z(n25642) );
    VMW_AO22 U1996 ( .A(matrixInput[1451]), .B(n25096), .C(matrixInput[1443]), 
        .D(n25081), .Z(n25813) );
    VMW_FD \matrixInput_reg[1412]  ( .D(n25844), .CP(Clk), .Q(matrixInput
        [1412]) );
    VMW_FD \matrixInput_reg[681]  ( .D(n26575), .CP(Clk), .Q(matrixInput[681])
         );
    VMW_FD \matrixInput_reg[205]  ( .D(n27051), .CP(Clk), .Q(matrixInput[205])
         );
    VMW_FD \matrixInput_reg[698]  ( .D(n26558), .CP(Clk), .Q(matrixInput[698])
         );
    VMW_AO22 U2165 ( .A(matrixInput[1299]), .B(n25096), .C(matrixInput[1291]), 
        .D(n25081), .Z(n25965) );
    VMW_FD \matrixInput_reg[1722]  ( .D(n25534), .CP(Clk), .Q(matrixInput
        [1722]) );
    VMW_FD \matrixInput_reg[1096]  ( .D(n26160), .CP(Clk), .Q(matrixInput
        [1096]) );
    VMW_FD \matrixInput_reg[135]  ( .D(n27121), .CP(Clk), .Q(matrixInput[135])
         );
    VMW_AO22 U975 ( .A(matrixInput[527]), .B(n25096), .C(matrixInput[519]), 
        .D(n25081), .Z(n26737) );
    VMW_AO22 U1069 ( .A(matrixInput[442]), .B(n25096), .C(matrixInput[434]), 
        .D(n25081), .Z(n26822) );
    VMW_AO22 U1155 ( .A(matrixInput[365]), .B(n25096), .C(matrixInput[357]), 
        .D(n25081), .Z(n26899) );
    VMW_FD \matrixInput_reg[1438]  ( .D(n25818), .CP(Clk), .Q(matrixInput
        [1438]) );
    VMW_FD \matrixInput_reg[236]  ( .D(n27020), .CP(Clk), .Q(matrixInput[236])
         );
    VMW_AO22 U1744 ( .A(matrixInput[1678]), .B(n25096), .C(matrixInput[1670]), 
        .D(n25081), .Z(n25586) );
    VMW_FD \matrixInput_reg[1421]  ( .D(n25835), .CP(Clk), .Q(matrixInput
        [1421]) );
    VMW_AO22 U1678 ( .A(matrixInput[180]), .B(n25096), .C(matrixInput[172]), 
        .D(n25081), .Z(n27084) );
    VMW_FD \matrixInput_reg[1855]  ( .D(n25401), .CP(Clk), .Q(matrixInput
        [1855]) );
    VMW_AO22 U316 ( .A(vectorInput[105]), .B(n25095), .C(vectorInput[97]), .D(
        n25080), .Z(n27287) );
    VMW_AO22 U497 ( .A(matrixInput[102]), .B(n25096), .C(matrixInput[94]), .D(
        n25081), .Z(n27162) );
    VMW_FD \vectorInput_reg[115]  ( .D(n27269), .CP(Clk), .Q(vectorInput[115])
         );
    VMW_AO22 U2059 ( .A(matrixInput[1395]), .B(n25096), .C(matrixInput[1387]), 
        .D(n25081), .Z(n25869) );
    VMW_AO22 U331 ( .A(vectorInput[91]), .B(n25095), .C(vectorInput[83]), .D(
        n25080), .Z(n27301) );
    VMW_AO22 U610 ( .A(matrixInput[856]), .B(n25096), .C(matrixInput[848]), 
        .D(n25081), .Z(n26408) );
    VMW_AO22 U637 ( .A(matrixInput[831]), .B(n25096), .C(matrixInput[823]), 
        .D(n25081), .Z(n26433) );
    VMW_AO22 U1359 ( .A(matrixInput[2024]), .B(n25096), .C(matrixInput[2016]), 
        .D(n25081), .Z(n25240) );
    VMW_FD \matrixInput_reg[1866]  ( .D(n25390), .CP(Clk), .Q(matrixInput
        [1866]) );
    VMW_FD \vectorInput_reg[96]  ( .D(n27288), .CP(Clk), .Q(vectorInput[96])
         );
    VMW_AO22 U1548 ( .A(matrixInput[1855]), .B(n25096), .C(matrixInput[1847]), 
        .D(n25081), .Z(n25409) );
    VMW_OAI21 U2578 ( .A(n25136), .B(n25137), .C(n25094), .Z(n25069) );
    VMW_AO22 U780 ( .A(matrixInput[703]), .B(n25096), .C(matrixInput[695]), 
        .D(n25081), .Z(n26561) );
    VMW_AO22 U2369 ( .A(matrixInput[1115]), .B(n25096), .C(matrixInput[1107]), 
        .D(n25081), .Z(n26149) );
    VMW_FD \matrixInput_reg[855]  ( .D(n26401), .CP(Clk), .Q(matrixInput[855])
         );
    VMW_FD \vectorInput_reg[126]  ( .D(n27258), .CP(Clk), .Q(vectorInput[126])
         );
    VMW_AO22 U952 ( .A(matrixInput[61]), .B(n25096), .C(matrixInput[53]), .D(
        n25081), .Z(n27203) );
    VMW_FD \matrixInput_reg[866]  ( .D(n26390), .CP(Clk), .Q(matrixInput[866])
         );
    VMW_FD \matrixInput_reg[15]  ( .D(n27241), .CP(Clk), .Q(matrixInput[15])
         );
    VMW_FD \matrixInput_reg[26]  ( .D(n27230), .CP(Clk), .Q(matrixInput[26])
         );
    VMW_AO22 U378 ( .A(vectorInput[48]), .B(n25095), .C(vectorInput[40]), .D(
        n25080), .Z(n27344) );
    VMW_AO22 U520 ( .A(matrixInput[937]), .B(n25096), .C(matrixInput[929]), 
        .D(n25081), .Z(n26327) );
    VMW_AO22 U1007 ( .A(matrixInput[498]), .B(n25096), .C(matrixInput[490]), 
        .D(n25081), .Z(n26766) );
    VMW_AO22 U1020 ( .A(matrixInput[487]), .B(n25096), .C(matrixInput[479]), 
        .D(n25081), .Z(n26777) );
    VMW_AO22 U1280 ( .A(matrixInput[252]), .B(n25096), .C(matrixInput[244]), 
        .D(n25081), .Z(n27012) );
    VMW_AO22 U1310 ( .A(matrixInput[225]), .B(n25096), .C(matrixInput[217]), 
        .D(n25081), .Z(n27039) );
    VMW_AO22 U1491 ( .A(matrixInput[1907]), .B(n25096), .C(matrixInput[1899]), 
        .D(n25081), .Z(n25357) );
    VMW_AO22 U1501 ( .A(matrixInput[196]), .B(n25096), .C(matrixInput[188]), 
        .D(n25081), .Z(n27068) );
    VMW_AO22 U1973 ( .A(matrixInput[1472]), .B(n25096), .C(matrixInput[1464]), 
        .D(n25081), .Z(n25792) );
    VMW_AO22 U2320 ( .A(matrixInput[1159]), .B(n25096), .C(matrixInput[1151]), 
        .D(n25081), .Z(n26105) );
    VMW_AO22 U2531 ( .A(cOutput[115]), .B(n25087), .C(cOutput[99]), .D(n25084), 
        .Z(n25147) );
    VMW_FD \matrixInput_reg[1679]  ( .D(n25577), .CP(Clk), .Q(matrixInput
        [1679]) );
    VMW_FD \matrixInput_reg[1660]  ( .D(n25596), .CP(Clk), .Q(matrixInput
        [1660]) );
    VMW_FD \matrixInput_reg[1563]  ( .D(n25693), .CP(Clk), .Q(matrixInput
        [1563]) );
    VMW_FD \matrixInput_reg[374]  ( .D(n26882), .CP(Clk), .Q(matrixInput[374])
         );
    VMW_FD \matrixInput_reg[2007]  ( .D(n25249), .CP(Clk), .Q(matrixInput
        [2007]) );
    VMW_FD \matrixInput_reg[1653]  ( .D(n25603), .CP(Clk), .Q(matrixInput
        [1653]) );
    VMW_AO22 U1197 ( .A(matrixInput[327]), .B(n25096), .C(matrixInput[319]), 
        .D(n25081), .Z(n26937) );
    VMW_AO22 U1616 ( .A(matrixInput[1794]), .B(n25096), .C(matrixInput[1786]), 
        .D(n25081), .Z(n25470) );
    VMW_AO22 U1631 ( .A(matrixInput[1780]), .B(n25096), .C(matrixInput[1772]), 
        .D(n25081), .Z(n25484) );
    VMW_AO22 U2010 ( .A(matrixInput[1438]), .B(n25096), .C(matrixInput[1430]), 
        .D(n25081), .Z(n25826) );
    VMW_AO22 U2180 ( .A(matrixInput[1286]), .B(n25096), .C(matrixInput[1278]), 
        .D(n25081), .Z(n25978) );
    VMW_INV U2601 ( .A(\holder[5] ), .Z(n25071) );
    VMW_FD \matrixInput_reg[2034]  ( .D(n25222), .CP(Clk), .Q(matrixInput
        [2034]) );
    VMW_FD \matrixInput_reg[1550]  ( .D(n25706), .CP(Clk), .Q(matrixInput
        [1550]) );
    VMW_FD \matrixInput_reg[1549]  ( .D(n25707), .CP(Clk), .Q(matrixInput
        [1549]) );
    VMW_FD \matrixInput_reg[679]  ( .D(n26577), .CP(Clk), .Q(matrixInput[679])
         );
    VMW_FD \matrixInput_reg[347]  ( .D(n26909), .CP(Clk), .Q(matrixInput[347])
         );
    VMW_AO22 U1786 ( .A(matrixInput[1640]), .B(n25096), .C(matrixInput[1632]), 
        .D(n25081), .Z(n25624) );
    VMW_FD \matrixInput_reg[660]  ( .D(n26596), .CP(Clk), .Q(matrixInput[660])
         );
    VMW_AO22 U2037 ( .A(matrixInput[1414]), .B(n25096), .C(matrixInput[1406]), 
        .D(n25081), .Z(n25850) );
    VMW_FD \matrixInput_reg[1077]  ( .D(n26179), .CP(Clk), .Q(matrixInput
        [1077]) );
    VMW_FD \matrixInput_reg[563]  ( .D(n26693), .CP(Clk), .Q(matrixInput[563])
         );
    VMW_AO22 U455 ( .A(matrixInput[996]), .B(n25096), .C(matrixInput[988]), 
        .D(n25081), .Z(n26268) );
    VMW_AO22 U569 ( .A(matrixInput[893]), .B(n25096), .C(matrixInput[885]), 
        .D(n25081), .Z(n26371) );
    VMW_BUFIZ U2626 ( .A(n25199), .E(RD), .Z(\DataOut[29]1 ) );
    VMW_AO22 U659 ( .A(matrixInput[811]), .B(n25096), .C(matrixInput[803]), 
        .D(n25081), .Z(n26453) );
    VMW_AO22 U1337 ( .A(matrixInput[2044]), .B(n25096), .C(matrixInput[2036]), 
        .D(n25081), .Z(n25220) );
    VMW_AO22 U1526 ( .A(matrixInput[1875]), .B(n25096), .C(matrixInput[1867]), 
        .D(n25081), .Z(n25389) );
    VMW_FD \matrixInput_reg[1374]  ( .D(n25882), .CP(Clk), .Q(matrixInput
        [1374]) );
    VMW_FD \matrixInput_reg[1044]  ( .D(n26212), .CP(Clk), .Q(matrixInput
        [1044]) );
    VMW_AO22 U1954 ( .A(matrixInput[1489]), .B(n25096), .C(matrixInput[1481]), 
        .D(n25081), .Z(n25775) );
    VMW_FD \matrixInput_reg[653]  ( .D(n26603), .CP(Clk), .Q(matrixInput[653])
         );
    VMW_AO22 U2297 ( .A(matrixInput[1180]), .B(n25096), .C(matrixInput[1172]), 
        .D(n25081), .Z(n26084) );
    VMW_AO22 U2307 ( .A(matrixInput[1171]), .B(n25096), .C(matrixInput[1163]), 
        .D(n25081), .Z(n26093) );
    VMW_FD \matrixInput_reg[1347]  ( .D(n25909), .CP(Clk), .Q(matrixInput
        [1347]) );
    VMW_AO22 U2486 ( .A(matrixInput[1009]), .B(n25096), .C(matrixInput[1001]), 
        .D(n25081), .Z(n26255) );
    VMW_FD \matrixInput_reg[550]  ( .D(n26706), .CP(Clk), .Q(matrixInput[550])
         );
    VMW_AO22 U2516 ( .A(cOutput[20]), .B(n25087), .C(cOutput[4]), .D(n25084), 
        .Z(n25130) );
    VMW_FD \matrixInput_reg[549]  ( .D(n26707), .CP(Clk), .Q(matrixInput[549])
         );
    VMW_AO22 U765 ( .A(matrixInput[716]), .B(n25096), .C(matrixInput[708]), 
        .D(n25081), .Z(n26548) );
    VMW_AO22 U827 ( .A(matrixInput[660]), .B(n25096), .C(matrixInput[652]), 
        .D(n25081), .Z(n26604) );
    VMW_AO22 U1868 ( .A(matrixInput[1567]), .B(n25096), .C(matrixInput[1559]), 
        .D(n25081), .Z(n25697) );
    VMW_FD \matrixInput_reg[924]  ( .D(n26332), .CP(Clk), .Q(matrixInput[924])
         );
    VMW_FD \matrixInput_reg[917]  ( .D(n26339), .CP(Clk), .Q(matrixInput[917])
         );
    VMW_FD \vectorInput_reg[44]  ( .D(n27340), .CP(Clk), .Q(vectorInput[44])
         );
    VMW_AO22 U469 ( .A(matrixInput[983]), .B(n25096), .C(matrixInput[975]), 
        .D(n25081), .Z(n26281) );
    VMW_AO22 U472 ( .A(matrixInput[980]), .B(n25096), .C(matrixInput[972]), 
        .D(n25081), .Z(n26284) );
    VMW_AO22 U800 ( .A(matrixInput[685]), .B(n25096), .C(matrixInput[677]), 
        .D(n25081), .Z(n26579) );
    VMW_FD \matrixInput_reg[1887]  ( .D(n25369), .CP(Clk), .Q(matrixInput
        [1887]) );
    VMW_FD \vectorInput_reg[77]  ( .D(n27307), .CP(Clk), .Q(vectorInput[77])
         );
    VMW_AO22 U990 ( .A(matrixInput[513]), .B(n25096), .C(matrixInput[505]), 
        .D(n25081), .Z(n26751) );
    VMW_AO22 U742 ( .A(matrixInput[737]), .B(n25096), .C(matrixInput[729]), 
        .D(n25081), .Z(n26527) );
    VMW_FD \matrixInput_reg[1924]  ( .D(n25332), .CP(Clk), .Q(matrixInput
        [1924]) );
    VMW_FD \matrixInput_reg[1917]  ( .D(n25339), .CP(Clk), .Q(matrixInput
        [1917]) );
    VMW_FD \matrixInput_reg[7]  ( .D(n27249), .CP(Clk), .Q(matrixInput[7]) );
    VMW_AO22 U759 ( .A(matrixInput[721]), .B(n25096), .C(matrixInput[713]), 
        .D(n25081), .Z(n26543) );
    VMW_AO22 U1237 ( .A(matrixInput[291]), .B(n25096), .C(matrixInput[283]), 
        .D(n25081), .Z(n26973) );
    VMW_FD \matrixInput_reg[887]  ( .D(n26369), .CP(Clk), .Q(matrixInput[887])
         );
    VMW_AO22 U1426 ( .A(matrixInput[1965]), .B(n25096), .C(matrixInput[1957]), 
        .D(n25081), .Z(n25299) );
    VMW_FD \matrixInput_reg[643]  ( .D(n26613), .CP(Clk), .Q(matrixInput[643])
         );
    VMW_AO22 U1854 ( .A(matrixInput[1579]), .B(n25096), .C(matrixInput[1571]), 
        .D(n25081), .Z(n25685) );
    VMW_FD \matrixInput_reg[1054]  ( .D(n26202), .CP(Clk), .Q(matrixInput
        [1054]) );
    VMW_AO22 U2397 ( .A(matrixInput[1090]), .B(n25096), .C(matrixInput[1082]), 
        .D(n25081), .Z(n26174) );
    VMW_AO22 U2416 ( .A(matrixInput[1073]), .B(n25096), .C(matrixInput[1065]), 
        .D(n25081), .Z(n26191) );
    VMW_AO22 U1097 ( .A(matrixInput[417]), .B(n25096), .C(matrixInput[409]), 
        .D(n25081), .Z(n26847) );
    VMW_AO22 U1107 ( .A(matrixInput[11]), .B(n25096), .C(matrixInput[3]), .D(
        n25081), .Z(n27253) );
    VMW_AO22 U1686 ( .A(matrixInput[1730]), .B(n25096), .C(matrixInput[1722]), 
        .D(n25081), .Z(n25534) );
    VMW_AO22 U2207 ( .A(matrixInput[1261]), .B(n25096), .C(matrixInput[1253]), 
        .D(n25081), .Z(n26003) );
    VMW_FD \matrixInput_reg[559]  ( .D(n26697), .CP(Clk), .Q(matrixInput[559])
         );
    VMW_OAI21 U2586 ( .A(n25158), .B(n25159), .C(n25094), .Z(n25063) );
    VMW_FD \matrixInput_reg[1357]  ( .D(n25899), .CP(Clk), .Q(matrixInput
        [1357]) );
    VMW_FD \matrixInput_reg[540]  ( .D(n26716), .CP(Clk), .Q(matrixInput[540])
         );
    VMW_FD \matrixInput_reg[1067]  ( .D(n26189), .CP(Clk), .Q(matrixInput
        [1067]) );
    VMW_FD \matrixInput_reg[670]  ( .D(n26586), .CP(Clk), .Q(matrixInput[670])
         );
    VMW_AO22 U1716 ( .A(matrixInput[1704]), .B(n25096), .C(matrixInput[1696]), 
        .D(n25081), .Z(n25560) );
    VMW_FD \matrixInput_reg[669]  ( .D(n26587), .CP(Clk), .Q(matrixInput[669])
         );
    VMW_FD \matrixInput_reg[1364]  ( .D(n25892), .CP(Clk), .Q(matrixInput
        [1364]) );
    VMW_AO22 U2137 ( .A(matrixInput[1324]), .B(n25096), .C(matrixInput[1316]), 
        .D(n25081), .Z(n25940) );
    VMW_FD \matrixInput_reg[573]  ( .D(n26683), .CP(Clk), .Q(matrixInput[573])
         );
    VMW_PULLDOWN U281 ( .Z(n25199) );
    VMW_NOR2 U311 ( .A(n25092), .B(Addr[2]), .Z(n25093) );
    VMW_AO22 U336 ( .A(vectorInput[87]), .B(n25095), .C(vectorInput[79]), .D(
        n25080), .Z(n27305) );
    VMW_AO22 U343 ( .A(vectorInput[80]), .B(n25095), .C(vectorInput[72]), .D(
        n25080), .Z(n27312) );
    VMW_AO22 U344 ( .A(vectorInput[79]), .B(n25095), .C(vectorInput[71]), .D(
        n25080), .Z(n27313) );
    VMW_AO22 U363 ( .A(vectorInput[62]), .B(n25095), .C(vectorInput[54]), .D(
        n25080), .Z(n27330) );
    VMW_AO22 U642 ( .A(matrixInput[827]), .B(n25096), .C(matrixInput[819]), 
        .D(n25081), .Z(n26437) );
    VMW_AO22 U1120 ( .A(matrixInput[397]), .B(n25096), .C(matrixInput[389]), 
        .D(n25081), .Z(n26867) );
    VMW_AO22 U1731 ( .A(matrixInput[1690]), .B(n25096), .C(matrixInput[1682]), 
        .D(n25081), .Z(n25574) );
    VMW_FD \matrixInput_reg[1643]  ( .D(n25613), .CP(Clk), .Q(matrixInput
        [1643]) );
    VMW_AO22 U1210 ( .A(matrixInput[315]), .B(n25096), .C(matrixInput[307]), 
        .D(n25081), .Z(n26949) );
    VMW_AO22 U1380 ( .A(matrixInput[2007]), .B(n25096), .C(matrixInput[1999]), 
        .D(n25081), .Z(n25257) );
    VMW_AO22 U2080 ( .A(matrixInput[1376]), .B(n25096), .C(matrixInput[1368]), 
        .D(n25081), .Z(n25888) );
    VMW_AO22 U2110 ( .A(matrixInput[1348]), .B(n25096), .C(matrixInput[1340]), 
        .D(n25081), .Z(n25916) );
    VMW_FD \matrixInput_reg[2024]  ( .D(n25232), .CP(Clk), .Q(matrixInput
        [2024]) );
    VMW_FD \matrixInput_reg[1559]  ( .D(n25697), .CP(Clk), .Q(matrixInput
        [1559]) );
    VMW_FD \matrixInput_reg[357]  ( .D(n26899), .CP(Clk), .Q(matrixInput[357])
         );
    VMW_FD \matrixInput_reg[1540]  ( .D(n25716), .CP(Clk), .Q(matrixInput
        [1540]) );
    VMW_AO22 U1401 ( .A(matrixInput[205]), .B(n25096), .C(matrixInput[197]), 
        .D(n25081), .Z(n27059) );
    VMW_AO22 U1591 ( .A(matrixInput[1816]), .B(n25096), .C(matrixInput[1808]), 
        .D(n25081), .Z(n25448) );
    VMW_AO22 U1873 ( .A(matrixInput[1562]), .B(n25096), .C(matrixInput[1554]), 
        .D(n25081), .Z(n25702) );
    VMW_FD \matrixInput_reg[1670]  ( .D(n25586), .CP(Clk), .Q(matrixInput
        [1670]) );
    VMW_FD \matrixInput_reg[1669]  ( .D(n25587), .CP(Clk), .Q(matrixInput
        [1669]) );
    VMW_AO22 U2220 ( .A(matrixInput[1249]), .B(n25096), .C(matrixInput[1241]), 
        .D(n25081), .Z(n26015) );
    VMW_FD \matrixInput_reg[2017]  ( .D(n25239), .CP(Clk), .Q(matrixInput
        [2017]) );
    VMW_FD \matrixInput_reg[1573]  ( .D(n25683), .CP(Clk), .Q(matrixInput
        [1573]) );
    VMW_FD \matrixInput_reg[364]  ( .D(n26892), .CP(Clk), .Q(matrixInput[364])
         );
    VMW_AO22 U2431 ( .A(matrixInput[1059]), .B(n25096), .C(matrixInput[1051]), 
        .D(n25081), .Z(n26205) );
    VMW_AO22 U890 ( .A(matrixInput[604]), .B(n25096), .C(matrixInput[596]), 
        .D(n25081), .Z(n26660) );
    VMW_FD \matrixInput_reg[1907]  ( .D(n25349), .CP(Clk), .Q(matrixInput
        [1907]) );
    VMW_FD \matrixInput_reg[897]  ( .D(n26359), .CP(Clk), .Q(matrixInput[897])
         );
    VMW_AO22 U900 ( .A(matrixInput[595]), .B(n25096), .C(matrixInput[587]), 
        .D(n25081), .Z(n26669) );
    VMW_FD \matrixInput_reg[1934]  ( .D(n25322), .CP(Clk), .Q(matrixInput
        [1934]) );
    VMW_AO22 U555 ( .A(matrixInput[906]), .B(n25096), .C(matrixInput[898]), 
        .D(n25081), .Z(n26358) );
    VMW_AO22 U572 ( .A(matrixInput[890]), .B(n25096), .C(matrixInput[882]), 
        .D(n25081), .Z(n26374) );
    VMW_AO22 U927 ( .A(matrixInput[570]), .B(n25096), .C(matrixInput[562]), 
        .D(n25081), .Z(n26694) );
    VMW_FD \matrixInput_reg[907]  ( .D(n26349), .CP(Clk), .Q(matrixInput[907])
         );
    VMW_AO22 U381 ( .A(vectorInput[46]), .B(n25095), .C(vectorInput[38]), .D(
        n25080), .Z(n27346) );
    VMW_AO22 U386 ( .A(vectorInput[41]), .B(n25095), .C(vectorInput[33]), .D(
        n25080), .Z(n27351) );
    VMW_AO22 U407 ( .A(vectorInput[22]), .B(n25095), .C(vectorInput[14]), .D(
        n25080), .Z(n27370) );
    VMW_AO22 U420 ( .A(vectorInput[126]), .B(n25095), .C(vectorInput[118]), 
        .D(n25080), .Z(n27266) );
    VMW_AO22 U665 ( .A(matrixInput[807]), .B(n25096), .C(matrixInput[799]), 
        .D(n25081), .Z(n26457) );
    VMW_FD \matrixInput_reg[1897]  ( .D(n25359), .CP(Clk), .Q(matrixInput
        [1897]) );
    VMW_FD \vectorInput_reg[67]  ( .D(n27317), .CP(Clk), .Q(vectorInput[67])
         );
    VMW_AO22 U852 ( .A(matrixInput[70]), .B(n25096), .C(matrixInput[62]), .D(
        n25081), .Z(n27194) );
    VMW_AO22 U949 ( .A(matrixInput[550]), .B(n25096), .C(matrixInput[542]), 
        .D(n25081), .Z(n26714) );
    VMW_AO22 U1968 ( .A(matrixInput[1477]), .B(n25096), .C(matrixInput[1469]), 
        .D(n25081), .Z(n25787) );
    VMW_FD \matrixInput_reg[934]  ( .D(n26322), .CP(Clk), .Q(matrixInput[934])
         );
    VMW_FD \vectorInput_reg[54]  ( .D(n27330), .CP(Clk), .Q(vectorInput[54])
         );
    VMW_AO22 U2065 ( .A(matrixInput[1389]), .B(n25096), .C(matrixInput[1381]), 
        .D(n25081), .Z(n25875) );
    VMW_FD \matrixInput_reg[1732]  ( .D(n25524), .CP(Clk), .Q(matrixInput
        [1732]) );
    VMW_FD \matrixInput_reg[125]  ( .D(n27131), .CP(Clk), .Q(matrixInput[125])
         );
    VMW_AO22 U1055 ( .A(matrixInput[455]), .B(n25096), .C(matrixInput[447]), 
        .D(n25081), .Z(n26809) );
    VMW_AO22 U1644 ( .A(matrixInput[1768]), .B(n25096), .C(matrixInput[1760]), 
        .D(n25081), .Z(n25496) );
    VMW_FD \matrixInput_reg[1431]  ( .D(n25825), .CP(Clk), .Q(matrixInput
        [1431]) );
    VMW_FD \matrixInput_reg[1428]  ( .D(n25828), .CP(Clk), .Q(matrixInput
        [1428]) );
    VMW_AO22 U1072 ( .A(matrixInput[439]), .B(n25096), .C(matrixInput[431]), 
        .D(n25081), .Z(n26825) );
    VMW_AO22 U1342 ( .A(matrixInput[2039]), .B(n25096), .C(matrixInput[2031]), 
        .D(n25081), .Z(n25225) );
    VMW_AO22 U1365 ( .A(matrixInput[2018]), .B(n25096), .C(matrixInput[2010]), 
        .D(n25081), .Z(n25246) );
    VMW_AO22 U1574 ( .A(matrixInput[1831]), .B(n25096), .C(matrixInput[1823]), 
        .D(n25081), .Z(n25433) );
    VMW_AO22 U2355 ( .A(matrixInput[119]), .B(n25096), .C(matrixInput[111]), 
        .D(n25081), .Z(n27145) );
    VMW_FD \matrixInput_reg[1385]  ( .D(n25871), .CP(Clk), .Q(matrixInput
        [1385]) );
    VMW_FD \matrixInput_reg[226]  ( .D(n27030), .CP(Clk), .Q(matrixInput[226])
         );
    VMW_FD \matrixInput_reg[592]  ( .D(n26664), .CP(Clk), .Q(matrixInput[592])
         );
    VMW_FD \matrixInput_reg[116]  ( .D(n27140), .CP(Clk), .Q(matrixInput[116])
         );
    VMW_AO22 U2544 ( .A(cOutput[25]), .B(n25089), .C(cOutput[9]), .D(n25088), 
        .Z(n25164) );
    VMW_FD \matrixInput_reg[1718]  ( .D(n25538), .CP(Clk), .Q(matrixInput
        [1718]) );
    VMW_FD \matrixInput_reg[1701]  ( .D(n25555), .CP(Clk), .Q(matrixInput
        [1701]) );
    VMW_FD \matrixInput_reg[215]  ( .D(n27041), .CP(Clk), .Q(matrixInput[215])
         );
    VMW_FD \matrixInput_reg[1402]  ( .D(n25854), .CP(Clk), .Q(matrixInput
        [1402]) );
    VMW_AO22 U1896 ( .A(matrixInput[1541]), .B(n25096), .C(matrixInput[1533]), 
        .D(n25081), .Z(n25723) );
    VMW_AO22 U1906 ( .A(matrixInput[1532]), .B(n25096), .C(matrixInput[1524]), 
        .D(n25081), .Z(n25732) );
    VMW_FD \matrixInput_reg[1086]  ( .D(n26170), .CP(Clk), .Q(matrixInput
        [1086]) );
    VMW_FD \matrixInput_reg[688]  ( .D(n26568), .CP(Clk), .Q(matrixInput[688])
         );
    VMW_FD \matrixInput_reg[691]  ( .D(n26565), .CP(Clk), .Q(matrixInput[691])
         );
    VMW_AO22 U2372 ( .A(matrixInput[1112]), .B(n25096), .C(matrixInput[1104]), 
        .D(n25081), .Z(n26152) );
    VMW_OAI21 U2563 ( .A(n25097), .B(n25098), .C(n25090), .Z(n25106) );
    VMW_FD \matrixInput_reg[1125]  ( .D(n26131), .CP(Clk), .Q(matrixInput
        [1125]) );
    VMW_FD \matrixInput_reg[732]  ( .D(n26524), .CP(Clk), .Q(matrixInput[732])
         );
    VMW_FD \vectorInput_reg[8]  ( .D(n27376), .CP(Clk), .Q(vectorInput[8]) );
    VMW_AO22 U1553 ( .A(matrixInput[1850]), .B(n25096), .C(matrixInput[1842]), 
        .D(n25081), .Z(n25414) );
    VMW_AO22 U1921 ( .A(matrixInput[1518]), .B(n25096), .C(matrixInput[1510]), 
        .D(n25081), .Z(n25746) );
    VMW_FD \matrixInput_reg[1226]  ( .D(n26030), .CP(Clk), .Q(matrixInput
        [1226]) );
    VMW_AO22 U2042 ( .A(matrixInput[1409]), .B(n25096), .C(matrixInput[1401]), 
        .D(n25081), .Z(n25855) );
    VMW_FD \matrixInput_reg[1592]  ( .D(n25664), .CP(Clk), .Q(matrixInput
        [1592]) );
    VMW_FD \matrixInput_reg[431]  ( .D(n26825), .CP(Clk), .Q(matrixInput[431])
         );
    VMW_FD \matrixInput_reg[428]  ( .D(n26828), .CP(Clk), .Q(matrixInput[428])
         );
    VMW_FD \matrixInput_reg[385]  ( .D(n26871), .CP(Clk), .Q(matrixInput[385])
         );
    VMW_FD \matrixInput_reg[1691]  ( .D(n25565), .CP(Clk), .Q(matrixInput
        [1691]) );
    VMW_FD \matrixInput_reg[1688]  ( .D(n25568), .CP(Clk), .Q(matrixInput
        [1688]) );
    VMW_FD \matrixInput_reg[1215]  ( .D(n26041), .CP(Clk), .Q(matrixInput
        [1215]) );
    VMW_FD \matrixInput_reg[1116]  ( .D(n26140), .CP(Clk), .Q(matrixInput
        [1116]) );
    VMW_FD \matrixInput_reg[718]  ( .D(n26538), .CP(Clk), .Q(matrixInput[718])
         );
    VMW_FD \matrixInput_reg[701]  ( .D(n26555), .CP(Clk), .Q(matrixInput[701])
         );
    VMW_FD \matrixInput_reg[402]  ( .D(n26854), .CP(Clk), .Q(matrixInput[402])
         );
    VMW_AO22 U1663 ( .A(matrixInput[1751]), .B(n25096), .C(matrixInput[1743]), 
        .D(n25081), .Z(n25513) );
    VMW_FD \matrixInput_reg[876]  ( .D(n26380), .CP(Clk), .Q(matrixInput[876])
         );
    VMW_FD \matrixInput_reg[36]  ( .D(n27220), .CP(Clk), .Q(matrixInput[36])
         );
    VMW_AO22 U597 ( .A(matrixInput[93]), .B(n25096), .C(matrixInput[85]), .D(
        n25081), .Z(n27171) );
    VMW_AO22 U680 ( .A(matrixInput[793]), .B(n25096), .C(matrixInput[785]), 
        .D(n25081), .Z(n26471) );
    VMW_AO22 U710 ( .A(matrixInput[766]), .B(n25096), .C(matrixInput[758]), 
        .D(n25081), .Z(n26498) );
    VMW_FD \matrixInput_reg[845]  ( .D(n26411), .CP(Clk), .Q(matrixInput[845])
         );
    VMW_AO22 U737 ( .A(matrixInput[741]), .B(n25096), .C(matrixInput[733]), 
        .D(n25081), .Z(n26523) );
    VMW_AO22 U1259 ( .A(matrixInput[271]), .B(n25096), .C(matrixInput[263]), 
        .D(n25081), .Z(n26993) );
    VMW_AO22 U1448 ( .A(matrixInput[1945]), .B(n25096), .C(matrixInput[1937]), 
        .D(n25081), .Z(n25319) );
    VMW_FD \matrixInput_reg[1876]  ( .D(n25380), .CP(Clk), .Q(matrixInput
        [1876]) );
    VMW_AO22 U2269 ( .A(matrixInput[1206]), .B(n25096), .C(matrixInput[1198]), 
        .D(n25081), .Z(n26058) );
    VMW_FD \vectorInput_reg[86]  ( .D(n27298), .CP(Clk), .Q(vectorInput[86])
         );
    VMW_AO22 U2478 ( .A(matrixInput[1017]), .B(n25096), .C(matrixInput[1009]), 
        .D(n25081), .Z(n26247) );
    VMW_AO22 U875 ( .A(matrixInput[617]), .B(n25096), .C(matrixInput[609]), 
        .D(n25081), .Z(n26647) );
    VMW_AO22 U1169 ( .A(matrixInput[352]), .B(n25096), .C(matrixInput[344]), 
        .D(n25081), .Z(n26912) );
    VMW_AO22 U1778 ( .A(matrixInput[171]), .B(n25096), .C(matrixInput[163]), 
        .D(n25081), .Z(n27093) );
    VMW_FD \matrixInput_reg[1845]  ( .D(n25411), .CP(Clk), .Q(matrixInput
        [1845]) );
    VMW_FD \vectorInput_reg[105]  ( .D(n27279), .CP(Clk), .Q(vectorInput[105])
         );
    VMW_AO22 U2159 ( .A(matrixInput[1305]), .B(n25096), .C(matrixInput[1297]), 
        .D(n25081), .Z(n25959) );
    VMW_AO22 U969 ( .A(matrixInput[532]), .B(n25096), .C(matrixInput[524]), 
        .D(n25081), .Z(n26732) );
    VMW_AO22 U1075 ( .A(matrixInput[437]), .B(n25096), .C(matrixInput[429]), 
        .D(n25081), .Z(n26827) );
    VMW_AO22 U1664 ( .A(matrixInput[1750]), .B(n25096), .C(matrixInput[1742]), 
        .D(n25081), .Z(n25514) );
    VMW_FD \matrixInput_reg[224]  ( .D(n27032), .CP(Clk), .Q(matrixInput[224])
         );
    VMW_FD \matrixInput_reg[1433]  ( .D(n25823), .CP(Clk), .Q(matrixInput
        [1433]) );
    VMW_AO22 U1052 ( .A(matrixInput[52]), .B(n25096), .C(matrixInput[44]), .D(
        n25081), .Z(n27212) );
    VMW_AO22 U1345 ( .A(matrixInput[2037]), .B(n25096), .C(matrixInput[2029]), 
        .D(n25081), .Z(n25227) );
    VMW_AO22 U1554 ( .A(matrixInput[1849]), .B(n25096), .C(matrixInput[1841]), 
        .D(n25081), .Z(n25415) );
    VMW_AO22 U1926 ( .A(matrixInput[1514]), .B(n25096), .C(matrixInput[1506]), 
        .D(n25081), .Z(n25750) );
    VMW_AO22 U2045 ( .A(matrixInput[147]), .B(n25096), .C(matrixInput[139]), 
        .D(n25081), .Z(n27117) );
    VMW_FD \matrixInput_reg[127]  ( .D(n27129), .CP(Clk), .Q(matrixInput[127])
         );
    VMW_FD \matrixInput_reg[1730]  ( .D(n25526), .CP(Clk), .Q(matrixInput
        [1730]) );
    VMW_FD \matrixInput_reg[1729]  ( .D(n25527), .CP(Clk), .Q(matrixInput
        [1729]) );
    VMW_FD \matrixInput_reg[1084]  ( .D(n26172), .CP(Clk), .Q(matrixInput
        [1084]) );
    VMW_FD \matrixInput_reg[693]  ( .D(n26563), .CP(Clk), .Q(matrixInput[693])
         );
    VMW_FD \matrixInput_reg[1419]  ( .D(n25837), .CP(Clk), .Q(matrixInput
        [1419]) );
    VMW_FD \matrixInput_reg[1400]  ( .D(n25856), .CP(Clk), .Q(matrixInput
        [1400]) );
    VMW_AO22 U1362 ( .A(matrixInput[2021]), .B(n25096), .C(matrixInput[2013]), 
        .D(n25081), .Z(n25243) );
    VMW_AO22 U1891 ( .A(matrixInput[1546]), .B(n25096), .C(matrixInput[1538]), 
        .D(n25081), .Z(n25718) );
    VMW_AO22 U2375 ( .A(matrixInput[1109]), .B(n25096), .C(matrixInput[1101]), 
        .D(n25081), .Z(n26155) );
    VMW_FD \matrixInput_reg[217]  ( .D(n27039), .CP(Clk), .Q(matrixInput[217])
         );
    VMW_OAI21 U2564 ( .A(n25099), .B(n25100), .C(n25091), .Z(n25105) );
    VMW_FD \matrixInput_reg[1703]  ( .D(n25553), .CP(Clk), .Q(matrixInput
        [1703]) );
    VMW_FD \matrixInput_reg[1387]  ( .D(n25869), .CP(Clk), .Q(matrixInput
        [1387]) );
    VMW_FD \matrixInput_reg[590]  ( .D(n26666), .CP(Clk), .Q(matrixInput[590])
         );
    VMW_FD \matrixInput_reg[114]  ( .D(n27142), .CP(Clk), .Q(matrixInput[114])
         );
    VMW_FD \matrixInput_reg[589]  ( .D(n26667), .CP(Clk), .Q(matrixInput[589])
         );
    VMW_FD \matrixInput_reg[433]  ( .D(n26823), .CP(Clk), .Q(matrixInput[433])
         );
    VMW_AO22 U1901 ( .A(matrixInput[1537]), .B(n25096), .C(matrixInput[1529]), 
        .D(n25081), .Z(n25727) );
    VMW_FD \matrixInput_reg[1224]  ( .D(n26032), .CP(Clk), .Q(matrixInput
        [1224]) );
    VMW_AO22 U1573 ( .A(matrixInput[1832]), .B(n25096), .C(matrixInput[1824]), 
        .D(n25081), .Z(n25432) );
    VMW_AO22 U2352 ( .A(matrixInput[1130]), .B(n25096), .C(matrixInput[1122]), 
        .D(n25081), .Z(n26134) );
    VMW_AO22 U2543 ( .A(cOutput[17]), .B(n25087), .C(cOutput[1]), .D(n25084), 
        .Z(n25163) );
    VMW_FD \matrixInput_reg[1127]  ( .D(n26129), .CP(Clk), .Q(matrixInput
        [1127]) );
    VMW_FD \matrixInput_reg[730]  ( .D(n26526), .CP(Clk), .Q(matrixInput[730])
         );
    VMW_FD \matrixInput_reg[729]  ( .D(n26527), .CP(Clk), .Q(matrixInput[729])
         );
    VMW_AO22 U1643 ( .A(matrixInput[1769]), .B(n25096), .C(matrixInput[1761]), 
        .D(n25081), .Z(n25495) );
    VMW_AO22 U2062 ( .A(matrixInput[1392]), .B(n25096), .C(matrixInput[1384]), 
        .D(n25081), .Z(n25872) );
    VMW_FD \matrixInput_reg[1693]  ( .D(n25563), .CP(Clk), .Q(matrixInput
        [1693]) );
    VMW_FD \matrixInput_reg[1217]  ( .D(n26039), .CP(Clk), .Q(matrixInput
        [1217]) );
    VMW_FD \matrixInput_reg[1114]  ( .D(n26142), .CP(Clk), .Q(matrixInput
        [1114]) );
    VMW_FD \matrixInput_reg[419]  ( .D(n26837), .CP(Clk), .Q(matrixInput[419])
         );
    VMW_FD \matrixInput_reg[400]  ( .D(n26856), .CP(Clk), .Q(matrixInput[400])
         );
    VMW_FD \matrixInput_reg[703]  ( .D(n26553), .CP(Clk), .Q(matrixInput[703])
         );
    VMW_FD \matrixInput_reg[387]  ( .D(n26869), .CP(Clk), .Q(matrixInput[387])
         );
    VMW_FD \matrixInput_reg[1590]  ( .D(n25666), .CP(Clk), .Q(matrixInput
        [1590]) );
    VMW_FD \matrixInput_reg[1589]  ( .D(n25667), .CP(Clk), .Q(matrixInput
        [1589]) );
    VMW_AO22 U400 ( .A(vectorInput[28]), .B(n25095), .C(vectorInput[20]), .D(
        n25080), .Z(n27364) );
    VMW_AO22 U427 ( .A(vectorInput[119]), .B(n25095), .C(vectorInput[111]), 
        .D(n25080), .Z(n27273) );
    VMW_AO22 U590 ( .A(matrixInput[874]), .B(n25096), .C(matrixInput[866]), 
        .D(n25081), .Z(n26390) );
    VMW_AO22 U687 ( .A(matrixInput[787]), .B(n25096), .C(matrixInput[779]), 
        .D(n25081), .Z(n26477) );
    VMW_AO22 U730 ( .A(matrixInput[81]), .B(n25096), .C(matrixInput[73]), .D(
        n25081), .Z(n27183) );
    VMW_AO22 U872 ( .A(matrixInput[619]), .B(n25096), .C(matrixInput[611]), 
        .D(n25081), .Z(n26645) );
    VMW_FD \matrixInput_reg[34]  ( .D(n27222), .CP(Clk), .Q(matrixInput[34])
         );
    VMW_FD \matrixInput_reg[874]  ( .D(n26382), .CP(Clk), .Q(matrixInput[874])
         );
    VMW_FD \matrixInput_reg[847]  ( .D(n26409), .CP(Clk), .Q(matrixInput[847])
         );
    VMW_AO22 U717 ( .A(matrixInput[759]), .B(n25096), .C(matrixInput[751]), 
        .D(n25081), .Z(n26505) );
    VMW_AO22 U2249 ( .A(matrixInput[1223]), .B(n25096), .C(matrixInput[1215]), 
        .D(n25081), .Z(n26041) );
    VMW_AO22 U2458 ( .A(matrixInput[1035]), .B(n25096), .C(matrixInput[1027]), 
        .D(n25081), .Z(n26229) );
    VMW_AO22 U1279 ( .A(matrixInput[253]), .B(n25096), .C(matrixInput[245]), 
        .D(n25081), .Z(n27011) );
    VMW_AO22 U1468 ( .A(matrixInput[1927]), .B(n25096), .C(matrixInput[1919]), 
        .D(n25081), .Z(n25337) );
    VMW_FD \vectorInput_reg[84]  ( .D(n27300), .CP(Clk), .Q(vectorInput[84])
         );
    VMW_AO22 U2179 ( .A(matrixInput[1287]), .B(n25096), .C(matrixInput[1279]), 
        .D(n25081), .Z(n25977) );
    VMW_FD \matrixInput_reg[1874]  ( .D(n25382), .CP(Clk), .Q(matrixInput
        [1874]) );
    VMW_FD \vectorInput_reg[107]  ( .D(n27277), .CP(Clk), .Q(vectorInput[107])
         );
    VMW_AO22 U449 ( .A(matrixInput[1001]), .B(n25096), .C(matrixInput[993]), 
        .D(n25081), .Z(n26263) );
    VMW_AO22 U779 ( .A(matrixInput[704]), .B(n25096), .C(matrixInput[696]), 
        .D(n25081), .Z(n26560) );
    VMW_AO22 U855 ( .A(matrixInput[635]), .B(n25096), .C(matrixInput[627]), 
        .D(n25081), .Z(n26629) );
    VMW_AO22 U1149 ( .A(matrixInput[370]), .B(n25096), .C(matrixInput[362]), 
        .D(n25081), .Z(n26894) );
    VMW_AO22 U1758 ( .A(matrixInput[1666]), .B(n25096), .C(matrixInput[1658]), 
        .D(n25081), .Z(n25598) );
    VMW_FD \matrixInput_reg[1847]  ( .D(n25409), .CP(Clk), .Q(matrixInput
        [1847]) );
    VMW_AO22 U2436 ( .A(matrixInput[1055]), .B(n25096), .C(matrixInput[1047]), 
        .D(n25081), .Z(n26209) );
    VMW_FD \matrixInput_reg[1355]  ( .D(n25901), .CP(Clk), .Q(matrixInput
        [1355]) );
    VMW_AO22 U1217 ( .A(matrixInput[308]), .B(n25096), .C(matrixInput[300]), 
        .D(n25081), .Z(n26956) );
    VMW_AO22 U1596 ( .A(matrixInput[1811]), .B(n25096), .C(matrixInput[1803]), 
        .D(n25081), .Z(n25453) );
    VMW_AO22 U1874 ( .A(matrixInput[1561]), .B(n25096), .C(matrixInput[1553]), 
        .D(n25081), .Z(n25703) );
    VMW_AO22 U2227 ( .A(matrixInput[1243]), .B(n25096), .C(matrixInput[1235]), 
        .D(n25081), .Z(n26021) );
    VMW_FD \matrixInput_reg[542]  ( .D(n26714), .CP(Clk), .Q(matrixInput[542])
         );
    VMW_FD \matrixInput_reg[1056]  ( .D(n26200), .CP(Clk), .Q(matrixInput
        [1056]) );
    VMW_FD \matrixInput_reg[641]  ( .D(n26615), .CP(Clk), .Q(matrixInput[641])
         );
    VMW_AO22 U1387 ( .A(matrixInput[2000]), .B(n25096), .C(matrixInput[1992]), 
        .D(n25081), .Z(n25264) );
    VMW_AO22 U1406 ( .A(matrixInput[1983]), .B(n25096), .C(matrixInput[1975]), 
        .D(n25081), .Z(n25281) );
    VMW_FD \matrixInput_reg[658]  ( .D(n26598), .CP(Clk), .Q(matrixInput[658])
         );
    VMW_AO22 U2087 ( .A(matrixInput[1369]), .B(n25096), .C(matrixInput[1361]), 
        .D(n25081), .Z(n25895) );
    VMW_AO22 U662 ( .A(matrixInput[808]), .B(n25096), .C(matrixInput[800]), 
        .D(n25081), .Z(n26456) );
    VMW_AO22 U1090 ( .A(matrixInput[423]), .B(n25096), .C(matrixInput[415]), 
        .D(n25081), .Z(n26841) );
    VMW_AO22 U1127 ( .A(matrixInput[390]), .B(n25096), .C(matrixInput[382]), 
        .D(n25081), .Z(n26874) );
    VMW_AO22 U2117 ( .A(matrixInput[1342]), .B(n25096), .C(matrixInput[1334]), 
        .D(n25081), .Z(n25922) );
    VMW_FD \matrixInput_reg[568]  ( .D(n26688), .CP(Clk), .Q(matrixInput[568])
         );
    VMW_FD \matrixInput_reg[1366]  ( .D(n25890), .CP(Clk), .Q(matrixInput
        [1366]) );
    VMW_FD \matrixInput_reg[571]  ( .D(n26685), .CP(Clk), .Q(matrixInput[571])
         );
    VMW_AO22 U1736 ( .A(matrixInput[1686]), .B(n25096), .C(matrixInput[1678]), 
        .D(n25081), .Z(n25578) );
    VMW_FD \matrixInput_reg[672]  ( .D(n26584), .CP(Clk), .Q(matrixInput[672])
         );
    VMW_AO22 U2130 ( .A(matrixInput[1330]), .B(n25096), .C(matrixInput[1322]), 
        .D(n25081), .Z(n25934) );
    VMW_FD \matrixInput_reg[2026]  ( .D(n25230), .CP(Clk), .Q(matrixInput
        [2026]) );
    VMW_FD \matrixInput_reg[1542]  ( .D(n25714), .CP(Clk), .Q(matrixInput
        [1542]) );
    VMW_FD \matrixInput_reg[1065]  ( .D(n26191), .CP(Clk), .Q(matrixInput
        [1065]) );
    VMW_FD \matrixInput_reg[355]  ( .D(n26901), .CP(Clk), .Q(matrixInput[355])
         );
    VMW_AO22 U1100 ( .A(matrixInput[414]), .B(n25096), .C(matrixInput[406]), 
        .D(n25081), .Z(n26850) );
    VMW_AO22 U1711 ( .A(matrixInput[24]), .B(n25096), .C(matrixInput[16]), .D(
        n25081), .Z(n27240) );
    VMW_AO22 U1230 ( .A(matrixInput[36]), .B(n25096), .C(matrixInput[28]), .D(
        n25081), .Z(n27228) );
    VMW_AO22 U1421 ( .A(matrixInput[1969]), .B(n25096), .C(matrixInput[1961]), 
        .D(n25081), .Z(n25295) );
    VMW_AO22 U1681 ( .A(matrixInput[1735]), .B(n25096), .C(matrixInput[1727]), 
        .D(n25081), .Z(n25529) );
    VMW_AO22 U1853 ( .A(matrixInput[1580]), .B(n25096), .C(matrixInput[1572]), 
        .D(n25081), .Z(n25684) );
    VMW_AO22 U2200 ( .A(matrixInput[133]), .B(n25096), .C(matrixInput[125]), 
        .D(n25081), .Z(n27131) );
    VMW_OAI21 U2581 ( .A(n25145), .B(n25146), .C(n25093), .Z(n25151) );
    VMW_FD \matrixInput_reg[1658]  ( .D(n25598), .CP(Clk), .Q(matrixInput
        [1658]) );
    VMW_FD \matrixInput_reg[1641]  ( .D(n25615), .CP(Clk), .Q(matrixInput
        [1641]) );
    VMW_AO22 U2390 ( .A(matrixInput[1097]), .B(n25096), .C(matrixInput[1089]), 
        .D(n25081), .Z(n26167) );
    VMW_AO22 U2411 ( .A(matrixInput[114]), .B(n25096), .C(matrixInput[106]), 
        .D(n25081), .Z(n27150) );
    VMW_FD \matrixInput_reg[2015]  ( .D(n25241), .CP(Clk), .Q(matrixInput
        [2015]) );
    VMW_FD \matrixInput_reg[1571]  ( .D(n25685), .CP(Clk), .Q(matrixInput
        [1571]) );
    VMW_FD \matrixInput_reg[1568]  ( .D(n25688), .CP(Clk), .Q(matrixInput
        [1568]) );
    VMW_FD \matrixInput_reg[366]  ( .D(n26890), .CP(Clk), .Q(matrixInput[366])
         );
    VMW_FD \matrixInput_reg[1672]  ( .D(n25584), .CP(Clk), .Q(matrixInput
        [1672]) );
    VMW_FD \matrixInput_reg[1905]  ( .D(n25351), .CP(Clk), .Q(matrixInput
        [1905]) );
    VMW_FD \matrixInput_reg[895]  ( .D(n26361), .CP(Clk), .Q(matrixInput[895])
         );
    VMW_AO22 U358 ( .A(vectorInput[67]), .B(n25095), .C(vectorInput[59]), .D(
        n25080), .Z(n27325) );
    VMW_AO22 U364 ( .A(vectorInput[61]), .B(n25095), .C(vectorInput[53]), .D(
        n25080), .Z(n27331) );
    VMW_AO22 U552 ( .A(matrixInput[16]), .B(n25096), .C(matrixInput[8]), .D(
        n25081), .Z(n27248) );
    VMW_AO22 U575 ( .A(matrixInput[95]), .B(n25096), .C(matrixInput[87]), .D(
        n25081), .Z(n27169) );
    VMW_AO22 U920 ( .A(matrixInput[577]), .B(n25096), .C(matrixInput[569]), 
        .D(n25081), .Z(n26687) );
    VMW_FD \matrixInput_reg[1936]  ( .D(n25320), .CP(Clk), .Q(matrixInput
        [1936]) );
    VMW_FD \matrixInput_reg[1895]  ( .D(n25361), .CP(Clk), .Q(matrixInput
        [1895]) );
    VMW_FD \vectorInput_reg[65]  ( .D(n27319), .CP(Clk), .Q(vectorInput[65])
         );
    VMW_AO22 U645 ( .A(matrixInput[824]), .B(n25096), .C(matrixInput[816]), 
        .D(n25081), .Z(n26440) );
    VMW_AO22 U897 ( .A(matrixInput[66]), .B(n25096), .C(matrixInput[58]), .D(
        n25081), .Z(n27198) );
    VMW_AO22 U907 ( .A(matrixInput[588]), .B(n25096), .C(matrixInput[580]), 
        .D(n25081), .Z(n26676) );
    VMW_FD \matrixInput_reg[905]  ( .D(n26351), .CP(Clk), .Q(matrixInput[905])
         );
    VMW_AO22 U1948 ( .A(matrixInput[1495]), .B(n25096), .C(matrixInput[1487]), 
        .D(n25081), .Z(n25769) );
    VMW_FD \matrixInput_reg[936]  ( .D(n26320), .CP(Clk), .Q(matrixInput[936])
         );
    VMW_FD \vectorInput_reg[56]  ( .D(n27328), .CP(Clk), .Q(vectorInput[56])
         );
    VMW_AO22 U1000 ( .A(matrixInput[505]), .B(n25096), .C(matrixInput[497]), 
        .D(n25081), .Z(n26759) );
    VMW_AO22 U1330 ( .A(DataIn[2]), .B(n25096), .C(matrixInput[2042]), .D(
        n25081), .Z(n25214) );
    VMW_AO22 U1953 ( .A(matrixInput[1490]), .B(n25096), .C(matrixInput[1482]), 
        .D(n25081), .Z(n25774) );
    VMW_AO22 U2290 ( .A(matrixInput[1187]), .B(n25096), .C(matrixInput[1179]), 
        .D(n25081), .Z(n26077) );
    VMW_AO22 U2511 ( .A(cOutput[85]), .B(n25087), .C(cOutput[69]), .D(n25084), 
        .Z(n25123) );
    VMW_FD \matrixInput_reg[2005]  ( .D(n25251), .CP(Clk), .Q(matrixInput
        [2005]) );
    VMW_AO22 U2300 ( .A(matrixInput[124]), .B(n25096), .C(matrixInput[116]), 
        .D(n25081), .Z(n27140) );
    VMW_AO22 U2481 ( .A(matrixInput[1014]), .B(n25096), .C(matrixInput[1006]), 
        .D(n25081), .Z(n26250) );
    VMW_FD \matrixInput_reg[1662]  ( .D(n25594), .CP(Clk), .Q(matrixInput
        [1662]) );
    VMW_FD \matrixInput_reg[1578]  ( .D(n25678), .CP(Clk), .Q(matrixInput
        [1578]) );
    VMW_FD \matrixInput_reg[1561]  ( .D(n25695), .CP(Clk), .Q(matrixInput
        [1561]) );
    VMW_FD \matrixInput_reg[376]  ( .D(n26880), .CP(Clk), .Q(matrixInput[376])
         );
    VMW_AO22 U1521 ( .A(matrixInput[1879]), .B(n25096), .C(matrixInput[1871]), 
        .D(n25081), .Z(n25385) );
    VMW_AO22 U2030 ( .A(matrixInput[1420]), .B(n25096), .C(matrixInput[1412]), 
        .D(n25081), .Z(n25844) );
    VMW_BUFIZ U2621 ( .A(\holder[6] ), .E(RD), .Z(\DataOut[6]1 ) );
    VMW_FD \matrixInput_reg[1552]  ( .D(n25704), .CP(Clk), .Q(matrixInput
        [1552]) );
    VMW_FD \matrixInput_reg[345]  ( .D(n26911), .CP(Clk), .Q(matrixInput[345])
         );
    VMW_FD \matrixInput_reg[2036]  ( .D(n25220), .CP(Clk), .Q(matrixInput
        [2036]) );
    VMW_AO22 U1190 ( .A(matrixInput[333]), .B(n25096), .C(matrixInput[325]), 
        .D(n25081), .Z(n26931) );
    VMW_AO22 U1781 ( .A(matrixInput[1645]), .B(n25096), .C(matrixInput[1637]), 
        .D(n25081), .Z(n25619) );
    VMW_AO22 U1611 ( .A(matrixInput[1798]), .B(n25096), .C(matrixInput[1790]), 
        .D(n25081), .Z(n25466) );
    VMW_AO22 U2017 ( .A(matrixInput[1432]), .B(n25096), .C(matrixInput[1424]), 
        .D(n25081), .Z(n25832) );
    VMW_FD \matrixInput_reg[1651]  ( .D(n25605), .CP(Clk), .Q(matrixInput
        [1651]) );
    VMW_FD \matrixInput_reg[1648]  ( .D(n25608), .CP(Clk), .Q(matrixInput
        [1648]) );
    VMW_FD \matrixInput_reg[1376]  ( .D(n25880), .CP(Clk), .Q(matrixInput
        [1376]) );
    VMW_AO22 U452 ( .A(matrixInput[998]), .B(n25096), .C(matrixInput[990]), 
        .D(n25081), .Z(n26266) );
    VMW_AO22 U475 ( .A(matrixInput[104]), .B(n25096), .C(matrixInput[96]), .D(
        n25081), .Z(n27160) );
    VMW_AO22 U549 ( .A(matrixInput[910]), .B(n25096), .C(matrixInput[902]), 
        .D(n25081), .Z(n26354) );
    VMW_AO22 U2187 ( .A(matrixInput[1279]), .B(n25096), .C(matrixInput[1271]), 
        .D(n25081), .Z(n25985) );
    VMW_FD \matrixInput_reg[561]  ( .D(n26695), .CP(Clk), .Q(matrixInput[561])
         );
    VMW_INV U2606 ( .A(\holder[4] ), .Z(n25068) );
    VMW_FD \matrixInput_reg[578]  ( .D(n26678), .CP(Clk), .Q(matrixInput[578])
         );
    VMW_AO22 U679 ( .A(matrixInput[794]), .B(n25096), .C(matrixInput[786]), 
        .D(n25081), .Z(n26470) );
    VMW_AO22 U1027 ( .A(matrixInput[480]), .B(n25096), .C(matrixInput[472]), 
        .D(n25081), .Z(n26784) );
    VMW_AO22 U1636 ( .A(matrixInput[1776]), .B(n25096), .C(matrixInput[1768]), 
        .D(n25081), .Z(n25488) );
    VMW_FD \matrixInput_reg[1075]  ( .D(n26181), .CP(Clk), .Q(matrixInput
        [1075]) );
    VMW_AO22 U2327 ( .A(matrixInput[1153]), .B(n25096), .C(matrixInput[1145]), 
        .D(n25081), .Z(n26111) );
    VMW_FD \matrixInput_reg[662]  ( .D(n26594), .CP(Clk), .Q(matrixInput[662])
         );
    VMW_FD \matrixInput_reg[552]  ( .D(n26704), .CP(Clk), .Q(matrixInput[552])
         );
    VMW_AO22 U2536 ( .A(cOutput[50]), .B(n25087), .C(cOutput[34]), .D(n25084), 
        .Z(n25154) );
    VMW_AO22 U745 ( .A(matrixInput[734]), .B(n25096), .C(matrixInput[726]), 
        .D(n25081), .Z(n26530) );
    VMW_AO22 U1287 ( .A(matrixInput[246]), .B(n25096), .C(matrixInput[238]), 
        .D(n25081), .Z(n27018) );
    VMW_AO22 U1506 ( .A(matrixInput[1893]), .B(n25096), .C(matrixInput[1885]), 
        .D(n25081), .Z(n25371) );
    VMW_AO22 U1974 ( .A(matrixInput[1471]), .B(n25096), .C(matrixInput[1463]), 
        .D(n25081), .Z(n25793) );
    VMW_FD \matrixInput_reg[1345]  ( .D(n25911), .CP(Clk), .Q(matrixInput
        [1345]) );
    VMW_FD \matrixInput_reg[648]  ( .D(n26608), .CP(Clk), .Q(matrixInput[648])
         );
    VMW_AO22 U1317 ( .A(matrixInput[218]), .B(n25096), .C(matrixInput[210]), 
        .D(n25081), .Z(n27046) );
    VMW_AO22 U1496 ( .A(matrixInput[1902]), .B(n25096), .C(matrixInput[1894]), 
        .D(n25081), .Z(n25362) );
    VMW_FD \matrixInput_reg[651]  ( .D(n26605), .CP(Clk), .Q(matrixInput[651])
         );
    VMW_AO22 U1848 ( .A(matrixInput[1585]), .B(n25096), .C(matrixInput[1577]), 
        .D(n25081), .Z(n25679) );
    VMW_FD \matrixInput_reg[1046]  ( .D(n26210), .CP(Clk), .Q(matrixInput
        [1046]) );
    VMW_FD \vectorInput_reg[46]  ( .D(n27338), .CP(Clk), .Q(vectorInput[46])
         );
    VMW_FD \matrixInput_reg[926]  ( .D(n26330), .CP(Clk), .Q(matrixInput[926])
         );
    VMW_FD \matrixInput_reg[1885]  ( .D(n25371), .CP(Clk), .Q(matrixInput
        [1885]) );
    VMW_FD \vectorInput_reg[75]  ( .D(n27309), .CP(Clk), .Q(vectorInput[75])
         );
    VMW_AO22 U807 ( .A(matrixInput[678]), .B(n25096), .C(matrixInput[670]), 
        .D(n25081), .Z(n26586) );
    VMW_AO22 U997 ( .A(matrixInput[57]), .B(n25096), .C(matrixInput[49]), .D(
        n25081), .Z(n27207) );
    VMW_FD \matrixInput_reg[915]  ( .D(n26341), .CP(Clk), .Q(matrixInput[915])
         );
    VMW_FD \matrixInput_reg[1926]  ( .D(n25330), .CP(Clk), .Q(matrixInput
        [1926]) );
    VMW_FD \matrixInput_reg[5]  ( .D(n27251), .CP(Clk), .Q(matrixInput[5]) );
    VMW_AO22 U527 ( .A(matrixInput[930]), .B(n25096), .C(matrixInput[922]), 
        .D(n25081), .Z(n26334) );
    VMW_AO22 U762 ( .A(matrixInput[718]), .B(n25096), .C(matrixInput[710]), 
        .D(n25081), .Z(n26546) );
    VMW_AO22 U820 ( .A(matrixInput[667]), .B(n25096), .C(matrixInput[659]), 
        .D(n25081), .Z(n26597) );
    VMW_FD \matrixInput_reg[885]  ( .D(n26371), .CP(Clk), .Q(matrixInput[885])
         );
    VMW_AO22 U869 ( .A(matrixInput[622]), .B(n25096), .C(matrixInput[614]), 
        .D(n25081), .Z(n26642) );
    VMW_AO22 U1152 ( .A(matrixInput[43]), .B(n25096), .C(matrixInput[35]), .D(
        n25081), .Z(n27221) );
    VMW_AO22 U1743 ( .A(matrixInput[1679]), .B(n25096), .C(matrixInput[1671]), 
        .D(n25081), .Z(n25585) );
    VMW_FD \matrixInput_reg[1915]  ( .D(n25341), .CP(Clk), .Q(matrixInput
        [1915]) );
    VMW_FD \matrixInput_reg[1683]  ( .D(n25573), .CP(Clk), .Q(matrixInput
        [1683]) );
    VMW_AO22 U1175 ( .A(matrixInput[347]), .B(n25096), .C(matrixInput[339]), 
        .D(n25081), .Z(n26917) );
    VMW_AO22 U1245 ( .A(matrixInput[284]), .B(n25096), .C(matrixInput[276]), 
        .D(n25081), .Z(n26980) );
    VMW_AO22 U1262 ( .A(matrixInput[268]), .B(n25096), .C(matrixInput[260]), 
        .D(n25081), .Z(n26996) );
    VMW_AO22 U1473 ( .A(matrixInput[1922]), .B(n25096), .C(matrixInput[1914]), 
        .D(n25081), .Z(n25342) );
    VMW_AO22 U1801 ( .A(matrixInput[1627]), .B(n25096), .C(matrixInput[1619]), 
        .D(n25081), .Z(n25637) );
    VMW_AO22 U2162 ( .A(matrixInput[1302]), .B(n25096), .C(matrixInput[1294]), 
        .D(n25081), .Z(n25962) );
    VMW_FD \matrixInput_reg[1599]  ( .D(n25657), .CP(Clk), .Q(matrixInput
        [1599]) );
    VMW_FD \matrixInput_reg[1207]  ( .D(n26049), .CP(Clk), .Q(matrixInput
        [1207]) );
    VMW_FD \matrixInput_reg[410]  ( .D(n26846), .CP(Clk), .Q(matrixInput[410])
         );
    VMW_FD \matrixInput_reg[409]  ( .D(n26847), .CP(Clk), .Q(matrixInput[409])
         );
    VMW_FD \matrixInput_reg[1104]  ( .D(n26152), .CP(Clk), .Q(matrixInput
        [1104]) );
    VMW_FD \matrixInput_reg[713]  ( .D(n26543), .CP(Clk), .Q(matrixInput[713])
         );
    VMW_FD \matrixInput_reg[1580]  ( .D(n25676), .CP(Clk), .Q(matrixInput
        [1580]) );
    VMW_FD \matrixInput_reg[397]  ( .D(n26859), .CP(Clk), .Q(matrixInput[397])
         );
    VMW_AO22 U1991 ( .A(matrixInput[1456]), .B(n25096), .C(matrixInput[1448]), 
        .D(n25081), .Z(n25808) );
    VMW_FD \matrixInput_reg[1234]  ( .D(n26022), .CP(Clk), .Q(matrixInput
        [1234]) );
    VMW_FD \matrixInput_reg[423]  ( .D(n26833), .CP(Clk), .Q(matrixInput[423])
         );
    VMW_AO22 U1826 ( .A(matrixInput[1605]), .B(n25096), .C(matrixInput[1597]), 
        .D(n25081), .Z(n25659) );
    VMW_AO22 U2252 ( .A(matrixInput[1220]), .B(n25096), .C(matrixInput[1212]), 
        .D(n25081), .Z(n26044) );
    VMW_AO22 U2443 ( .A(matrixInput[1048]), .B(n25096), .C(matrixInput[1040]), 
        .D(n25081), .Z(n26216) );
    VMW_FD \matrixInput_reg[1137]  ( .D(n26119), .CP(Clk), .Q(matrixInput
        [1137]) );
    VMW_FD \matrixInput_reg[1094]  ( .D(n26162), .CP(Clk), .Q(matrixInput
        [1094]) );
    VMW_FD \matrixInput_reg[739]  ( .D(n26517), .CP(Clk), .Q(matrixInput[739])
         );
    VMW_FD \matrixInput_reg[720]  ( .D(n26536), .CP(Clk), .Q(matrixInput[720])
         );
    VMW_FD \vectorInput_reg[3]  ( .D(n27381), .CP(Clk), .Q(vectorInput[3]) );
    VMW_FD \matrixInput_reg[683]  ( .D(n26573), .CP(Clk), .Q(matrixInput[683])
         );
    VMW_FD \matrixInput_reg[1409]  ( .D(n25847), .CP(Clk), .Q(matrixInput
        [1409]) );
    VMW_FD \matrixInput_reg[207]  ( .D(n27049), .CP(Clk), .Q(matrixInput[207])
         );
    VMW_AO22 U1454 ( .A(matrixInput[1939]), .B(n25096), .C(matrixInput[1931]), 
        .D(n25081), .Z(n25325) );
    VMW_AO22 U2275 ( .A(matrixInput[1200]), .B(n25096), .C(matrixInput[1192]), 
        .D(n25081), .Z(n26064) );
    VMW_AO22 U2464 ( .A(matrixInput[1029]), .B(n25096), .C(matrixInput[1021]), 
        .D(n25081), .Z(n26235) );
    VMW_FD \matrixInput_reg[1713]  ( .D(n25543), .CP(Clk), .Q(matrixInput
        [1713]) );
    VMW_FD \matrixInput_reg[1410]  ( .D(n25846), .CP(Clk), .Q(matrixInput
        [1410]) );
    VMW_FD \matrixInput_reg[104]  ( .D(n27152), .CP(Clk), .Q(matrixInput[104])
         );
    VMW_FD \matrixInput_reg[1397]  ( .D(n25859), .CP(Clk), .Q(matrixInput
        [1397]) );
    VMW_FD \matrixInput_reg[599]  ( .D(n26657), .CP(Clk), .Q(matrixInput[599])
         );
    VMW_FD \matrixInput_reg[580]  ( .D(n26676), .CP(Clk), .Q(matrixInput[580])
         );
    VMW_AO22 U1764 ( .A(matrixInput[1660]), .B(n25096), .C(matrixInput[1652]), 
        .D(n25081), .Z(n25604) );
    VMW_FD \matrixInput_reg[1423]  ( .D(n25833), .CP(Clk), .Q(matrixInput
        [1423]) );
    VMW_FD \matrixInput_reg[234]  ( .D(n27022), .CP(Clk), .Q(matrixInput[234])
         );
    VMW_AO22 U2145 ( .A(matrixInput[1317]), .B(n25096), .C(matrixInput[1309]), 
        .D(n25081), .Z(n25947) );
    VMW_FD \matrixInput_reg[1720]  ( .D(n25536), .CP(Clk), .Q(matrixInput
        [1720]) );
    VMW_FD \matrixInput_reg[1739]  ( .D(n25517), .CP(Clk), .Q(matrixInput
        [1739]) );
    VMW_FD \matrixInput_reg[137]  ( .D(n27119), .CP(Clk), .Q(matrixInput[137])
         );
    VMW_AO22 U2079 ( .A(matrixInput[1377]), .B(n25096), .C(matrixInput[1369]), 
        .D(n25081), .Z(n25887) );
    VMW_AO22 U617 ( .A(matrixInput[849]), .B(n25096), .C(matrixInput[841]), 
        .D(n25081), .Z(n26415) );
    VMW_AO22 U955 ( .A(matrixInput[545]), .B(n25096), .C(matrixInput[537]), 
        .D(n25081), .Z(n26719) );
    VMW_FD \vectorInput_reg[117]  ( .D(n27267), .CP(Clk), .Q(vectorInput[117])
         );
    VMW_AO22 U1049 ( .A(matrixInput[460]), .B(n25096), .C(matrixInput[452]), 
        .D(n25081), .Z(n26804) );
    VMW_FD \matrixInput_reg[1857]  ( .D(n25399), .CP(Clk), .Q(matrixInput
        [1857]) );
    VMW_AO22 U1658 ( .A(matrixInput[1756]), .B(n25096), .C(matrixInput[1748]), 
        .D(n25081), .Z(n25508) );
    VMW_AO22 U2558 ( .A(cOutput[112]), .B(n25087), .C(cOutput[96]), .D(n25084), 
        .Z(n25180) );
    VMW_AO22 U630 ( .A(matrixInput[90]), .B(n25096), .C(matrixInput[82]), .D(
        n25081), .Z(n27174) );
    VMW_AO22 U787 ( .A(matrixInput[697]), .B(n25096), .C(matrixInput[689]), 
        .D(n25081), .Z(n26567) );
    VMW_FD \vectorInput_reg[124]  ( .D(n27260), .CP(Clk), .Q(vectorInput[124])
         );
    VMW_AO22 U1379 ( .A(matrixInput[207]), .B(n25096), .C(matrixInput[199]), 
        .D(n25081), .Z(n27057) );
    VMW_AO22 U2349 ( .A(matrixInput[1133]), .B(n25096), .C(matrixInput[1125]), 
        .D(n25081), .Z(n26131) );
    VMW_AO22 U1568 ( .A(matrixInput[1837]), .B(n25096), .C(matrixInput[1829]), 
        .D(n25081), .Z(n25427) );
    VMW_FD \matrixInput_reg[1864]  ( .D(n25392), .CP(Clk), .Q(matrixInput
        [1864]) );
    VMW_FD \vectorInput_reg[94]  ( .D(n27290), .CP(Clk), .Q(vectorInput[94])
         );
    VMW_FD \matrixInput_reg[17]  ( .D(n27239), .CP(Clk), .Q(matrixInput[17])
         );
    VMW_FD \matrixInput_reg[857]  ( .D(n26399), .CP(Clk), .Q(matrixInput[857])
         );
    VMW_AO22 U490 ( .A(matrixInput[964]), .B(n25096), .C(matrixInput[956]), 
        .D(n25081), .Z(n26300) );
    VMW_PULLDOWN U293 ( .Z(Logic01) );
    VMW_AO22 U324 ( .A(vectorInput[16]), .B(n25095), .C(vectorInput[8]), .D(
        n25080), .Z(n27376) );
    VMW_AO22 U500 ( .A(matrixInput[955]), .B(n25096), .C(matrixInput[947]), 
        .D(n25081), .Z(n26309) );
    VMW_AO22 U947 ( .A(matrixInput[552]), .B(n25096), .C(matrixInput[544]), 
        .D(n25081), .Z(n26712) );
    VMW_AO22 U972 ( .A(matrixInput[529]), .B(n25096), .C(matrixInput[521]), 
        .D(n25081), .Z(n26735) );
    VMW_FD \matrixInput_reg[918]  ( .D(n26338), .CP(Clk), .Q(matrixInput[918])
         );
    VMW_FD \matrixInput_reg[901]  ( .D(n26355), .CP(Clk), .Q(matrixInput[901])
         );
    VMW_FD \matrixInput_reg[864]  ( .D(n26392), .CP(Clk), .Q(matrixInput[864])
         );
    VMW_FD \matrixInput_reg[24]  ( .D(n27232), .CP(Clk), .Q(matrixInput[24])
         );
    VMW_AO22 U535 ( .A(matrixInput[923]), .B(n25096), .C(matrixInput[915]), 
        .D(n25081), .Z(n26341) );
    VMW_AO22 U605 ( .A(matrixInput[860]), .B(n25096), .C(matrixInput[852]), 
        .D(n25081), .Z(n26404) );
    VMW_AO22 U795 ( .A(matrixInput[689]), .B(n25096), .C(matrixInput[681]), 
        .D(n25081), .Z(n26575) );
    VMW_FD \matrixInput_reg[1891]  ( .D(n25365), .CP(Clk), .Q(matrixInput
        [1891]) );
    VMW_FD \matrixInput_reg[1888]  ( .D(n25368), .CP(Clk), .Q(matrixInput
        [1888]) );
    VMW_FD \vectorInput_reg[78]  ( .D(n27306), .CP(Clk), .Q(vectorInput[78])
         );
    VMW_FD \vectorInput_reg[61]  ( .D(n27323), .CP(Clk), .Q(vectorInput[61])
         );
    VMW_AO22 U622 ( .A(matrixInput[845]), .B(n25096), .C(matrixInput[837]), 
        .D(n25081), .Z(n26419) );
    VMW_AO22 U1898 ( .A(matrixInput[1539]), .B(n25096), .C(matrixInput[1531]), 
        .D(n25081), .Z(n25725) );
    VMW_AO22 U1908 ( .A(matrixInput[1530]), .B(n25096), .C(matrixInput[1522]), 
        .D(n25081), .Z(n25734) );
    VMW_FD \matrixInput_reg[932]  ( .D(n26324), .CP(Clk), .Q(matrixInput[932])
         );
    VMW_FD \vectorInput_reg[52]  ( .D(n27332), .CP(Clk), .Q(vectorInput[52])
         );
    IntMatMul_Control_pVectorSize16_pWordSize8_pScan1_DW01_cmp2_15_0 lt_130 ( 
        .A({Addr[14], Addr[13], Addr[12], Addr[11], Addr[10], Addr[9], Addr[8], 
        Addr[7], Addr[6], Addr[5], Addr[4], UNCONNECTED_1, UNCONNECTED_2, 
        UNCONNECTED_3, UNCONNECTED_4}), .B({Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic11, Logic01, 
        Logic01, Logic01, Logic01}), .LEQ(n27393), .TC(n27393), .LT_LE(n164)
         );
    VMW_AO22 U960 ( .A(matrixInput[540]), .B(n25096), .C(matrixInput[532]), 
        .D(n25081), .Z(n26724) );
    VMW_FD \matrixInput_reg[1918]  ( .D(n25338), .CP(Clk), .Q(matrixInput
        [1918]) );
    VMW_FD \matrixInput_reg[1901]  ( .D(n25355), .CP(Clk), .Q(matrixInput
        [1901]) );
    VMW_FD \matrixInput_reg[891]  ( .D(n26365), .CP(Clk), .Q(matrixInput[891])
         );
    VMW_FD \matrixInput_reg[888]  ( .D(n26368), .CP(Clk), .Q(matrixInput[888])
         );
    VMW_FD \matrixInput_reg[1932]  ( .D(n25324), .CP(Clk), .Q(matrixInput
        [1932]) );
    VMW_FD \matrixInput_reg[8]  ( .D(n27248), .CP(Clk), .Q(matrixInput[8]) );
    VMW_AND2 U303 ( .A(n25083), .B(n25055), .Z(n25082) );
    VMW_AO22 U512 ( .A(matrixInput[944]), .B(n25096), .C(matrixInput[936]), 
        .D(n25081), .Z(n26320) );
    VMW_AO22 U388 ( .A(vectorInput[39]), .B(n25095), .C(vectorInput[31]), .D(
        n25080), .Z(n27353) );
    VMW_AO22 U482 ( .A(matrixInput[971]), .B(n25096), .C(matrixInput[963]), 
        .D(n25081), .Z(n26293) );
    VMW_AO22 U599 ( .A(matrixInput[866]), .B(n25096), .C(matrixInput[858]), 
        .D(n25081), .Z(n26398) );
    VMW_AO22 U739 ( .A(matrixInput[739]), .B(n25096), .C(matrixInput[731]), 
        .D(n25081), .Z(n26525) );
    VMW_AO22 U1140 ( .A(matrixInput[378]), .B(n25096), .C(matrixInput[370]), 
        .D(n25081), .Z(n26886) );
    VMW_FD \matrixInput_reg[1645]  ( .D(n25611), .CP(Clk), .Q(matrixInput
        [1645]) );
    VMW_AO22 U1257 ( .A(matrixInput[273]), .B(n25096), .C(matrixInput[265]), 
        .D(n25081), .Z(n26991) );
    VMW_AO22 U1270 ( .A(matrixInput[261]), .B(n25096), .C(matrixInput[253]), 
        .D(n25081), .Z(n27003) );
    VMW_AO22 U1751 ( .A(matrixInput[1672]), .B(n25096), .C(matrixInput[1664]), 
        .D(n25081), .Z(n25592) );
    VMW_AO22 U2170 ( .A(matrixInput[1295]), .B(n25096), .C(matrixInput[1287]), 
        .D(n25081), .Z(n25969) );
    VMW_FD \matrixInput_reg[2022]  ( .D(n25234), .CP(Clk), .Q(matrixInput
        [2022]) );
    VMW_FD \matrixInput_reg[1546]  ( .D(n25710), .CP(Clk), .Q(matrixInput
        [1546]) );
    VMW_FD \matrixInput_reg[351]  ( .D(n26905), .CP(Clk), .Q(matrixInput[351])
         );
    VMW_FD \matrixInput_reg[348]  ( .D(n26908), .CP(Clk), .Q(matrixInput[348])
         );
    VMW_AO22 U1446 ( .A(matrixInput[1947]), .B(n25096), .C(matrixInput[1939]), 
        .D(n25081), .Z(n25317) );
    VMW_AO22 U1461 ( .A(matrixInput[1933]), .B(n25096), .C(matrixInput[1925]), 
        .D(n25081), .Z(n25331) );
    VMW_AO22 U1813 ( .A(matrixInput[1616]), .B(n25096), .C(matrixInput[1608]), 
        .D(n25081), .Z(n25648) );
    VMW_AO22 U1983 ( .A(matrixInput[1463]), .B(n25096), .C(matrixInput[1455]), 
        .D(n25081), .Z(n25801) );
    VMW_FD \matrixInput_reg[1676]  ( .D(n25580), .CP(Clk), .Q(matrixInput
        [1676]) );
    VMW_AO22 U2240 ( .A(matrixInput[1231]), .B(n25096), .C(matrixInput[1223]), 
        .D(n25081), .Z(n26033) );
    VMW_AO22 U2451 ( .A(matrixInput[1041]), .B(n25096), .C(matrixInput[1033]), 
        .D(n25081), .Z(n26223) );
    VMW_FD \matrixInput_reg[2011]  ( .D(n25245), .CP(Clk), .Q(matrixInput
        [2011]) );
    VMW_FD \matrixInput_reg[1575]  ( .D(n25681), .CP(Clk), .Q(matrixInput
        [1575]) );
    VMW_FD \matrixInput_reg[362]  ( .D(n26894), .CP(Clk), .Q(matrixInput[362])
         );
    VMW_FD \matrixInput_reg[2008]  ( .D(n25248), .CP(Clk), .Q(matrixInput
        [2008]) );
    VMW_FD \matrixInput_reg[645]  ( .D(n26611), .CP(Clk), .Q(matrixInput[645])
         );
    VMW_AO22 U1834 ( .A(matrixInput[166]), .B(n25096), .C(matrixInput[158]), 
        .D(n25081), .Z(n27098) );
    VMW_FD \matrixInput_reg[1052]  ( .D(n26204), .CP(Clk), .Q(matrixInput
        [1052]) );
    VMW_AO22 U2267 ( .A(matrixInput[127]), .B(n25096), .C(matrixInput[119]), 
        .D(n25081), .Z(n27137) );
    VMW_FD \matrixInput_reg[546]  ( .D(n26710), .CP(Clk), .Q(matrixInput[546])
         );
    VMW_AO22 U2476 ( .A(matrixInput[1018]), .B(n25096), .C(matrixInput[1010]), 
        .D(n25081), .Z(n26246) );
    VMW_AO22 U1167 ( .A(matrixInput[354]), .B(n25096), .C(matrixInput[346]), 
        .D(n25081), .Z(n26910) );
    VMW_AO22 U1776 ( .A(matrixInput[1649]), .B(n25096), .C(matrixInput[1641]), 
        .D(n25081), .Z(n25615) );
    VMW_FD \matrixInput_reg[1351]  ( .D(n25905), .CP(Clk), .Q(matrixInput
        [1351]) );
    VMW_FD \matrixInput_reg[1348]  ( .D(n25908), .CP(Clk), .Q(matrixInput
        [1348]) );
    VMW_FD \matrixInput_reg[1078]  ( .D(n26178), .CP(Clk), .Q(matrixInput
        [1078]) );
    VMW_FD \matrixInput_reg[1061]  ( .D(n26195), .CP(Clk), .Q(matrixInput
        [1061]) );
    VMW_AO22 U2157 ( .A(matrixInput[1307]), .B(n25096), .C(matrixInput[1299]), 
        .D(n25081), .Z(n25957) );
    VMW_FD \matrixInput_reg[1362]  ( .D(n25894), .CP(Clk), .Q(matrixInput
        [1362]) );
    VMW_FD \matrixInput_reg[676]  ( .D(n26580), .CP(Clk), .Q(matrixInput[676])
         );
    VMW_FD \matrixInput_reg[575]  ( .D(n26681), .CP(Clk), .Q(matrixInput[575])
         );
    VMW_AO22 U409 ( .A(vectorInput[20]), .B(n25095), .C(vectorInput[12]), .D(
        n25080), .Z(n27372) );
    VMW_AO22 U467 ( .A(matrixInput[985]), .B(n25096), .C(matrixInput[977]), 
        .D(n25081), .Z(n26279) );
    VMW_AO22 U757 ( .A(matrixInput[723]), .B(n25096), .C(matrixInput[715]), 
        .D(n25081), .Z(n26541) );
    VMW_AO22 U1239 ( .A(matrixInput[289]), .B(n25096), .C(matrixInput[281]), 
        .D(n25081), .Z(n26975) );
    VMW_FD \matrixInput_reg[1870]  ( .D(n25386), .CP(Clk), .Q(matrixInput
        [1870]) );
    VMW_FD \matrixInput_reg[1869]  ( .D(n25387), .CP(Clk), .Q(matrixInput
        [1869]) );
    VMW_AO22 U1428 ( .A(matrixInput[1963]), .B(n25096), .C(matrixInput[1955]), 
        .D(n25081), .Z(n25301) );
    VMW_AO22 U2418 ( .A(matrixInput[1071]), .B(n25096), .C(matrixInput[1063]), 
        .D(n25081), .Z(n26193) );
    VMW_FD \vectorInput_reg[99]  ( .D(n27285), .CP(Clk), .Q(vectorInput[99])
         );
    VMW_FD \vectorInput_reg[80]  ( .D(n27304), .CP(Clk), .Q(vectorInput[80])
         );
    VMW_AO22 U815 ( .A(matrixInput[671]), .B(n25096), .C(matrixInput[663]), 
        .D(n25081), .Z(n26593) );
    VMW_AO22 U1099 ( .A(matrixInput[415]), .B(n25096), .C(matrixInput[407]), 
        .D(n25081), .Z(n26849) );
    VMW_AO22 U1109 ( .A(matrixInput[407]), .B(n25096), .C(matrixInput[399]), 
        .D(n25081), .Z(n26857) );
    VMW_AO22 U2209 ( .A(matrixInput[1259]), .B(n25096), .C(matrixInput[1251]), 
        .D(n25081), .Z(n26005) );
    VMW_AO22 U2399 ( .A(matrixInput[1088]), .B(n25096), .C(matrixInput[1080]), 
        .D(n25081), .Z(n26176) );
    VMW_OAI21 U2588 ( .A(n25165), .B(n25166), .C(n25091), .Z(n25171) );
    VMW_AO22 U1688 ( .A(matrixInput[1728]), .B(n25096), .C(matrixInput[1720]), 
        .D(n25081), .Z(n25536) );
    VMW_AO22 U1718 ( .A(matrixInput[1702]), .B(n25096), .C(matrixInput[1694]), 
        .D(n25081), .Z(n25562) );
    VMW_FD \matrixInput_reg[1843]  ( .D(n25413), .CP(Clk), .Q(matrixInput
        [1843]) );
    VMW_AO22 U985 ( .A(matrixInput[58]), .B(n25096), .C(matrixInput[50]), .D(
        n25081), .Z(n27206) );
    VMW_AO22 U2139 ( .A(matrixInput[1322]), .B(n25096), .C(matrixInput[1314]), 
        .D(n25081), .Z(n25942) );
    VMW_PULLDOWN U280 ( .Z(n25198) );
    VMW_PULLDOWN U288 ( .Z(n25206) );
    VMW_AO22 U351 ( .A(vectorInput[73]), .B(n25095), .C(vectorInput[65]), .D(
        n25080), .Z(n27319) );
    VMW_AO22 U440 ( .A(vectorInput[8]), .B(n25095), .C(vectorInput[0]), .D(
        n25080), .Z(n27384) );
    VMW_AO22 U832 ( .A(matrixInput[656]), .B(n25096), .C(matrixInput[648]), 
        .D(n25081), .Z(n26608) );
    VMW_FD \matrixInput_reg[870]  ( .D(n26386), .CP(Clk), .Q(matrixInput[870])
         );
    VMW_FD \matrixInput_reg[869]  ( .D(n26387), .CP(Clk), .Q(matrixInput[869])
         );
    VMW_FD \vectorInput_reg[103]  ( .D(n27281), .CP(Clk), .Q(vectorInput[103])
         );
    VMW_FD \matrixInput_reg[30]  ( .D(n27226), .CP(Clk), .Q(matrixInput[30])
         );
    VMW_FD \matrixInput_reg[29]  ( .D(n27227), .CP(Clk), .Q(matrixInput[29])
         );
    VMW_AO22 U540 ( .A(matrixInput[918]), .B(n25096), .C(matrixInput[910]), 
        .D(n25081), .Z(n26346) );
    VMW_AO22 U670 ( .A(matrixInput[802]), .B(n25096), .C(matrixInput[794]), 
        .D(n25081), .Z(n26462) );
    VMW_AO22 U770 ( .A(matrixInput[711]), .B(n25096), .C(matrixInput[703]), 
        .D(n25081), .Z(n26553) );
    VMW_FD \matrixInput_reg[843]  ( .D(n26413), .CP(Clk), .Q(matrixInput[843])
         );
    VMW_AO22 U929 ( .A(matrixInput[568]), .B(n25096), .C(matrixInput[560]), 
        .D(n25081), .Z(n26696) );
    VMW_AO22 U1012 ( .A(matrixInput[494]), .B(n25096), .C(matrixInput[486]), 
        .D(n25081), .Z(n26770) );
    VMW_AO22 U1182 ( .A(matrixInput[340]), .B(n25096), .C(matrixInput[332]), 
        .D(n25081), .Z(n26924) );
    VMW_AO22 U1322 ( .A(matrixInput[214]), .B(n25096), .C(matrixInput[206]), 
        .D(n25081), .Z(n27050) );
    VMW_AO22 U1533 ( .A(matrixInput[1868]), .B(n25096), .C(matrixInput[1860]), 
        .D(n25081), .Z(n25396) );
    VMW_AO22 U2282 ( .A(matrixInput[1194]), .B(n25096), .C(matrixInput[1186]), 
        .D(n25081), .Z(n26070) );
    VMW_AO22 U2312 ( .A(matrixInput[1167]), .B(n25096), .C(matrixInput[1159]), 
        .D(n25081), .Z(n26097) );
    VMW_AO22 U2493 ( .A(cOutput[87]), .B(n25087), .C(cOutput[71]), .D(n25084), 
        .Z(n25101) );
    VMW_FD \matrixInput_reg[1123]  ( .D(n26133), .CP(Clk), .Q(matrixInput
        [1123]) );
    VMW_FD \matrixInput_reg[734]  ( .D(n26522), .CP(Clk), .Q(matrixInput[734])
         );
    VMW_AO22 U2503 ( .A(cOutput[94]), .B(n25089), .C(cOutput[78]), .D(n25088), 
        .Z(n25113) );
    VMW_AO22 U1941 ( .A(matrixInput[1501]), .B(n25096), .C(matrixInput[1493]), 
        .D(n25081), .Z(n25763) );
    VMW_AO22 U2022 ( .A(matrixInput[149]), .B(n25096), .C(matrixInput[141]), 
        .D(n25081), .Z(n27115) );
    VMW_FD \matrixInput_reg[1594]  ( .D(n25662), .CP(Clk), .Q(matrixInput
        [1594]) );
    VMW_FD \matrixInput_reg[1239]  ( .D(n26017), .CP(Clk), .Q(matrixInput
        [1239]) );
    VMW_FD \matrixInput_reg[1220]  ( .D(n26036), .CP(Clk), .Q(matrixInput
        [1220]) );
    VMW_FD \matrixInput_reg[437]  ( .D(n26819), .CP(Clk), .Q(matrixInput[437])
         );
    VMW_BUFIZ U2633 ( .A(\holder[7] ), .E(RD), .Z(\DataOut[7]1 ) );
    VMW_FD \matrixInput_reg[383]  ( .D(n26873), .CP(Clk), .Q(matrixInput[383])
         );
    VMW_FD \matrixInput_reg[1697]  ( .D(n25559), .CP(Clk), .Q(matrixInput
        [1697]) );
    VMW_FD \matrixInput_reg[1213]  ( .D(n26043), .CP(Clk), .Q(matrixInput
        [1213]) );
    VMW_FD \matrixInput_reg[1110]  ( .D(n26146), .CP(Clk), .Q(matrixInput
        [1110]) );
    VMW_FD \matrixInput_reg[707]  ( .D(n26549), .CP(Clk), .Q(matrixInput[707])
         );
    VMW_FD \matrixInput_reg[1109]  ( .D(n26147), .CP(Clk), .Q(matrixInput
        [1109]) );
    VMW_FD \matrixInput_reg[404]  ( .D(n26852), .CP(Clk), .Q(matrixInput[404])
         );
    VMW_AO22 U1603 ( .A(matrixInput[1806]), .B(n25096), .C(matrixInput[1798]), 
        .D(n25081), .Z(n25458) );
    VMW_AO22 U1793 ( .A(matrixInput[1634]), .B(n25096), .C(matrixInput[1626]), 
        .D(n25081), .Z(n25630) );
    VMW_AO22 U2005 ( .A(matrixInput[1443]), .B(n25096), .C(matrixInput[1435]), 
        .D(n25081), .Z(n25821) );
    VMW_AO22 U2195 ( .A(matrixInput[1272]), .B(n25096), .C(matrixInput[1264]), 
        .D(n25081), .Z(n25992) );
    VMW_BUFIZ U2614 ( .A(n25190), .E(RD), .Z(\DataOut[9]1 ) );
    VMW_FD \matrixInput_reg[1734]  ( .D(n25522), .CP(Clk), .Q(matrixInput
        [1734]) );
    VMW_FD \matrixInput_reg[123]  ( .D(n27133), .CP(Clk), .Q(matrixInput[123])
         );
    VMW_AO22 U1035 ( .A(matrixInput[473]), .B(n25096), .C(matrixInput[465]), 
        .D(n25081), .Z(n26791) );
    VMW_AO22 U1295 ( .A(matrixInput[238]), .B(n25096), .C(matrixInput[230]), 
        .D(n25081), .Z(n27026) );
    VMW_AO22 U1305 ( .A(matrixInput[229]), .B(n25096), .C(matrixInput[221]), 
        .D(n25081), .Z(n27035) );
    VMW_AO22 U1484 ( .A(matrixInput[1912]), .B(n25096), .C(matrixInput[1904]), 
        .D(n25081), .Z(n25352) );
    VMW_AO22 U1624 ( .A(matrixInput[1787]), .B(n25096), .C(matrixInput[1779]), 
        .D(n25081), .Z(n25477) );
    VMW_AO22 U2335 ( .A(matrixInput[1146]), .B(n25096), .C(matrixInput[1138]), 
        .D(n25081), .Z(n26118) );
    VMW_AND3 U2524 ( .A(n25138), .B(n25139), .C(n25140), .Z(n25070) );
    VMW_FD \matrixInput_reg[1707]  ( .D(n25549), .CP(Clk), .Q(matrixInput
        [1707]) );
    VMW_FD \matrixInput_reg[1437]  ( .D(n25819), .CP(Clk), .Q(matrixInput
        [1437]) );
    VMW_FD \matrixInput_reg[1383]  ( .D(n25873), .CP(Clk), .Q(matrixInput
        [1383]) );
    VMW_FD \matrixInput_reg[239]  ( .D(n27017), .CP(Clk), .Q(matrixInput[239])
         );
    VMW_FD \matrixInput_reg[220]  ( .D(n27036), .CP(Clk), .Q(matrixInput[220])
         );
    VMW_FD \matrixInput_reg[594]  ( .D(n26662), .CP(Clk), .Q(matrixInput[594])
         );
    VMW_FD \matrixInput_reg[110]  ( .D(n27146), .CP(Clk), .Q(matrixInput[110])
         );
    VMW_FD \matrixInput_reg[109]  ( .D(n27147), .CP(Clk), .Q(matrixInput[109])
         );
    VMW_FD \matrixInput_reg[213]  ( .D(n27043), .CP(Clk), .Q(matrixInput[213])
         );
    VMW_AO22 U1514 ( .A(matrixInput[1886]), .B(n25096), .C(matrixInput[1878]), 
        .D(n25081), .Z(n25378) );
    VMW_FD \matrixInput_reg[1404]  ( .D(n25852), .CP(Clk), .Q(matrixInput
        [1404]) );
    VMW_AO22 U1966 ( .A(matrixInput[1478]), .B(n25096), .C(matrixInput[1470]), 
        .D(n25081), .Z(n25786) );
    VMW_FD \matrixInput_reg[1099]  ( .D(n26157), .CP(Clk), .Q(matrixInput
        [1099]) );
    VMW_FD \matrixInput_reg[1080]  ( .D(n26176), .CP(Clk), .Q(matrixInput
        [1080]) );
    VMW_FD \matrixInput_reg[697]  ( .D(n26559), .CP(Clk), .Q(matrixInput[697])
         );
    VMW_FD \matrixInput_reg[853]  ( .D(n26403), .CP(Clk), .Q(matrixInput[853])
         );
    VMW_AO22 U932 ( .A(matrixInput[566]), .B(n25096), .C(matrixInput[558]), 
        .D(n25081), .Z(n26698) );
    VMW_FD \matrixInput_reg[879]  ( .D(n26377), .CP(Clk), .Q(matrixInput[879])
         );
    VMW_FD \matrixInput_reg[860]  ( .D(n26396), .CP(Clk), .Q(matrixInput[860])
         );
    VMW_FD \matrixInput_reg[13]  ( .D(n27243), .CP(Clk), .Q(matrixInput[13])
         );
    VMW_FD \matrixInput_reg[39]  ( .D(n27217), .CP(Clk), .Q(matrixInput[39])
         );
    VMW_FD \matrixInput_reg[20]  ( .D(n27236), .CP(Clk), .Q(matrixInput[20])
         );
    VMW_AO22 U376 ( .A(vectorInput[50]), .B(n25095), .C(vectorInput[42]), .D(
        n25080), .Z(n27342) );
    VMW_AO22 U885 ( .A(matrixInput[13]), .B(n25096), .C(matrixInput[5]), .D(
        n25081), .Z(n27251) );
    VMW_AO22 U1009 ( .A(matrixInput[497]), .B(n25096), .C(matrixInput[489]), 
        .D(n25081), .Z(n26767) );
    VMW_AO22 U1199 ( .A(matrixInput[325]), .B(n25096), .C(matrixInput[317]), 
        .D(n25081), .Z(n26939) );
    VMW_AO22 U1618 ( .A(matrixInput[1792]), .B(n25096), .C(matrixInput[1784]), 
        .D(n25081), .Z(n25472) );
    VMW_AO22 U1788 ( .A(matrixInput[1638]), .B(n25096), .C(matrixInput[1630]), 
        .D(n25081), .Z(n25626) );
    VMW_FD \matrixInput_reg[1853]  ( .D(n25403), .CP(Clk), .Q(matrixInput
        [1853]) );
    VMW_AO22 U915 ( .A(matrixInput[581]), .B(n25096), .C(matrixInput[573]), 
        .D(n25081), .Z(n26683) );
    VMW_AO22 U2039 ( .A(matrixInput[1412]), .B(n25096), .C(matrixInput[1404]), 
        .D(n25081), .Z(n25852) );
    VMW_AO22 U393 ( .A(vectorInput[35]), .B(n25095), .C(vectorInput[27]), .D(
        n25080), .Z(n27357) );
    VMW_AO22 U567 ( .A(matrixInput[895]), .B(n25096), .C(matrixInput[887]), 
        .D(n25081), .Z(n26369) );
    VMW_BUFIZ U2628 ( .A(n25201), .E(RD), .Z(\DataOut[26]1 ) );
    VMW_FD \vectorInput_reg[113]  ( .D(n27271), .CP(Clk), .Q(vectorInput[113])
         );
    VMW_AO22 U582 ( .A(matrixInput[881]), .B(n25096), .C(matrixInput[873]), 
        .D(n25081), .Z(n26383) );
    VMW_AO22 U657 ( .A(matrixInput[813]), .B(n25096), .C(matrixInput[805]), 
        .D(n25081), .Z(n26451) );
    VMW_AO22 U1339 ( .A(matrixInput[2042]), .B(n25096), .C(matrixInput[2034]), 
        .D(n25081), .Z(n25222) );
    VMW_AO22 U1528 ( .A(matrixInput[1873]), .B(n25096), .C(matrixInput[1865]), 
        .D(n25081), .Z(n25391) );
    VMW_FD \matrixInput_reg[1879]  ( .D(n25377), .CP(Clk), .Q(matrixInput
        [1879]) );
    VMW_FD \matrixInput_reg[1860]  ( .D(n25396), .CP(Clk), .Q(matrixInput
        [1860]) );
    VMW_FD \vectorInput_reg[90]  ( .D(n27294), .CP(Clk), .Q(vectorInput[90])
         );
    VMW_FD \vectorInput_reg[89]  ( .D(n27295), .CP(Clk), .Q(vectorInput[89])
         );
    VMW_AO22 U2309 ( .A(matrixInput[1169]), .B(n25096), .C(matrixInput[1161]), 
        .D(n25081), .Z(n26095) );
    VMW_AO22 U2488 ( .A(matrixInput[8]), .B(n25096), .C(matrixInput[0]), .D(
        n25081), .Z(n27256) );
    VMW_FD \vectorInput_reg[120]  ( .D(n27264), .CP(Clk), .Q(vectorInput[120])
         );
    VMW_AO22 U2518 ( .A(cOutput[52]), .B(n25087), .C(cOutput[36]), .D(n25084), 
        .Z(n25132) );
    VMW_AO22 U829 ( .A(matrixInput[658]), .B(n25096), .C(matrixInput[650]), 
        .D(n25081), .Z(n26606) );
    VMW_AO22 U1205 ( .A(matrixInput[319]), .B(n25096), .C(matrixInput[311]), 
        .D(n25081), .Z(n26945) );
    VMW_AO22 U1395 ( .A(matrixInput[1993]), .B(n25096), .C(matrixInput[1985]), 
        .D(n25081), .Z(n25271) );
    VMW_AO22 U1414 ( .A(matrixInput[1976]), .B(n25096), .C(matrixInput[1968]), 
        .D(n25081), .Z(n25288) );
    VMW_AO22 U2235 ( .A(matrixInput[1236]), .B(n25096), .C(matrixInput[1228]), 
        .D(n25081), .Z(n26028) );
    VMW_AO22 U2299 ( .A(matrixInput[1178]), .B(n25096), .C(matrixInput[1170]), 
        .D(n25081), .Z(n26086) );
    VMW_FD \matrixInput_reg[1393]  ( .D(n25863), .CP(Clk), .Q(matrixInput
        [1393]) );
    VMW_FD \matrixInput_reg[584]  ( .D(n26672), .CP(Clk), .Q(matrixInput[584])
         );
    VMW_AO22 U2424 ( .A(matrixInput[1066]), .B(n25096), .C(matrixInput[1058]), 
        .D(n25081), .Z(n26198) );
    VMW_FD \matrixInput_reg[1717]  ( .D(n25539), .CP(Clk), .Q(matrixInput
        [1717]) );
    VMW_FD \matrixInput_reg[119]  ( .D(n27137), .CP(Clk), .Q(matrixInput[119])
         );
    VMW_FD \matrixInput_reg[100]  ( .D(n27156), .CP(Clk), .Q(matrixInput[100])
         );
    VMW_FD \matrixInput_reg[1414]  ( .D(n25842), .CP(Clk), .Q(matrixInput
        [1414]) );
    VMW_AO22 U1584 ( .A(matrixInput[1822]), .B(n25096), .C(matrixInput[1814]), 
        .D(n25081), .Z(n25442) );
    VMW_AO22 U1866 ( .A(matrixInput[1568]), .B(n25096), .C(matrixInput[1560]), 
        .D(n25081), .Z(n25696) );
    VMW_FD \matrixInput_reg[203]  ( .D(n27053), .CP(Clk), .Q(matrixInput[203])
         );
    VMW_AO22 U2095 ( .A(matrixInput[1362]), .B(n25096), .C(matrixInput[1354]), 
        .D(n25081), .Z(n25902) );
    VMW_AO22 U2105 ( .A(matrixInput[1353]), .B(n25096), .C(matrixInput[1345]), 
        .D(n25081), .Z(n25911) );
    VMW_FD \matrixInput_reg[1090]  ( .D(n26166), .CP(Clk), .Q(matrixInput
        [1090]) );
    VMW_FD \matrixInput_reg[1089]  ( .D(n26167), .CP(Clk), .Q(matrixInput
        [1089]) );
    VMW_FD \matrixInput_reg[687]  ( .D(n26569), .CP(Clk), .Q(matrixInput[687])
         );
    VMW_FD \matrixInput_reg[133]  ( .D(n27123), .CP(Clk), .Q(matrixInput[133])
         );
    VMW_FD \matrixInput_reg[1724]  ( .D(n25532), .CP(Clk), .Q(matrixInput
        [1724]) );
    VMW_AO22 U860 ( .A(matrixInput[630]), .B(n25096), .C(matrixInput[622]), 
        .D(n25081), .Z(n26634) );
    VMW_AO22 U1082 ( .A(matrixInput[430]), .B(n25096), .C(matrixInput[422]), 
        .D(n25081), .Z(n26834) );
    VMW_AO22 U1112 ( .A(matrixInput[404]), .B(n25096), .C(matrixInput[396]), 
        .D(n25081), .Z(n26860) );
    VMW_AO22 U1135 ( .A(matrixInput[383]), .B(n25096), .C(matrixInput[375]), 
        .D(n25081), .Z(n26881) );
    VMW_AO22 U1724 ( .A(matrixInput[1697]), .B(n25096), .C(matrixInput[1689]), 
        .D(n25081), .Z(n25567) );
    VMW_FD \matrixInput_reg[230]  ( .D(n27026), .CP(Clk), .Q(matrixInput[230])
         );
    VMW_FD \matrixInput_reg[229]  ( .D(n27027), .CP(Clk), .Q(matrixInput[229])
         );
    VMW_FD \matrixInput_reg[1427]  ( .D(n25829), .CP(Clk), .Q(matrixInput
        [1427]) );
    VMW_AO22 U2122 ( .A(matrixInput[140]), .B(n25096), .C(matrixInput[132]), 
        .D(n25081), .Z(n27124) );
    VMW_FD \matrixInput_reg[393]  ( .D(n26863), .CP(Clk), .Q(matrixInput[393])
         );
    VMW_FD \matrixInput_reg[1584]  ( .D(n25672), .CP(Clk), .Q(matrixInput
        [1584]) );
    VMW_FD \matrixInput_reg[1203]  ( .D(n26053), .CP(Clk), .Q(matrixInput
        [1203]) );
    VMW_FD \matrixInput_reg[1119]  ( .D(n26137), .CP(Clk), .Q(matrixInput
        [1119]) );
    VMW_FD \matrixInput_reg[1100]  ( .D(n26156), .CP(Clk), .Q(matrixInput
        [1100]) );
    VMW_FD \matrixInput_reg[717]  ( .D(n26539), .CP(Clk), .Q(matrixInput[717])
         );
    VMW_FD \matrixInput_reg[414]  ( .D(n26842), .CP(Clk), .Q(matrixInput[414])
         );
    VMW_AO22 U1693 ( .A(matrixInput[1724]), .B(n25096), .C(matrixInput[1716]), 
        .D(n25081), .Z(n25540) );
    VMW_AO22 U1222 ( .A(matrixInput[305]), .B(n25096), .C(matrixInput[297]), 
        .D(n25081), .Z(n26959) );
    VMW_AO22 U1703 ( .A(matrixInput[1715]), .B(n25096), .C(matrixInput[1707]), 
        .D(n25081), .Z(n25549) );
    VMW_AO22 U2212 ( .A(matrixInput[1257]), .B(n25096), .C(matrixInput[1249]), 
        .D(n25081), .Z(n26007) );
    VMW_AO22 U2382 ( .A(matrixInput[1104]), .B(n25096), .C(matrixInput[1096]), 
        .D(n25081), .Z(n26160) );
    VMW_AO22 U2403 ( .A(matrixInput[1085]), .B(n25096), .C(matrixInput[1077]), 
        .D(n25081), .Z(n26179) );
    VMW_FD \matrixInput_reg[1687]  ( .D(n25569), .CP(Clk), .Q(matrixInput
        [1687]) );
    VMW_FD \matrixInput_reg[1133]  ( .D(n26123), .CP(Clk), .Q(matrixInput
        [1133]) );
    VMW_FD \matrixInput_reg[724]  ( .D(n26532), .CP(Clk), .Q(matrixInput[724])
         );
    VMW_FD \vectorInput_reg[7]  ( .D(n27377), .CP(Clk), .Q(vectorInput[7]) );
    VMW_OAI21 U2593 ( .A(n25178), .B(n25179), .C(n25093), .Z(n25184) );
    VMW_AO22 U1433 ( .A(matrixInput[1958]), .B(n25096), .C(matrixInput[1950]), 
        .D(n25081), .Z(n25306) );
    VMW_AO22 U1841 ( .A(matrixInput[1591]), .B(n25096), .C(matrixInput[1583]), 
        .D(n25081), .Z(n25673) );
    VMW_FD \matrixInput_reg[1230]  ( .D(n26026), .CP(Clk), .Q(matrixInput
        [1230]) );
    VMW_FD \matrixInput_reg[427]  ( .D(n26829), .CP(Clk), .Q(matrixInput[427])
         );
    VMW_FD \matrixInput_reg[1229]  ( .D(n26027), .CP(Clk), .Q(matrixInput
        [1229]) );
    VMW_AO22 U412 ( .A(DataIn[5]), .B(n25095), .C(vectorInput[125]), .D(n25080
        ), .Z(n27259) );
    VMW_AO22 U435 ( .A(vectorInput[112]), .B(n25095), .C(vectorInput[104]), 
        .D(n25080), .Z(n27280) );
    VMW_AO22 U695 ( .A(matrixInput[779]), .B(n25096), .C(matrixInput[771]), 
        .D(n25081), .Z(n26485) );
    VMW_AO22 U705 ( .A(matrixInput[770]), .B(n25096), .C(matrixInput[762]), 
        .D(n25081), .Z(n26494) );
    VMW_AO22 U722 ( .A(matrixInput[755]), .B(n25096), .C(matrixInput[747]), 
        .D(n25081), .Z(n26509) );
    VMW_FD \matrixInput_reg[1922]  ( .D(n25334), .CP(Clk), .Q(matrixInput
        [1922]) );
    VMW_FD \matrixInput_reg[1]  ( .D(n27255), .CP(Clk), .Q(matrixInput[1]) );
    VMW_FD \matrixInput_reg[1911]  ( .D(n25345), .CP(Clk), .Q(matrixInput
        [1911]) );
    VMW_FD \matrixInput_reg[1908]  ( .D(n25348), .CP(Clk), .Q(matrixInput
        [1908]) );
    VMW_FD \matrixInput_reg[898]  ( .D(n26358), .CP(Clk), .Q(matrixInput[898])
         );
    VMW_FD \matrixInput_reg[881]  ( .D(n26375), .CP(Clk), .Q(matrixInput[881])
         );
    VMW_AO22 U847 ( .A(matrixInput[642]), .B(n25096), .C(matrixInput[634]), 
        .D(n25081), .Z(n26622) );
    VMW_AO22 U1808 ( .A(matrixInput[1620]), .B(n25096), .C(matrixInput[1612]), 
        .D(n25081), .Z(n25644) );
    VMW_AO22 U1998 ( .A(matrixInput[1449]), .B(n25096), .C(matrixInput[1441]), 
        .D(n25081), .Z(n25815) );
    VMW_FD \matrixInput_reg[922]  ( .D(n26334), .CP(Clk), .Q(matrixInput[922])
         );
    VMW_FD \vectorInput_reg[42]  ( .D(n27342), .CP(Clk), .Q(vectorInput[42])
         );
    VMW_FD \matrixInput_reg[911]  ( .D(n26345), .CP(Clk), .Q(matrixInput[911])
         );
    VMW_FD \matrixInput_reg[908]  ( .D(n26348), .CP(Clk), .Q(matrixInput[908])
         );
    VMW_AO22 U1067 ( .A(matrixInput[444]), .B(n25096), .C(matrixInput[436]), 
        .D(n25081), .Z(n26820) );
    VMW_FD \matrixInput_reg[1898]  ( .D(n25358), .CP(Clk), .Q(matrixInput
        [1898]) );
    VMW_FD \matrixInput_reg[1881]  ( .D(n25375), .CP(Clk), .Q(matrixInput
        [1881]) );
    VMW_FD \vectorInput_reg[71]  ( .D(n27313), .CP(Clk), .Q(vectorInput[71])
         );
    VMW_FD \vectorInput_reg[68]  ( .D(n27316), .CP(Clk), .Q(vectorInput[68])
         );
    VMW_AO22 U1676 ( .A(matrixInput[1739]), .B(n25096), .C(matrixInput[1731]), 
        .D(n25081), .Z(n25525) );
    VMW_FD \matrixInput_reg[666]  ( .D(n26590), .CP(Clk), .Q(matrixInput[666])
         );
    VMW_FD \matrixInput_reg[1071]  ( .D(n26185), .CP(Clk), .Q(matrixInput
        [1071]) );
    VMW_FD \matrixInput_reg[1068]  ( .D(n26188), .CP(Clk), .Q(matrixInput
        [1068]) );
    VMW_AO22 U318 ( .A(vectorInput[103]), .B(n25095), .C(vectorInput[95]), .D(
        n25080), .Z(n27289) );
    VMW_AO22 U509 ( .A(matrixInput[947]), .B(n25096), .C(matrixInput[939]), 
        .D(n25081), .Z(n26317) );
    VMW_AO22 U2057 ( .A(matrixInput[1397]), .B(n25096), .C(matrixInput[1389]), 
        .D(n25081), .Z(n25867) );
    VMW_AO22 U337 ( .A(vectorInput[86]), .B(n25095), .C(vectorInput[78]), .D(
        n25080), .Z(n27306) );
    VMW_AO22 U499 ( .A(matrixInput[956]), .B(n25096), .C(matrixInput[948]), 
        .D(n25081), .Z(n26308) );
    VMW_FD \matrixInput_reg[565]  ( .D(n26691), .CP(Clk), .Q(matrixInput[565])
         );
    VMW_AO22 U639 ( .A(matrixInput[829]), .B(n25096), .C(matrixInput[821]), 
        .D(n25081), .Z(n26435) );
    VMW_AO22 U1357 ( .A(matrixInput[2026]), .B(n25096), .C(matrixInput[2018]), 
        .D(n25081), .Z(n25238) );
    VMW_FD \matrixInput_reg[1372]  ( .D(n25884), .CP(Clk), .Q(matrixInput
        [1372]) );
    VMW_FD \matrixInput_reg[1042]  ( .D(n26214), .CP(Clk), .Q(matrixInput
        [1042]) );
    VMW_FD \matrixInput_reg[655]  ( .D(n26601), .CP(Clk), .Q(matrixInput[655])
         );
    VMW_AO22 U1546 ( .A(matrixInput[1857]), .B(n25096), .C(matrixInput[1849]), 
        .D(n25081), .Z(n25407) );
    VMW_AO22 U1934 ( .A(matrixInput[157]), .B(n25096), .C(matrixInput[149]), 
        .D(n25081), .Z(n27107) );
    VMW_OAI21 U2576 ( .A(n25132), .B(n25133), .C(n25091), .Z(n25138) );
    VMW_FD \matrixInput_reg[1358]  ( .D(n25898), .CP(Clk), .Q(matrixInput
        [1358]) );
    VMW_FD \matrixInput_reg[1341]  ( .D(n25915), .CP(Clk), .Q(matrixInput
        [1341]) );
    VMW_AO22 U868 ( .A(matrixInput[623]), .B(n25096), .C(matrixInput[615]), 
        .D(n25081), .Z(n26641) );
    VMW_AO22 U1040 ( .A(matrixInput[468]), .B(n25096), .C(matrixInput[460]), 
        .D(n25081), .Z(n26796) );
    VMW_AO22 U1370 ( .A(matrixInput[2014]), .B(n25096), .C(matrixInput[2006]), 
        .D(n25081), .Z(n25250) );
    VMW_AO22 U1561 ( .A(matrixInput[1843]), .B(n25096), .C(matrixInput[1835]), 
        .D(n25081), .Z(n25421) );
    VMW_AO22 U2367 ( .A(matrixInput[1117]), .B(n25096), .C(matrixInput[1109]), 
        .D(n25081), .Z(n26147) );
    VMW_FD \matrixInput_reg[556]  ( .D(n26700), .CP(Clk), .Q(matrixInput[556])
         );
    VMW_AO22 U1651 ( .A(matrixInput[1762]), .B(n25096), .C(matrixInput[1754]), 
        .D(n25081), .Z(n25502) );
    VMW_AO22 U1883 ( .A(matrixInput[1553]), .B(n25096), .C(matrixInput[1545]), 
        .D(n25081), .Z(n25711) );
    VMW_AO22 U1913 ( .A(matrixInput[1526]), .B(n25096), .C(matrixInput[1518]), 
        .D(n25081), .Z(n25738) );
    VMW_AO22 U2340 ( .A(matrixInput[1141]), .B(n25096), .C(matrixInput[1133]), 
        .D(n25081), .Z(n26123) );
    VMW_FD \matrixInput_reg[1666]  ( .D(n25590), .CP(Clk), .Q(matrixInput
        [1666]) );
    VMW_FD \matrixInput_reg[1565]  ( .D(n25691), .CP(Clk), .Q(matrixInput
        [1565]) );
    VMW_FD \matrixInput_reg[372]  ( .D(n26884), .CP(Clk), .Q(matrixInput[372])
         );
    VMW_AND3 U2551 ( .A(n25171), .B(n25172), .C(n25173), .Z(n25061) );
    VMW_FD \matrixInput_reg[2018]  ( .D(n25238), .CP(Clk), .Q(matrixInput
        [2018]) );
    VMW_FD \matrixInput_reg[2001]  ( .D(n25255), .CP(Clk), .Q(matrixInput
        [2001]) );
    VMW_FD \matrixInput_reg[1655]  ( .D(n25601), .CP(Clk), .Q(matrixInput
        [1655]) );
    VMW_AO22 U1153 ( .A(matrixInput[367]), .B(n25096), .C(matrixInput[359]), 
        .D(n25081), .Z(n26897) );
    VMW_AO22 U2070 ( .A(matrixInput[1385]), .B(n25096), .C(matrixInput[1377]), 
        .D(n25081), .Z(n25879) );
    VMW_FD \matrixInput_reg[2032]  ( .D(n25224), .CP(Clk), .Q(matrixInput
        [2032]) );
    VMW_AO22 U2163 ( .A(matrixInput[1301]), .B(n25096), .C(matrixInput[1293]), 
        .D(n25081), .Z(n25963) );
    VMW_FD \matrixInput_reg[1556]  ( .D(n25700), .CP(Clk), .Q(matrixInput
        [1556]) );
    VMW_FD \matrixInput_reg[1165]  ( .D(n26091), .CP(Clk), .Q(matrixInput
        [1165]) );
    VMW_FD \matrixInput_reg[772]  ( .D(n26484), .CP(Clk), .Q(matrixInput[772])
         );
    VMW_FD \matrixInput_reg[358]  ( .D(n26898), .CP(Clk), .Q(matrixInput[358])
         );
    VMW_FD \matrixInput_reg[341]  ( .D(n26915), .CP(Clk), .Q(matrixInput[341])
         );
    VMW_AO22 U1244 ( .A(matrixInput[285]), .B(n25096), .C(matrixInput[277]), 
        .D(n25081), .Z(n26979) );
    VMW_AO22 U1263 ( .A(matrixInput[33]), .B(n25096), .C(matrixInput[25]), .D(
        n25081), .Z(n27231) );
    VMW_AO22 U1742 ( .A(matrixInput[1680]), .B(n25096), .C(matrixInput[1672]), 
        .D(n25081), .Z(n25584) );
    VMW_AO22 U1800 ( .A(matrixInput[169]), .B(n25096), .C(matrixInput[161]), 
        .D(n25081), .Z(n27095) );
    VMW_AO22 U1990 ( .A(matrixInput[1457]), .B(n25096), .C(matrixInput[1449]), 
        .D(n25081), .Z(n25807) );
    VMW_AO22 U2253 ( .A(matrixInput[1219]), .B(n25096), .C(matrixInput[1211]), 
        .D(n25081), .Z(n26045) );
    VMW_AO22 U2442 ( .A(matrixInput[1049]), .B(n25096), .C(matrixInput[1041]), 
        .D(n25081), .Z(n26215) );
    VMW_FD \matrixInput_reg[1266]  ( .D(n25990), .CP(Clk), .Q(matrixInput
        [1266]) );
    VMW_FD \matrixInput_reg[471]  ( .D(n26785), .CP(Clk), .Q(matrixInput[471])
         );
    VMW_FD \matrixInput_reg[468]  ( .D(n26788), .CP(Clk), .Q(matrixInput[468])
         );
    VMW_FD \matrixInput_reg[1156]  ( .D(n26100), .CP(Clk), .Q(matrixInput
        [1156]) );
    VMW_FD \matrixInput_reg[758]  ( .D(n26498), .CP(Clk), .Q(matrixInput[758])
         );
    VMW_FD \matrixInput_reg[741]  ( .D(n26515), .CP(Clk), .Q(matrixInput[741])
         );
    VMW_FD \matrixInput_reg[1255]  ( .D(n26001), .CP(Clk), .Q(matrixInput
        [1255]) );
    VMW_FD \matrixInput_reg[442]  ( .D(n26814), .CP(Clk), .Q(matrixInput[442])
         );
    VMW_AO22 U1455 ( .A(matrixInput[1938]), .B(n25096), .C(matrixInput[1930]), 
        .D(n25081), .Z(n25326) );
    VMW_AO22 U1472 ( .A(matrixInput[1923]), .B(n25096), .C(matrixInput[1915]), 
        .D(n25081), .Z(n25341) );
    VMW_AO22 U1827 ( .A(matrixInput[1604]), .B(n25096), .C(matrixInput[1596]), 
        .D(n25081), .Z(n25660) );
    VMW_AO22 U2274 ( .A(matrixInput[1201]), .B(n25096), .C(matrixInput[1193]), 
        .D(n25081), .Z(n26063) );
    VMW_FD \matrixInput_reg[165]  ( .D(n27091), .CP(Clk), .Q(matrixInput[165])
         );
    VMW_AO22 U2465 ( .A(matrixInput[1028]), .B(n25096), .C(matrixInput[1020]), 
        .D(n25081), .Z(n26236) );
    VMW_FD \matrixInput_reg[1772]  ( .D(n25484), .CP(Clk), .Q(matrixInput
        [1772]) );
    VMW_FD \matrixInput_reg[1468]  ( .D(n25788), .CP(Clk), .Q(matrixInput
        [1468]) );
    VMW_FD \matrixInput_reg[266]  ( .D(n26990), .CP(Clk), .Q(matrixInput[266])
         );
    VMW_FD \matrixInput_reg[1471]  ( .D(n25785), .CP(Clk), .Q(matrixInput
        [1471]) );
    VMW_AO22 U1048 ( .A(matrixInput[461]), .B(n25096), .C(matrixInput[453]), 
        .D(n25081), .Z(n26803) );
    VMW_AO22 U1174 ( .A(matrixInput[41]), .B(n25096), .C(matrixInput[33]), .D(
        n25081), .Z(n27223) );
    VMW_AO22 U1765 ( .A(matrixInput[1659]), .B(n25096), .C(matrixInput[1651]), 
        .D(n25081), .Z(n25605) );
    VMW_AO22 U2144 ( .A(matrixInput[138]), .B(n25096), .C(matrixInput[130]), 
        .D(n25081), .Z(n27126) );
    VMW_FD \matrixInput_reg[1758]  ( .D(n25498), .CP(Clk), .Q(matrixInput
        [1758]) );
    VMW_FD \matrixInput_reg[1741]  ( .D(n25515), .CP(Clk), .Q(matrixInput
        [1741]) );
    VMW_FD \matrixInput_reg[156]  ( .D(n27100), .CP(Clk), .Q(matrixInput[156])
         );
    VMW_FD \matrixInput_reg[1442]  ( .D(n25814), .CP(Clk), .Q(matrixInput
        [1442]) );
    VMW_AO22 U1659 ( .A(matrixInput[1755]), .B(n25096), .C(matrixInput[1747]), 
        .D(n25081), .Z(n25509) );
    VMW_FD \matrixInput_reg[1836]  ( .D(n25420), .CP(Clk), .Q(matrixInput
        [1836]) );
    VMW_FD \matrixInput_reg[255]  ( .D(n27001), .CP(Clk), .Q(matrixInput[255])
         );
    VMW_AO22 U501 ( .A(matrixInput[954]), .B(n25096), .C(matrixInput[946]), 
        .D(n25081), .Z(n26310) );
    VMW_AO22 U526 ( .A(matrixInput[931]), .B(n25096), .C(matrixInput[923]), 
        .D(n25081), .Z(n26333) );
    VMW_AO22 U2078 ( .A(matrixInput[144]), .B(n25096), .C(matrixInput[136]), 
        .D(n25081), .Z(n27120) );
    VMW_AO22 U616 ( .A(matrixInput[850]), .B(n25096), .C(matrixInput[842]), 
        .D(n25081), .Z(n26414) );
    VMW_AO22 U786 ( .A(matrixInput[76]), .B(n25096), .C(matrixInput[68]), .D(
        n25081), .Z(n27188) );
    VMW_AO22 U954 ( .A(matrixInput[546]), .B(n25096), .C(matrixInput[538]), 
        .D(n25081), .Z(n26718) );
    VMW_AO22 U1378 ( .A(matrixInput[27]), .B(n25096), .C(matrixInput[19]), .D(
        n25081), .Z(n27237) );
    VMW_AO22 U1569 ( .A(matrixInput[1836]), .B(n25096), .C(matrixInput[1828]), 
        .D(n25081), .Z(n25428) );
    VMW_AO22 U2348 ( .A(matrixInput[1134]), .B(n25096), .C(matrixInput[1126]), 
        .D(n25081), .Z(n26130) );
    VMW_FD \matrixInput_reg[1805]  ( .D(n25451), .CP(Clk), .Q(matrixInput
        [1805]) );
    VMW_FD \matrixInput_reg[995]  ( .D(n26261), .CP(Clk), .Q(matrixInput[995])
         );
    VMW_AO22 U631 ( .A(matrixInput[837]), .B(n25096), .C(matrixInput[829]), 
        .D(n25081), .Z(n26427) );
    VMW_AO22 U2559 ( .A(cOutput[120]), .B(n25089), .C(cOutput[104]), .D(n25088
        ), .Z(n25181) );
    VMW_FD \matrixInput_reg[836]  ( .D(n26420), .CP(Clk), .Q(matrixInput[836])
         );
    VMW_FD \matrixInput_reg[76]  ( .D(n27180), .CP(Clk), .Q(matrixInput[76])
         );
    VMW_FD \matrixInput_reg[805]  ( .D(n26451), .CP(Clk), .Q(matrixInput[805])
         );
    VMW_AND2 U310 ( .A(Addr[2]), .B(n25092), .Z(n25091) );
    VMW_AO22 U491 ( .A(matrixInput[963]), .B(n25096), .C(matrixInput[955]), 
        .D(n25081), .Z(n26301) );
    VMW_AO22 U359 ( .A(vectorInput[66]), .B(n25095), .C(vectorInput[58]), .D(
        n25080), .Z(n27326) );
    VMW_AO22 U548 ( .A(matrixInput[911]), .B(n25096), .C(matrixInput[903]), 
        .D(n25081), .Z(n26353) );
    VMW_AO22 U973 ( .A(matrixInput[528]), .B(n25096), .C(matrixInput[520]), 
        .D(n25081), .Z(n26736) );
    VMW_AO22 U1001 ( .A(matrixInput[504]), .B(n25096), .C(matrixInput[496]), 
        .D(n25081), .Z(n26760) );
    VMW_AO22 U1191 ( .A(matrixInput[332]), .B(n25096), .C(matrixInput[324]), 
        .D(n25081), .Z(n26932) );
    VMW_AO22 U1331 ( .A(DataIn[1]), .B(n25096), .C(matrixInput[2041]), .D(
        n25081), .Z(n25215) );
    VMW_AO22 U1520 ( .A(matrixInput[1880]), .B(n25096), .C(matrixInput[1872]), 
        .D(n25081), .Z(n25384) );
    VMW_AO22 U1952 ( .A(matrixInput[1491]), .B(n25096), .C(matrixInput[1483]), 
        .D(n25081), .Z(n25773) );
    VMW_FD \matrixInput_reg[1995]  ( .D(n25261), .CP(Clk), .Q(matrixInput
        [1995]) );
    VMW_FD \matrixInput_reg[45]  ( .D(n27211), .CP(Clk), .Q(matrixInput[45])
         );
    VMW_FD \matrixInput_reg[1603]  ( .D(n25653), .CP(Clk), .Q(matrixInput
        [1603]) );
    VMW_FD \matrixInput_reg[1287]  ( .D(n25969), .CP(Clk), .Q(matrixInput
        [1287]) );
    VMW_FD \matrixInput_reg[490]  ( .D(n26766), .CP(Clk), .Q(matrixInput[490])
         );
    VMW_FD \matrixInput_reg[489]  ( .D(n26767), .CP(Clk), .Q(matrixInput[489])
         );
    VMW_AO22 U1610 ( .A(matrixInput[1799]), .B(n25096), .C(matrixInput[1791]), 
        .D(n25081), .Z(n25465) );
    VMW_AO22 U2291 ( .A(matrixInput[1186]), .B(n25096), .C(matrixInput[1178]), 
        .D(n25081), .Z(n26078) );
    VMW_AO22 U2301 ( .A(matrixInput[1177]), .B(n25096), .C(matrixInput[1169]), 
        .D(n25081), .Z(n26087) );
    VMW_FD \matrixInput_reg[793]  ( .D(n26463), .CP(Clk), .Q(matrixInput[793])
         );
    VMW_AO22 U2480 ( .A(matrixInput[1015]), .B(n25096), .C(matrixInput[1007]), 
        .D(n25081), .Z(n26249) );
    VMW_AO22 U2510 ( .A(cOutput[61]), .B(n25089), .C(cOutput[45]), .D(n25088), 
        .Z(n25122) );
    VMW_FD \matrixInput_reg[1519]  ( .D(n25737), .CP(Clk), .Q(matrixInput
        [1519]) );
    VMW_FD \matrixInput_reg[1500]  ( .D(n25756), .CP(Clk), .Q(matrixInput
        [1500]) );
    VMW_FD \matrixInput_reg[1184]  ( .D(n26072), .CP(Clk), .Q(matrixInput
        [1184]) );
    VMW_FD \matrixInput_reg[317]  ( .D(n26939), .CP(Clk), .Q(matrixInput[317])
         );
    VMW_AO22 U1780 ( .A(matrixInput[1646]), .B(n25096), .C(matrixInput[1638]), 
        .D(n25081), .Z(n25618) );
    VMW_AO22 U1026 ( .A(matrixInput[481]), .B(n25096), .C(matrixInput[473]), 
        .D(n25081), .Z(n26783) );
    VMW_AO22 U2031 ( .A(matrixInput[1419]), .B(n25096), .C(matrixInput[1411]), 
        .D(n25081), .Z(n25845) );
    VMW_FD \matrixInput_reg[1630]  ( .D(n25626), .CP(Clk), .Q(matrixInput
        [1630]) );
    VMW_FD \matrixInput_reg[1629]  ( .D(n25627), .CP(Clk), .Q(matrixInput
        [1629]) );
    VMW_FD \matrixInput_reg[1533]  ( .D(n25723), .CP(Clk), .Q(matrixInput
        [1533]) );
    VMW_FD \matrixInput_reg[324]  ( .D(n26932), .CP(Clk), .Q(matrixInput[324])
         );
    VMW_BUFIZ U2620 ( .A(n25195), .E(RD), .Z(\DataOut[12]1 ) );
    VMW_FD \matrixInput_reg[1014]  ( .D(n26242), .CP(Clk), .Q(matrixInput
        [1014]) );
    VMW_AO22 U1637 ( .A(matrixInput[1775]), .B(n25096), .C(matrixInput[1767]), 
        .D(n25081), .Z(n25489) );
    VMW_FD \matrixInput_reg[1793]  ( .D(n25463), .CP(Clk), .Q(matrixInput
        [1793]) );
    VMW_FD \matrixInput_reg[1490]  ( .D(n25766), .CP(Clk), .Q(matrixInput
        [1490]) );
    VMW_FD \matrixInput_reg[603]  ( .D(n26653), .CP(Clk), .Q(matrixInput[603])
         );
    VMW_FD \matrixInput_reg[287]  ( .D(n26969), .CP(Clk), .Q(matrixInput[287])
         );
    VMW_FD \matrixInput_reg[1489]  ( .D(n25767), .CP(Clk), .Q(matrixInput
        [1489]) );
    VMW_FD \matrixInput_reg[184]  ( .D(n27072), .CP(Clk), .Q(matrixInput[184])
         );
    VMW_FD \matrixInput_reg[1317]  ( .D(n25939), .CP(Clk), .Q(matrixInput
        [1317]) );
    VMW_AO22 U2186 ( .A(matrixInput[1280]), .B(n25096), .C(matrixInput[1272]), 
        .D(n25081), .Z(n25984) );
    VMW_INV U2607 ( .A(\holder[0] ), .Z(n25056) );
    VMW_FD \matrixInput_reg[500]  ( .D(n26756), .CP(Clk), .Q(matrixInput[500])
         );
    VMW_AO22 U453 ( .A(matrixInput[106]), .B(n25096), .C(matrixInput[98]), .D(
        n25081), .Z(n27158) );
    VMW_AO22 U474 ( .A(matrixInput[978]), .B(n25096), .C(matrixInput[970]), 
        .D(n25081), .Z(n26286) );
    VMW_AO22 U678 ( .A(matrixInput[795]), .B(n25096), .C(matrixInput[787]), 
        .D(n25081), .Z(n26469) );
    VMW_AO22 U1286 ( .A(matrixInput[247]), .B(n25096), .C(matrixInput[239]), 
        .D(n25081), .Z(n27017) );
    VMW_AO22 U1316 ( .A(matrixInput[219]), .B(n25096), .C(matrixInput[211]), 
        .D(n25081), .Z(n27045) );
    VMW_AO22 U1975 ( .A(matrixInput[1470]), .B(n25096), .C(matrixInput[1462]), 
        .D(n25081), .Z(n25794) );
    VMW_AO22 U2016 ( .A(matrixInput[1433]), .B(n25096), .C(matrixInput[1425]), 
        .D(n25081), .Z(n25831) );
    VMW_FD \matrixInput_reg[519]  ( .D(n26737), .CP(Clk), .Q(matrixInput[519])
         );
    VMW_AO22 U1497 ( .A(matrixInput[1901]), .B(n25096), .C(matrixInput[1893]), 
        .D(n25081), .Z(n25363) );
    VMW_FD \matrixInput_reg[629]  ( .D(n26627), .CP(Clk), .Q(matrixInput[629])
         );
    VMW_AO22 U1507 ( .A(matrixInput[1892]), .B(n25096), .C(matrixInput[1884]), 
        .D(n25081), .Z(n25372) );
    VMW_FD \matrixInput_reg[630]  ( .D(n26626), .CP(Clk), .Q(matrixInput[630])
         );
    VMW_FD \matrixInput_reg[1027]  ( .D(n26229), .CP(Clk), .Q(matrixInput
        [1027]) );
    VMW_FD \matrixInput_reg[533]  ( .D(n26723), .CP(Clk), .Q(matrixInput[533])
         );
    VMW_AO22 U744 ( .A(matrixInput[735]), .B(n25096), .C(matrixInput[727]), 
        .D(n25081), .Z(n26529) );
    VMW_AO22 U2326 ( .A(matrixInput[1154]), .B(n25096), .C(matrixInput[1146]), 
        .D(n25081), .Z(n26110) );
    VMW_AO22 U2537 ( .A(cOutput[58]), .B(n25089), .C(cOutput[42]), .D(n25088), 
        .Z(n25155) );
    VMW_FD \matrixInput_reg[1324]  ( .D(n25932), .CP(Clk), .Q(matrixInput
        [1324]) );
    VMW_FD \matrixInput_reg[947]  ( .D(n26309), .CP(Clk), .Q(matrixInput[947])
         );
    VMW_AO22 U1849 ( .A(matrixInput[1584]), .B(n25096), .C(matrixInput[1576]), 
        .D(n25081), .Z(n25680) );
    VMW_FD \vectorInput_reg[27]  ( .D(n27357), .CP(Clk), .Q(vectorInput[27])
         );
    VMW_AO22 U806 ( .A(matrixInput[679]), .B(n25096), .C(matrixInput[671]), 
        .D(n25081), .Z(n26585) );
    VMW_AO22 U996 ( .A(matrixInput[12]), .B(n25096), .C(matrixInput[4]), .D(
        n25081), .Z(n27252) );
    VMW_FD \matrixInput_reg[974]  ( .D(n26282), .CP(Clk), .Q(matrixInput[974])
         );
    VMW_FD \matrixInput_reg[1947]  ( .D(n25309), .CP(Clk), .Q(matrixInput
        [1947]) );
    VMW_FD \vectorInput_reg[14]  ( .D(n27370), .CP(Clk), .Q(vectorInput[14])
         );
    VMW_FD \matrixInput_reg[97]  ( .D(n27159), .CP(Clk), .Q(matrixInput[97])
         );
    VMW_AO22 U763 ( .A(matrixInput[78]), .B(n25096), .C(matrixInput[70]), .D(
        n25081), .Z(n27186) );
    VMW_AO22 U821 ( .A(matrixInput[666]), .B(n25096), .C(matrixInput[658]), 
        .D(n25081), .Z(n26598) );
    VMW_AO22 U1216 ( .A(matrixInput[309]), .B(n25096), .C(matrixInput[301]), 
        .D(n25081), .Z(n26955) );
    VMW_AO22 U1386 ( .A(matrixInput[2001]), .B(n25096), .C(matrixInput[1993]), 
        .D(n25081), .Z(n25263) );
    VMW_AO22 U1875 ( .A(matrixInput[1560]), .B(n25096), .C(matrixInput[1552]), 
        .D(n25081), .Z(n25704) );
    VMW_FD \matrixInput_reg[1974]  ( .D(n25282), .CP(Clk), .Q(matrixInput
        [1974]) );
    VMW_FD \matrixInput_reg[1037]  ( .D(n26219), .CP(Clk), .Q(matrixInput
        [1037]) );
    VMW_AO22 U1407 ( .A(matrixInput[1982]), .B(n25096), .C(matrixInput[1974]), 
        .D(n25081), .Z(n25282) );
    VMW_FD \matrixInput_reg[620]  ( .D(n26636), .CP(Clk), .Q(matrixInput[620])
         );
    VMW_AO22 U1597 ( .A(matrixInput[1810]), .B(n25096), .C(matrixInput[1802]), 
        .D(n25081), .Z(n25454) );
    VMW_FD \matrixInput_reg[639]  ( .D(n26617), .CP(Clk), .Q(matrixInput[639])
         );
    VMW_FD \matrixInput_reg[1334]  ( .D(n25922), .CP(Clk), .Q(matrixInput
        [1334]) );
    VMW_FD \holder_reg[1]  ( .D(n27391), .CP(Clk), .Q(\holder[1] ) );
    VMW_PULLDOWN U270 ( .Z(n25188) );
    VMW_PULLDOWN U277 ( .Z(n25195) );
    VMW_PULLDOWN U289 ( .Z(n25207) );
    VMW_AO22 U319 ( .A(vectorInput[102]), .B(n25095), .C(vectorInput[94]), .D(
        n25080), .Z(n27290) );
    VMW_AO22 U342 ( .A(vectorInput[81]), .B(n25095), .C(vectorInput[73]), .D(
        n25080), .Z(n27311) );
    VMW_AO22 U448 ( .A(matrixInput[1002]), .B(n25096), .C(matrixInput[994]), 
        .D(n25081), .Z(n26262) );
    VMW_AO22 U778 ( .A(matrixInput[705]), .B(n25096), .C(matrixInput[697]), 
        .D(n25081), .Z(n26559) );
    VMW_AO22 U2226 ( .A(matrixInput[1244]), .B(n25096), .C(matrixInput[1236]), 
        .D(n25081), .Z(n26020) );
    VMW_FD \matrixInput_reg[523]  ( .D(n26733), .CP(Clk), .Q(matrixInput[523])
         );
    VMW_AO22 U1126 ( .A(matrixInput[391]), .B(n25096), .C(matrixInput[383]), 
        .D(n25081), .Z(n26873) );
    VMW_AO22 U1737 ( .A(matrixInput[1685]), .B(n25096), .C(matrixInput[1677]), 
        .D(n25081), .Z(n25579) );
    VMW_AO22 U2437 ( .A(matrixInput[1054]), .B(n25096), .C(matrixInput[1046]), 
        .D(n25081), .Z(n26210) );
    VMW_FD \matrixInput_reg[613]  ( .D(n26643), .CP(Clk), .Q(matrixInput[613])
         );
    VMW_AO22 U2116 ( .A(matrixInput[1343]), .B(n25096), .C(matrixInput[1335]), 
        .D(n25081), .Z(n25921) );
    VMW_FD \matrixInput_reg[1783]  ( .D(n25473), .CP(Clk), .Q(matrixInput
        [1783]) );
    VMW_FD \matrixInput_reg[1499]  ( .D(n25757), .CP(Clk), .Q(matrixInput
        [1499]) );
    VMW_FD \matrixInput_reg[1004]  ( .D(n26252), .CP(Clk), .Q(matrixInput
        [1004]) );
    VMW_FD \matrixInput_reg[1480]  ( .D(n25776), .CP(Clk), .Q(matrixInput
        [1480]) );
    VMW_FD \matrixInput_reg[297]  ( .D(n26959), .CP(Clk), .Q(matrixInput[297])
         );
    VMW_FD \matrixInput_reg[509]  ( .D(n26747), .CP(Clk), .Q(matrixInput[509])
         );
    VMW_FD \matrixInput_reg[194]  ( .D(n27062), .CP(Clk), .Q(matrixInput[194])
         );
    VMW_AO22 U553 ( .A(matrixInput[97]), .B(n25096), .C(matrixInput[89]), .D(
        n25081), .Z(n27167) );
    VMW_AO22 U663 ( .A(matrixInput[15]), .B(n25096), .C(matrixInput[7]), .D(
        n25081), .Z(n27249) );
    VMW_AO22 U1091 ( .A(matrixInput[422]), .B(n25096), .C(matrixInput[414]), 
        .D(n25081), .Z(n26842) );
    VMW_AO22 U1101 ( .A(matrixInput[413]), .B(n25096), .C(matrixInput[405]), 
        .D(n25081), .Z(n26851) );
    VMW_AO22 U1680 ( .A(matrixInput[1736]), .B(n25096), .C(matrixInput[1728]), 
        .D(n25081), .Z(n25528) );
    VMW_AO22 U2086 ( .A(matrixInput[1370]), .B(n25096), .C(matrixInput[1362]), 
        .D(n25081), .Z(n25894) );
    VMW_FD \matrixInput_reg[510]  ( .D(n26746), .CP(Clk), .Q(matrixInput[510])
         );
    VMW_FD \matrixInput_reg[1307]  ( .D(n25949), .CP(Clk), .Q(matrixInput
        [1307]) );
    VMW_AO22 U1710 ( .A(matrixInput[1708]), .B(n25096), .C(matrixInput[1700]), 
        .D(n25081), .Z(n25556) );
    VMW_AO22 U1231 ( .A(matrixInput[297]), .B(n25096), .C(matrixInput[289]), 
        .D(n25081), .Z(n26967) );
    VMW_AO22 U1852 ( .A(matrixInput[1581]), .B(n25096), .C(matrixInput[1573]), 
        .D(n25081), .Z(n25683) );
    VMW_AO22 U2131 ( .A(matrixInput[1329]), .B(n25096), .C(matrixInput[1321]), 
        .D(n25081), .Z(n25935) );
    VMW_FD \matrixInput_reg[2047]  ( .D(n25209), .CP(Clk), .Q(matrixInput
        [2047]) );
    VMW_FD \matrixInput_reg[1639]  ( .D(n25617), .CP(Clk), .Q(matrixInput
        [1639]) );
    VMW_FD \matrixInput_reg[1620]  ( .D(n25636), .CP(Clk), .Q(matrixInput
        [1620]) );
    VMW_FD \matrixInput_reg[1523]  ( .D(n25733), .CP(Clk), .Q(matrixInput
        [1523]) );
    VMW_FD \matrixInput_reg[334]  ( .D(n26922), .CP(Clk), .Q(matrixInput[334])
         );
    VMW_FD \matrixInput_reg[1613]  ( .D(n25643), .CP(Clk), .Q(matrixInput
        [1613]) );
    VMW_AO22 U1420 ( .A(matrixInput[1970]), .B(n25096), .C(matrixInput[1962]), 
        .D(n25081), .Z(n25294) );
    VMW_AO22 U2201 ( .A(matrixInput[1267]), .B(n25096), .C(matrixInput[1259]), 
        .D(n25081), .Z(n25997) );
    VMW_AO22 U2391 ( .A(matrixInput[1096]), .B(n25096), .C(matrixInput[1088]), 
        .D(n25081), .Z(n26168) );
    VMW_FD \matrixInput_reg[1297]  ( .D(n25959), .CP(Clk), .Q(matrixInput
        [1297]) );
    VMW_FD \matrixInput_reg[499]  ( .D(n26757), .CP(Clk), .Q(matrixInput[499])
         );
    VMW_FD \matrixInput_reg[480]  ( .D(n26776), .CP(Clk), .Q(matrixInput[480])
         );
    VMW_AO22 U2410 ( .A(matrixInput[1078]), .B(n25096), .C(matrixInput[1070]), 
        .D(n25081), .Z(n26186) );
    VMW_FD \matrixInput_reg[1194]  ( .D(n26062), .CP(Clk), .Q(matrixInput
        [1194]) );
    VMW_OAI21 U2580 ( .A(n25143), .B(n25144), .C(n25091), .Z(n25149) );
    VMW_FD \matrixInput_reg[1964]  ( .D(n25292), .CP(Clk), .Q(matrixInput
        [1964]) );
    VMW_FD \matrixInput_reg[1510]  ( .D(n25746), .CP(Clk), .Q(matrixInput
        [1510]) );
    VMW_FD \matrixInput_reg[1509]  ( .D(n25747), .CP(Clk), .Q(matrixInput
        [1509]) );
    VMW_FD \matrixInput_reg[783]  ( .D(n26473), .CP(Clk), .Q(matrixInput[783])
         );
    VMW_FD \matrixInput_reg[307]  ( .D(n26949), .CP(Clk), .Q(matrixInput[307])
         );
    VMW_AO22 U365 ( .A(vectorInput[60]), .B(n25095), .C(vectorInput[52]), .D(
        n25080), .Z(n27332) );
    VMW_AO22 U921 ( .A(matrixInput[576]), .B(n25096), .C(matrixInput[568]), 
        .D(n25081), .Z(n26688) );
    VMW_FD \matrixInput_reg[1957]  ( .D(n25299), .CP(Clk), .Q(matrixInput
        [1957]) );
    VMW_FD \matrixInput_reg[87]  ( .D(n27169), .CP(Clk), .Q(matrixInput[87])
         );
    VMW_AO22 U380 ( .A(vectorInput[47]), .B(n25095), .C(vectorInput[39]), .D(
        n25080), .Z(n27345) );
    VMW_AO22 U401 ( .A(vectorInput[9]), .B(n25095), .C(vectorInput[1]), .D(
        n25080), .Z(n27383) );
    VMW_AO22 U574 ( .A(matrixInput[888]), .B(n25096), .C(matrixInput[880]), 
        .D(n25081), .Z(n26376) );
    VMW_AO22 U591 ( .A(matrixInput[873]), .B(n25096), .C(matrixInput[865]), 
        .D(n25081), .Z(n26391) );
    VMW_AO22 U644 ( .A(matrixInput[825]), .B(n25096), .C(matrixInput[817]), 
        .D(n25081), .Z(n26439) );
    VMW_AO22 U896 ( .A(matrixInput[598]), .B(n25096), .C(matrixInput[590]), 
        .D(n25081), .Z(n26666) );
    VMW_AO22 U906 ( .A(matrixInput[589]), .B(n25096), .C(matrixInput[581]), 
        .D(n25081), .Z(n26675) );
    VMW_FD \matrixInput_reg[964]  ( .D(n26292), .CP(Clk), .Q(matrixInput[964])
         );
    VMW_FD \matrixInput_reg[957]  ( .D(n26299), .CP(Clk), .Q(matrixInput[957])
         );
    VMW_AO22 U968 ( .A(matrixInput[533]), .B(n25096), .C(matrixInput[525]), 
        .D(n25081), .Z(n26731) );
    VMW_AO22 U1949 ( .A(matrixInput[1494]), .B(n25096), .C(matrixInput[1486]), 
        .D(n25081), .Z(n25770) );
    VMW_FD \vectorInput_reg[37]  ( .D(n27347), .CP(Clk), .Q(vectorInput[37])
         );
    VMW_AO22 U1053 ( .A(matrixInput[457]), .B(n25096), .C(matrixInput[449]), 
        .D(n25081), .Z(n26807) );
    VMW_AO22 U1074 ( .A(matrixInput[50]), .B(n25096), .C(matrixInput[42]), .D(
        n25081), .Z(n27214) );
    VMW_AO22 U2044 ( .A(matrixInput[21]), .B(n25096), .C(matrixInput[13]), .D(
        n25081), .Z(n27243) );
    VMW_FD \matrixInput_reg[1748]  ( .D(n25508), .CP(Clk), .Q(matrixInput
        [1748]) );
    VMW_FD \matrixInput_reg[146]  ( .D(n27110), .CP(Clk), .Q(matrixInput[146])
         );
    VMW_FD \matrixInput_reg[1751]  ( .D(n25505), .CP(Clk), .Q(matrixInput
        [1751]) );
    VMW_FD \matrixInput_reg[1452]  ( .D(n25804), .CP(Clk), .Q(matrixInput
        [1452]) );
    VMW_FD \matrixInput_reg[245]  ( .D(n27011), .CP(Clk), .Q(matrixInput[245])
         );
    VMW_AO22 U1344 ( .A(matrixInput[210]), .B(n25096), .C(matrixInput[202]), 
        .D(n25081), .Z(n27054) );
    VMW_AO22 U1665 ( .A(matrixInput[1749]), .B(n25096), .C(matrixInput[1741]), 
        .D(n25081), .Z(n25515) );
    VMW_AO22 U1927 ( .A(matrixInput[1513]), .B(n25096), .C(matrixInput[1505]), 
        .D(n25081), .Z(n25751) );
    VMW_AO22 U2374 ( .A(matrixInput[1110]), .B(n25096), .C(matrixInput[1102]), 
        .D(n25081), .Z(n26154) );
    VMW_OAI21 U2565 ( .A(n25101), .B(n25102), .C(n25093), .Z(n25107) );
    VMW_FD \matrixInput_reg[1762]  ( .D(n25494), .CP(Clk), .Q(matrixInput
        [1762]) );
    VMW_FD \matrixInput_reg[175]  ( .D(n27081), .CP(Clk), .Q(matrixInput[175])
         );
    VMW_FD \matrixInput_reg[1461]  ( .D(n25795), .CP(Clk), .Q(matrixInput
        [1461]) );
    VMW_AO22 U1363 ( .A(matrixInput[2020]), .B(n25096), .C(matrixInput[2012]), 
        .D(n25081), .Z(n25244) );
    VMW_AO22 U1555 ( .A(matrixInput[1848]), .B(n25096), .C(matrixInput[1840]), 
        .D(n25081), .Z(n25416) );
    VMW_FD \matrixInput_reg[1478]  ( .D(n25778), .CP(Clk), .Q(matrixInput
        [1478]) );
    VMW_AO22 U1572 ( .A(matrixInput[1833]), .B(n25096), .C(matrixInput[1825]), 
        .D(n25081), .Z(n25431) );
    VMW_AO22 U1890 ( .A(matrixInput[1547]), .B(n25096), .C(matrixInput[1539]), 
        .D(n25081), .Z(n25717) );
    VMW_AO22 U1900 ( .A(matrixInput[160]), .B(n25096), .C(matrixInput[152]), 
        .D(n25081), .Z(n27104) );
    VMW_AO22 U2353 ( .A(matrixInput[1129]), .B(n25096), .C(matrixInput[1121]), 
        .D(n25081), .Z(n26135) );
    VMW_FD \matrixInput_reg[276]  ( .D(n26980), .CP(Clk), .Q(matrixInput[276])
         );
    VMW_AND3 U2542 ( .A(n25160), .B(n25161), .C(n25162), .Z(n25064) );
    VMW_FD \matrixInput_reg[1245]  ( .D(n26011), .CP(Clk), .Q(matrixInput
        [1245]) );
    VMW_FD \matrixInput_reg[1146]  ( .D(n26110), .CP(Clk), .Q(matrixInput
        [1146]) );
    VMW_FD \matrixInput_reg[751]  ( .D(n26505), .CP(Clk), .Q(matrixInput[751])
         );
    VMW_FD \matrixInput_reg[748]  ( .D(n26508), .CP(Clk), .Q(matrixInput[748])
         );
    VMW_FD \matrixInput_reg[452]  ( .D(n26804), .CP(Clk), .Q(matrixInput[452])
         );
    VMW_AO22 U1642 ( .A(matrixInput[1770]), .B(n25096), .C(matrixInput[1762]), 
        .D(n25081), .Z(n25494) );
    VMW_AO22 U2063 ( .A(matrixInput[1391]), .B(n25096), .C(matrixInput[1383]), 
        .D(n25081), .Z(n25873) );
    VMW_FD \matrixInput_reg[1175]  ( .D(n26081), .CP(Clk), .Q(matrixInput
        [1175]) );
    VMW_FD \matrixInput_reg[762]  ( .D(n26494), .CP(Clk), .Q(matrixInput[762])
         );
    VMW_FD \matrixInput_reg[1276]  ( .D(n25980), .CP(Clk), .Q(matrixInput
        [1276]) );
    VMW_FD \matrixInput_reg[815]  ( .D(n26441), .CP(Clk), .Q(matrixInput[815])
         );
    VMW_FD \matrixInput_reg[478]  ( .D(n26778), .CP(Clk), .Q(matrixInput[478])
         );
    VMW_FD \matrixInput_reg[461]  ( .D(n26795), .CP(Clk), .Q(matrixInput[461])
         );
    VMW_AO22 U392 ( .A(vectorInput[36]), .B(n25095), .C(vectorInput[28]), .D(
        n25080), .Z(n27356) );
    VMW_AO22 U413 ( .A(DataIn[4]), .B(n25095), .C(vectorInput[124]), .D(n25080
        ), .Z(n27260) );
    VMW_AO22 U426 ( .A(vectorInput[120]), .B(n25095), .C(vectorInput[112]), 
        .D(n25080), .Z(n27272) );
    VMW_AO22 U686 ( .A(matrixInput[85]), .B(n25096), .C(matrixInput[77]), .D(
        n25081), .Z(n27179) );
    VMW_AO22 U716 ( .A(matrixInput[760]), .B(n25096), .C(matrixInput[752]), 
        .D(n25081), .Z(n26504) );
    VMW_AO22 U731 ( .A(matrixInput[747]), .B(n25096), .C(matrixInput[739]), 
        .D(n25081), .Z(n26517) );
    VMW_AO22 U873 ( .A(matrixInput[618]), .B(n25096), .C(matrixInput[610]), 
        .D(n25081), .Z(n26646) );
    VMW_FD \matrixInput_reg[1985]  ( .D(n25271), .CP(Clk), .Q(matrixInput
        [1985]) );
    VMW_FD \matrixInput_reg[55]  ( .D(n27201), .CP(Clk), .Q(matrixInput[55])
         );
    VMW_FD \matrixInput_reg[826]  ( .D(n26430), .CP(Clk), .Q(matrixInput[826])
         );
    VMW_FD \matrixInput_reg[66]  ( .D(n27190), .CP(Clk), .Q(matrixInput[66])
         );
    VMW_AO22 U1278 ( .A(matrixInput[254]), .B(n25096), .C(matrixInput[246]), 
        .D(n25081), .Z(n27010) );
    VMW_AO22 U1469 ( .A(matrixInput[1926]), .B(n25096), .C(matrixInput[1918]), 
        .D(n25081), .Z(n25338) );
    VMW_FD \matrixInput_reg[1815]  ( .D(n25441), .CP(Clk), .Q(matrixInput
        [1815]) );
    VMW_FD \matrixInput_reg[985]  ( .D(n26271), .CP(Clk), .Q(matrixInput[985])
         );
    VMW_AO22 U2248 ( .A(matrixInput[1224]), .B(n25096), .C(matrixInput[1216]), 
        .D(n25081), .Z(n26040) );
    VMW_AO22 U2459 ( .A(matrixInput[1034]), .B(n25096), .C(matrixInput[1026]), 
        .D(n25081), .Z(n26230) );
    VMW_AO22 U1148 ( .A(matrixInput[371]), .B(n25096), .C(matrixInput[363]), 
        .D(n25081), .Z(n26893) );
    VMW_FD \matrixInput_reg[1826]  ( .D(n25430), .CP(Clk), .Q(matrixInput
        [1826]) );
    VMW_AO22 U1759 ( .A(matrixInput[1665]), .B(n25096), .C(matrixInput[1657]), 
        .D(n25081), .Z(n25599) );
    VMW_AO22 U854 ( .A(matrixInput[636]), .B(n25096), .C(matrixInput[628]), 
        .D(n25081), .Z(n26628) );
    VMW_AO22 U2178 ( .A(matrixInput[135]), .B(n25096), .C(matrixInput[127]), 
        .D(n25081), .Z(n27129) );
    VMW_AO22 U861 ( .A(matrixInput[629]), .B(n25096), .C(matrixInput[621]), 
        .D(n25081), .Z(n26635) );
    VMW_AO22 U434 ( .A(vectorInput[113]), .B(n25095), .C(vectorInput[105]), 
        .D(n25080), .Z(n27279) );
    VMW_AO22 U583 ( .A(matrixInput[880]), .B(n25096), .C(matrixInput[872]), 
        .D(n25081), .Z(n26384) );
    VMW_AO22 U694 ( .A(matrixInput[780]), .B(n25096), .C(matrixInput[772]), 
        .D(n25081), .Z(n26484) );
    VMW_AO22 U723 ( .A(matrixInput[754]), .B(n25096), .C(matrixInput[746]), 
        .D(n25081), .Z(n26510) );
    VMW_FD \matrixInput_reg[1970]  ( .D(n25286), .CP(Clk), .Q(matrixInput
        [1970]) );
    VMW_FD \matrixInput_reg[1969]  ( .D(n25287), .CP(Clk), .Q(matrixInput
        [1969]) );
    VMW_FD \matrixInput_reg[1943]  ( .D(n25313), .CP(Clk), .Q(matrixInput
        [1943]) );
    VMW_FD \matrixInput_reg[93]  ( .D(n27163), .CP(Clk), .Q(matrixInput[93])
         );
    VMW_AO22 U1809 ( .A(matrixInput[1619]), .B(n25096), .C(matrixInput[1611]), 
        .D(n25081), .Z(n25645) );
    VMW_AO22 U1999 ( .A(matrixInput[1448]), .B(n25096), .C(matrixInput[1440]), 
        .D(n25081), .Z(n25816) );
    VMW_FD \vectorInput_reg[23]  ( .D(n27361), .CP(Clk), .Q(vectorInput[23])
         );
    VMW_AO22 U704 ( .A(matrixInput[771]), .B(n25096), .C(matrixInput[763]), 
        .D(n25081), .Z(n26493) );
    VMW_AO22 U846 ( .A(matrixInput[643]), .B(n25096), .C(matrixInput[635]), 
        .D(n25081), .Z(n26621) );
    VMW_FD \matrixInput_reg[969]  ( .D(n26287), .CP(Clk), .Q(matrixInput[969])
         );
    VMW_FD \matrixInput_reg[943]  ( .D(n26313), .CP(Clk), .Q(matrixInput[943])
         );
    VMW_FD \vectorInput_reg[10]  ( .D(n27374), .CP(Clk), .Q(vectorInput[10])
         );
    VMW_FD \matrixInput_reg[970]  ( .D(n26286), .CP(Clk), .Q(matrixInput[970])
         );
    VMW_AO22 U498 ( .A(matrixInput[957]), .B(n25096), .C(matrixInput[949]), 
        .D(n25081), .Z(n26307) );
    VMW_AO22 U508 ( .A(matrixInput[101]), .B(n25096), .C(matrixInput[93]), .D(
        n25081), .Z(n27163) );
    VMW_AO22 U2056 ( .A(matrixInput[146]), .B(n25096), .C(matrixInput[138]), 
        .D(n25081), .Z(n27118) );
    VMW_AO22 U350 ( .A(vectorInput[74]), .B(n25095), .C(vectorInput[66]), .D(
        n25080), .Z(n27318) );
    VMW_AO22 U638 ( .A(matrixInput[830]), .B(n25096), .C(matrixInput[822]), 
        .D(n25081), .Z(n26434) );
    VMW_AO22 U1066 ( .A(matrixInput[445]), .B(n25096), .C(matrixInput[437]), 
        .D(n25081), .Z(n26819) );
    VMW_AO22 U1677 ( .A(matrixInput[1738]), .B(n25096), .C(matrixInput[1730]), 
        .D(n25081), .Z(n25526) );
    VMW_FD \matrixInput_reg[1797]  ( .D(n25459), .CP(Clk), .Q(matrixInput
        [1797]) );
    VMW_FD \matrixInput_reg[1313]  ( .D(n25943), .CP(Clk), .Q(matrixInput
        [1313]) );
    VMW_FD \matrixInput_reg[504]  ( .D(n26752), .CP(Clk), .Q(matrixInput[504])
         );
    VMW_FD \matrixInput_reg[1494]  ( .D(n25762), .CP(Clk), .Q(matrixInput
        [1494]) );
    VMW_FD \matrixInput_reg[199]  ( .D(n27057), .CP(Clk), .Q(matrixInput[199])
         );
    VMW_FD \matrixInput_reg[180]  ( .D(n27076), .CP(Clk), .Q(matrixInput[180])
         );
    VMW_FD \matrixInput_reg[283]  ( .D(n26973), .CP(Clk), .Q(matrixInput[283])
         );
    VMW_FD \matrixInput_reg[607]  ( .D(n26649), .CP(Clk), .Q(matrixInput[607])
         );
    VMW_AO22 U2366 ( .A(matrixInput[118]), .B(n25096), .C(matrixInput[110]), 
        .D(n25081), .Z(n27146) );
    VMW_FD \matrixInput_reg[1339]  ( .D(n25917), .CP(Clk), .Q(matrixInput
        [1339]) );
    VMW_FD \matrixInput_reg[1010]  ( .D(n26246), .CP(Clk), .Q(matrixInput
        [1010]) );
    VMW_FD \matrixInput_reg[1009]  ( .D(n26247), .CP(Clk), .Q(matrixInput
        [1009]) );
    VMW_FD \matrixInput_reg[1320]  ( .D(n25936), .CP(Clk), .Q(matrixInput
        [1320]) );
    VMW_FD \matrixInput_reg[537]  ( .D(n26719), .CP(Clk), .Q(matrixInput[537])
         );
    VMW_AO22 U671 ( .A(matrixInput[801]), .B(n25096), .C(matrixInput[793]), 
        .D(n25081), .Z(n26463) );
    VMW_AO22 U1041 ( .A(matrixInput[53]), .B(n25096), .C(matrixInput[45]), .D(
        n25081), .Z(n27211) );
    VMW_AO22 U1356 ( .A(matrixInput[2027]), .B(n25096), .C(matrixInput[2019]), 
        .D(n25081), .Z(n25237) );
    VMW_AO22 U1547 ( .A(matrixInput[1856]), .B(n25096), .C(matrixInput[1848]), 
        .D(n25081), .Z(n25408) );
    VMW_OAI21 U2577 ( .A(n25134), .B(n25135), .C(n25093), .Z(n25140) );
    VMW_FD \matrixInput_reg[1023]  ( .D(n26233), .CP(Clk), .Q(matrixInput
        [1023]) );
    VMW_FD \matrixInput_reg[634]  ( .D(n26622), .CP(Clk), .Q(matrixInput[634])
         );
    VMW_AO22 U1371 ( .A(matrixInput[2013]), .B(n25096), .C(matrixInput[2005]), 
        .D(n25081), .Z(n25251) );
    VMW_AO22 U1935 ( .A(matrixInput[1507]), .B(n25096), .C(matrixInput[1499]), 
        .D(n25081), .Z(n25757) );
    VMW_AO22 U2341 ( .A(matrixInput[1140]), .B(n25096), .C(matrixInput[1132]), 
        .D(n25081), .Z(n26124) );
    VMW_AO22 U2550 ( .A(cOutput[121]), .B(n25089), .C(cOutput[105]), .D(n25088
        ), .Z(n25170) );
    VMW_FD \matrixInput_reg[1504]  ( .D(n25752), .CP(Clk), .Q(matrixInput
        [1504]) );
    VMW_FD \matrixInput_reg[313]  ( .D(n26943), .CP(Clk), .Q(matrixInput[313])
         );
    VMW_FD \matrixInput_reg[1180]  ( .D(n26076), .CP(Clk), .Q(matrixInput
        [1180]) );
    VMW_FD \matrixInput_reg[1199]  ( .D(n26057), .CP(Clk), .Q(matrixInput
        [1199]) );
    VMW_FD \matrixInput_reg[797]  ( .D(n26459), .CP(Clk), .Q(matrixInput[797])
         );
    VMW_AO22 U1560 ( .A(matrixInput[1844]), .B(n25096), .C(matrixInput[1836]), 
        .D(n25081), .Z(n25420) );
    VMW_AO22 U1882 ( .A(matrixInput[1554]), .B(n25096), .C(matrixInput[1546]), 
        .D(n25081), .Z(n25710) );
    VMW_FD \matrixInput_reg[1283]  ( .D(n25973), .CP(Clk), .Q(matrixInput
        [1283]) );
    VMW_FD \matrixInput_reg[494]  ( .D(n26762), .CP(Clk), .Q(matrixInput[494])
         );
    VMW_AO22 U1912 ( .A(matrixInput[1527]), .B(n25096), .C(matrixInput[1519]), 
        .D(n25081), .Z(n25737) );
    VMW_AO22 U2071 ( .A(matrixInput[1384]), .B(n25096), .C(matrixInput[1376]), 
        .D(n25081), .Z(n25880) );
    VMW_FD \matrixInput_reg[1607]  ( .D(n25649), .CP(Clk), .Q(matrixInput
        [1607]) );
    VMW_FD \matrixInput_reg[1634]  ( .D(n25622), .CP(Clk), .Q(matrixInput
        [1634]) );
    VMW_FD \matrixInput_reg[1537]  ( .D(n25719), .CP(Clk), .Q(matrixInput
        [1537]) );
    VMW_FD \matrixInput_reg[339]  ( .D(n26917), .CP(Clk), .Q(matrixInput[339])
         );
    VMW_FD \matrixInput_reg[320]  ( .D(n26936), .CP(Clk), .Q(matrixInput[320])
         );
    VMW_AO22 U1650 ( .A(matrixInput[1763]), .B(n25096), .C(matrixInput[1755]), 
        .D(n25081), .Z(n25501) );
    VMW_AO22 U933 ( .A(matrixInput[565]), .B(n25096), .C(matrixInput[557]), 
        .D(n25081), .Z(n26699) );
    VMW_FD \matrixInput_reg[1991]  ( .D(n25265), .CP(Clk), .Q(matrixInput
        [1991]) );
    VMW_FD \matrixInput_reg[832]  ( .D(n26424), .CP(Clk), .Q(matrixInput[832])
         );
    VMW_FD \matrixInput_reg[72]  ( .D(n27184), .CP(Clk), .Q(matrixInput[72])
         );
    VMW_FD \matrixInput_reg[58]  ( .D(n27198), .CP(Clk), .Q(matrixInput[58])
         );
    VMW_FD \matrixInput_reg[1988]  ( .D(n25268), .CP(Clk), .Q(matrixInput
        [1988]) );
    VMW_FD \matrixInput_reg[41]  ( .D(n27215), .CP(Clk), .Q(matrixInput[41])
         );
    VMW_AO22 U377 ( .A(vectorInput[49]), .B(n25095), .C(vectorInput[41]), .D(
        n25080), .Z(n27343) );
    VMW_AO22 U541 ( .A(matrixInput[98]), .B(n25096), .C(matrixInput[90]), .D(
        n25081), .Z(n27166) );
    VMW_AO22 U566 ( .A(matrixInput[896]), .B(n25096), .C(matrixInput[888]), 
        .D(n25081), .Z(n26368) );
    VMW_AO22 U884 ( .A(matrixInput[608]), .B(n25096), .C(matrixInput[600]), 
        .D(n25081), .Z(n26656) );
    VMW_AO22 U914 ( .A(matrixInput[582]), .B(n25096), .C(matrixInput[574]), 
        .D(n25081), .Z(n26682) );
    VMW_FD \matrixInput_reg[818]  ( .D(n26438), .CP(Clk), .Q(matrixInput[818])
         );
    VMW_FD \matrixInput_reg[801]  ( .D(n26455), .CP(Clk), .Q(matrixInput[801])
         );
    VMW_BUFIZ U2629 ( .A(n25202), .E(RD), .Z(\DataOut[24]1 ) );
    VMW_AO22 U656 ( .A(matrixInput[814]), .B(n25096), .C(matrixInput[806]), 
        .D(n25081), .Z(n26450) );
    VMW_AO22 U1008 ( .A(matrixInput[56]), .B(n25096), .C(matrixInput[48]), .D(
        n25081), .Z(n27208) );
    VMW_AO22 U1789 ( .A(matrixInput[170]), .B(n25096), .C(matrixInput[162]), 
        .D(n25081), .Z(n27094) );
    VMW_AO22 U2038 ( .A(matrixInput[1413]), .B(n25096), .C(matrixInput[1405]), 
        .D(n25081), .Z(n25851) );
    VMW_AO22 U1198 ( .A(matrixInput[326]), .B(n25096), .C(matrixInput[318]), 
        .D(n25081), .Z(n26938) );
    VMW_AO22 U1619 ( .A(matrixInput[1791]), .B(n25096), .C(matrixInput[1783]), 
        .D(n25081), .Z(n25473) );
    VMW_AO22 U2298 ( .A(matrixInput[1179]), .B(n25096), .C(matrixInput[1171]), 
        .D(n25081), .Z(n26085) );
    VMW_FD \matrixInput_reg[1832]  ( .D(n25424), .CP(Clk), .Q(matrixInput
        [1832]) );
    VMW_FD \matrixInput_reg[991]  ( .D(n26265), .CP(Clk), .Q(matrixInput[991])
         );
    VMW_AO22 U756 ( .A(matrixInput[724]), .B(n25096), .C(matrixInput[716]), 
        .D(n25081), .Z(n26540) );
    VMW_AO22 U828 ( .A(matrixInput[659]), .B(n25096), .C(matrixInput[651]), 
        .D(n25081), .Z(n26605) );
    VMW_AO22 U1134 ( .A(matrixInput[384]), .B(n25096), .C(matrixInput[376]), 
        .D(n25081), .Z(n26880) );
    VMW_AO22 U1204 ( .A(matrixInput[320]), .B(n25096), .C(matrixInput[312]), 
        .D(n25081), .Z(n26944) );
    VMW_AO22 U1338 ( .A(matrixInput[2043]), .B(n25096), .C(matrixInput[2035]), 
        .D(n25081), .Z(n25221) );
    VMW_AO22 U2308 ( .A(matrixInput[1170]), .B(n25096), .C(matrixInput[1162]), 
        .D(n25081), .Z(n26094) );
    VMW_AO22 U2519 ( .A(cOutput[60]), .B(n25089), .C(cOutput[44]), .D(n25088), 
        .Z(n25133) );
    VMW_FD \matrixInput_reg[988]  ( .D(n26268), .CP(Clk), .Q(matrixInput[988])
         );
    VMW_AO22 U2489 ( .A(cOutput[23]), .B(n25087), .C(cOutput[7]), .D(n25084), 
        .Z(n25097) );
    VMW_FD \matrixInput_reg[1818]  ( .D(n25438), .CP(Clk), .Q(matrixInput
        [1818]) );
    VMW_FD \matrixInput_reg[1801]  ( .D(n25455), .CP(Clk), .Q(matrixInput
        [1801]) );
    VMW_AO22 U1529 ( .A(matrixInput[1872]), .B(n25096), .C(matrixInput[1864]), 
        .D(n25081), .Z(n25392) );
    VMW_FD \matrixInput_reg[1475]  ( .D(n25781), .CP(Clk), .Q(matrixInput
        [1475]) );
    VMW_AO22 U1394 ( .A(matrixInput[1994]), .B(n25096), .C(matrixInput[1986]), 
        .D(n25081), .Z(n25270) );
    VMW_AO22 U1585 ( .A(matrixInput[1821]), .B(n25096), .C(matrixInput[1813]), 
        .D(n25081), .Z(n25443) );
    VMW_AO22 U1415 ( .A(matrixInput[1975]), .B(n25096), .C(matrixInput[1967]), 
        .D(n25081), .Z(n25289) );
    VMW_AO22 U1867 ( .A(matrixInput[163]), .B(n25096), .C(matrixInput[155]), 
        .D(n25081), .Z(n27101) );
    VMW_FD \matrixInput_reg[262]  ( .D(n26994), .CP(Clk), .Q(matrixInput[262])
         );
    VMW_AO22 U2234 ( .A(matrixInput[1237]), .B(n25096), .C(matrixInput[1229]), 
        .D(n25081), .Z(n26027) );
    VMW_AO22 U2425 ( .A(matrixInput[1065]), .B(n25096), .C(matrixInput[1057]), 
        .D(n25081), .Z(n26199) );
    VMW_FD \matrixInput_reg[1776]  ( .D(n25480), .CP(Clk), .Q(matrixInput
        [1776]) );
    VMW_FD \matrixInput_reg[1446]  ( .D(n25810), .CP(Clk), .Q(matrixInput
        [1446]) );
    VMW_FD \matrixInput_reg[251]  ( .D(n27005), .CP(Clk), .Q(matrixInput[251])
         );
    VMW_FD \matrixInput_reg[178]  ( .D(n27078), .CP(Clk), .Q(matrixInput[178])
         );
    VMW_FD \matrixInput_reg[161]  ( .D(n27095), .CP(Clk), .Q(matrixInput[161])
         );
    VMW_FD \matrixInput_reg[248]  ( .D(n27008), .CP(Clk), .Q(matrixInput[248])
         );
    VMW_AO22 U1725 ( .A(matrixInput[1696]), .B(n25096), .C(matrixInput[1688]), 
        .D(n25081), .Z(n25568) );
    VMW_AO22 U2094 ( .A(matrixInput[1363]), .B(n25096), .C(matrixInput[1355]), 
        .D(n25081), .Z(n25901) );
    VMW_FD \matrixInput_reg[152]  ( .D(n27104), .CP(Clk), .Q(matrixInput[152])
         );
    VMW_AO22 U2104 ( .A(matrixInput[1354]), .B(n25096), .C(matrixInput[1346]), 
        .D(n25081), .Z(n25910) );
    VMW_FD \matrixInput_reg[1745]  ( .D(n25511), .CP(Clk), .Q(matrixInput
        [1745]) );
    VMW_AO22 U1083 ( .A(matrixInput[429]), .B(n25096), .C(matrixInput[421]), 
        .D(n25081), .Z(n26835) );
    VMW_AO22 U1702 ( .A(matrixInput[1716]), .B(n25096), .C(matrixInput[1708]), 
        .D(n25081), .Z(n25548) );
    VMW_FD \matrixInput_reg[1262]  ( .D(n25994), .CP(Clk), .Q(matrixInput
        [1262]) );
    VMW_FD \matrixInput_reg[475]  ( .D(n26781), .CP(Clk), .Q(matrixInput[475])
         );
    VMW_AO22 U1113 ( .A(matrixInput[403]), .B(n25096), .C(matrixInput[395]), 
        .D(n25081), .Z(n26861) );
    VMW_AO22 U1692 ( .A(matrixInput[1725]), .B(n25096), .C(matrixInput[1717]), 
        .D(n25081), .Z(n25539) );
    VMW_AO22 U1223 ( .A(matrixInput[304]), .B(n25096), .C(matrixInput[296]), 
        .D(n25081), .Z(n26960) );
    VMW_AO22 U1432 ( .A(matrixInput[1959]), .B(n25096), .C(matrixInput[1951]), 
        .D(n25081), .Z(n25305) );
    VMW_AO22 U2123 ( .A(matrixInput[1337]), .B(n25096), .C(matrixInput[1329]), 
        .D(n25081), .Z(n25927) );
    VMW_FD \matrixInput_reg[1178]  ( .D(n26078), .CP(Clk), .Q(matrixInput
        [1178]) );
    VMW_FD \matrixInput_reg[1161]  ( .D(n26095), .CP(Clk), .Q(matrixInput
        [1161]) );
    VMW_FD \matrixInput_reg[776]  ( .D(n26480), .CP(Clk), .Q(matrixInput[776])
         );
    VMW_AO22 U1840 ( .A(matrixInput[1592]), .B(n25096), .C(matrixInput[1584]), 
        .D(n25081), .Z(n25672) );
    VMW_FD \matrixInput_reg[1251]  ( .D(n26005), .CP(Clk), .Q(matrixInput
        [1251]) );
    VMW_FD \matrixInput_reg[446]  ( .D(n26810), .CP(Clk), .Q(matrixInput[446])
         );
    VMW_AO22 U2208 ( .A(matrixInput[1260]), .B(n25096), .C(matrixInput[1252]), 
        .D(n25081), .Z(n26004) );
    VMW_AO22 U2213 ( .A(matrixInput[1256]), .B(n25096), .C(matrixInput[1248]), 
        .D(n25081), .Z(n26008) );
    VMW_FD \matrixInput_reg[1248]  ( .D(n26008), .CP(Clk), .Q(matrixInput
        [1248]) );
    VMW_FD \matrixInput_reg[1152]  ( .D(n26104), .CP(Clk), .Q(matrixInput
        [1152]) );
    VMW_FD \matrixInput_reg[745]  ( .D(n26511), .CP(Clk), .Q(matrixInput[745])
         );
    VMW_AO22 U2383 ( .A(matrixInput[1103]), .B(n25096), .C(matrixInput[1095]), 
        .D(n25081), .Z(n26161) );
    VMW_OAI21 U2592 ( .A(n25176), .B(n25177), .C(n25091), .Z(n25182) );
    VMW_AO22 U2402 ( .A(matrixInput[1086]), .B(n25096), .C(matrixInput[1078]), 
        .D(n25081), .Z(n26178) );
    VMW_FD \matrixInput_reg[998]  ( .D(n26258), .CP(Clk), .Q(matrixInput[998])
         );
    VMW_AO22 U2398 ( .A(matrixInput[1089]), .B(n25096), .C(matrixInput[1081]), 
        .D(n25081), .Z(n26175) );
    VMW_OAI21 U2589 ( .A(n25167), .B(n25168), .C(n25093), .Z(n25173) );
    VMW_FD \matrixInput_reg[981]  ( .D(n26275), .CP(Clk), .Q(matrixInput[981])
         );
    VMW_AO22 U814 ( .A(matrixInput[672]), .B(n25096), .C(matrixInput[664]), 
        .D(n25081), .Z(n26592) );
    VMW_AO22 U984 ( .A(matrixInput[518]), .B(n25096), .C(matrixInput[510]), 
        .D(n25081), .Z(n26746) );
    VMW_AO22 U1238 ( .A(matrixInput[290]), .B(n25096), .C(matrixInput[282]), 
        .D(n25081), .Z(n26974) );
    VMW_AO22 U1429 ( .A(matrixInput[1962]), .B(n25096), .C(matrixInput[1954]), 
        .D(n25081), .Z(n25302) );
    VMW_AO22 U2419 ( .A(matrixInput[1070]), .B(n25096), .C(matrixInput[1062]), 
        .D(n25081), .Z(n26194) );
    VMW_FD \matrixInput_reg[1811]  ( .D(n25445), .CP(Clk), .Q(matrixInput
        [1811]) );
    VMW_FD \matrixInput_reg[1808]  ( .D(n25448), .CP(Clk), .Q(matrixInput
        [1808]) );
    VMW_PULLUP U292 ( .Z(Logic11) );
    VMW_AND4 U302 ( .A(RD), .B(n164), .C(n25080), .D(n25081), .Z(n25055) );
    VMW_AO22 U325 ( .A(vectorInput[97]), .B(n25095), .C(vectorInput[89]), .D(
        n25080), .Z(n27295) );
    VMW_AO22 U441 ( .A(matrixInput[17]), .B(n25096), .C(matrixInput[9]), .D(
        n25081), .Z(n27247) );
    VMW_AO22 U466 ( .A(matrixInput[986]), .B(n25096), .C(matrixInput[978]), 
        .D(n25081), .Z(n26278) );
    VMW_AO22 U2138 ( .A(matrixInput[1323]), .B(n25096), .C(matrixInput[1315]), 
        .D(n25081), .Z(n25941) );
    VMW_AO22 U833 ( .A(matrixInput[655]), .B(n25096), .C(matrixInput[647]), 
        .D(n25081), .Z(n26609) );
    VMW_AO22 U1098 ( .A(matrixInput[416]), .B(n25096), .C(matrixInput[408]), 
        .D(n25081), .Z(n26848) );
    VMW_AO22 U1719 ( .A(matrixInput[1701]), .B(n25096), .C(matrixInput[1693]), 
        .D(n25081), .Z(n25563) );
    VMW_AO22 U1108 ( .A(matrixInput[47]), .B(n25096), .C(matrixInput[39]), .D(
        n25081), .Z(n27217) );
    VMW_AO22 U1689 ( .A(matrixInput[179]), .B(n25096), .C(matrixInput[171]), 
        .D(n25081), .Z(n27085) );
    VMW_FD \matrixInput_reg[1822]  ( .D(n25434), .CP(Clk), .Q(matrixInput
        [1822]) );
    VMW_FD \matrixInput_reg[1998]  ( .D(n25258), .CP(Clk), .Q(matrixInput
        [1998]) );
    VMW_FD \matrixInput_reg[1981]  ( .D(n25275), .CP(Clk), .Q(matrixInput
        [1981]) );
    VMW_FD \matrixInput_reg[51]  ( .D(n27205), .CP(Clk), .Q(matrixInput[51])
         );
    VMW_FD \matrixInput_reg[48]  ( .D(n27208), .CP(Clk), .Q(matrixInput[48])
         );
    VMW_AO22 U534 ( .A(matrixInput[924]), .B(n25096), .C(matrixInput[916]), 
        .D(n25081), .Z(n26340) );
    VMW_AO22 U771 ( .A(matrixInput[710]), .B(n25096), .C(matrixInput[702]), 
        .D(n25081), .Z(n26554) );
    VMW_FD \matrixInput_reg[811]  ( .D(n26445), .CP(Clk), .Q(matrixInput[811])
         );
    VMW_FD \matrixInput_reg[808]  ( .D(n26448), .CP(Clk), .Q(matrixInput[808])
         );
    VMW_AO22 U928 ( .A(matrixInput[569]), .B(n25096), .C(matrixInput[561]), 
        .D(n25081), .Z(n26695) );
    VMW_AO22 U1013 ( .A(matrixInput[493]), .B(n25096), .C(matrixInput[485]), 
        .D(n25081), .Z(n26771) );
    VMW_AO22 U1323 ( .A(matrixInput[213]), .B(n25096), .C(matrixInput[205]), 
        .D(n25081), .Z(n27051) );
    VMW_FD \matrixInput_reg[822]  ( .D(n26434), .CP(Clk), .Q(matrixInput[822])
         );
    VMW_FD \matrixInput_reg[62]  ( .D(n27194), .CP(Clk), .Q(matrixInput[62])
         );
    VMW_AO22 U1532 ( .A(matrixInput[1869]), .B(n25096), .C(matrixInput[1861]), 
        .D(n25081), .Z(n25395) );
    VMW_AO22 U1792 ( .A(matrixInput[1635]), .B(n25096), .C(matrixInput[1627]), 
        .D(n25081), .Z(n25629) );
    VMW_AO22 U1940 ( .A(matrixInput[1502]), .B(n25096), .C(matrixInput[1494]), 
        .D(n25081), .Z(n25762) );
    VMW_FD \matrixInput_reg[1258]  ( .D(n25998), .CP(Clk), .Q(matrixInput
        [1258]) );
    VMW_AO22 U2283 ( .A(matrixInput[1193]), .B(n25096), .C(matrixInput[1185]), 
        .D(n25081), .Z(n26071) );
    VMW_FD \matrixInput_reg[1241]  ( .D(n26015), .CP(Clk), .Q(matrixInput
        [1241]) );
    VMW_FD \matrixInput_reg[1142]  ( .D(n26114), .CP(Clk), .Q(matrixInput
        [1142]) );
    VMW_FD \matrixInput_reg[456]  ( .D(n26800), .CP(Clk), .Q(matrixInput[456])
         );
    VMW_FD \matrixInput_reg[755]  ( .D(n26501), .CP(Clk), .Q(matrixInput[755])
         );
    VMW_AO22 U2313 ( .A(matrixInput[1166]), .B(n25096), .C(matrixInput[1158]), 
        .D(n25081), .Z(n26098) );
    VMW_AO22 U2502 ( .A(cOutput[86]), .B(n25087), .C(cOutput[70]), .D(n25084), 
        .Z(n25112) );
    VMW_AO22 U2492 ( .A(cOutput[63]), .B(n25089), .C(cOutput[47]), .D(n25088), 
        .Z(n25100) );
    VMW_FD \matrixInput_reg[1272]  ( .D(n25984), .CP(Clk), .Q(matrixInput
        [1272]) );
    VMW_FD \matrixInput_reg[465]  ( .D(n26791), .CP(Clk), .Q(matrixInput[465])
         );
    VMW_AO22 U1034 ( .A(matrixInput[474]), .B(n25096), .C(matrixInput[466]), 
        .D(n25081), .Z(n26790) );
    VMW_AO22 U1183 ( .A(matrixInput[339]), .B(n25096), .C(matrixInput[331]), 
        .D(n25081), .Z(n26925) );
    VMW_AO22 U1602 ( .A(matrixInput[1807]), .B(n25096), .C(matrixInput[1799]), 
        .D(n25081), .Z(n25457) );
    VMW_AO22 U1625 ( .A(matrixInput[1786]), .B(n25096), .C(matrixInput[1778]), 
        .D(n25081), .Z(n25478) );
    VMW_AO22 U2023 ( .A(matrixInput[1427]), .B(n25096), .C(matrixInput[1419]), 
        .D(n25081), .Z(n25837) );
    VMW_BUFIZ U2632 ( .A(n25204), .E(RD), .Z(\DataOut[15]1 ) );
    VMW_FD \matrixInput_reg[1171]  ( .D(n26085), .CP(Clk), .Q(matrixInput
        [1171]) );
    VMW_FD \matrixInput_reg[766]  ( .D(n26490), .CP(Clk), .Q(matrixInput[766])
         );
    VMW_FD \matrixInput_reg[1168]  ( .D(n26088), .CP(Clk), .Q(matrixInput
        [1168]) );
    VMW_FD \matrixInput_reg[1456]  ( .D(n25800), .CP(Clk), .Q(matrixInput
        [1456]) );
    VMW_AO22 U2004 ( .A(matrixInput[1444]), .B(n25096), .C(matrixInput[1436]), 
        .D(n25081), .Z(n25820) );
    VMW_FD \matrixInput_reg[258]  ( .D(n26998), .CP(Clk), .Q(matrixInput[258])
         );
    VMW_FD \matrixInput_reg[241]  ( .D(n27015), .CP(Clk), .Q(matrixInput[241])
         );
    VMW_AO22 U2194 ( .A(matrixInput[1273]), .B(n25096), .C(matrixInput[1265]), 
        .D(n25081), .Z(n25991) );
    VMW_BUFIZ U2615 ( .A(\holder[4] ), .E(RD), .Z(\DataOut[4]1 ) );
    VMW_FD \matrixInput_reg[1755]  ( .D(n25501), .CP(Clk), .Q(matrixInput
        [1755]) );
    VMW_FD \matrixInput_reg[142]  ( .D(n27114), .CP(Clk), .Q(matrixInput[142])
         );
    VMW_AO22 U946 ( .A(matrixInput[553]), .B(n25096), .C(matrixInput[545]), 
        .D(n25081), .Z(n26711) );
    VMW_AO22 U1294 ( .A(matrixInput[239]), .B(n25096), .C(matrixInput[231]), 
        .D(n25081), .Z(n27025) );
    VMW_FD \matrixInput_reg[272]  ( .D(n26984), .CP(Clk), .Q(matrixInput[272])
         );
    VMW_AO22 U1304 ( .A(matrixInput[230]), .B(n25096), .C(matrixInput[222]), 
        .D(n25081), .Z(n27034) );
    VMW_AO22 U1515 ( .A(matrixInput[1885]), .B(n25096), .C(matrixInput[1877]), 
        .D(n25081), .Z(n25379) );
    VMW_FD \matrixInput_reg[1465]  ( .D(n25791), .CP(Clk), .Q(matrixInput
        [1465]) );
    VMW_AO22 U1485 ( .A(matrixInput[1911]), .B(n25096), .C(matrixInput[1903]), 
        .D(n25081), .Z(n25353) );
    VMW_AO22 U1967 ( .A(matrixInput[154]), .B(n25096), .C(matrixInput[146]), 
        .D(n25081), .Z(n27110) );
    VMW_AO22 U2334 ( .A(matrixInput[1147]), .B(n25096), .C(matrixInput[1139]), 
        .D(n25081), .Z(n26117) );
    VMW_FD \matrixInput_reg[171]  ( .D(n27085), .CP(Clk), .Q(matrixInput[171])
         );
    VMW_FD \matrixInput_reg[168]  ( .D(n27088), .CP(Clk), .Q(matrixInput[168])
         );
    VMW_AO22 U2525 ( .A(cOutput[19]), .B(n25087), .C(cOutput[3]), .D(n25084), 
        .Z(n25141) );
    VMW_FD \matrixInput_reg[1766]  ( .D(n25490), .CP(Clk), .Q(matrixInput
        [1766]) );
    VMW_FD \vectorInput_reg[19]  ( .D(n27365), .CP(Clk), .Q(vectorInput[19])
         );
    VMW_FD \matrixInput_reg[979]  ( .D(n26277), .CP(Clk), .Q(matrixInput[979])
         );
    VMW_FD \matrixInput_reg[960]  ( .D(n26296), .CP(Clk), .Q(matrixInput[960])
         );
    VMW_AO22 U483 ( .A(matrixInput[970]), .B(n25096), .C(matrixInput[962]), 
        .D(n25081), .Z(n26294) );
    VMW_AO22 U604 ( .A(matrixInput[861]), .B(n25096), .C(matrixInput[853]), 
        .D(n25081), .Z(n26403) );
    VMW_AO22 U1899 ( .A(matrixInput[1538]), .B(n25096), .C(matrixInput[1530]), 
        .D(n25081), .Z(n25726) );
    VMW_FD \vectorInput_reg[33]  ( .D(n27351), .CP(Clk), .Q(vectorInput[33])
         );
    VMW_AO22 U1909 ( .A(matrixInput[1529]), .B(n25096), .C(matrixInput[1521]), 
        .D(n25081), .Z(n25735) );
    VMW_AO22 U623 ( .A(matrixInput[844]), .B(n25096), .C(matrixInput[836]), 
        .D(n25081), .Z(n26420) );
    VMW_AO22 U794 ( .A(matrixInput[690]), .B(n25096), .C(matrixInput[682]), 
        .D(n25081), .Z(n26574) );
    VMW_FD \matrixInput_reg[953]  ( .D(n26303), .CP(Clk), .Q(matrixInput[953])
         );
    VMW_AO22 U961 ( .A(matrixInput[539]), .B(n25096), .C(matrixInput[531]), 
        .D(n25081), .Z(n26725) );
    VMW_FD \matrixInput_reg[1979]  ( .D(n25277), .CP(Clk), .Q(matrixInput
        [1979]) );
    VMW_FD \matrixInput_reg[1960]  ( .D(n25296), .CP(Clk), .Q(matrixInput
        [1960]) );
    VMW_FD \matrixInput_reg[1953]  ( .D(n25303), .CP(Clk), .Q(matrixInput
        [1953]) );
    VMW_FD \matrixInput_reg[83]  ( .D(n27173), .CP(Clk), .Q(matrixInput[83])
         );
    VMW_AO22 U513 ( .A(matrixInput[943]), .B(n25096), .C(matrixInput[935]), 
        .D(n25081), .Z(n26321) );
    VMW_OAI211 U295 ( .A(n25055), .B(n25059), .C(n25060), .D(n25061), .Z(
        n27391) );
    VMW_AO22 U389 ( .A(vectorInput[38]), .B(n25095), .C(vectorInput[30]), .D(
        n25080), .Z(n27354) );
    VMW_AO22 U408 ( .A(vectorInput[21]), .B(n25095), .C(vectorInput[13]), .D(
        n25080), .Z(n27371) );
    VMW_AO22 U738 ( .A(matrixInput[740]), .B(n25096), .C(matrixInput[732]), 
        .D(n25081), .Z(n26524) );
    VMW_AO22 U1141 ( .A(matrixInput[44]), .B(n25096), .C(matrixInput[36]), .D(
        n25081), .Z(n27220) );
    VMW_AO22 U1750 ( .A(matrixInput[1673]), .B(n25096), .C(matrixInput[1665]), 
        .D(n25081), .Z(n25591) );
    VMW_AO22 U2171 ( .A(matrixInput[1294]), .B(n25096), .C(matrixInput[1286]), 
        .D(n25081), .Z(n25970) );
    VMW_FD \matrixInput_reg[2043]  ( .D(n25213), .CP(Clk), .Q(matrixInput
        [2043]) );
    VMW_FD \matrixInput_reg[1624]  ( .D(n25632), .CP(Clk), .Q(matrixInput
        [1624]) );
    VMW_FD \matrixInput_reg[1527]  ( .D(n25729), .CP(Clk), .Q(matrixInput
        [1527]) );
    VMW_FD \matrixInput_reg[330]  ( .D(n26926), .CP(Clk), .Q(matrixInput[330])
         );
    VMW_FD \matrixInput_reg[329]  ( .D(n26927), .CP(Clk), .Q(matrixInput[329])
         );
    VMW_AO22 U1271 ( .A(matrixInput[260]), .B(n25096), .C(matrixInput[252]), 
        .D(n25081), .Z(n27004) );
    VMW_AO22 U1460 ( .A(matrixInput[1934]), .B(n25096), .C(matrixInput[1926]), 
        .D(n25081), .Z(n25330) );
    VMW_AO22 U2241 ( .A(matrixInput[1230]), .B(n25096), .C(matrixInput[1222]), 
        .D(n25081), .Z(n26034) );
    VMW_FD \matrixInput_reg[1514]  ( .D(n25742), .CP(Clk), .Q(matrixInput
        [1514]) );
    VMW_FD \matrixInput_reg[787]  ( .D(n26469), .CP(Clk), .Q(matrixInput[787])
         );
    VMW_FD \matrixInput_reg[303]  ( .D(n26953), .CP(Clk), .Q(matrixInput[303])
         );
    VMW_AO22 U2450 ( .A(matrixInput[1042]), .B(n25096), .C(matrixInput[1034]), 
        .D(n25081), .Z(n26222) );
    VMW_FD \matrixInput_reg[1189]  ( .D(n26067), .CP(Clk), .Q(matrixInput
        [1189]) );
    VMW_FD \matrixInput_reg[1293]  ( .D(n25963), .CP(Clk), .Q(matrixInput
        [1293]) );
    VMW_FD \matrixInput_reg[1190]  ( .D(n26066), .CP(Clk), .Q(matrixInput
        [1190]) );
    VMW_FD \matrixInput_reg[484]  ( .D(n26772), .CP(Clk), .Q(matrixInput[484])
         );
    VMW_AO22 U1812 ( .A(matrixInput[1617]), .B(n25096), .C(matrixInput[1609]), 
        .D(n25081), .Z(n25647) );
    VMW_FD \matrixInput_reg[1617]  ( .D(n25639), .CP(Clk), .Q(matrixInput
        [1617]) );
    VMW_AO22 U1982 ( .A(matrixInput[1464]), .B(n25096), .C(matrixInput[1456]), 
        .D(n25081), .Z(n25800) );
    VMW_FD \matrixInput_reg[527]  ( .D(n26729), .CP(Clk), .Q(matrixInput[527])
         );
    VMW_AO22 U1256 ( .A(matrixInput[274]), .B(n25096), .C(matrixInput[266]), 
        .D(n25081), .Z(n26990) );
    VMW_AO22 U2266 ( .A(matrixInput[19]), .B(n25096), .C(matrixInput[11]), .D(
        n25081), .Z(n27245) );
    VMW_AO22 U2477 ( .A(matrixInput[108]), .B(n25096), .C(matrixInput[100]), 
        .D(n25081), .Z(n27156) );
    VMW_FD \matrixInput_reg[1330]  ( .D(n25926), .CP(Clk), .Q(matrixInput
        [1330]) );
    VMW_FD \matrixInput_reg[1329]  ( .D(n25927), .CP(Clk), .Q(matrixInput
        [1329]) );
    VMW_FD \holder_reg[5]  ( .D(n27387), .CP(Clk), .Q(\holder[5] ) );
    VMW_AO22 U1447 ( .A(matrixInput[1946]), .B(n25096), .C(matrixInput[1938]), 
        .D(n25081), .Z(n25318) );
    VMW_FD \matrixInput_reg[624]  ( .D(n26632), .CP(Clk), .Q(matrixInput[624])
         );
    VMW_AO22 U1835 ( .A(matrixInput[1597]), .B(n25096), .C(matrixInput[1589]), 
        .D(n25081), .Z(n25667) );
    VMW_FD \matrixInput_reg[1033]  ( .D(n26223), .CP(Clk), .Q(matrixInput
        [1033]) );
    VMW_FD \matrixInput_reg[1303]  ( .D(n25953), .CP(Clk), .Q(matrixInput
        [1303]) );
    VMW_FD \matrixInput_reg[514]  ( .D(n26742), .CP(Clk), .Q(matrixInput[514])
         );
    VMW_AO22 U598 ( .A(matrixInput[867]), .B(n25096), .C(matrixInput[859]), 
        .D(n25081), .Z(n26397) );
    VMW_AO22 U1166 ( .A(matrixInput[355]), .B(n25096), .C(matrixInput[347]), 
        .D(n25081), .Z(n26909) );
    VMW_AO22 U2156 ( .A(matrixInput[137]), .B(n25096), .C(matrixInput[129]), 
        .D(n25081), .Z(n27127) );
    VMW_FD \matrixInput_reg[1787]  ( .D(n25469), .CP(Clk), .Q(matrixInput
        [1787]) );
    VMW_FD \matrixInput_reg[190]  ( .D(n27066), .CP(Clk), .Q(matrixInput[190])
         );
    VMW_FD \matrixInput_reg[189]  ( .D(n27067), .CP(Clk), .Q(matrixInput[189])
         );
    VMW_FD \matrixInput_reg[1484]  ( .D(n25772), .CP(Clk), .Q(matrixInput
        [1484]) );
    VMW_FD \matrixInput_reg[293]  ( .D(n26963), .CP(Clk), .Q(matrixInput[293])
         );
    VMW_FD \matrixInput_reg[1019]  ( .D(n26237), .CP(Clk), .Q(matrixInput
        [1019]) );
    VMW_FD \matrixInput_reg[1000]  ( .D(n26256), .CP(Clk), .Q(matrixInput
        [1000]) );
    VMW_AO22 U1777 ( .A(matrixInput[1648]), .B(n25096), .C(matrixInput[1640]), 
        .D(n25081), .Z(n25616) );
    VMW_FD \matrixInput_reg[617]  ( .D(n26639), .CP(Clk), .Q(matrixInput[617])
         );
    VMW_AND2 U305 ( .A(n25055), .B(Addr[1]), .Z(n25086) );
    VMW_AO22 U514 ( .A(matrixInput[942]), .B(n25096), .C(matrixInput[934]), 
        .D(n25081), .Z(n26322) );
    VMW_AO22 U322 ( .A(vectorInput[99]), .B(n25095), .C(vectorInput[91]), .D(
        n25080), .Z(n27293) );
    VMW_AO22 U484 ( .A(matrixInput[969]), .B(n25096), .C(matrixInput[961]), 
        .D(n25081), .Z(n26295) );
    VMW_AO22 U603 ( .A(matrixInput[862]), .B(n25096), .C(matrixInput[854]), 
        .D(n25081), .Z(n26402) );
    VMW_AO22 U624 ( .A(matrixInput[843]), .B(n25096), .C(matrixInput[835]), 
        .D(n25081), .Z(n26421) );
    VMW_AO22 U966 ( .A(matrixInput[535]), .B(n25096), .C(matrixInput[527]), 
        .D(n25081), .Z(n26729) );
    VMW_FD \matrixInput_reg[962]  ( .D(n26294), .CP(Clk), .Q(matrixInput[962])
         );
    VMW_FD \matrixInput_reg[951]  ( .D(n26305), .CP(Clk), .Q(matrixInput[951])
         );
    VMW_FD \matrixInput_reg[948]  ( .D(n26308), .CP(Clk), .Q(matrixInput[948])
         );
    VMW_AO22 U793 ( .A(matrixInput[691]), .B(n25096), .C(matrixInput[683]), 
        .D(n25081), .Z(n26573) );
    VMW_AO22 U1929 ( .A(matrixInput[1511]), .B(n25096), .C(matrixInput[1503]), 
        .D(n25081), .Z(n25753) );
    VMW_FD \matrixInput_reg[1962]  ( .D(n25294), .CP(Clk), .Q(matrixInput
        [1962]) );
    VMW_FD \vectorInput_reg[31]  ( .D(n27353), .CP(Clk), .Q(vectorInput[31])
         );
    VMW_FD \vectorInput_reg[28]  ( .D(n27356), .CP(Clk), .Q(vectorInput[28])
         );
    VMW_AO22 U428 ( .A(vectorInput[118]), .B(n25095), .C(vectorInput[110]), 
        .D(n25080), .Z(n27274) );
    VMW_AO22 U533 ( .A(matrixInput[925]), .B(n25096), .C(matrixInput[917]), 
        .D(n25081), .Z(n26339) );
    VMW_AO22 U688 ( .A(matrixInput[786]), .B(n25096), .C(matrixInput[778]), 
        .D(n25081), .Z(n26478) );
    VMW_AO22 U718 ( .A(matrixInput[758]), .B(n25096), .C(matrixInput[750]), 
        .D(n25081), .Z(n26506) );
    VMW_AO22 U941 ( .A(matrixInput[62]), .B(n25096), .C(matrixInput[54]), .D(
        n25081), .Z(n27202) );
    VMW_FD \matrixInput_reg[1951]  ( .D(n25305), .CP(Clk), .Q(matrixInput
        [1951]) );
    VMW_FD \matrixInput_reg[1948]  ( .D(n25308), .CP(Clk), .Q(matrixInput
        [1948]) );
    VMW_FD \matrixInput_reg[98]  ( .D(n27158), .CP(Clk), .Q(matrixInput[98])
         );
    VMW_FD \matrixInput_reg[81]  ( .D(n27175), .CP(Clk), .Q(matrixInput[81])
         );
    VMW_AO22 U1161 ( .A(matrixInput[359]), .B(n25096), .C(matrixInput[351]), 
        .D(n25081), .Z(n26905) );
    VMW_AO22 U1770 ( .A(matrixInput[1655]), .B(n25096), .C(matrixInput[1647]), 
        .D(n25081), .Z(n25609) );
    VMW_AO22 U1251 ( .A(matrixInput[278]), .B(n25096), .C(matrixInput[270]), 
        .D(n25081), .Z(n26986) );
    VMW_AO22 U1440 ( .A(matrixInput[1952]), .B(n25096), .C(matrixInput[1944]), 
        .D(n25081), .Z(n25312) );
    VMW_AO22 U1832 ( .A(matrixInput[1599]), .B(n25096), .C(matrixInput[1591]), 
        .D(n25081), .Z(n25665) );
    VMW_AO22 U2151 ( .A(matrixInput[1311]), .B(n25096), .C(matrixInput[1303]), 
        .D(n25081), .Z(n25953) );
    VMW_FD \matrixInput_reg[2041]  ( .D(n25215), .CP(Clk), .Q(matrixInput
        [2041]) );
    VMW_FD \matrixInput_reg[1626]  ( .D(n25630), .CP(Clk), .Q(matrixInput
        [1626]) );
    VMW_FD \matrixInput_reg[1525]  ( .D(n25731), .CP(Clk), .Q(matrixInput
        [1525]) );
    VMW_FD \matrixInput_reg[332]  ( .D(n26924), .CP(Clk), .Q(matrixInput[332])
         );
    VMW_FD \matrixInput_reg[1615]  ( .D(n25641), .CP(Clk), .Q(matrixInput
        [1615]) );
    VMW_FD \matrixInput_reg[1291]  ( .D(n25965), .CP(Clk), .Q(matrixInput
        [1291]) );
    VMW_FD \matrixInput_reg[1288]  ( .D(n25968), .CP(Clk), .Q(matrixInput
        [1288]) );
    VMW_AO22 U1276 ( .A(matrixInput[256]), .B(n25096), .C(matrixInput[248]), 
        .D(n25081), .Z(n27008) );
    VMW_AO22 U1815 ( .A(matrixInput[1614]), .B(n25096), .C(matrixInput[1606]), 
        .D(n25081), .Z(n25650) );
    VMW_AO22 U1985 ( .A(matrixInput[1461]), .B(n25096), .C(matrixInput[1453]), 
        .D(n25081), .Z(n25803) );
    VMW_AO22 U2261 ( .A(matrixInput[1212]), .B(n25096), .C(matrixInput[1204]), 
        .D(n25081), .Z(n26052) );
    VMW_FD \matrixInput_reg[486]  ( .D(n26770), .CP(Clk), .Q(matrixInput[486])
         );
    VMW_AO22 U2470 ( .A(matrixInput[1024]), .B(n25096), .C(matrixInput[1016]), 
        .D(n25081), .Z(n26240) );
    VMW_FD \matrixInput_reg[1192]  ( .D(n26064), .CP(Clk), .Q(matrixInput
        [1192]) );
    VMW_FD \matrixInput_reg[1516]  ( .D(n25740), .CP(Clk), .Q(matrixInput
        [1516]) );
    VMW_FD \matrixInput_reg[785]  ( .D(n26471), .CP(Clk), .Q(matrixInput[785])
         );
    VMW_FD \matrixInput_reg[318]  ( .D(n26938), .CP(Clk), .Q(matrixInput[318])
         );
    VMW_FD \matrixInput_reg[301]  ( .D(n26955), .CP(Clk), .Q(matrixInput[301])
         );
    VMW_FD \matrixInput_reg[1031]  ( .D(n26225), .CP(Clk), .Q(matrixInput
        [1031]) );
    VMW_FD \matrixInput_reg[1028]  ( .D(n26228), .CP(Clk), .Q(matrixInput
        [1028]) );
    VMW_AO22 U1467 ( .A(matrixInput[199]), .B(n25096), .C(matrixInput[191]), 
        .D(n25081), .Z(n27065) );
    VMW_FD \matrixInput_reg[1332]  ( .D(n25924), .CP(Clk), .Q(matrixInput
        [1332]) );
    VMW_FD \matrixInput_reg[626]  ( .D(n26630), .CP(Clk), .Q(matrixInput[626])
         );
    VMW_FD \holder_reg[7]  ( .D(n27385), .CP(Clk), .Q(\holder[7] ) );
    VMW_AO22 U2457 ( .A(matrixInput[1036]), .B(n25096), .C(matrixInput[1028]), 
        .D(n25081), .Z(n26228) );
    VMW_FD \matrixInput_reg[525]  ( .D(n26731), .CP(Clk), .Q(matrixInput[525])
         );
    VMW_AO22 U1146 ( .A(matrixInput[373]), .B(n25096), .C(matrixInput[365]), 
        .D(n25081), .Z(n26891) );
    VMW_AO22 U2246 ( .A(matrixInput[1226]), .B(n25096), .C(matrixInput[1218]), 
        .D(n25081), .Z(n26038) );
    VMW_AO22 U1757 ( .A(matrixInput[1667]), .B(n25096), .C(matrixInput[1659]), 
        .D(n25081), .Z(n25597) );
    VMW_FD \matrixInput_reg[615]  ( .D(n26641), .CP(Clk), .Q(matrixInput[615])
         );
    VMW_FD \matrixInput_reg[1785]  ( .D(n25471), .CP(Clk), .Q(matrixInput
        [1785]) );
    VMW_FD \matrixInput_reg[1486]  ( .D(n25770), .CP(Clk), .Q(matrixInput
        [1486]) );
    VMW_FD \matrixInput_reg[1002]  ( .D(n26254), .CP(Clk), .Q(matrixInput
        [1002]) );
    VMW_FD \matrixInput_reg[291]  ( .D(n26965), .CP(Clk), .Q(matrixInput[291])
         );
    VMW_FD \matrixInput_reg[288]  ( .D(n26968), .CP(Clk), .Q(matrixInput[288])
         );
    VMW_FD \matrixInput_reg[516]  ( .D(n26740), .CP(Clk), .Q(matrixInput[516])
         );
    VMW_FD \matrixInput_reg[192]  ( .D(n27064), .CP(Clk), .Q(matrixInput[192])
         );
    VMW_AO22 U446 ( .A(matrixInput[1004]), .B(n25096), .C(matrixInput[996]), 
        .D(n25081), .Z(n26260) );
    VMW_AO22 U776 ( .A(matrixInput[707]), .B(n25096), .C(matrixInput[699]), 
        .D(n25081), .Z(n26557) );
    VMW_AO22 U1218 ( .A(matrixInput[10]), .B(n25096), .C(matrixInput[2]), .D(
        n25081), .Z(n27254) );
    VMW_AO22 U1388 ( .A(matrixInput[1999]), .B(n25096), .C(matrixInput[1991]), 
        .D(n25081), .Z(n25265) );
    VMW_AO22 U1409 ( .A(matrixInput[1980]), .B(n25096), .C(matrixInput[1972]), 
        .D(n25081), .Z(n25284) );
    VMW_AO22 U2176 ( .A(matrixInput[1289]), .B(n25096), .C(matrixInput[1281]), 
        .D(n25081), .Z(n25975) );
    VMW_FD \matrixInput_reg[1318]  ( .D(n25938), .CP(Clk), .Q(matrixInput
        [1318]) );
    VMW_FD \matrixInput_reg[1301]  ( .D(n25955), .CP(Clk), .Q(matrixInput
        [1301]) );
    VMW_AO22 U1599 ( .A(matrixInput[1808]), .B(n25096), .C(matrixInput[1800]), 
        .D(n25081), .Z(n25456) );
    VMW_AO22 U2228 ( .A(matrixInput[1242]), .B(n25096), .C(matrixInput[1234]), 
        .D(n25081), .Z(n26022) );
    VMW_FD \matrixInput_reg[1813]  ( .D(n25443), .CP(Clk), .Q(matrixInput
        [1813]) );
    VMW_AO22 U1128 ( .A(matrixInput[389]), .B(n25096), .C(matrixInput[381]), 
        .D(n25081), .Z(n26875) );
    VMW_AO22 U1739 ( .A(matrixInput[1683]), .B(n25096), .C(matrixInput[1675]), 
        .D(n25081), .Z(n25581) );
    VMW_AO22 U2439 ( .A(matrixInput[1052]), .B(n25096), .C(matrixInput[1044]), 
        .D(n25081), .Z(n26212) );
    VMW_FD \matrixInput_reg[1839]  ( .D(n25417), .CP(Clk), .Q(matrixInput
        [1839]) );
    VMW_FD \matrixInput_reg[983]  ( .D(n26273), .CP(Clk), .Q(matrixInput[983])
         );
    VMW_FD \matrixInput_reg[1820]  ( .D(n25436), .CP(Clk), .Q(matrixInput
        [1820]) );
    VMW_AO22 U2088 ( .A(matrixInput[1368]), .B(n25096), .C(matrixInput[1360]), 
        .D(n25081), .Z(n25896) );
    VMW_AO22 U2118 ( .A(matrixInput[1341]), .B(n25096), .C(matrixInput[1333]), 
        .D(n25081), .Z(n25923) );
    VMW_AO22 U461 ( .A(matrixInput[990]), .B(n25096), .C(matrixInput[982]), 
        .D(n25081), .Z(n26274) );
    VMW_AO22 U834 ( .A(matrixInput[654]), .B(n25096), .C(matrixInput[646]), 
        .D(n25081), .Z(n26610) );
    VMW_FD \matrixInput_reg[813]  ( .D(n26443), .CP(Clk), .Q(matrixInput[813])
         );
    VMW_PULLDOWN U279 ( .Z(n25197) );
    VMW_AO22 U339 ( .A(vectorInput[84]), .B(n25095), .C(vectorInput[76]), .D(
        n25080), .Z(n27308) );
    VMW_AO22 U357 ( .A(vectorInput[13]), .B(n25095), .C(vectorInput[5]), .D(
        n25080), .Z(n27379) );
    VMW_AO22 U370 ( .A(vectorInput[56]), .B(n25095), .C(vectorInput[48]), .D(
        n25080), .Z(n27336) );
    VMW_AO22 U651 ( .A(matrixInput[818]), .B(n25096), .C(matrixInput[810]), 
        .D(n25081), .Z(n26446) );
    VMW_AO22 U751 ( .A(matrixInput[728]), .B(n25096), .C(matrixInput[720]), 
        .D(n25081), .Z(n26536) );
    VMW_AO22 U813 ( .A(matrixInput[673]), .B(n25096), .C(matrixInput[665]), 
        .D(n25081), .Z(n26591) );
    VMW_FD \matrixInput_reg[1983]  ( .D(n25273), .CP(Clk), .Q(matrixInput
        [1983]) );
    VMW_FD \matrixInput_reg[53]  ( .D(n27203), .CP(Clk), .Q(matrixInput[53])
         );
    VMW_AO22 U983 ( .A(matrixInput[519]), .B(n25096), .C(matrixInput[511]), 
        .D(n25081), .Z(n26745) );
    VMW_FD \matrixInput_reg[839]  ( .D(n26417), .CP(Clk), .Q(matrixInput[839])
         );
    VMW_FD \matrixInput_reg[820]  ( .D(n26436), .CP(Clk), .Q(matrixInput[820])
         );
    VMW_FD \matrixInput_reg[79]  ( .D(n27177), .CP(Clk), .Q(matrixInput[79])
         );
    VMW_FD \matrixInput_reg[60]  ( .D(n27196), .CP(Clk), .Q(matrixInput[60])
         );
    VMW_AO22 U898 ( .A(matrixInput[597]), .B(n25096), .C(matrixInput[589]), 
        .D(n25081), .Z(n26667) );
    VMW_AO22 U1033 ( .A(matrixInput[475]), .B(n25096), .C(matrixInput[467]), 
        .D(n25081), .Z(n26789) );
    VMW_AO22 U1293 ( .A(matrixInput[240]), .B(n25096), .C(matrixInput[232]), 
        .D(n25081), .Z(n27024) );
    VMW_AO22 U1303 ( .A(matrixInput[231]), .B(n25096), .C(matrixInput[223]), 
        .D(n25081), .Z(n27033) );
    VMW_AO22 U1482 ( .A(matrixInput[1914]), .B(n25096), .C(matrixInput[1906]), 
        .D(n25081), .Z(n25350) );
    VMW_AO22 U1960 ( .A(matrixInput[1484]), .B(n25096), .C(matrixInput[1476]), 
        .D(n25081), .Z(n25780) );
    VMW_AO22 U2333 ( .A(matrixInput[121]), .B(n25096), .C(matrixInput[113]), 
        .D(n25081), .Z(n27143) );
    VMW_AO22 U2522 ( .A(cOutput[116]), .B(n25087), .C(cOutput[100]), .D(n25084
        ), .Z(n25136) );
    VMW_FD \matrixInput_reg[1243]  ( .D(n26013), .CP(Clk), .Q(matrixInput
        [1243]) );
    VMW_FD \matrixInput_reg[1159]  ( .D(n26097), .CP(Clk), .Q(matrixInput
        [1159]) );
    VMW_FD \matrixInput_reg[1140]  ( .D(n26116), .CP(Clk), .Q(matrixInput
        [1140]) );
    VMW_FD \matrixInput_reg[757]  ( .D(n26499), .CP(Clk), .Q(matrixInput[757])
         );
    VMW_FD \matrixInput_reg[454]  ( .D(n26802), .CP(Clk), .Q(matrixInput[454])
         );
    VMW_AO22 U1512 ( .A(matrixInput[195]), .B(n25096), .C(matrixInput[187]), 
        .D(n25081), .Z(n27069) );
    VMW_AO22 U2003 ( .A(matrixInput[1445]), .B(n25096), .C(matrixInput[1437]), 
        .D(n25081), .Z(n25819) );
    VMW_AO22 U2193 ( .A(matrixInput[1274]), .B(n25096), .C(matrixInput[1266]), 
        .D(n25081), .Z(n25990) );
    VMW_FD \matrixInput_reg[1173]  ( .D(n26083), .CP(Clk), .Q(matrixInput
        [1173]) );
    VMW_FD \matrixInput_reg[764]  ( .D(n26492), .CP(Clk), .Q(matrixInput[764])
         );
    VMW_BUFIZ U2612 ( .A(\holder[0] ), .E(RD), .Z(\DataOut[0]1 ) );
    VMW_AO22 U1622 ( .A(matrixInput[1788]), .B(n25096), .C(matrixInput[1780]), 
        .D(n25081), .Z(n25476) );
    VMW_FD \matrixInput_reg[1270]  ( .D(n25986), .CP(Clk), .Q(matrixInput
        [1270]) );
    VMW_FD \matrixInput_reg[1269]  ( .D(n25987), .CP(Clk), .Q(matrixInput
        [1269]) );
    VMW_FD \matrixInput_reg[467]  ( .D(n26789), .CP(Clk), .Q(matrixInput[467])
         );
    VMW_AO22 U908 ( .A(matrixInput[65]), .B(n25096), .C(matrixInput[57]), .D(
        n25081), .Z(n27199) );
    VMW_AO22 U1014 ( .A(matrixInput[492]), .B(n25096), .C(matrixInput[484]), 
        .D(n25081), .Z(n26772) );
    VMW_AO22 U1184 ( .A(matrixInput[338]), .B(n25096), .C(matrixInput[330]), 
        .D(n25081), .Z(n26926) );
    VMW_AO22 U2024 ( .A(matrixInput[1426]), .B(n25096), .C(matrixInput[1418]), 
        .D(n25081), .Z(n25838) );
    VMW_FD \matrixInput_reg[159]  ( .D(n27097), .CP(Clk), .Q(matrixInput[159])
         );
    VMW_FD \matrixInput_reg[140]  ( .D(n27116), .CP(Clk), .Q(matrixInput[140])
         );
    VMW_BUFIZ U2635 ( .A(n25205), .E(RD), .Z(\DataOut[22]1 ) );
    VMW_FD \matrixInput_reg[1757]  ( .D(n25499), .CP(Clk), .Q(matrixInput
        [1757]) );
    VMW_FD \matrixInput_reg[243]  ( .D(n27013), .CP(Clk), .Q(matrixInput[243])
         );
    VMW_AO22 U1605 ( .A(matrixInput[1804]), .B(n25096), .C(matrixInput[1796]), 
        .D(n25081), .Z(n25460) );
    VMW_FD \matrixInput_reg[1454]  ( .D(n25802), .CP(Clk), .Q(matrixInput
        [1454]) );
    VMW_AO22 U1324 ( .A(matrixInput[212]), .B(n25096), .C(matrixInput[204]), 
        .D(n25081), .Z(n27052) );
    VMW_AO22 U1535 ( .A(matrixInput[1867]), .B(n25096), .C(matrixInput[1859]), 
        .D(n25081), .Z(n25397) );
    VMW_AO22 U1795 ( .A(matrixInput[1632]), .B(n25096), .C(matrixInput[1624]), 
        .D(n25081), .Z(n25632) );
    VMW_AO22 U1947 ( .A(matrixInput[1496]), .B(n25096), .C(matrixInput[1488]), 
        .D(n25081), .Z(n25768) );
    VMW_AO22 U2284 ( .A(matrixInput[1192]), .B(n25096), .C(matrixInput[1184]), 
        .D(n25081), .Z(n26072) );
    VMW_AO22 U2314 ( .A(matrixInput[1165]), .B(n25096), .C(matrixInput[1157]), 
        .D(n25081), .Z(n26099) );
    VMW_AO22 U2495 ( .A(cOutput[119]), .B(n25087), .C(cOutput[103]), .D(n25084
        ), .Z(n25103) );
    VMW_AO22 U2505 ( .A(cOutput[126]), .B(n25089), .C(cOutput[110]), .D(n25088
        ), .Z(n25115) );
    VMW_FD \matrixInput_reg[1764]  ( .D(n25492), .CP(Clk), .Q(matrixInput
        [1764]) );
    VMW_FD \matrixInput_reg[173]  ( .D(n27083), .CP(Clk), .Q(matrixInput[173])
         );
    VMW_FD \matrixInput_reg[1467]  ( .D(n25789), .CP(Clk), .Q(matrixInput
        [1467]) );
    VMW_FD \matrixInput_reg[830]  ( .D(n26426), .CP(Clk), .Q(matrixInput[830])
         );
    VMW_FD \matrixInput_reg[270]  ( .D(n26986), .CP(Clk), .Q(matrixInput[270])
         );
    VMW_FD \matrixInput_reg[269]  ( .D(n26987), .CP(Clk), .Q(matrixInput[269])
         );
    VMW_FD \matrixInput_reg[829]  ( .D(n26427), .CP(Clk), .Q(matrixInput[829])
         );
    VMW_FD \matrixInput_reg[70]  ( .D(n27186), .CP(Clk), .Q(matrixInput[70])
         );
    VMW_FD \matrixInput_reg[69]  ( .D(n27187), .CP(Clk), .Q(matrixInput[69])
         );
    VMW_FD \matrixInput_reg[803]  ( .D(n26453), .CP(Clk), .Q(matrixInput[803])
         );
    VMW_AO22 U546 ( .A(matrixInput[913]), .B(n25096), .C(matrixInput[905]), 
        .D(n25081), .Z(n26351) );
    VMW_AO22 U561 ( .A(matrixInput[900]), .B(n25096), .C(matrixInput[892]), 
        .D(n25081), .Z(n26364) );
    VMW_AO22 U883 ( .A(matrixInput[609]), .B(n25096), .C(matrixInput[601]), 
        .D(n25081), .Z(n26655) );
    VMW_AO22 U913 ( .A(matrixInput[583]), .B(n25096), .C(matrixInput[575]), 
        .D(n25081), .Z(n26681) );
    VMW_AO22 U1028 ( .A(matrixInput[479]), .B(n25096), .C(matrixInput[471]), 
        .D(n25081), .Z(n26785) );
    VMW_FD \matrixInput_reg[1993]  ( .D(n25263), .CP(Clk), .Q(matrixInput
        [1993]) );
    VMW_FD \matrixInput_reg[1830]  ( .D(n25426), .CP(Clk), .Q(matrixInput
        [1830]) );
    VMW_FD \matrixInput_reg[43]  ( .D(n27213), .CP(Clk), .Q(matrixInput[43])
         );
    VMW_FD \matrixInput_reg[1829]  ( .D(n25427), .CP(Clk), .Q(matrixInput
        [1829]) );
    VMW_AO22 U1639 ( .A(matrixInput[1773]), .B(n25096), .C(matrixInput[1765]), 
        .D(n25081), .Z(n25491) );
    VMW_AO22 U2188 ( .A(matrixInput[1278]), .B(n25096), .C(matrixInput[1270]), 
        .D(n25081), .Z(n25986) );
    VMW_BUFIZ U2609 ( .A(n25186), .E(RD), .Z(\DataOut[23]1 ) );
    VMW_AO22 U395 ( .A(vectorInput[33]), .B(n25095), .C(vectorInput[25]), .D(
        n25080), .Z(n27359) );
    VMW_AO22 U433 ( .A(vectorInput[114]), .B(n25095), .C(vectorInput[106]), 
        .D(n25080), .Z(n27278) );
    VMW_AO22 U676 ( .A(matrixInput[797]), .B(n25096), .C(matrixInput[789]), 
        .D(n25081), .Z(n26467) );
    VMW_AO22 U934 ( .A(matrixInput[564]), .B(n25096), .C(matrixInput[556]), 
        .D(n25081), .Z(n26700) );
    VMW_AO22 U2018 ( .A(matrixInput[1431]), .B(n25096), .C(matrixInput[1423]), 
        .D(n25081), .Z(n25833) );
    VMW_AO22 U1288 ( .A(matrixInput[245]), .B(n25096), .C(matrixInput[237]), 
        .D(n25081), .Z(n27019) );
    VMW_AO22 U1318 ( .A(matrixInput[28]), .B(n25096), .C(matrixInput[20]), .D(
        n25081), .Z(n27236) );
    VMW_AO22 U1499 ( .A(matrixInput[1899]), .B(n25096), .C(matrixInput[1891]), 
        .D(n25081), .Z(n25365) );
    VMW_AO22 U1509 ( .A(matrixInput[1890]), .B(n25096), .C(matrixInput[1882]), 
        .D(n25081), .Z(n25374) );
    VMW_FD \matrixInput_reg[1803]  ( .D(n25453), .CP(Clk), .Q(matrixInput
        [1803]) );
    VMW_AO22 U808 ( .A(matrixInput[74]), .B(n25096), .C(matrixInput[66]), .D(
        n25081), .Z(n27190) );
    VMW_AO22 U1224 ( .A(matrixInput[303]), .B(n25096), .C(matrixInput[295]), 
        .D(n25081), .Z(n26961) );
    VMW_AO22 U1847 ( .A(matrixInput[1586]), .B(n25096), .C(matrixInput[1578]), 
        .D(n25081), .Z(n25678) );
    VMW_AO22 U2214 ( .A(matrixInput[1255]), .B(n25096), .C(matrixInput[1247]), 
        .D(n25081), .Z(n26009) );
    VMW_AO22 U2328 ( .A(matrixInput[1152]), .B(n25096), .C(matrixInput[1144]), 
        .D(n25081), .Z(n26112) );
    VMW_AO22 U2539 ( .A(cOutput[90]), .B(n25089), .C(cOutput[74]), .D(n25088), 
        .Z(n25157) );
    VMW_FD \matrixInput_reg[993]  ( .D(n26263), .CP(Clk), .Q(matrixInput[993])
         );
    VMW_AO22 U2384 ( .A(matrixInput[1102]), .B(n25096), .C(matrixInput[1094]), 
        .D(n25081), .Z(n26162) );
    VMW_AO22 U2405 ( .A(matrixInput[1083]), .B(n25096), .C(matrixInput[1075]), 
        .D(n25081), .Z(n26181) );
    VMW_FD \matrixInput_reg[163]  ( .D(n27093), .CP(Clk), .Q(matrixInput[163])
         );
    VMW_INV U2595 ( .A(n25080), .Z(n25095) );
    VMW_FD \matrixInput_reg[1774]  ( .D(n25482), .CP(Clk), .Q(matrixInput
        [1774]) );
    VMW_FD \matrixInput_reg[1477]  ( .D(n25779), .CP(Clk), .Q(matrixInput
        [1477]) );
    VMW_FD \matrixInput_reg[279]  ( .D(n26977), .CP(Clk), .Q(matrixInput[279])
         );
    VMW_FD \matrixInput_reg[260]  ( .D(n26996), .CP(Clk), .Q(matrixInput[260])
         );
    VMW_AO22 U1435 ( .A(matrixInput[1957]), .B(n25096), .C(matrixInput[1949]), 
        .D(n25081), .Z(n25307) );
    VMW_AO22 U998 ( .A(matrixInput[507]), .B(n25096), .C(matrixInput[499]), 
        .D(n25081), .Z(n26757) );
    VMW_AO22 U1084 ( .A(matrixInput[428]), .B(n25096), .C(matrixInput[420]), 
        .D(n25081), .Z(n26836) );
    VMW_AO22 U1114 ( .A(matrixInput[402]), .B(n25096), .C(matrixInput[394]), 
        .D(n25081), .Z(n26862) );
    VMW_AO22 U2124 ( .A(matrixInput[1336]), .B(n25096), .C(matrixInput[1328]), 
        .D(n25081), .Z(n25928) );
    VMW_FD \matrixInput_reg[1747]  ( .D(n25509), .CP(Clk), .Q(matrixInput
        [1747]) );
    VMW_FD \matrixInput_reg[1444]  ( .D(n25812), .CP(Clk), .Q(matrixInput
        [1444]) );
    VMW_FD \matrixInput_reg[150]  ( .D(n27106), .CP(Clk), .Q(matrixInput[150])
         );
    VMW_FD \matrixInput_reg[149]  ( .D(n27107), .CP(Clk), .Q(matrixInput[149])
         );
    VMW_AO22 U1695 ( .A(matrixInput[1722]), .B(n25096), .C(matrixInput[1714]), 
        .D(n25081), .Z(n25542) );
    VMW_AO22 U1133 ( .A(matrixInput[385]), .B(n25096), .C(matrixInput[377]), 
        .D(n25081), .Z(n26879) );
    VMW_AO22 U1705 ( .A(matrixInput[1713]), .B(n25096), .C(matrixInput[1705]), 
        .D(n25081), .Z(n25551) );
    VMW_AO22 U1722 ( .A(matrixInput[1698]), .B(n25096), .C(matrixInput[1690]), 
        .D(n25081), .Z(n25566) );
    VMW_AO22 U2093 ( .A(matrixInput[1364]), .B(n25096), .C(matrixInput[1356]), 
        .D(n25081), .Z(n25900) );
    VMW_AO22 U2103 ( .A(matrixInput[1355]), .B(n25096), .C(matrixInput[1347]), 
        .D(n25081), .Z(n25909) );
    VMW_FD \matrixInput_reg[1163]  ( .D(n26093), .CP(Clk), .Q(matrixInput
        [1163]) );
    VMW_FD \matrixInput_reg[774]  ( .D(n26482), .CP(Clk), .Q(matrixInput[774])
         );
    VMW_FD \matrixInput_reg[253]  ( .D(n27003), .CP(Clk), .Q(matrixInput[253])
         );
    VMW_AO22 U1203 ( .A(matrixInput[321]), .B(n25096), .C(matrixInput[313]), 
        .D(n25081), .Z(n26943) );
    VMW_AO22 U1393 ( .A(matrixInput[1995]), .B(n25096), .C(matrixInput[1987]), 
        .D(n25081), .Z(n25269) );
    VMW_AO22 U1412 ( .A(matrixInput[204]), .B(n25096), .C(matrixInput[196]), 
        .D(n25081), .Z(n27060) );
    VMW_AO22 U1860 ( .A(matrixInput[1574]), .B(n25096), .C(matrixInput[1566]), 
        .D(n25081), .Z(n25690) );
    VMW_AO22 U2233 ( .A(matrixInput[130]), .B(n25096), .C(matrixInput[122]), 
        .D(n25081), .Z(n27134) );
    VMW_FD \matrixInput_reg[1279]  ( .D(n25977), .CP(Clk), .Q(matrixInput
        [1279]) );
    VMW_FD \matrixInput_reg[1260]  ( .D(n25996), .CP(Clk), .Q(matrixInput
        [1260]) );
    VMW_FD \matrixInput_reg[477]  ( .D(n26779), .CP(Clk), .Q(matrixInput[477])
         );
    VMW_AO22 U2422 ( .A(matrixInput[113]), .B(n25096), .C(matrixInput[105]), 
        .D(n25081), .Z(n27151) );
    VMW_FD \matrixInput_reg[1150]  ( .D(n26106), .CP(Clk), .Q(matrixInput
        [1150]) );
    VMW_FD \matrixInput_reg[1149]  ( .D(n26107), .CP(Clk), .Q(matrixInput
        [1149]) );
    VMW_FD \matrixInput_reg[747]  ( .D(n26509), .CP(Clk), .Q(matrixInput[747])
         );
    VMW_FD \matrixInput_reg[1253]  ( .D(n26003), .CP(Clk), .Q(matrixInput
        [1253]) );
    VMW_FD \matrixInput_reg[444]  ( .D(n26812), .CP(Clk), .Q(matrixInput[444])
         );
    VMW_AO22 U1582 ( .A(matrixInput[1824]), .B(n25096), .C(matrixInput[1816]), 
        .D(n25081), .Z(n25440) );
    VMW_FD \matrixInput_reg[1958]  ( .D(n25298), .CP(Clk), .Q(matrixInput
        [1958]) );
    VMW_FD \matrixInput_reg[91]  ( .D(n27165), .CP(Clk), .Q(matrixInput[91])
         );
    VMW_FD \matrixInput_reg[1941]  ( .D(n25315), .CP(Clk), .Q(matrixInput
        [1941]) );
    VMW_FD \matrixInput_reg[88]  ( .D(n27168), .CP(Clk), .Q(matrixInput[88])
         );
    VMW_AO22 U584 ( .A(matrixInput[879]), .B(n25096), .C(matrixInput[871]), 
        .D(n25081), .Z(n26385) );
    VMW_AO22 U693 ( .A(matrixInput[781]), .B(n25096), .C(matrixInput[773]), 
        .D(n25081), .Z(n26483) );
    VMW_AO22 U703 ( .A(matrixInput[772]), .B(n25096), .C(matrixInput[764]), 
        .D(n25081), .Z(n26492) );
    VMW_AO22 U841 ( .A(matrixInput[71]), .B(n25096), .C(matrixInput[63]), .D(
        n25081), .Z(n27193) );
    VMW_AO22 U724 ( .A(matrixInput[753]), .B(n25096), .C(matrixInput[745]), 
        .D(n25081), .Z(n26511) );
    VMW_FD \matrixInput_reg[1972]  ( .D(n25284), .CP(Clk), .Q(matrixInput
        [1972]) );
    VMW_FD \matrixInput_reg[958]  ( .D(n26298), .CP(Clk), .Q(matrixInput[958])
         );
    VMW_FD \matrixInput_reg[941]  ( .D(n26315), .CP(Clk), .Q(matrixInput[941])
         );
    VMW_AO22 U1829 ( .A(matrixInput[1602]), .B(n25096), .C(matrixInput[1594]), 
        .D(n25081), .Z(n25662) );
    VMW_FD \vectorInput_reg[38]  ( .D(n27346), .CP(Clk), .Q(vectorInput[38])
         );
    VMW_FD \vectorInput_reg[21]  ( .D(n27363), .CP(Clk), .Q(vectorInput[21])
         );
    VMW_AO22 U414 ( .A(DataIn[3]), .B(n25095), .C(vectorInput[123]), .D(n25080
        ), .Z(n27261) );
    VMW_AO22 U866 ( .A(matrixInput[625]), .B(n25096), .C(matrixInput[617]), 
        .D(n25081), .Z(n26639) );
    VMW_FD \matrixInput_reg[972]  ( .D(n26284), .CP(Clk), .Q(matrixInput[972])
         );
    VMW_AO22 U1046 ( .A(matrixInput[463]), .B(n25096), .C(matrixInput[455]), 
        .D(n25081), .Z(n26801) );
    VMW_AO22 U1657 ( .A(matrixInput[1757]), .B(n25096), .C(matrixInput[1749]), 
        .D(n25081), .Z(n25507) );
    VMW_FD \matrixInput_reg[1012]  ( .D(n26244), .CP(Clk), .Q(matrixInput
        [1012]) );
    VMW_FD \vectorInput_reg[12]  ( .D(n27372), .CP(Clk), .Q(vectorInput[12])
         );
    VMW_FD \matrixInput_reg[605]  ( .D(n26651), .CP(Clk), .Q(matrixInput[605])
         );
    VMW_FD \matrixInput_reg[1795]  ( .D(n25461), .CP(Clk), .Q(matrixInput
        [1795]) );
    VMW_FD \matrixInput_reg[1496]  ( .D(n25760), .CP(Clk), .Q(matrixInput
        [1496]) );
    VMW_FD \matrixInput_reg[298]  ( .D(n26958), .CP(Clk), .Q(matrixInput[298])
         );
    VMW_FD \matrixInput_reg[281]  ( .D(n26975), .CP(Clk), .Q(matrixInput[281])
         );
    VMW_FD \matrixInput_reg[182]  ( .D(n27074), .CP(Clk), .Q(matrixInput[182])
         );
    VMW_FD \matrixInput_reg[1311]  ( .D(n25945), .CP(Clk), .Q(matrixInput
        [1311]) );
    VMW_FD \matrixInput_reg[1308]  ( .D(n25948), .CP(Clk), .Q(matrixInput
        [1308]) );
    VMW_AO22 U387 ( .A(vectorInput[40]), .B(n25095), .C(vectorInput[32]), .D(
        n25080), .Z(n27352) );
    VMW_AO22 U421 ( .A(vectorInput[125]), .B(n25095), .C(vectorInput[117]), 
        .D(n25080), .Z(n27267) );
    VMW_AO22 U528 ( .A(matrixInput[929]), .B(n25096), .C(matrixInput[921]), 
        .D(n25081), .Z(n26335) );
    VMW_AO22 U2076 ( .A(matrixInput[1379]), .B(n25096), .C(matrixInput[1371]), 
        .D(n25081), .Z(n25885) );
    VMW_FD \matrixInput_reg[506]  ( .D(n26750), .CP(Clk), .Q(matrixInput[506])
         );
    VMW_AO22 U618 ( .A(matrixInput[848]), .B(n25096), .C(matrixInput[840]), 
        .D(n25081), .Z(n26416) );
    VMW_AO22 U788 ( .A(matrixInput[696]), .B(n25096), .C(matrixInput[688]), 
        .D(n25081), .Z(n26568) );
    VMW_AO22 U1376 ( .A(matrixInput[2008]), .B(n25096), .C(matrixInput[2000]), 
        .D(n25081), .Z(n25256) );
    VMW_AO22 U1567 ( .A(matrixInput[190]), .B(n25096), .C(matrixInput[182]), 
        .D(n25081), .Z(n27074) );
    VMW_AO22 U1885 ( .A(matrixInput[1551]), .B(n25096), .C(matrixInput[1543]), 
        .D(n25081), .Z(n25713) );
    VMW_AO22 U1915 ( .A(matrixInput[1524]), .B(n25096), .C(matrixInput[1516]), 
        .D(n25081), .Z(n25740) );
    VMW_FD \matrixInput_reg[636]  ( .D(n26620), .CP(Clk), .Q(matrixInput[636])
         );
    VMW_FD \matrixInput_reg[1038]  ( .D(n26218), .CP(Clk), .Q(matrixInput
        [1038]) );
    VMW_FD \matrixInput_reg[1021]  ( .D(n26235), .CP(Clk), .Q(matrixInput
        [1021]) );
    VMW_AO22 U2346 ( .A(matrixInput[1136]), .B(n25096), .C(matrixInput[1128]), 
        .D(n25081), .Z(n26128) );
    VMW_AO22 U853 ( .A(matrixInput[637]), .B(n25096), .C(matrixInput[629]), 
        .D(n25081), .Z(n26627) );
    VMW_AO22 U948 ( .A(matrixInput[551]), .B(n25096), .C(matrixInput[543]), 
        .D(n25081), .Z(n26713) );
    VMW_AO22 U1054 ( .A(matrixInput[456]), .B(n25096), .C(matrixInput[448]), 
        .D(n25081), .Z(n26808) );
    VMW_AO22 U1061 ( .A(matrixInput[449]), .B(n25096), .C(matrixInput[441]), 
        .D(n25081), .Z(n26815) );
    VMW_AO22 U1351 ( .A(matrixInput[2031]), .B(n25096), .C(matrixInput[2023]), 
        .D(n25081), .Z(n25233) );
    VMW_AO22 U1932 ( .A(matrixInput[1508]), .B(n25096), .C(matrixInput[1500]), 
        .D(n25081), .Z(n25756) );
    VMW_AO22 U2557 ( .A(cOutput[88]), .B(n25089), .C(cOutput[72]), .D(n25088), 
        .Z(n25179) );
    VMW_FD \matrixInput_reg[1605]  ( .D(n25651), .CP(Clk), .Q(matrixInput
        [1605]) );
    VMW_FD \matrixInput_reg[1322]  ( .D(n25934), .CP(Clk), .Q(matrixInput
        [1322]) );
    VMW_FD \matrixInput_reg[535]  ( .D(n26721), .CP(Clk), .Q(matrixInput[535])
         );
    VMW_FD \matrixInput_reg[1298]  ( .D(n25958), .CP(Clk), .Q(matrixInput
        [1298]) );
    VMW_FD \matrixInput_reg[496]  ( .D(n26760), .CP(Clk), .Q(matrixInput[496])
         );
    VMW_AO22 U1540 ( .A(matrixInput[1862]), .B(n25096), .C(matrixInput[1854]), 
        .D(n25081), .Z(n25402) );
    VMW_FD \matrixInput_reg[1281]  ( .D(n25975), .CP(Clk), .Q(matrixInput
        [1281]) );
    VMW_AO22 U2361 ( .A(matrixInput[1122]), .B(n25096), .C(matrixInput[1114]), 
        .D(n25081), .Z(n26142) );
    VMW_OAI21 U2570 ( .A(n25114), .B(n25115), .C(n25094), .Z(n25075) );
    VMW_FD \matrixInput_reg[795]  ( .D(n26461), .CP(Clk), .Q(matrixInput[795])
         );
    VMW_FD \matrixInput_reg[1182]  ( .D(n26074), .CP(Clk), .Q(matrixInput
        [1182]) );
    VMW_FD \matrixInput_reg[1506]  ( .D(n25750), .CP(Clk), .Q(matrixInput
        [1506]) );
    VMW_FD \matrixInput_reg[311]  ( .D(n26945), .CP(Clk), .Q(matrixInput[311])
         );
    VMW_FD \matrixInput_reg[308]  ( .D(n26948), .CP(Clk), .Q(matrixInput[308])
         );
    VMW_AO22 U1670 ( .A(matrixInput[1745]), .B(n25096), .C(matrixInput[1737]), 
        .D(n25081), .Z(n25519) );
    VMW_AO22 U2051 ( .A(matrixInput[1402]), .B(n25096), .C(matrixInput[1394]), 
        .D(n25081), .Z(n25862) );
    VMW_FD \matrixInput_reg[1636]  ( .D(n25620), .CP(Clk), .Q(matrixInput
        [1636]) );
    VMW_FD \matrixInput_reg[1535]  ( .D(n25721), .CP(Clk), .Q(matrixInput
        [1535]) );
    VMW_FD \matrixInput_reg[322]  ( .D(n26934), .CP(Clk), .Q(matrixInput[322])
         );
    VMW_FD \matrixInput_reg[1450]  ( .D(n25806), .CP(Clk), .Q(matrixInput
        [1450]) );
    VMW_AO22 U1645 ( .A(matrixInput[183]), .B(n25096), .C(matrixInput[175]), 
        .D(n25081), .Z(n27081) );
    VMW_FD \matrixInput_reg[1449]  ( .D(n25807), .CP(Clk), .Q(matrixInput
        [1449]) );
    VMW_AO22 U2064 ( .A(matrixInput[1390]), .B(n25096), .C(matrixInput[1382]), 
        .D(n25081), .Z(n25874) );
    VMW_FD \matrixInput_reg[247]  ( .D(n27009), .CP(Clk), .Q(matrixInput[247])
         );
    VMW_FD \matrixInput_reg[1753]  ( .D(n25503), .CP(Clk), .Q(matrixInput
        [1753]) );
    VMW_FD \matrixInput_reg[144]  ( .D(n27112), .CP(Clk), .Q(matrixInput[144])
         );
    VMW_AO22 U1073 ( .A(matrixInput[438]), .B(n25096), .C(matrixInput[430]), 
        .D(n25081), .Z(n26826) );
    VMW_AO22 U1343 ( .A(matrixInput[2038]), .B(n25096), .C(matrixInput[2030]), 
        .D(n25081), .Z(n25226) );
    VMW_AO22 U1364 ( .A(matrixInput[2019]), .B(n25096), .C(matrixInput[2011]), 
        .D(n25081), .Z(n25245) );
    VMW_FD \matrixInput_reg[1463]  ( .D(n25793), .CP(Clk), .Q(matrixInput
        [1463]) );
    VMW_FD \matrixInput_reg[274]  ( .D(n26982), .CP(Clk), .Q(matrixInput[274])
         );
    VMW_AO22 U1552 ( .A(matrixInput[1851]), .B(n25096), .C(matrixInput[1843]), 
        .D(n25081), .Z(n25413) );
    VMW_AO22 U1575 ( .A(matrixInput[1830]), .B(n25096), .C(matrixInput[1822]), 
        .D(n25081), .Z(n25434) );
    VMW_AO22 U1897 ( .A(matrixInput[1540]), .B(n25096), .C(matrixInput[1532]), 
        .D(n25081), .Z(n25724) );
    VMW_AO22 U1907 ( .A(matrixInput[1531]), .B(n25096), .C(matrixInput[1523]), 
        .D(n25081), .Z(n25733) );
    VMW_AO22 U2354 ( .A(matrixInput[1128]), .B(n25096), .C(matrixInput[1120]), 
        .D(n25081), .Z(n26136) );
    VMW_AO22 U2545 ( .A(cOutput[49]), .B(n25087), .C(cOutput[33]), .D(n25084), 
        .Z(n25165) );
    VMW_FD \matrixInput_reg[177]  ( .D(n27079), .CP(Clk), .Q(matrixInput[177])
         );
    VMW_FD \matrixInput_reg[1779]  ( .D(n25477), .CP(Clk), .Q(matrixInput
        [1779]) );
    VMW_FD \matrixInput_reg[1760]  ( .D(n25496), .CP(Clk), .Q(matrixInput
        [1760]) );
    VMW_AO22 U1662 ( .A(matrixInput[1752]), .B(n25096), .C(matrixInput[1744]), 
        .D(n25081), .Z(n25512) );
    VMW_AO22 U1920 ( .A(matrixInput[1519]), .B(n25096), .C(matrixInput[1511]), 
        .D(n25081), .Z(n25745) );
    VMW_AO22 U2373 ( .A(matrixInput[1111]), .B(n25096), .C(matrixInput[1103]), 
        .D(n25081), .Z(n26153) );
    VMW_FD \matrixInput_reg[1247]  ( .D(n26009), .CP(Clk), .Q(matrixInput
        [1247]) );
    VMW_FD \matrixInput_reg[1144]  ( .D(n26112), .CP(Clk), .Q(matrixInput
        [1144]) );
    VMW_FD \matrixInput_reg[450]  ( .D(n26806), .CP(Clk), .Q(matrixInput[450])
         );
    VMW_FD \matrixInput_reg[449]  ( .D(n26807), .CP(Clk), .Q(matrixInput[449])
         );
    VMW_FD \matrixInput_reg[753]  ( .D(n26503), .CP(Clk), .Q(matrixInput[753])
         );
    VMW_NAND3 U2562 ( .A(WR), .B(n25083), .C(Addr[0]), .Z(n25080) );
    VMW_FD \matrixInput_reg[1274]  ( .D(n25982), .CP(Clk), .Q(matrixInput
        [1274]) );
    VMW_FD \matrixInput_reg[463]  ( .D(n26793), .CP(Clk), .Q(matrixInput[463])
         );
    VMW_AO22 U2043 ( .A(matrixInput[1408]), .B(n25096), .C(matrixInput[1400]), 
        .D(n25081), .Z(n25856) );
    VMW_FD \matrixInput_reg[1177]  ( .D(n26079), .CP(Clk), .Q(matrixInput
        [1177]) );
    VMW_FD \matrixInput_reg[779]  ( .D(n26477), .CP(Clk), .Q(matrixInput[779])
         );
    VMW_FD \matrixInput_reg[760]  ( .D(n26496), .CP(Clk), .Q(matrixInput[760])
         );
    VMW_FD \matrixInput_reg[1987]  ( .D(n25269), .CP(Clk), .Q(matrixInput
        [1987]) );
    VMW_FD \matrixInput_reg[57]  ( .D(n27199), .CP(Clk), .Q(matrixInput[57])
         );
    VMW_AO22 U681 ( .A(matrixInput[792]), .B(n25096), .C(matrixInput[784]), 
        .D(n25081), .Z(n26472) );
    VMW_FD \matrixInput_reg[817]  ( .D(n26439), .CP(Clk), .Q(matrixInput[817])
         );
    VMW_AO22 U711 ( .A(matrixInput[765]), .B(n25096), .C(matrixInput[757]), 
        .D(n25081), .Z(n26499) );
    VMW_AO22 U736 ( .A(matrixInput[742]), .B(n25096), .C(matrixInput[734]), 
        .D(n25081), .Z(n26522) );
    VMW_FD \matrixInput_reg[824]  ( .D(n26432), .CP(Clk), .Q(matrixInput[824])
         );
    VMW_FD \matrixInput_reg[64]  ( .D(n27192), .CP(Clk), .Q(matrixInput[64])
         );
    VMW_AO22 U874 ( .A(matrixInput[68]), .B(n25096), .C(matrixInput[60]), .D(
        n25081), .Z(n27196) );
    VMW_AO22 U1258 ( .A(matrixInput[272]), .B(n25096), .C(matrixInput[264]), 
        .D(n25081), .Z(n26992) );
    VMW_AO22 U2268 ( .A(matrixInput[1207]), .B(n25096), .C(matrixInput[1199]), 
        .D(n25081), .Z(n26057) );
    VMW_AO22 U2479 ( .A(matrixInput[1016]), .B(n25096), .C(matrixInput[1008]), 
        .D(n25081), .Z(n26248) );
    VMW_FD \matrixInput_reg[987]  ( .D(n26269), .CP(Clk), .Q(matrixInput[987])
         );
    VMW_FD \matrixInput_reg[1817]  ( .D(n25439), .CP(Clk), .Q(matrixInput
        [1817]) );
    VMW_AO22 U1449 ( .A(matrixInput[1944]), .B(n25096), .C(matrixInput[1936]), 
        .D(n25081), .Z(n25320) );
    VMW_AO22 U406 ( .A(vectorInput[23]), .B(n25095), .C(vectorInput[15]), .D(
        n25080), .Z(n27369) );
    VMW_AO22 U596 ( .A(matrixInput[868]), .B(n25096), .C(matrixInput[860]), 
        .D(n25081), .Z(n26396) );
    VMW_AO22 U2158 ( .A(matrixInput[1306]), .B(n25096), .C(matrixInput[1298]), 
        .D(n25081), .Z(n25958) );
    VMW_AO22 U758 ( .A(matrixInput[722]), .B(n25096), .C(matrixInput[714]), 
        .D(n25081), .Z(n26542) );
    VMW_AO22 U1168 ( .A(matrixInput[353]), .B(n25096), .C(matrixInput[345]), 
        .D(n25081), .Z(n26911) );
    VMW_AO22 U1779 ( .A(matrixInput[1647]), .B(n25096), .C(matrixInput[1639]), 
        .D(n25081), .Z(n25617) );
    VMW_AO22 U2206 ( .A(matrixInput[1262]), .B(n25096), .C(matrixInput[1254]), 
        .D(n25081), .Z(n26002) );
    VMW_OAI21 U2587 ( .A(n25163), .B(n25164), .C(n25090), .Z(n25172) );
    VMW_FD \matrixInput_reg[1824]  ( .D(n25432), .CP(Clk), .Q(matrixInput
        [1824]) );
    VMW_FD \matrixInput_reg[538]  ( .D(n26718), .CP(Clk), .Q(matrixInput[538])
         );
    VMW_AO22 U1236 ( .A(matrixInput[292]), .B(n25096), .C(matrixInput[284]), 
        .D(n25081), .Z(n26972) );
    VMW_AO22 U1427 ( .A(matrixInput[1964]), .B(n25096), .C(matrixInput[1956]), 
        .D(n25081), .Z(n25300) );
    VMW_AO22 U2396 ( .A(matrixInput[1091]), .B(n25096), .C(matrixInput[1083]), 
        .D(n25081), .Z(n26173) );
    VMW_AO22 U2417 ( .A(matrixInput[1072]), .B(n25096), .C(matrixInput[1064]), 
        .D(n25081), .Z(n26192) );
    VMW_FD \matrixInput_reg[521]  ( .D(n26735), .CP(Clk), .Q(matrixInput[521])
         );
    VMW_FD \matrixInput_reg[1336]  ( .D(n25920), .CP(Clk), .Q(matrixInput
        [1336]) );
    VMW_FD \holder_reg[3]  ( .D(n27389), .CP(Clk), .Q(\holder[3] ) );
    VMW_FD \matrixInput_reg[622]  ( .D(n26634), .CP(Clk), .Q(matrixInput[622])
         );
    VMW_AO22 U1855 ( .A(matrixInput[1578]), .B(n25096), .C(matrixInput[1570]), 
        .D(n25081), .Z(n25686) );
    VMW_FD \matrixInput_reg[1035]  ( .D(n26221), .CP(Clk), .Q(matrixInput
        [1035]) );
    VMW_FD \matrixInput_reg[1305]  ( .D(n25951), .CP(Clk), .Q(matrixInput
        [1305]) );
    VMW_AO22 U345 ( .A(vectorInput[78]), .B(n25095), .C(vectorInput[70]), .D(
        n25080), .Z(n27314) );
    VMW_AO22 U362 ( .A(vectorInput[63]), .B(n25095), .C(vectorInput[55]), .D(
        n25080), .Z(n27329) );
    VMW_AO22 U468 ( .A(matrixInput[984]), .B(n25096), .C(matrixInput[976]), 
        .D(n25081), .Z(n26280) );
    VMW_AO22 U2136 ( .A(matrixInput[1325]), .B(n25096), .C(matrixInput[1317]), 
        .D(n25081), .Z(n25939) );
    VMW_FD \matrixInput_reg[512]  ( .D(n26744), .CP(Clk), .Q(matrixInput[512])
         );
    VMW_AO22 U573 ( .A(matrixInput[889]), .B(n25096), .C(matrixInput[881]), 
        .D(n25081), .Z(n26375) );
    VMW_AO22 U643 ( .A(matrixInput[826]), .B(n25096), .C(matrixInput[818]), 
        .D(n25081), .Z(n26438) );
    VMW_AO22 U1096 ( .A(matrixInput[48]), .B(n25096), .C(matrixInput[40]), .D(
        n25081), .Z(n27216) );
    VMW_FD \matrixInput_reg[1798]  ( .D(n25458), .CP(Clk), .Q(matrixInput
        [1798]) );
    VMW_FD \matrixInput_reg[1781]  ( .D(n25475), .CP(Clk), .Q(matrixInput
        [1781]) );
    VMW_FD \matrixInput_reg[196]  ( .D(n27060), .CP(Clk), .Q(matrixInput[196])
         );
    VMW_FD \matrixInput_reg[1482]  ( .D(n25774), .CP(Clk), .Q(matrixInput
        [1482]) );
    VMW_FD \matrixInput_reg[295]  ( .D(n26961), .CP(Clk), .Q(matrixInput[295])
         );
    VMW_FD \matrixInput_reg[1006]  ( .D(n26250), .CP(Clk), .Q(matrixInput
        [1006]) );
    VMW_AO22 U1106 ( .A(matrixInput[408]), .B(n25096), .C(matrixInput[400]), 
        .D(n25081), .Z(n26856) );
    VMW_AO22 U1717 ( .A(matrixInput[1703]), .B(n25096), .C(matrixInput[1695]), 
        .D(n25081), .Z(n25561) );
    VMW_FD \matrixInput_reg[611]  ( .D(n26645), .CP(Clk), .Q(matrixInput[611])
         );
    VMW_AO22 U1121 ( .A(matrixInput[396]), .B(n25096), .C(matrixInput[388]), 
        .D(n25081), .Z(n26868) );
    VMW_AO22 U1687 ( .A(matrixInput[1729]), .B(n25096), .C(matrixInput[1721]), 
        .D(n25081), .Z(n25535) );
    VMW_FD \matrixInput_reg[608]  ( .D(n26648), .CP(Clk), .Q(matrixInput[608])
         );
    VMW_AO22 U2081 ( .A(matrixInput[1375]), .B(n25096), .C(matrixInput[1367]), 
        .D(n25081), .Z(n25889) );
    VMW_AO22 U2111 ( .A(matrixInput[141]), .B(n25096), .C(matrixInput[133]), 
        .D(n25081), .Z(n27123) );
    VMW_FD \matrixInput_reg[2045]  ( .D(n25211), .CP(Clk), .Q(matrixInput
        [2045]) );
    VMW_FD \matrixInput_reg[1622]  ( .D(n25634), .CP(Clk), .Q(matrixInput
        [1622]) );
    VMW_FD \matrixInput_reg[1538]  ( .D(n25718), .CP(Clk), .Q(matrixInput
        [1538]) );
    VMW_FD \matrixInput_reg[336]  ( .D(n26920), .CP(Clk), .Q(matrixInput[336])
         );
    VMW_FD \matrixInput_reg[1521]  ( .D(n25735), .CP(Clk), .Q(matrixInput
        [1521]) );
    VMW_AO22 U1211 ( .A(matrixInput[314]), .B(n25096), .C(matrixInput[306]), 
        .D(n25081), .Z(n26950) );
    VMW_AO22 U1590 ( .A(matrixInput[1817]), .B(n25096), .C(matrixInput[1809]), 
        .D(n25081), .Z(n25447) );
    VMW_AO22 U1730 ( .A(matrixInput[1691]), .B(n25096), .C(matrixInput[1683]), 
        .D(n25081), .Z(n25573) );
    VMW_AO22 U2221 ( .A(matrixInput[1248]), .B(n25096), .C(matrixInput[1240]), 
        .D(n25081), .Z(n26016) );
    VMW_AO22 U2430 ( .A(matrixInput[1060]), .B(n25096), .C(matrixInput[1052]), 
        .D(n25081), .Z(n26204) );
    VMW_FD \matrixInput_reg[1512]  ( .D(n25744), .CP(Clk), .Q(matrixInput
        [1512]) );
    VMW_FD \matrixInput_reg[798]  ( .D(n26458), .CP(Clk), .Q(matrixInput[798])
         );
    VMW_FD \matrixInput_reg[781]  ( .D(n26475), .CP(Clk), .Q(matrixInput[781])
         );
    VMW_FD \matrixInput_reg[305]  ( .D(n26951), .CP(Clk), .Q(matrixInput[305])
         );
    VMW_FD \matrixInput_reg[1196]  ( .D(n26060), .CP(Clk), .Q(matrixInput
        [1196]) );
    VMW_FD \matrixInput_reg[482]  ( .D(n26774), .CP(Clk), .Q(matrixInput[482])
         );
    VMW_AO22 U1381 ( .A(matrixInput[2006]), .B(n25096), .C(matrixInput[1998]), 
        .D(n25081), .Z(n25258) );
    VMW_AO22 U1400 ( .A(matrixInput[1988]), .B(n25096), .C(matrixInput[1980]), 
        .D(n25081), .Z(n25276) );
    VMW_FD \matrixInput_reg[1295]  ( .D(n25961), .CP(Clk), .Q(matrixInput
        [1295]) );
    VMW_AO22 U1872 ( .A(matrixInput[1563]), .B(n25096), .C(matrixInput[1555]), 
        .D(n25081), .Z(n25701) );
    VMW_FD \matrixInput_reg[1611]  ( .D(n25645), .CP(Clk), .Q(matrixInput
        [1611]) );
    VMW_FD \matrixInput_reg[1608]  ( .D(n25648), .CP(Clk), .Q(matrixInput
        [1608]) );
    VMW_AO22 U891 ( .A(matrixInput[603]), .B(n25096), .C(matrixInput[595]), 
        .D(n25081), .Z(n26661) );
    VMW_AO22 U901 ( .A(matrixInput[594]), .B(n25096), .C(matrixInput[586]), 
        .D(n25081), .Z(n26670) );
    VMW_FD \matrixInput_reg[1966]  ( .D(n25290), .CP(Clk), .Q(matrixInput
        [1966]) );
    VMW_FD \matrixInput_reg[1955]  ( .D(n25301), .CP(Clk), .Q(matrixInput
        [1955]) );
    VMW_FD \matrixInput_reg[85]  ( .D(n27171), .CP(Clk), .Q(matrixInput[85])
         );
    VMW_AO22 U926 ( .A(matrixInput[571]), .B(n25096), .C(matrixInput[563]), 
        .D(n25081), .Z(n26693) );
    VMW_FD \matrixInput_reg[966]  ( .D(n26290), .CP(Clk), .Q(matrixInput[966])
         );
    VMW_AO22 U379 ( .A(vectorInput[11]), .B(n25095), .C(vectorInput[3]), .D(
        n25080), .Z(n27381) );
    VMW_AO22 U554 ( .A(matrixInput[907]), .B(n25096), .C(matrixInput[899]), 
        .D(n25081), .Z(n26357) );
    VMW_AO22 U568 ( .A(matrixInput[894]), .B(n25096), .C(matrixInput[886]), 
        .D(n25081), .Z(n26370) );
    VMW_AO22 U664 ( .A(matrixInput[87]), .B(n25096), .C(matrixInput[79]), .D(
        n25081), .Z(n27177) );
    VMW_AO22 U1969 ( .A(matrixInput[1476]), .B(n25096), .C(matrixInput[1468]), 
        .D(n25081), .Z(n25788) );
    VMW_FD \vectorInput_reg[35]  ( .D(n27349), .CP(Clk), .Q(vectorInput[35])
         );
    VMW_AO22 U1021 ( .A(matrixInput[486]), .B(n25096), .C(matrixInput[478]), 
        .D(n25081), .Z(n26778) );
    VMW_AO22 U1281 ( .A(matrixInput[251]), .B(n25096), .C(matrixInput[243]), 
        .D(n25081), .Z(n27013) );
    VMW_AO22 U1500 ( .A(matrixInput[1898]), .B(n25096), .C(matrixInput[1890]), 
        .D(n25081), .Z(n25366) );
    VMW_AO22 U2321 ( .A(matrixInput[1158]), .B(n25096), .C(matrixInput[1150]), 
        .D(n25081), .Z(n26106) );
    VMW_FD \matrixInput_reg[1502]  ( .D(n25754), .CP(Clk), .Q(matrixInput
        [1502]) );
    VMW_FD \matrixInput_reg[955]  ( .D(n26301), .CP(Clk), .Q(matrixInput[955])
         );
    VMW_FD \matrixInput_reg[315]  ( .D(n26941), .CP(Clk), .Q(matrixInput[315])
         );
    VMW_AO22 U2530 ( .A(cOutput[91]), .B(n25089), .C(cOutput[75]), .D(n25088), 
        .Z(n25146) );
    VMW_FD \matrixInput_reg[1186]  ( .D(n26070), .CP(Clk), .Q(matrixInput
        [1186]) );
    VMW_FD \matrixInput_reg[791]  ( .D(n26465), .CP(Clk), .Q(matrixInput[791])
         );
    VMW_FD \matrixInput_reg[788]  ( .D(n26468), .CP(Clk), .Q(matrixInput[788])
         );
    VMW_FD \matrixInput_reg[1285]  ( .D(n25971), .CP(Clk), .Q(matrixInput
        [1285]) );
    VMW_AO22 U1311 ( .A(matrixInput[224]), .B(n25096), .C(matrixInput[216]), 
        .D(n25081), .Z(n27040) );
    VMW_AO22 U1490 ( .A(matrixInput[197]), .B(n25096), .C(matrixInput[189]), 
        .D(n25081), .Z(n27067) );
    VMW_AO22 U1630 ( .A(matrixInput[1781]), .B(n25096), .C(matrixInput[1773]), 
        .D(n25081), .Z(n25483) );
    VMW_AO22 U1972 ( .A(matrixInput[1473]), .B(n25096), .C(matrixInput[1465]), 
        .D(n25081), .Z(n25791) );
    VMW_FD \matrixInput_reg[492]  ( .D(n26764), .CP(Clk), .Q(matrixInput[492])
         );
    VMW_AO22 U2011 ( .A(matrixInput[150]), .B(n25096), .C(matrixInput[142]), 
        .D(n25081), .Z(n27114) );
    VMW_FD \matrixInput_reg[1618]  ( .D(n25638), .CP(Clk), .Q(matrixInput
        [1618]) );
    VMW_FD \matrixInput_reg[1601]  ( .D(n25655), .CP(Clk), .Q(matrixInput
        [1601]) );
    VMW_AO22 U2181 ( .A(matrixInput[1285]), .B(n25096), .C(matrixInput[1277]), 
        .D(n25081), .Z(n25979) );
    VMW_INV U2600 ( .A(\holder[1] ), .Z(n25059) );
    VMW_FD \matrixInput_reg[1632]  ( .D(n25624), .CP(Clk), .Q(matrixInput
        [1632]) );
    VMW_FD \matrixInput_reg[1531]  ( .D(n25725), .CP(Clk), .Q(matrixInput
        [1531]) );
    VMW_FD \matrixInput_reg[1528]  ( .D(n25728), .CP(Clk), .Q(matrixInput
        [1528]) );
    VMW_FD \matrixInput_reg[326]  ( .D(n26930), .CP(Clk), .Q(matrixInput[326])
         );
    VMW_FD \matrixInput_reg[502]  ( .D(n26754), .CP(Clk), .Q(matrixInput[502])
         );
    VMW_BUFIZ U2627 ( .A(n25200), .E(RD), .Z(\DataOut[20]1 ) );
    VMW_AO22 U454 ( .A(matrixInput[997]), .B(n25096), .C(matrixInput[989]), 
        .D(n25081), .Z(n26267) );
    VMW_AO22 U658 ( .A(matrixInput[812]), .B(n25096), .C(matrixInput[804]), 
        .D(n25081), .Z(n26452) );
    VMW_AO22 U1006 ( .A(matrixInput[499]), .B(n25096), .C(matrixInput[491]), 
        .D(n25081), .Z(n26765) );
    VMW_AO22 U2036 ( .A(matrixInput[1415]), .B(n25096), .C(matrixInput[1407]), 
        .D(n25081), .Z(n25849) );
    VMW_FD \matrixInput_reg[1791]  ( .D(n25465), .CP(Clk), .Q(matrixInput
        [1791]) );
    VMW_FD \matrixInput_reg[1788]  ( .D(n25468), .CP(Clk), .Q(matrixInput
        [1788]) );
    VMW_FD \matrixInput_reg[1315]  ( .D(n25941), .CP(Clk), .Q(matrixInput
        [1315]) );
    VMW_FD \matrixInput_reg[1492]  ( .D(n25764), .CP(Clk), .Q(matrixInput
        [1492]) );
    VMW_FD \matrixInput_reg[186]  ( .D(n27070), .CP(Clk), .Q(matrixInput[186])
         );
    VMW_FD \matrixInput_reg[285]  ( .D(n26971), .CP(Clk), .Q(matrixInput[285])
         );
    VMW_AO22 U1196 ( .A(matrixInput[39]), .B(n25096), .C(matrixInput[31]), .D(
        n25081), .Z(n27225) );
    VMW_AO22 U1787 ( .A(matrixInput[1639]), .B(n25096), .C(matrixInput[1631]), 
        .D(n25081), .Z(n25625) );
    VMW_FD \matrixInput_reg[618]  ( .D(n26638), .CP(Clk), .Q(matrixInput[618])
         );
    VMW_AO22 U1617 ( .A(matrixInput[1793]), .B(n25096), .C(matrixInput[1785]), 
        .D(n25081), .Z(n25471) );
    VMW_FD \matrixInput_reg[601]  ( .D(n26655), .CP(Clk), .Q(matrixInput[601])
         );
    VMW_FD \matrixInput_reg[1326]  ( .D(n25930), .CP(Clk), .Q(matrixInput
        [1326]) );
    VMW_FD \matrixInput_reg[1016]  ( .D(n26240), .CP(Clk), .Q(matrixInput
        [1016]) );
    VMW_AO22 U764 ( .A(matrixInput[717]), .B(n25096), .C(matrixInput[709]), 
        .D(n25081), .Z(n26547) );
    VMW_AO22 U1336 ( .A(matrixInput[2045]), .B(n25096), .C(matrixInput[2037]), 
        .D(n25081), .Z(n25219) );
    VMW_AO22 U2296 ( .A(matrixInput[1181]), .B(n25096), .C(matrixInput[1173]), 
        .D(n25081), .Z(n26083) );
    VMW_AO22 U2517 ( .A(cOutput[28]), .B(n25089), .C(cOutput[12]), .D(n25088), 
        .Z(n25131) );
    VMW_FD \matrixInput_reg[531]  ( .D(n26725), .CP(Clk), .Q(matrixInput[531])
         );
    VMW_AO22 U2306 ( .A(matrixInput[1172]), .B(n25096), .C(matrixInput[1164]), 
        .D(n25081), .Z(n26092) );
    VMW_AO22 U2487 ( .A(matrixInput[1008]), .B(n25096), .C(matrixInput[1000]), 
        .D(n25081), .Z(n26256) );
    VMW_FD \matrixInput_reg[528]  ( .D(n26728), .CP(Clk), .Q(matrixInput[528])
         );
    VMW_FD \matrixInput_reg[1025]  ( .D(n26231), .CP(Clk), .Q(matrixInput
        [1025]) );
    VMW_AO22 U1527 ( .A(matrixInput[1874]), .B(n25096), .C(matrixInput[1866]), 
        .D(n25081), .Z(n25390) );
    VMW_AO22 U1869 ( .A(matrixInput[1566]), .B(n25096), .C(matrixInput[1558]), 
        .D(n25081), .Z(n25698) );
    VMW_AO22 U1955 ( .A(matrixInput[1488]), .B(n25096), .C(matrixInput[1480]), 
        .D(n25081), .Z(n25776) );
    VMW_FD \matrixInput_reg[632]  ( .D(n26624), .CP(Clk), .Q(matrixInput[632])
         );
    VMW_FD \vectorInput_reg[25]  ( .D(n27359), .CP(Clk), .Q(vectorInput[25])
         );
    VMW_AO22 U826 ( .A(matrixInput[661]), .B(n25096), .C(matrixInput[653]), 
        .D(n25081), .Z(n26603) );
    VMW_FD \matrixInput_reg[976]  ( .D(n26280), .CP(Clk), .Q(matrixInput[976])
         );
    VMW_FD \matrixInput_reg[945]  ( .D(n26311), .CP(Clk), .Q(matrixInput[945])
         );
    VMW_FD \vectorInput_reg[16]  ( .D(n27368), .CP(Clk), .Q(vectorInput[16])
         );
    VMW_AO22 U473 ( .A(matrixInput[979]), .B(n25096), .C(matrixInput[971]), 
        .D(n25081), .Z(n26285) );
    VMW_AO22 U801 ( .A(matrixInput[684]), .B(n25096), .C(matrixInput[676]), 
        .D(n25081), .Z(n26580) );
    VMW_AO22 U991 ( .A(matrixInput[512]), .B(n25096), .C(matrixInput[504]), 
        .D(n25081), .Z(n26752) );
    VMW_AO22 U743 ( .A(matrixInput[736]), .B(n25096), .C(matrixInput[728]), 
        .D(n25081), .Z(n26528) );
    VMW_FD \matrixInput_reg[1976]  ( .D(n25280), .CP(Clk), .Q(matrixInput
        [1976]) );
    VMW_FD \matrixInput_reg[1945]  ( .D(n25311), .CP(Clk), .Q(matrixInput
        [1945]) );
    VMW_FD \matrixInput_reg[95]  ( .D(n27161), .CP(Clk), .Q(matrixInput[95])
         );
    VMW_AO22 U1173 ( .A(matrixInput[348]), .B(n25096), .C(matrixInput[340]), 
        .D(n25081), .Z(n26916) );
    VMW_FD \matrixInput_reg[1264]  ( .D(n25992), .CP(Clk), .Q(matrixInput
        [1264]) );
    VMW_FD \matrixInput_reg[473]  ( .D(n26783), .CP(Clk), .Q(matrixInput[473])
         );
    VMW_AO22 U1243 ( .A(matrixInput[286]), .B(n25096), .C(matrixInput[278]), 
        .D(n25081), .Z(n26978) );
    VMW_AO22 U1762 ( .A(matrixInput[1662]), .B(n25096), .C(matrixInput[1654]), 
        .D(n25081), .Z(n25602) );
    VMW_AO22 U2143 ( .A(matrixInput[1318]), .B(n25096), .C(matrixInput[1310]), 
        .D(n25081), .Z(n25946) );
    VMW_FD \matrixInput_reg[1167]  ( .D(n26089), .CP(Clk), .Q(matrixInput
        [1167]) );
    VMW_FD \matrixInput_reg[770]  ( .D(n26486), .CP(Clk), .Q(matrixInput[770])
         );
    VMW_FD \matrixInput_reg[769]  ( .D(n26487), .CP(Clk), .Q(matrixInput[769])
         );
    VMW_AO22 U1264 ( .A(matrixInput[267]), .B(n25096), .C(matrixInput[259]), 
        .D(n25081), .Z(n26997) );
    VMW_AO22 U1452 ( .A(matrixInput[1941]), .B(n25096), .C(matrixInput[1933]), 
        .D(n25081), .Z(n25323) );
    VMW_AO22 U1475 ( .A(matrixInput[1920]), .B(n25096), .C(matrixInput[1912]), 
        .D(n25081), .Z(n25344) );
    VMW_AO22 U1820 ( .A(matrixInput[1609]), .B(n25096), .C(matrixInput[1601]), 
        .D(n25081), .Z(n25655) );
    VMW_FD \matrixInput_reg[1257]  ( .D(n25999), .CP(Clk), .Q(matrixInput
        [1257]) );
    VMW_FD \matrixInput_reg[459]  ( .D(n26797), .CP(Clk), .Q(matrixInput[459])
         );
    VMW_FD \matrixInput_reg[440]  ( .D(n26816), .CP(Clk), .Q(matrixInput[440])
         );
    VMW_AO22 U2273 ( .A(matrixInput[1202]), .B(n25096), .C(matrixInput[1194]), 
        .D(n25081), .Z(n26062) );
    VMW_AO22 U2462 ( .A(matrixInput[1031]), .B(n25096), .C(matrixInput[1023]), 
        .D(n25081), .Z(n26233) );
    VMW_FD \matrixInput_reg[1154]  ( .D(n26102), .CP(Clk), .Q(matrixInput
        [1154]) );
    VMW_FD \matrixInput_reg[743]  ( .D(n26513), .CP(Clk), .Q(matrixInput[743])
         );
    VMW_FD \matrixInput_reg[1473]  ( .D(n25783), .CP(Clk), .Q(matrixInput
        [1473]) );
    VMW_AO22 U1807 ( .A(matrixInput[1621]), .B(n25096), .C(matrixInput[1613]), 
        .D(n25081), .Z(n25643) );
    VMW_FD \matrixInput_reg[264]  ( .D(n26992), .CP(Clk), .Q(matrixInput[264])
         );
    VMW_AO22 U1997 ( .A(matrixInput[1450]), .B(n25096), .C(matrixInput[1442]), 
        .D(n25081), .Z(n25814) );
    VMW_PULLDOWN U267 ( .Z(n25185) );
    VMW_PULLDOWN U269 ( .Z(n25187) );
    VMW_PULLDOWN U287 ( .Z(n25205) );
    VMW_AO22 U317 ( .A(vectorInput[104]), .B(n25095), .C(vectorInput[96]), .D(
        n25080), .Z(n27288) );
    VMW_AO22 U848 ( .A(matrixInput[641]), .B(n25096), .C(matrixInput[633]), 
        .D(n25081), .Z(n26623) );
    VMW_AO22 U1154 ( .A(matrixInput[366]), .B(n25096), .C(matrixInput[358]), 
        .D(n25081), .Z(n26898) );
    VMW_AO22 U1745 ( .A(matrixInput[174]), .B(n25096), .C(matrixInput[166]), 
        .D(n25081), .Z(n27090) );
    VMW_AO22 U2254 ( .A(matrixInput[1218]), .B(n25096), .C(matrixInput[1210]), 
        .D(n25081), .Z(n26046) );
    VMW_AO22 U2445 ( .A(matrixInput[1047]), .B(n25096), .C(matrixInput[1039]), 
        .D(n25081), .Z(n26217) );
    VMW_FD \matrixInput_reg[1770]  ( .D(n25486), .CP(Clk), .Q(matrixInput
        [1770]) );
    VMW_FD \matrixInput_reg[1769]  ( .D(n25487), .CP(Clk), .Q(matrixInput
        [1769]) );
    VMW_FD \matrixInput_reg[1459]  ( .D(n25797), .CP(Clk), .Q(matrixInput
        [1459]) );
    VMW_FD \matrixInput_reg[257]  ( .D(n26999), .CP(Clk), .Q(matrixInput[257])
         );
    VMW_FD \matrixInput_reg[167]  ( .D(n27089), .CP(Clk), .Q(matrixInput[167])
         );
    VMW_FD \matrixInput_reg[1440]  ( .D(n25816), .CP(Clk), .Q(matrixInput
        [1440]) );
    VMW_AO22 U2164 ( .A(matrixInput[1300]), .B(n25096), .C(matrixInput[1292]), 
        .D(n25081), .Z(n25964) );
    VMW_FD \matrixInput_reg[154]  ( .D(n27102), .CP(Clk), .Q(matrixInput[154])
         );
    VMW_FD \matrixInput_reg[1743]  ( .D(n25513), .CP(Clk), .Q(matrixInput
        [1743]) );
    VMW_AO22 U974 ( .A(matrixInput[59]), .B(n25096), .C(matrixInput[51]), .D(
        n25081), .Z(n27205) );
    VMW_AO22 U496 ( .A(matrixInput[958]), .B(n25096), .C(matrixInput[950]), 
        .D(n25081), .Z(n26306) );
    VMW_AO22 U2058 ( .A(matrixInput[1396]), .B(n25096), .C(matrixInput[1388]), 
        .D(n25081), .Z(n25868) );
    VMW_AO22 U330 ( .A(vectorInput[92]), .B(n25095), .C(vectorInput[84]), .D(
        n25080), .Z(n27300) );
    VMW_AO22 U506 ( .A(matrixInput[949]), .B(n25096), .C(matrixInput[941]), 
        .D(n25081), .Z(n26315) );
    VMW_AO22 U521 ( .A(matrixInput[936]), .B(n25096), .C(matrixInput[928]), 
        .D(n25081), .Z(n26328) );
    VMW_AO22 U611 ( .A(matrixInput[855]), .B(n25096), .C(matrixInput[847]), 
        .D(n25081), .Z(n26409) );
    VMW_AO22 U636 ( .A(matrixInput[832]), .B(n25096), .C(matrixInput[824]), 
        .D(n25081), .Z(n26432) );
    VMW_AO22 U1068 ( .A(matrixInput[443]), .B(n25096), .C(matrixInput[435]), 
        .D(n25081), .Z(n26821) );
    VMW_AO22 U1679 ( .A(matrixInput[1737]), .B(n25096), .C(matrixInput[1729]), 
        .D(n25081), .Z(n25527) );
    VMW_AO22 U2368 ( .A(matrixInput[1116]), .B(n25096), .C(matrixInput[1108]), 
        .D(n25081), .Z(n26148) );
    VMW_FD \matrixInput_reg[1834]  ( .D(n25422), .CP(Clk), .Q(matrixInput
        [1834]) );
    VMW_AO22 U1358 ( .A(matrixInput[2025]), .B(n25096), .C(matrixInput[2017]), 
        .D(n25081), .Z(n25239) );
    VMW_AO22 U1549 ( .A(matrixInput[1854]), .B(n25096), .C(matrixInput[1846]), 
        .D(n25081), .Z(n25410) );
    VMW_OAI21 U2579 ( .A(n25141), .B(n25142), .C(n25090), .Z(n25150) );
    VMW_FD \matrixInput_reg[1807]  ( .D(n25449), .CP(Clk), .Q(matrixInput
        [1807]) );
    VMW_FD \matrixInput_reg[997]  ( .D(n26259), .CP(Clk), .Q(matrixInput[997])
         );
    VMW_AO22 U781 ( .A(matrixInput[702]), .B(n25096), .C(matrixInput[694]), 
        .D(n25081), .Z(n26562) );
    VMW_AO22 U953 ( .A(matrixInput[547]), .B(n25096), .C(matrixInput[539]), 
        .D(n25081), .Z(n26717) );
    VMW_FD \matrixInput_reg[1997]  ( .D(n25259), .CP(Clk), .Q(matrixInput
        [1997]) );
    VMW_FD \matrixInput_reg[834]  ( .D(n26422), .CP(Clk), .Q(matrixInput[834])
         );
    VMW_FD \matrixInput_reg[74]  ( .D(n27182), .CP(Clk), .Q(matrixInput[74])
         );
    VMW_FD \matrixInput_reg[47]  ( .D(n27209), .CP(Clk), .Q(matrixInput[47])
         );
    VMW_AO22 U397 ( .A(vectorInput[31]), .B(n25095), .C(vectorInput[23]), .D(
        n25080), .Z(n27361) );
    VMW_AO22 U586 ( .A(matrixInput[94]), .B(n25096), .C(matrixInput[86]), .D(
        n25081), .Z(n27170) );
    VMW_AO22 U726 ( .A(matrixInput[751]), .B(n25096), .C(matrixInput[743]), 
        .D(n25081), .Z(n26513) );
    VMW_AO22 U958 ( .A(matrixInput[542]), .B(n25096), .C(matrixInput[534]), 
        .D(n25081), .Z(n26722) );
    VMW_AO22 U1063 ( .A(matrixInput[51]), .B(n25096), .C(matrixInput[43]), .D(
        n25081), .Z(n27213) );
    VMW_AO22 U1353 ( .A(matrixInput[2029]), .B(n25096), .C(matrixInput[2021]), 
        .D(n25081), .Z(n25235) );
    VMW_AO22 U2363 ( .A(matrixInput[1120]), .B(n25096), .C(matrixInput[1112]), 
        .D(n25081), .Z(n26144) );
    VMW_OAI21 U2572 ( .A(n25121), .B(n25122), .C(n25091), .Z(n25127) );
    VMW_FD \matrixInput_reg[1145]  ( .D(n26111), .CP(Clk), .Q(matrixInput
        [1145]) );
    VMW_FD \matrixInput_reg[807]  ( .D(n26449), .CP(Clk), .Q(matrixInput[807])
         );
    VMW_FD \matrixInput_reg[752]  ( .D(n26504), .CP(Clk), .Q(matrixInput[752])
         );
    VMW_AO22 U1542 ( .A(matrixInput[1860]), .B(n25096), .C(matrixInput[1852]), 
        .D(n25081), .Z(n25404) );
    VMW_AO22 U1930 ( .A(matrixInput[1510]), .B(n25096), .C(matrixInput[1502]), 
        .D(n25081), .Z(n25754) );
    VMW_FD \matrixInput_reg[1246]  ( .D(n26010), .CP(Clk), .Q(matrixInput
        [1246]) );
    VMW_FD \matrixInput_reg[451]  ( .D(n26805), .CP(Clk), .Q(matrixInput[451])
         );
    VMW_FD \matrixInput_reg[448]  ( .D(n26808), .CP(Clk), .Q(matrixInput[448])
         );
    VMW_AO22 U2053 ( .A(matrixInput[1400]), .B(n25096), .C(matrixInput[1392]), 
        .D(n25081), .Z(n25864) );
    VMW_FD \matrixInput_reg[1275]  ( .D(n25981), .CP(Clk), .Q(matrixInput
        [1275]) );
    VMW_FD \matrixInput_reg[1176]  ( .D(n26080), .CP(Clk), .Q(matrixInput
        [1176]) );
    VMW_FD \matrixInput_reg[778]  ( .D(n26478), .CP(Clk), .Q(matrixInput[778])
         );
    VMW_FD \matrixInput_reg[761]  ( .D(n26495), .CP(Clk), .Q(matrixInput[761])
         );
    VMW_FD \matrixInput_reg[462]  ( .D(n26794), .CP(Clk), .Q(matrixInput[462])
         );
    VMW_AO22 U1672 ( .A(matrixInput[1743]), .B(n25096), .C(matrixInput[1735]), 
        .D(n25081), .Z(n25521) );
    VMW_AO22 U2074 ( .A(matrixInput[1381]), .B(n25096), .C(matrixInput[1373]), 
        .D(n25081), .Z(n25883) );
    VMW_FD \matrixInput_reg[1752]  ( .D(n25504), .CP(Clk), .Q(matrixInput
        [1752]) );
    VMW_FD \matrixInput_reg[145]  ( .D(n27111), .CP(Clk), .Q(matrixInput[145])
         );
    VMW_AO22 U1044 ( .A(matrixInput[465]), .B(n25096), .C(matrixInput[457]), 
        .D(n25081), .Z(n26799) );
    VMW_AO22 U1655 ( .A(matrixInput[1758]), .B(n25096), .C(matrixInput[1750]), 
        .D(n25081), .Z(n25506) );
    VMW_FD \matrixInput_reg[1448]  ( .D(n25808), .CP(Clk), .Q(matrixInput
        [1448]) );
    VMW_FD \matrixInput_reg[246]  ( .D(n27010), .CP(Clk), .Q(matrixInput[246])
         );
    VMW_AO22 U1248 ( .A(matrixInput[281]), .B(n25096), .C(matrixInput[273]), 
        .D(n25081), .Z(n26983) );
    VMW_AO22 U1374 ( .A(matrixInput[2010]), .B(n25096), .C(matrixInput[2002]), 
        .D(n25081), .Z(n25254) );
    VMW_AO22 U1565 ( .A(matrixInput[1839]), .B(n25096), .C(matrixInput[1831]), 
        .D(n25081), .Z(n25425) );
    VMW_AO22 U2344 ( .A(matrixInput[120]), .B(n25096), .C(matrixInput[112]), 
        .D(n25081), .Z(n27144) );
    VMW_FD \matrixInput_reg[1761]  ( .D(n25495), .CP(Clk), .Q(matrixInput
        [1761]) );
    VMW_FD \matrixInput_reg[1451]  ( .D(n25805), .CP(Clk), .Q(matrixInput
        [1451]) );
    VMW_AO22 U2555 ( .A(cOutput[56]), .B(n25089), .C(cOutput[40]), .D(n25088), 
        .Z(n25177) );
    VMW_FD \matrixInput_reg[1778]  ( .D(n25478), .CP(Clk), .Q(matrixInput
        [1778]) );
    VMW_FD \matrixInput_reg[176]  ( .D(n27080), .CP(Clk), .Q(matrixInput[176])
         );
    VMW_AO22 U1459 ( .A(matrixInput[1935]), .B(n25096), .C(matrixInput[1927]), 
        .D(n25081), .Z(n25329) );
    VMW_AO22 U1887 ( .A(matrixInput[1549]), .B(n25096), .C(matrixInput[1541]), 
        .D(n25081), .Z(n25715) );
    VMW_AO22 U1917 ( .A(matrixInput[1522]), .B(n25096), .C(matrixInput[1514]), 
        .D(n25081), .Z(n25742) );
    VMW_FD \matrixInput_reg[1462]  ( .D(n25794), .CP(Clk), .Q(matrixInput
        [1462]) );
    VMW_FD \matrixInput_reg[275]  ( .D(n26981), .CP(Clk), .Q(matrixInput[275])
         );
    VMW_FD \matrixInput_reg[1816]  ( .D(n25440), .CP(Clk), .Q(matrixInput
        [1816]) );
    VMW_AO22 U2278 ( .A(matrixInput[126]), .B(n25096), .C(matrixInput[118]), 
        .D(n25081), .Z(n27138) );
    VMW_AO22 U2469 ( .A(matrixInput[1025]), .B(n25096), .C(matrixInput[1017]), 
        .D(n25081), .Z(n26239) );
    VMW_AO22 U864 ( .A(matrixInput[627]), .B(n25096), .C(matrixInput[619]), 
        .D(n25081), .Z(n26637) );
    VMW_AO22 U1178 ( .A(matrixInput[344]), .B(n25096), .C(matrixInput[336]), 
        .D(n25081), .Z(n26920) );
    VMW_AO22 U1769 ( .A(matrixInput[1656]), .B(n25096), .C(matrixInput[1648]), 
        .D(n25081), .Z(n25608) );
    VMW_FD \matrixInput_reg[986]  ( .D(n26270), .CP(Clk), .Q(matrixInput[986])
         );
    VMW_FD \matrixInput_reg[1825]  ( .D(n25431), .CP(Clk), .Q(matrixInput
        [1825]) );
    VMW_AO22 U2148 ( .A(matrixInput[1314]), .B(n25096), .C(matrixInput[1306]), 
        .D(n25081), .Z(n25950) );
    VMW_AO22 U416 ( .A(DataIn[1]), .B(n25095), .C(vectorInput[121]), .D(n25080
        ), .Z(n27263) );
    VMW_AO22 U431 ( .A(vectorInput[116]), .B(n25095), .C(vectorInput[108]), 
        .D(n25080), .Z(n27276) );
    VMW_AO22 U843 ( .A(matrixInput[646]), .B(n25096), .C(matrixInput[638]), 
        .D(n25081), .Z(n26618) );
    VMW_FD \matrixInput_reg[1986]  ( .D(n25270), .CP(Clk), .Q(matrixInput
        [1986]) );
    VMW_FD \matrixInput_reg[816]  ( .D(n26440), .CP(Clk), .Q(matrixInput[816])
         );
    VMW_FD \matrixInput_reg[56]  ( .D(n27200), .CP(Clk), .Q(matrixInput[56])
         );
    VMW_AO22 U478 ( .A(matrixInput[975]), .B(n25096), .C(matrixInput[967]), 
        .D(n25081), .Z(n26289) );
    VMW_AO22 U691 ( .A(matrixInput[783]), .B(n25096), .C(matrixInput[775]), 
        .D(n25081), .Z(n26481) );
    VMW_AO22 U701 ( .A(matrixInput[774]), .B(n25096), .C(matrixInput[766]), 
        .D(n25081), .Z(n26490) );
    VMW_FD \matrixInput_reg[825]  ( .D(n26431), .CP(Clk), .Q(matrixInput[825])
         );
    VMW_AO22 U748 ( .A(matrixInput[731]), .B(n25096), .C(matrixInput[723]), 
        .D(n25081), .Z(n26533) );
    VMW_AO22 U1131 ( .A(matrixInput[387]), .B(n25096), .C(matrixInput[379]), 
        .D(n25081), .Z(n26877) );
    VMW_AO22 U1720 ( .A(matrixInput[1700]), .B(n25096), .C(matrixInput[1692]), 
        .D(n25081), .Z(n25564) );
    VMW_FD \matrixInput_reg[1623]  ( .D(n25633), .CP(Clk), .Q(matrixInput
        [1623]) );
    VMW_FD \matrixInput_reg[65]  ( .D(n27191), .CP(Clk), .Q(matrixInput[65])
         );
    VMW_AO22 U1201 ( .A(matrixInput[323]), .B(n25096), .C(matrixInput[315]), 
        .D(n25081), .Z(n26941) );
    VMW_AO22 U1391 ( .A(matrixInput[1997]), .B(n25096), .C(matrixInput[1989]), 
        .D(n25081), .Z(n25267) );
    VMW_AO22 U1410 ( .A(matrixInput[1979]), .B(n25096), .C(matrixInput[1971]), 
        .D(n25081), .Z(n25285) );
    VMW_AO22 U2091 ( .A(matrixInput[1366]), .B(n25096), .C(matrixInput[1358]), 
        .D(n25081), .Z(n25898) );
    VMW_AO22 U2101 ( .A(matrixInput[1357]), .B(n25096), .C(matrixInput[1349]), 
        .D(n25081), .Z(n25907) );
    VMW_FD \matrixInput_reg[2044]  ( .D(n25212), .CP(Clk), .Q(matrixInput
        [2044]) );
    VMW_FD \matrixInput_reg[1539]  ( .D(n25717), .CP(Clk), .Q(matrixInput
        [1539]) );
    VMW_FD \matrixInput_reg[1520]  ( .D(n25736), .CP(Clk), .Q(matrixInput
        [1520]) );
    VMW_FD \matrixInput_reg[337]  ( .D(n26919), .CP(Clk), .Q(matrixInput[337])
         );
    VMW_FD \matrixInput_reg[1294]  ( .D(n25962), .CP(Clk), .Q(matrixInput
        [1294]) );
    VMW_AO22 U1580 ( .A(matrixInput[1826]), .B(n25096), .C(matrixInput[1818]), 
        .D(n25081), .Z(n25438) );
    VMW_AO22 U1226 ( .A(matrixInput[301]), .B(n25096), .C(matrixInput[293]), 
        .D(n25081), .Z(n26963) );
    VMW_AO22 U1862 ( .A(matrixInput[1572]), .B(n25096), .C(matrixInput[1564]), 
        .D(n25081), .Z(n25692) );
    VMW_FD \matrixInput_reg[483]  ( .D(n26773), .CP(Clk), .Q(matrixInput[483])
         );
    VMW_AO22 U2231 ( .A(matrixInput[1239]), .B(n25096), .C(matrixInput[1231]), 
        .D(n25081), .Z(n26025) );
    VMW_FD \matrixInput_reg[1610]  ( .D(n25646), .CP(Clk), .Q(matrixInput
        [1610]) );
    VMW_FD \matrixInput_reg[1609]  ( .D(n25647), .CP(Clk), .Q(matrixInput
        [1609]) );
    VMW_FD \matrixInput_reg[1513]  ( .D(n25743), .CP(Clk), .Q(matrixInput
        [1513]) );
    VMW_FD \matrixInput_reg[304]  ( .D(n26952), .CP(Clk), .Q(matrixInput[304])
         );
    VMW_AO22 U2420 ( .A(matrixInput[1069]), .B(n25096), .C(matrixInput[1061]), 
        .D(n25081), .Z(n26195) );
    VMW_FD \matrixInput_reg[1197]  ( .D(n26059), .CP(Clk), .Q(matrixInput
        [1197]) );
    VMW_FD \matrixInput_reg[1034]  ( .D(n26222), .CP(Clk), .Q(matrixInput
        [1034]) );
    VMW_FD \matrixInput_reg[799]  ( .D(n26457), .CP(Clk), .Q(matrixInput[799])
         );
    VMW_FD \matrixInput_reg[780]  ( .D(n26476), .CP(Clk), .Q(matrixInput[780])
         );
    VMW_AO22 U1437 ( .A(matrixInput[1955]), .B(n25096), .C(matrixInput[1947]), 
        .D(n25081), .Z(n25309) );
    VMW_AO22 U1845 ( .A(matrixInput[165]), .B(n25096), .C(matrixInput[157]), 
        .D(n25081), .Z(n27099) );
    VMW_FD \matrixInput_reg[623]  ( .D(n26633), .CP(Clk), .Q(matrixInput[623])
         );
    VMW_AO22 U2407 ( .A(matrixInput[1081]), .B(n25096), .C(matrixInput[1073]), 
        .D(n25081), .Z(n26183) );
    VMW_FD \matrixInput_reg[1337]  ( .D(n25919), .CP(Clk), .Q(matrixInput
        [1337]) );
    VMW_FD \holder_reg[2]  ( .D(n27390), .CP(Clk), .Q(\holder[2] ) );
    VMW_AO22 U1086 ( .A(matrixInput[427]), .B(n25096), .C(matrixInput[419]), 
        .D(n25081), .Z(n26837) );
    VMW_AO22 U1116 ( .A(matrixInput[400]), .B(n25096), .C(matrixInput[392]), 
        .D(n25081), .Z(n26864) );
    VMW_AO22 U2216 ( .A(matrixInput[1253]), .B(n25096), .C(matrixInput[1245]), 
        .D(n25081), .Z(n26011) );
    VMW_AO22 U2386 ( .A(matrixInput[1100]), .B(n25096), .C(matrixInput[1092]), 
        .D(n25081), .Z(n26164) );
    VMW_INV U2597 ( .A(Addr[1]), .Z(n25083) );
    VMW_FD \matrixInput_reg[520]  ( .D(n26736), .CP(Clk), .Q(matrixInput[520])
         );
    VMW_FD \matrixInput_reg[1483]  ( .D(n25773), .CP(Clk), .Q(matrixInput
        [1483]) );
    VMW_FD \matrixInput_reg[539]  ( .D(n26717), .CP(Clk), .Q(matrixInput[539])
         );
    VMW_FD \matrixInput_reg[609]  ( .D(n26647), .CP(Clk), .Q(matrixInput[609])
         );
    VMW_FD \matrixInput_reg[294]  ( .D(n26962), .CP(Clk), .Q(matrixInput[294])
         );
    VMW_AO22 U1697 ( .A(matrixInput[1720]), .B(n25096), .C(matrixInput[1712]), 
        .D(n25081), .Z(n25544) );
    VMW_FD \matrixInput_reg[610]  ( .D(n26646), .CP(Clk), .Q(matrixInput[610])
         );
    VMW_AO22 U1707 ( .A(matrixInput[1711]), .B(n25096), .C(matrixInput[1703]), 
        .D(n25081), .Z(n25553) );
    VMW_FD \matrixInput_reg[1007]  ( .D(n26249), .CP(Clk), .Q(matrixInput
        [1007]) );
    VMW_FD \matrixInput_reg[513]  ( .D(n26743), .CP(Clk), .Q(matrixInput[513])
         );
    VMW_AO22 U2126 ( .A(matrixInput[1334]), .B(n25096), .C(matrixInput[1326]), 
        .D(n25081), .Z(n25930) );
    VMW_PULLDOWN U272 ( .Z(n25190) );
    VMW_AO22 U355 ( .A(vectorInput[69]), .B(n25095), .C(vectorInput[61]), .D(
        n25080), .Z(n27323) );
    VMW_AO22 U544 ( .A(matrixInput[915]), .B(n25096), .C(matrixInput[907]), 
        .D(n25081), .Z(n26349) );
    VMW_AO22 U936 ( .A(matrixInput[562]), .B(n25096), .C(matrixInput[554]), 
        .D(n25081), .Z(n26702) );
    VMW_FD \matrixInput_reg[1799]  ( .D(n25457), .CP(Clk), .Q(matrixInput
        [1799]) );
    VMW_FD \matrixInput_reg[1304]  ( .D(n25952), .CP(Clk), .Q(matrixInput
        [1304]) );
    VMW_FD \matrixInput_reg[1780]  ( .D(n25476), .CP(Clk), .Q(matrixInput
        [1780]) );
    VMW_FD \matrixInput_reg[967]  ( .D(n26289), .CP(Clk), .Q(matrixInput[967])
         );
    VMW_FD \matrixInput_reg[197]  ( .D(n27059), .CP(Clk), .Q(matrixInput[197])
         );
    VMW_AO22 U369 ( .A(vectorInput[57]), .B(n25095), .C(vectorInput[49]), .D(
        n25080), .Z(n27335) );
    VMW_AO22 U372 ( .A(vectorInput[54]), .B(n25095), .C(vectorInput[46]), .D(
        n25080), .Z(n27338) );
    VMW_AO22 U653 ( .A(matrixInput[817]), .B(n25096), .C(matrixInput[809]), 
        .D(n25081), .Z(n26447) );
    VMW_AO22 U674 ( .A(matrixInput[798]), .B(n25096), .C(matrixInput[790]), 
        .D(n25081), .Z(n26466) );
    VMW_AO22 U1979 ( .A(matrixInput[1467]), .B(n25096), .C(matrixInput[1459]), 
        .D(n25081), .Z(n25797) );
    VMW_FD \matrixInput_reg[954]  ( .D(n26302), .CP(Clk), .Q(matrixInput[954])
         );
    VMW_FD \matrixInput_reg[1967]  ( .D(n25289), .CP(Clk), .Q(matrixInput
        [1967]) );
    VMW_FD \vectorInput_reg[34]  ( .D(n27350), .CP(Clk), .Q(vectorInput[34])
         );
    VMW_AO22 U881 ( .A(matrixInput[611]), .B(n25096), .C(matrixInput[603]), 
        .D(n25081), .Z(n26653) );
    VMW_AO22 U911 ( .A(matrixInput[585]), .B(n25096), .C(matrixInput[577]), 
        .D(n25081), .Z(n26679) );
    VMW_AO22 U563 ( .A(matrixInput[898]), .B(n25096), .C(matrixInput[890]), 
        .D(n25081), .Z(n26366) );
    VMW_AO22 U1016 ( .A(matrixInput[490]), .B(n25096), .C(matrixInput[482]), 
        .D(n25081), .Z(n26774) );
    VMW_AO22 U1186 ( .A(matrixInput[337]), .B(n25096), .C(matrixInput[329]), 
        .D(n25081), .Z(n26927) );
    VMW_FD \matrixInput_reg[1954]  ( .D(n25302), .CP(Clk), .Q(matrixInput
        [1954]) );
    VMW_FD \matrixInput_reg[1493]  ( .D(n25763), .CP(Clk), .Q(matrixInput
        [1493]) );
    VMW_FD \matrixInput_reg[284]  ( .D(n26972), .CP(Clk), .Q(matrixInput[284])
         );
    VMW_FD \matrixInput_reg[84]  ( .D(n27172), .CP(Clk), .Q(matrixInput[84])
         );
    VMW_FD \matrixInput_reg[1017]  ( .D(n26239), .CP(Clk), .Q(matrixInput
        [1017]) );
    VMW_FD \matrixInput_reg[600]  ( .D(n26656), .CP(Clk), .Q(matrixInput[600])
         );
    VMW_AO22 U1607 ( .A(matrixInput[1802]), .B(n25096), .C(matrixInput[1794]), 
        .D(n25081), .Z(n25462) );
    VMW_FD \matrixInput_reg[619]  ( .D(n26637), .CP(Clk), .Q(matrixInput[619])
         );
    VMW_AO22 U1797 ( .A(matrixInput[1630]), .B(n25096), .C(matrixInput[1622]), 
        .D(n25081), .Z(n25634) );
    VMW_AO22 U2026 ( .A(matrixInput[1424]), .B(n25096), .C(matrixInput[1416]), 
        .D(n25081), .Z(n25840) );
    VMW_FD \matrixInput_reg[1314]  ( .D(n25942), .CP(Clk), .Q(matrixInput
        [1314]) );
    VMW_AO22 U463 ( .A(matrixInput[988]), .B(n25096), .C(matrixInput[980]), 
        .D(n25081), .Z(n26276) );
    VMW_AO22 U578 ( .A(matrixInput[885]), .B(n25096), .C(matrixInput[877]), 
        .D(n25081), .Z(n26379) );
    VMW_BUFIZ U2637 ( .A(n25207), .E(RD), .Z(\DataOut[11]1 ) );
    VMW_FD \matrixInput_reg[503]  ( .D(n26753), .CP(Clk), .Q(matrixInput[503])
         );
    VMW_AO22 U648 ( .A(matrixInput[821]), .B(n25096), .C(matrixInput[813]), 
        .D(n25081), .Z(n26443) );
    VMW_AO22 U1326 ( .A(DataIn[6]), .B(n25096), .C(matrixInput[2046]), .D(
        n25081), .Z(n25210) );
    VMW_AO22 U1537 ( .A(matrixInput[1865]), .B(n25096), .C(matrixInput[1857]), 
        .D(n25081), .Z(n25399) );
    VMW_FD \matrixInput_reg[1790]  ( .D(n25466), .CP(Clk), .Q(matrixInput
        [1790]) );
    VMW_FD \matrixInput_reg[187]  ( .D(n27069), .CP(Clk), .Q(matrixInput[187])
         );
    VMW_FD \matrixInput_reg[1789]  ( .D(n25467), .CP(Clk), .Q(matrixInput
        [1789]) );
    VMW_FD \matrixInput_reg[633]  ( .D(n26623), .CP(Clk), .Q(matrixInput[633])
         );
    VMW_AO22 U1945 ( .A(matrixInput[156]), .B(n25096), .C(matrixInput[148]), 
        .D(n25081), .Z(n27108) );
    VMW_FD \matrixInput_reg[1024]  ( .D(n26232), .CP(Clk), .Q(matrixInput
        [1024]) );
    VMW_AO22 U2316 ( .A(matrixInput[1163]), .B(n25096), .C(matrixInput[1155]), 
        .D(n25081), .Z(n26101) );
    VMW_AND3 U2497 ( .A(n25105), .B(n25106), .C(n25107), .Z(n25079) );
    VMW_AO22 U2507 ( .A(cOutput[21]), .B(n25087), .C(cOutput[5]), .D(n25084), 
        .Z(n25119) );
    VMW_FD \matrixInput_reg[529]  ( .D(n26727), .CP(Clk), .Q(matrixInput[529])
         );
    VMW_AO22 U811 ( .A(matrixInput[675]), .B(n25096), .C(matrixInput[667]), 
        .D(n25081), .Z(n26589) );
    VMW_AO22 U1031 ( .A(matrixInput[477]), .B(n25096), .C(matrixInput[469]), 
        .D(n25081), .Z(n26787) );
    VMW_AO22 U1291 ( .A(matrixInput[242]), .B(n25096), .C(matrixInput[234]), 
        .D(n25081), .Z(n27022) );
    VMW_AO22 U1301 ( .A(matrixInput[233]), .B(n25096), .C(matrixInput[225]), 
        .D(n25081), .Z(n27031) );
    VMW_AO22 U1480 ( .A(matrixInput[1916]), .B(n25096), .C(matrixInput[1908]), 
        .D(n25081), .Z(n25348) );
    VMW_AO22 U2286 ( .A(matrixInput[1190]), .B(n25096), .C(matrixInput[1182]), 
        .D(n25081), .Z(n26074) );
    VMW_FD \matrixInput_reg[1327]  ( .D(n25929), .CP(Clk), .Q(matrixInput
        [1327]) );
    VMW_FD \matrixInput_reg[530]  ( .D(n26726), .CP(Clk), .Q(matrixInput[530])
         );
    VMW_FD \matrixInput_reg[493]  ( .D(n26763), .CP(Clk), .Q(matrixInput[493])
         );
    VMW_AO22 U1510 ( .A(matrixInput[1889]), .B(n25096), .C(matrixInput[1881]), 
        .D(n25081), .Z(n25375) );
    VMW_FD \matrixInput_reg[1284]  ( .D(n25972), .CP(Clk), .Q(matrixInput
        [1284]) );
    VMW_AO22 U1962 ( .A(matrixInput[1482]), .B(n25096), .C(matrixInput[1474]), 
        .D(n25081), .Z(n25782) );
    VMW_FD \matrixInput_reg[1619]  ( .D(n25637), .CP(Clk), .Q(matrixInput
        [1619]) );
    VMW_FD \matrixInput_reg[1600]  ( .D(n25656), .CP(Clk), .Q(matrixInput
        [1600]) );
    VMW_AO22 U2331 ( .A(matrixInput[1149]), .B(n25096), .C(matrixInput[1141]), 
        .D(n25081), .Z(n26115) );
    VMW_AO22 U2520 ( .A(cOutput[84]), .B(n25087), .C(cOutput[68]), .D(n25084), 
        .Z(n25134) );
    VMW_FD \matrixInput_reg[1503]  ( .D(n25753), .CP(Clk), .Q(matrixInput
        [1503]) );
    VMW_FD \matrixInput_reg[790]  ( .D(n26466), .CP(Clk), .Q(matrixInput[790])
         );
    VMW_FD \matrixInput_reg[314]  ( .D(n26942), .CP(Clk), .Q(matrixInput[314])
         );
    VMW_FD \matrixInput_reg[789]  ( .D(n26467), .CP(Clk), .Q(matrixInput[789])
         );
    VMW_FD \matrixInput_reg[1187]  ( .D(n26069), .CP(Clk), .Q(matrixInput
        [1187]) );
    VMW_FD \matrixInput_reg[1633]  ( .D(n25623), .CP(Clk), .Q(matrixInput
        [1633]) );
    VMW_AO22 U1620 ( .A(matrixInput[1790]), .B(n25096), .C(matrixInput[1782]), 
        .D(n25081), .Z(n25474) );
    VMW_AO22 U2001 ( .A(matrixInput[1447]), .B(n25096), .C(matrixInput[1439]), 
        .D(n25081), .Z(n25817) );
    VMW_AO22 U2191 ( .A(matrixInput[1276]), .B(n25096), .C(matrixInput[1268]), 
        .D(n25081), .Z(n25988) );
    VMW_BUFIZ U2610 ( .A(n25187), .E(RD), .Z(\DataOut[19]1 ) );
    VMW_FD \matrixInput_reg[1530]  ( .D(n25726), .CP(Clk), .Q(matrixInput
        [1530]) );
    VMW_FD \matrixInput_reg[1529]  ( .D(n25727), .CP(Clk), .Q(matrixInput
        [1529]) );
    VMW_FD \matrixInput_reg[327]  ( .D(n26929), .CP(Clk), .Q(matrixInput[327])
         );
    VMW_AO22 U981 ( .A(matrixInput[521]), .B(n25096), .C(matrixInput[513]), 
        .D(n25081), .Z(n26743) );
    VMW_FD \matrixInput_reg[1944]  ( .D(n25312), .CP(Clk), .Q(matrixInput
        [1944]) );
    VMW_FD \matrixInput_reg[94]  ( .D(n27162), .CP(Clk), .Q(matrixInput[94])
         );
    VMW_PULLDOWN U285 ( .Z(n25203) );
    VMW_OAI211 U297 ( .A(n25055), .B(n25065), .C(n25066), .D(n25067), .Z(
        n27389) );
    VMW_AO22 U320 ( .A(vectorInput[101]), .B(n25095), .C(vectorInput[93]), .D(
        n25080), .Z(n27291) );
    VMW_AO22 U444 ( .A(matrixInput[1006]), .B(n25096), .C(matrixInput[998]), 
        .D(n25081), .Z(n26258) );
    VMW_AO22 U753 ( .A(matrixInput[727]), .B(n25096), .C(matrixInput[719]), 
        .D(n25081), .Z(n26537) );
    VMW_AO22 U774 ( .A(matrixInput[14]), .B(n25096), .C(matrixInput[6]), .D(
        n25081), .Z(n27250) );
    VMW_FD \matrixInput_reg[1977]  ( .D(n25279), .CP(Clk), .Q(matrixInput
        [1977]) );
    VMW_AO22 U836 ( .A(matrixInput[652]), .B(n25096), .C(matrixInput[644]), 
        .D(n25081), .Z(n26612) );
    VMW_AO22 U1879 ( .A(matrixInput[1557]), .B(n25096), .C(matrixInput[1549]), 
        .D(n25081), .Z(n25707) );
    VMW_FD \matrixInput_reg[944]  ( .D(n26312), .CP(Clk), .Q(matrixInput[944])
         );
    VMW_FD \vectorInput_reg[24]  ( .D(n27360), .CP(Clk), .Q(vectorInput[24])
         );
    VMW_FD \matrixInput_reg[977]  ( .D(n26279), .CP(Clk), .Q(matrixInput[977])
         );
    VMW_AO22 U601 ( .A(matrixInput[864]), .B(n25096), .C(matrixInput[856]), 
        .D(n25081), .Z(n26400) );
    VMW_AO22 U791 ( .A(matrixInput[693]), .B(n25096), .C(matrixInput[685]), 
        .D(n25081), .Z(n26571) );
    VMW_AO22 U858 ( .A(matrixInput[632]), .B(n25096), .C(matrixInput[624]), 
        .D(n25081), .Z(n26632) );
    VMW_AO22 U1274 ( .A(matrixInput[32]), .B(n25096), .C(matrixInput[24]), .D(
        n25081), .Z(n27232) );
    VMW_AO22 U2244 ( .A(matrixInput[129]), .B(n25096), .C(matrixInput[121]), 
        .D(n25081), .Z(n27135) );
    VMW_AO22 U2455 ( .A(matrixInput[110]), .B(n25096), .C(matrixInput[102]), 
        .D(n25081), .Z(n27154) );
    VMW_FD \matrixInput_reg[166]  ( .D(n27090), .CP(Clk), .Q(matrixInput[166])
         );
    VMW_FD \vectorInput_reg[17]  ( .D(n27367), .CP(Clk), .Q(vectorInput[17])
         );
    VMW_FD \matrixInput_reg[1771]  ( .D(n25485), .CP(Clk), .Q(matrixInput
        [1771]) );
    VMW_FD \matrixInput_reg[1768]  ( .D(n25488), .CP(Clk), .Q(matrixInput
        [1768]) );
    VMW_FD \matrixInput_reg[265]  ( .D(n26991), .CP(Clk), .Q(matrixInput[265])
         );
    VMW_AO22 U1465 ( .A(matrixInput[1929]), .B(n25096), .C(matrixInput[1921]), 
        .D(n25081), .Z(n25335) );
    VMW_FD \matrixInput_reg[1472]  ( .D(n25784), .CP(Clk), .Q(matrixInput
        [1472]) );
    VMW_AO22 U1817 ( .A(matrixInput[1612]), .B(n25096), .C(matrixInput[1604]), 
        .D(n25081), .Z(n25652) );
    VMW_AO22 U1987 ( .A(matrixInput[1459]), .B(n25096), .C(matrixInput[1451]), 
        .D(n25081), .Z(n25805) );
    VMW_AO22 U2174 ( .A(matrixInput[1291]), .B(n25096), .C(matrixInput[1283]), 
        .D(n25081), .Z(n25973) );
    VMW_FD \matrixInput_reg[1742]  ( .D(n25514), .CP(Clk), .Q(matrixInput
        [1742]) );
    VMW_FD \matrixInput_reg[155]  ( .D(n27101), .CP(Clk), .Q(matrixInput[155])
         );
    VMW_AO22 U1144 ( .A(matrixInput[375]), .B(n25096), .C(matrixInput[367]), 
        .D(n25081), .Z(n26889) );
    VMW_AO22 U1163 ( .A(matrixInput[42]), .B(n25096), .C(matrixInput[34]), .D(
        n25081), .Z(n27222) );
    VMW_AO22 U1755 ( .A(matrixInput[1668]), .B(n25096), .C(matrixInput[1660]), 
        .D(n25081), .Z(n25596) );
    VMW_FD \matrixInput_reg[1458]  ( .D(n25798), .CP(Clk), .Q(matrixInput
        [1458]) );
    VMW_FD \matrixInput_reg[1441]  ( .D(n25815), .CP(Clk), .Q(matrixInput
        [1441]) );
    VMW_AO22 U1772 ( .A(matrixInput[1653]), .B(n25096), .C(matrixInput[1645]), 
        .D(n25081), .Z(n25611) );
    VMW_AO22 U2153 ( .A(matrixInput[1309]), .B(n25096), .C(matrixInput[1301]), 
        .D(n25081), .Z(n25955) );
    VMW_FD \matrixInput_reg[256]  ( .D(n27000), .CP(Clk), .Q(matrixInput[256])
         );
    VMW_FD \matrixInput_reg[1265]  ( .D(n25991), .CP(Clk), .Q(matrixInput
        [1265]) );
    VMW_FD \matrixInput_reg[1166]  ( .D(n26090), .CP(Clk), .Q(matrixInput
        [1166]) );
    VMW_FD \matrixInput_reg[771]  ( .D(n26485), .CP(Clk), .Q(matrixInput[771])
         );
    VMW_FD \matrixInput_reg[768]  ( .D(n26488), .CP(Clk), .Q(matrixInput[768])
         );
    VMW_FD \matrixInput_reg[472]  ( .D(n26784), .CP(Clk), .Q(matrixInput[472])
         );
    VMW_AO22 U1253 ( .A(matrixInput[277]), .B(n25096), .C(matrixInput[269]), 
        .D(n25081), .Z(n26987) );
    VMW_AO22 U1442 ( .A(matrixInput[1950]), .B(n25096), .C(matrixInput[1942]), 
        .D(n25081), .Z(n25314) );
    VMW_AO22 U2263 ( .A(matrixInput[1210]), .B(n25096), .C(matrixInput[1202]), 
        .D(n25081), .Z(n26054) );
    VMW_FD \matrixInput_reg[1155]  ( .D(n26101), .CP(Clk), .Q(matrixInput
        [1155]) );
    VMW_FD \matrixInput_reg[742]  ( .D(n26514), .CP(Clk), .Q(matrixInput[742])
         );
    VMW_AO22 U2472 ( .A(matrixInput[1022]), .B(n25096), .C(matrixInput[1014]), 
        .D(n25081), .Z(n26242) );
    VMW_AO22 U1830 ( .A(matrixInput[1601]), .B(n25096), .C(matrixInput[1593]), 
        .D(n25081), .Z(n25663) );
    VMW_FD \matrixInput_reg[1256]  ( .D(n26000), .CP(Clk), .Q(matrixInput
        [1256]) );
    VMW_FD \matrixInput_reg[835]  ( .D(n26421), .CP(Clk), .Q(matrixInput[835])
         );
    VMW_FD \matrixInput_reg[458]  ( .D(n26798), .CP(Clk), .Q(matrixInput[458])
         );
    VMW_FD \matrixInput_reg[441]  ( .D(n26815), .CP(Clk), .Q(matrixInput[441])
         );
    VMW_AO22 U943 ( .A(matrixInput[556]), .B(n25096), .C(matrixInput[548]), 
        .D(n25081), .Z(n26708) );
    VMW_FD \matrixInput_reg[806]  ( .D(n26450), .CP(Clk), .Q(matrixInput[806])
         );
    VMW_FD \matrixInput_reg[75]  ( .D(n27181), .CP(Clk), .Q(matrixInput[75])
         );
    VMW_FD \matrixInput_reg[1996]  ( .D(n25260), .CP(Clk), .Q(matrixInput
        [1996]) );
    VMW_FD \matrixInput_reg[46]  ( .D(n27210), .CP(Clk), .Q(matrixInput[46])
         );
    VMW_AO22 U531 ( .A(matrixInput[927]), .B(n25096), .C(matrixInput[919]), 
        .D(n25081), .Z(n26337) );
    VMW_AO22 U964 ( .A(matrixInput[537]), .B(n25096), .C(matrixInput[529]), 
        .D(n25081), .Z(n26727) );
    VMW_AO22 U1078 ( .A(matrixInput[434]), .B(n25096), .C(matrixInput[426]), 
        .D(n25081), .Z(n26830) );
    VMW_AO22 U1669 ( .A(matrixInput[1746]), .B(n25096), .C(matrixInput[1738]), 
        .D(n25081), .Z(n25518) );
    VMW_FD \matrixInput_reg[1835]  ( .D(n25421), .CP(Clk), .Q(matrixInput
        [1835]) );
    VMW_AND2 U307 ( .A(n25082), .B(Addr[0]), .Z(n25088) );
    VMW_AO22 U516 ( .A(matrixInput[940]), .B(n25096), .C(matrixInput[932]), 
        .D(n25081), .Z(n26324) );
    VMW_AO22 U2048 ( .A(matrixInput[1405]), .B(n25096), .C(matrixInput[1397]), 
        .D(n25081), .Z(n25859) );
    VMW_AO22 U315 ( .A(vectorInput[106]), .B(n25095), .C(vectorInput[98]), .D(
        n25080), .Z(n27286) );
    VMW_AO22 U332 ( .A(vectorInput[90]), .B(n25095), .C(vectorInput[82]), .D(
        n25080), .Z(n27302) );
    VMW_AO22 U486 ( .A(matrixInput[103]), .B(n25096), .C(matrixInput[95]), .D(
        n25081), .Z(n27161) );
    VMW_AO22 U523 ( .A(matrixInput[934]), .B(n25096), .C(matrixInput[926]), 
        .D(n25081), .Z(n26330) );
    VMW_AO22 U613 ( .A(matrixInput[853]), .B(n25096), .C(matrixInput[845]), 
        .D(n25081), .Z(n26411) );
    VMW_AO22 U626 ( .A(matrixInput[841]), .B(n25096), .C(matrixInput[833]), 
        .D(n25081), .Z(n26423) );
    VMW_AO22 U1348 ( .A(matrixInput[2034]), .B(n25096), .C(matrixInput[2026]), 
        .D(n25081), .Z(n25230) );
    VMW_FD \matrixInput_reg[1806]  ( .D(n25450), .CP(Clk), .Q(matrixInput
        [1806]) );
    VMW_AO22 U1559 ( .A(matrixInput[1845]), .B(n25096), .C(matrixInput[1837]), 
        .D(n25081), .Z(n25419) );
    VMW_OAI21 U2569 ( .A(n25112), .B(n25113), .C(n25093), .Z(n25118) );
    VMW_AO22 U2378 ( .A(matrixInput[117]), .B(n25096), .C(matrixInput[109]), 
        .D(n25081), .Z(n27147) );
    VMW_FD \matrixInput_reg[996]  ( .D(n26260), .CP(Clk), .Q(matrixInput[996])
         );
    VMW_AO22 U783 ( .A(matrixInput[700]), .B(n25096), .C(matrixInput[692]), 
        .D(n25081), .Z(n26564) );
    VMW_FD \matrixInput_reg[1963]  ( .D(n25293), .CP(Clk), .Q(matrixInput
        [1963]) );
    VMW_FD \matrixInput_reg[1950]  ( .D(n25306), .CP(Clk), .Q(matrixInput
        [1950]) );
    VMW_FD \matrixInput_reg[1949]  ( .D(n25307), .CP(Clk), .Q(matrixInput
        [1949]) );
    VMW_FD \matrixInput_reg[80]  ( .D(n27176), .CP(Clk), .Q(matrixInput[80])
         );
    VMW_FD \matrixInput_reg[99]  ( .D(n27157), .CP(Clk), .Q(matrixInput[99])
         );
    VMW_AO22 U951 ( .A(matrixInput[548]), .B(n25096), .C(matrixInput[540]), 
        .D(n25081), .Z(n26716) );
    VMW_AO22 U494 ( .A(matrixInput[960]), .B(n25096), .C(matrixInput[952]), 
        .D(n25081), .Z(n26304) );
    VMW_OAI211 U299 ( .A(n25055), .B(n25071), .C(n25072), .D(n25073), .Z(
        n27387) );
    VMW_AO22 U329 ( .A(vectorInput[93]), .B(n25095), .C(vectorInput[85]), .D(
        n25080), .Z(n27299) );
    VMW_AO22 U347 ( .A(vectorInput[77]), .B(n25095), .C(vectorInput[69]), .D(
        n25080), .Z(n27315) );
    VMW_AO22 U438 ( .A(vectorInput[109]), .B(n25095), .C(vectorInput[101]), 
        .D(n25080), .Z(n27283) );
    VMW_AO22 U504 ( .A(matrixInput[951]), .B(n25096), .C(matrixInput[943]), 
        .D(n25081), .Z(n26313) );
    VMW_AO22 U634 ( .A(matrixInput[834]), .B(n25096), .C(matrixInput[826]), 
        .D(n25081), .Z(n26430) );
    VMW_AO22 U976 ( .A(matrixInput[526]), .B(n25096), .C(matrixInput[518]), 
        .D(n25081), .Z(n26738) );
    VMW_FD \matrixInput_reg[963]  ( .D(n26293), .CP(Clk), .Q(matrixInput[963])
         );
    VMW_AO22 U1939 ( .A(matrixInput[1503]), .B(n25096), .C(matrixInput[1495]), 
        .D(n25081), .Z(n25761) );
    VMW_FD \vectorInput_reg[30]  ( .D(n27354), .CP(Clk), .Q(vectorInput[30])
         );
    VMW_FD \vectorInput_reg[29]  ( .D(n27355), .CP(Clk), .Q(vectorInput[29])
         );
    VMW_FD \matrixInput_reg[950]  ( .D(n26306), .CP(Clk), .Q(matrixInput[950])
         );
    VMW_FD \matrixInput_reg[949]  ( .D(n26307), .CP(Clk), .Q(matrixInput[949])
         );
    VMW_AO22 U698 ( .A(matrixInput[777]), .B(n25096), .C(matrixInput[769]), 
        .D(n25081), .Z(n26487) );
    VMW_AO22 U708 ( .A(matrixInput[83]), .B(n25096), .C(matrixInput[75]), .D(
        n25081), .Z(n27181) );
    VMW_AO22 U2256 ( .A(matrixInput[1217]), .B(n25096), .C(matrixInput[1209]), 
        .D(n25081), .Z(n26047) );
    VMW_AO22 U2447 ( .A(matrixInput[1045]), .B(n25096), .C(matrixInput[1037]), 
        .D(n25081), .Z(n26219) );
    VMW_AO22 U1266 ( .A(matrixInput[265]), .B(n25096), .C(matrixInput[257]), 
        .D(n25081), .Z(n26999) );
    VMW_AO22 U1477 ( .A(matrixInput[1918]), .B(n25096), .C(matrixInput[1910]), 
        .D(n25081), .Z(n25346) );
    VMW_AO22 U1805 ( .A(matrixInput[1623]), .B(n25096), .C(matrixInput[1615]), 
        .D(n25081), .Z(n25641) );
    VMW_FD \matrixInput_reg[1333]  ( .D(n25923), .CP(Clk), .Q(matrixInput
        [1333]) );
    VMW_FD \matrixInput_reg[524]  ( .D(n26732), .CP(Clk), .Q(matrixInput[524])
         );
    VMW_FD \holder_reg[6]  ( .D(n27386), .CP(Clk), .Q(\holder[6] ) );
    VMW_AO22 U1995 ( .A(matrixInput[1452]), .B(n25096), .C(matrixInput[1444]), 
        .D(n25081), .Z(n25812) );
    VMW_FD \matrixInput_reg[627]  ( .D(n26629), .CP(Clk), .Q(matrixInput[627])
         );
    VMW_AO22 U2166 ( .A(matrixInput[1298]), .B(n25096), .C(matrixInput[1290]), 
        .D(n25081), .Z(n25966) );
    VMW_FD \matrixInput_reg[1784]  ( .D(n25472), .CP(Clk), .Q(matrixInput
        [1784]) );
    VMW_FD \matrixInput_reg[1030]  ( .D(n26226), .CP(Clk), .Q(matrixInput
        [1030]) );
    VMW_FD \matrixInput_reg[1029]  ( .D(n26227), .CP(Clk), .Q(matrixInput
        [1029]) );
    VMW_FD \matrixInput_reg[193]  ( .D(n27063), .CP(Clk), .Q(matrixInput[193])
         );
    VMW_FD \matrixInput_reg[1319]  ( .D(n25937), .CP(Clk), .Q(matrixInput
        [1319]) );
    VMW_FD \matrixInput_reg[1300]  ( .D(n25956), .CP(Clk), .Q(matrixInput
        [1300]) );
    VMW_FD \matrixInput_reg[517]  ( .D(n26739), .CP(Clk), .Q(matrixInput[517])
         );
    VMW_AO22 U456 ( .A(matrixInput[995]), .B(n25096), .C(matrixInput[987]), 
        .D(n25081), .Z(n26269) );
    VMW_AO22 U471 ( .A(matrixInput[981]), .B(n25096), .C(matrixInput[973]), 
        .D(n25081), .Z(n26283) );
    VMW_AO22 U1156 ( .A(matrixInput[364]), .B(n25096), .C(matrixInput[356]), 
        .D(n25081), .Z(n26900) );
    VMW_AO22 U1747 ( .A(matrixInput[1676]), .B(n25096), .C(matrixInput[1668]), 
        .D(n25081), .Z(n25588) );
    VMW_FD \matrixInput_reg[1003]  ( .D(n26253), .CP(Clk), .Q(matrixInput
        [1003]) );
    VMW_FD \matrixInput_reg[614]  ( .D(n26642), .CP(Clk), .Q(matrixInput[614])
         );
    VMW_AO22 U1171 ( .A(matrixInput[350]), .B(n25096), .C(matrixInput[342]), 
        .D(n25081), .Z(n26914) );
    VMW_AO22 U2141 ( .A(matrixInput[1320]), .B(n25096), .C(matrixInput[1312]), 
        .D(n25081), .Z(n25944) );
    VMW_FD \matrixInput_reg[1524]  ( .D(n25732), .CP(Clk), .Q(matrixInput
        [1524]) );
    VMW_FD \matrixInput_reg[1487]  ( .D(n25769), .CP(Clk), .Q(matrixInput
        [1487]) );
    VMW_FD \matrixInput_reg[290]  ( .D(n26966), .CP(Clk), .Q(matrixInput[290])
         );
    VMW_FD \matrixInput_reg[289]  ( .D(n26967), .CP(Clk), .Q(matrixInput[289])
         );
    VMW_FD \matrixInput_reg[333]  ( .D(n26923), .CP(Clk), .Q(matrixInput[333])
         );
    VMW_FD \matrixInput_reg[2040]  ( .D(n25216), .CP(Clk), .Q(matrixInput
        [2040]) );
    VMW_AO22 U1241 ( .A(matrixInput[35]), .B(n25096), .C(matrixInput[27]), .D(
        n25081), .Z(n27229) );
    VMW_AO22 U1760 ( .A(matrixInput[1664]), .B(n25096), .C(matrixInput[1656]), 
        .D(n25081), .Z(n25600) );
    VMW_AO22 U1822 ( .A(matrixInput[23]), .B(n25096), .C(matrixInput[15]), .D(
        n25081), .Z(n27241) );
    VMW_AO22 U2271 ( .A(matrixInput[1204]), .B(n25096), .C(matrixInput[1196]), 
        .D(n25081), .Z(n26060) );
    VMW_AO22 U2460 ( .A(matrixInput[1033]), .B(n25096), .C(matrixInput[1025]), 
        .D(n25081), .Z(n26231) );
    VMW_FD \matrixInput_reg[1627]  ( .D(n25629), .CP(Clk), .Q(matrixInput
        [1627]) );
    VMW_FD \matrixInput_reg[784]  ( .D(n26472), .CP(Clk), .Q(matrixInput[784])
         );
    VMW_FD \matrixInput_reg[1193]  ( .D(n26063), .CP(Clk), .Q(matrixInput
        [1193]) );
    VMW_FD \matrixInput_reg[1614]  ( .D(n25642), .CP(Clk), .Q(matrixInput
        [1614]) );
    VMW_FD \matrixInput_reg[1517]  ( .D(n25739), .CP(Clk), .Q(matrixInput
        [1517]) );
    VMW_FD \matrixInput_reg[319]  ( .D(n26937), .CP(Clk), .Q(matrixInput[319])
         );
    VMW_FD \matrixInput_reg[300]  ( .D(n26956), .CP(Clk), .Q(matrixInput[300])
         );
    VMW_FD \matrixInput_reg[1289]  ( .D(n25967), .CP(Clk), .Q(matrixInput
        [1289]) );
    VMW_FD \matrixInput_reg[487]  ( .D(n26769), .CP(Clk), .Q(matrixInput[487])
         );
    VMW_AO22 U1450 ( .A(matrixInput[1943]), .B(n25096), .C(matrixInput[1935]), 
        .D(n25081), .Z(n25321) );
    VMW_FD \matrixInput_reg[1290]  ( .D(n25966), .CP(Clk), .Q(matrixInput
        [1290]) );
    VMW_AO22 U741 ( .A(matrixInput[80]), .B(n25096), .C(matrixInput[72]), .D(
        n25081), .Z(n27184) );
    VMW_AO22 U803 ( .A(matrixInput[682]), .B(n25096), .C(matrixInput[674]), 
        .D(n25081), .Z(n26582) );
    VMW_AO22 U993 ( .A(matrixInput[510]), .B(n25096), .C(matrixInput[502]), 
        .D(n25081), .Z(n26754) );
    VMW_FD \matrixInput_reg[1982]  ( .D(n25274), .CP(Clk), .Q(matrixInput
        [1982]) );
    VMW_FD \matrixInput_reg[812]  ( .D(n26444), .CP(Clk), .Q(matrixInput[812])
         );
    VMW_FD \matrixInput_reg[52]  ( .D(n27204), .CP(Clk), .Q(matrixInput[52])
         );
    VMW_FD \matrixInput_reg[78]  ( .D(n27178), .CP(Clk), .Q(matrixInput[78])
         );
    VMW_FD \matrixInput_reg[61]  ( .D(n27195), .CP(Clk), .Q(matrixInput[61])
         );
    VMW_AO22 U766 ( .A(matrixInput[715]), .B(n25096), .C(matrixInput[707]), 
        .D(n25081), .Z(n26549) );
    VMW_AO22 U2429 ( .A(matrixInput[1061]), .B(n25096), .C(matrixInput[1053]), 
        .D(n25081), .Z(n26203) );
    VMW_FD \matrixInput_reg[838]  ( .D(n26418), .CP(Clk), .Q(matrixInput[838])
         );
    VMW_FD \matrixInput_reg[821]  ( .D(n26435), .CP(Clk), .Q(matrixInput[821])
         );
    VMW_AO22 U1208 ( .A(matrixInput[317]), .B(n25096), .C(matrixInput[309]), 
        .D(n25081), .Z(n26947) );
    VMW_AO22 U1589 ( .A(matrixInput[188]), .B(n25096), .C(matrixInput[180]), 
        .D(n25081), .Z(n27076) );
    VMW_AO22 U2238 ( .A(matrixInput[1233]), .B(n25096), .C(matrixInput[1225]), 
        .D(n25081), .Z(n26031) );
    VMW_FD \matrixInput_reg[982]  ( .D(n26274), .CP(Clk), .Q(matrixInput[982])
         );
    VMW_AO22 U1398 ( .A(matrixInput[1990]), .B(n25096), .C(matrixInput[1982]), 
        .D(n25081), .Z(n25274) );
    VMW_AO22 U1419 ( .A(matrixInput[1971]), .B(n25096), .C(matrixInput[1963]), 
        .D(n25081), .Z(n25293) );
    VMW_AO22 U2098 ( .A(matrixInput[1359]), .B(n25096), .C(matrixInput[1351]), 
        .D(n25081), .Z(n25905) );
    VMW_FD \matrixInput_reg[1812]  ( .D(n25444), .CP(Clk), .Q(matrixInput
        [1812]) );
    VMW_AO22 U824 ( .A(matrixInput[663]), .B(n25096), .C(matrixInput[655]), 
        .D(n25081), .Z(n26601) );
    VMW_AO22 U2108 ( .A(matrixInput[1350]), .B(n25096), .C(matrixInput[1342]), 
        .D(n25081), .Z(n25914) );
    VMW_AO22 U888 ( .A(matrixInput[606]), .B(n25096), .C(matrixInput[598]), 
        .D(n25081), .Z(n26658) );
    VMW_AO22 U918 ( .A(matrixInput[578]), .B(n25096), .C(matrixInput[570]), 
        .D(n25081), .Z(n26686) );
    VMW_AO22 U1004 ( .A(matrixInput[501]), .B(n25096), .C(matrixInput[493]), 
        .D(n25081), .Z(n26763) );
    VMW_AO22 U1138 ( .A(matrixInput[380]), .B(n25096), .C(matrixInput[372]), 
        .D(n25081), .Z(n26884) );
    VMW_FD \matrixInput_reg[1838]  ( .D(n25418), .CP(Clk), .Q(matrixInput
        [1838]) );
    VMW_FD \matrixInput_reg[1821]  ( .D(n25435), .CP(Clk), .Q(matrixInput
        [1821]) );
    VMW_AO22 U1729 ( .A(matrixInput[1692]), .B(n25096), .C(matrixInput[1684]), 
        .D(n25081), .Z(n25572) );
    VMW_AO22 U1194 ( .A(matrixInput[329]), .B(n25096), .C(matrixInput[321]), 
        .D(n25081), .Z(n26935) );
    VMW_AO22 U1785 ( .A(matrixInput[1641]), .B(n25096), .C(matrixInput[1633]), 
        .D(n25081), .Z(n25623) );
    VMW_FD \matrixInput_reg[1455]  ( .D(n25801), .CP(Clk), .Q(matrixInput
        [1455]) );
    VMW_AO22 U1615 ( .A(matrixInput[1795]), .B(n25096), .C(matrixInput[1787]), 
        .D(n25081), .Z(n25469) );
    VMW_FD \matrixInput_reg[242]  ( .D(n27014), .CP(Clk), .Q(matrixInput[242])
         );
    VMW_AO22 U1023 ( .A(matrixInput[484]), .B(n25096), .C(matrixInput[476]), 
        .D(n25081), .Z(n26780) );
    VMW_AO22 U1283 ( .A(matrixInput[249]), .B(n25096), .C(matrixInput[241]), 
        .D(n25081), .Z(n27015) );
    VMW_AO22 U1334 ( .A(matrixInput[2047]), .B(n25096), .C(matrixInput[2039]), 
        .D(n25081), .Z(n25217) );
    VMW_AO22 U1957 ( .A(matrixInput[1487]), .B(n25096), .C(matrixInput[1479]), 
        .D(n25081), .Z(n25777) );
    VMW_AO22 U2034 ( .A(matrixInput[1417]), .B(n25096), .C(matrixInput[1409]), 
        .D(n25081), .Z(n25847) );
    VMW_BUFIZ U2625 ( .A(n25198), .E(RD), .Z(\DataOut[30]1 ) );
    VMW_FD \matrixInput_reg[1756]  ( .D(n25500), .CP(Clk), .Q(matrixInput
        [1756]) );
    VMW_FD \matrixInput_reg[158]  ( .D(n27098), .CP(Clk), .Q(matrixInput[158])
         );
    VMW_FD \matrixInput_reg[141]  ( .D(n27115), .CP(Clk), .Q(matrixInput[141])
         );
    VMW_FD \matrixInput_reg[271]  ( .D(n26985), .CP(Clk), .Q(matrixInput[271])
         );
    VMW_FD \matrixInput_reg[268]  ( .D(n26988), .CP(Clk), .Q(matrixInput[268])
         );
    VMW_AO22 U1502 ( .A(matrixInput[1897]), .B(n25096), .C(matrixInput[1889]), 
        .D(n25081), .Z(n25367) );
    VMW_AO22 U1525 ( .A(matrixInput[1876]), .B(n25096), .C(matrixInput[1868]), 
        .D(n25081), .Z(n25388) );
    VMW_FD \matrixInput_reg[1466]  ( .D(n25790), .CP(Clk), .Q(matrixInput
        [1466]) );
    VMW_AO22 U1970 ( .A(matrixInput[1475]), .B(n25096), .C(matrixInput[1467]), 
        .D(n25081), .Z(n25789) );
    VMW_AO22 U2294 ( .A(matrixInput[1183]), .B(n25096), .C(matrixInput[1175]), 
        .D(n25081), .Z(n26081) );
    VMW_AND3 U2515 ( .A(n25127), .B(n25128), .C(n25129), .Z(n25073) );
    VMW_FD \matrixInput_reg[172]  ( .D(n27084), .CP(Clk), .Q(matrixInput[172])
         );
    VMW_AO22 U2304 ( .A(matrixInput[1174]), .B(n25096), .C(matrixInput[1166]), 
        .D(n25081), .Z(n26090) );
    VMW_AO22 U2485 ( .A(matrixInput[1010]), .B(n25096), .C(matrixInput[1002]), 
        .D(n25081), .Z(n26254) );
    VMW_FD \matrixInput_reg[1765]  ( .D(n25491), .CP(Clk), .Q(matrixInput
        [1765]) );
    VMW_FD \matrixInput_reg[1242]  ( .D(n26014), .CP(Clk), .Q(matrixInput
        [1242]) );
    VMW_FD \matrixInput_reg[455]  ( .D(n26801), .CP(Clk), .Q(matrixInput[455])
         );
    VMW_AO22 U1313 ( .A(matrixInput[222]), .B(n25096), .C(matrixInput[214]), 
        .D(n25081), .Z(n27042) );
    VMW_AO22 U1492 ( .A(matrixInput[1906]), .B(n25096), .C(matrixInput[1898]), 
        .D(n25081), .Z(n25358) );
    VMW_AO22 U1632 ( .A(matrixInput[1779]), .B(n25096), .C(matrixInput[1771]), 
        .D(n25081), .Z(n25485) );
    VMW_AO22 U2323 ( .A(matrixInput[1157]), .B(n25096), .C(matrixInput[1149]), 
        .D(n25081), .Z(n26107) );
    VMW_AO22 U2532 ( .A(cOutput[123]), .B(n25089), .C(cOutput[107]), .D(n25088
        ), .Z(n25148) );
    VMW_FD \matrixInput_reg[1158]  ( .D(n26098), .CP(Clk), .Q(matrixInput
        [1158]) );
    VMW_FD \matrixInput_reg[1141]  ( .D(n26115), .CP(Clk), .Q(matrixInput
        [1141]) );
    VMW_FD \matrixInput_reg[756]  ( .D(n26500), .CP(Clk), .Q(matrixInput[756])
         );
    VMW_AO22 U2008 ( .A(matrixInput[1440]), .B(n25096), .C(matrixInput[1432]), 
        .D(n25081), .Z(n25824) );
    VMW_AO22 U2013 ( .A(matrixInput[1436]), .B(n25096), .C(matrixInput[1428]), 
        .D(n25081), .Z(n25828) );
    VMW_FD \matrixInput_reg[1271]  ( .D(n25985), .CP(Clk), .Q(matrixInput
        [1271]) );
    VMW_FD \matrixInput_reg[466]  ( .D(n26790), .CP(Clk), .Q(matrixInput[466])
         );
    VMW_FD \matrixInput_reg[1268]  ( .D(n25988), .CP(Clk), .Q(matrixInput
        [1268]) );
    VMW_FD \matrixInput_reg[1172]  ( .D(n26084), .CP(Clk), .Q(matrixInput
        [1172]) );
    VMW_FD \matrixInput_reg[765]  ( .D(n26491), .CP(Clk), .Q(matrixInput[765])
         );
    VMW_AO22 U2183 ( .A(matrixInput[1283]), .B(n25096), .C(matrixInput[1275]), 
        .D(n25081), .Z(n25981) );
    VMW_INV U2602 ( .A(\holder[7] ), .Z(n25077) );
    VMW_AO22 U360 ( .A(vectorInput[65]), .B(n25095), .C(vectorInput[57]), .D(
        n25080), .Z(n27327) );
    VMW_AO22 U556 ( .A(matrixInput[905]), .B(n25096), .C(matrixInput[897]), 
        .D(n25081), .Z(n26359) );
    VMW_AO22 U2198 ( .A(matrixInput[1269]), .B(n25096), .C(matrixInput[1261]), 
        .D(n25081), .Z(n25995) );
    VMW_BUFIZ U2619 ( .A(n25194), .E(RD), .Z(\DataOut[21]1 ) );
    VMW_AO22 U571 ( .A(matrixInput[891]), .B(n25096), .C(matrixInput[883]), 
        .D(n25081), .Z(n26373) );
    VMW_AO22 U641 ( .A(matrixInput[89]), .B(n25096), .C(matrixInput[81]), .D(
        n25081), .Z(n27175) );
    VMW_AO22 U666 ( .A(matrixInput[806]), .B(n25096), .C(matrixInput[798]), 
        .D(n25081), .Z(n26458) );
    VMW_AO22 U924 ( .A(matrixInput[573]), .B(n25096), .C(matrixInput[565]), 
        .D(n25081), .Z(n26691) );
    VMW_AO22 U1038 ( .A(matrixInput[470]), .B(n25096), .C(matrixInput[462]), 
        .D(n25081), .Z(n26794) );
    VMW_AO22 U1629 ( .A(matrixInput[1782]), .B(n25096), .C(matrixInput[1774]), 
        .D(n25081), .Z(n25482) );
    VMW_FD \matrixInput_reg[1831]  ( .D(n25425), .CP(Clk), .Q(matrixInput
        [1831]) );
    VMW_FD \matrixInput_reg[1828]  ( .D(n25428), .CP(Clk), .Q(matrixInput
        [1828]) );
    VMW_AO22 U2338 ( .A(matrixInput[1143]), .B(n25096), .C(matrixInput[1135]), 
        .D(n25081), .Z(n26121) );
    VMW_AO22 U2529 ( .A(cOutput[83]), .B(n25087), .C(cOutput[67]), .D(n25084), 
        .Z(n25145) );
    VMW_AO22 U1298 ( .A(matrixInput[236]), .B(n25096), .C(matrixInput[228]), 
        .D(n25081), .Z(n27028) );
    VMW_AO22 U1519 ( .A(matrixInput[1881]), .B(n25096), .C(matrixInput[1873]), 
        .D(n25081), .Z(n25383) );
    VMW_FD \matrixInput_reg[992]  ( .D(n26264), .CP(Clk), .Q(matrixInput[992])
         );
    VMW_AO22 U1308 ( .A(matrixInput[227]), .B(n25096), .C(matrixInput[219]), 
        .D(n25081), .Z(n27037) );
    VMW_AO22 U1489 ( .A(matrixInput[26]), .B(n25096), .C(matrixInput[18]), .D(
        n25081), .Z(n27238) );
    VMW_FD \matrixInput_reg[1802]  ( .D(n25454), .CP(Clk), .Q(matrixInput
        [1802]) );
    VMW_FD \matrixInput_reg[71]  ( .D(n27185), .CP(Clk), .Q(matrixInput[71])
         );
    VMW_FD \matrixInput_reg[68]  ( .D(n27188), .CP(Clk), .Q(matrixInput[68])
         );
    VMW_FD \matrixInput_reg[831]  ( .D(n26425), .CP(Clk), .Q(matrixInput[831])
         );
    VMW_FD \matrixInput_reg[828]  ( .D(n26428), .CP(Clk), .Q(matrixInput[828])
         );
    VMW_AO22 U385 ( .A(vectorInput[42]), .B(n25095), .C(vectorInput[34]), .D(
        n25080), .Z(n27350) );
    VMW_AO22 U734 ( .A(matrixInput[744]), .B(n25096), .C(matrixInput[736]), 
        .D(n25081), .Z(n26520) );
    VMW_AO22 U818 ( .A(matrixInput[668]), .B(n25096), .C(matrixInput[660]), 
        .D(n25081), .Z(n26596) );
    VMW_AO22 U893 ( .A(matrixInput[601]), .B(n25096), .C(matrixInput[593]), 
        .D(n25081), .Z(n26663) );
    VMW_AO22 U903 ( .A(matrixInput[592]), .B(n25096), .C(matrixInput[584]), 
        .D(n25081), .Z(n26672) );
    VMW_FD \matrixInput_reg[1992]  ( .D(n25264), .CP(Clk), .Q(matrixInput
        [1992]) );
    VMW_FD \matrixInput_reg[42]  ( .D(n27214), .CP(Clk), .Q(matrixInput[42])
         );
    VMW_AO22 U988 ( .A(matrixInput[515]), .B(n25096), .C(matrixInput[507]), 
        .D(n25081), .Z(n26749) );
    VMW_AO22 U1094 ( .A(matrixInput[419]), .B(n25096), .C(matrixInput[411]), 
        .D(n25081), .Z(n26845) );
    VMW_AO22 U1123 ( .A(matrixInput[394]), .B(n25096), .C(matrixInput[386]), 
        .D(n25081), .Z(n26870) );
    VMW_FD \matrixInput_reg[802]  ( .D(n26454), .CP(Clk), .Q(matrixInput[802])
         );
    VMW_AO22 U1213 ( .A(matrixInput[312]), .B(n25096), .C(matrixInput[304]), 
        .D(n25081), .Z(n26952) );
    VMW_AO22 U1592 ( .A(matrixInput[1815]), .B(n25096), .C(matrixInput[1807]), 
        .D(n25081), .Z(n25449) );
    VMW_AO22 U1732 ( .A(matrixInput[1689]), .B(n25096), .C(matrixInput[1681]), 
        .D(n25081), .Z(n25575) );
    VMW_AO22 U1870 ( .A(matrixInput[1565]), .B(n25096), .C(matrixInput[1557]), 
        .D(n25081), .Z(n25699) );
    VMW_AO22 U2083 ( .A(matrixInput[1373]), .B(n25096), .C(matrixInput[1365]), 
        .D(n25081), .Z(n25891) );
    VMW_FD \matrixInput_reg[1278]  ( .D(n25978), .CP(Clk), .Q(matrixInput
        [1278]) );
    VMW_FD \matrixInput_reg[1261]  ( .D(n25995), .CP(Clk), .Q(matrixInput
        [1261]) );
    VMW_FD \matrixInput_reg[1162]  ( .D(n26094), .CP(Clk), .Q(matrixInput
        [1162]) );
    VMW_FD \matrixInput_reg[476]  ( .D(n26780), .CP(Clk), .Q(matrixInput[476])
         );
    VMW_FD \matrixInput_reg[775]  ( .D(n26481), .CP(Clk), .Q(matrixInput[775])
         );
    VMW_AO22 U2113 ( .A(matrixInput[1346]), .B(n25096), .C(matrixInput[1338]), 
        .D(n25081), .Z(n25918) );
    VMW_FD \matrixInput_reg[1252]  ( .D(n26004), .CP(Clk), .Q(matrixInput
        [1252]) );
    VMW_FD \matrixInput_reg[445]  ( .D(n26811), .CP(Clk), .Q(matrixInput[445])
         );
    VMW_AO22 U1234 ( .A(matrixInput[294]), .B(n25096), .C(matrixInput[286]), 
        .D(n25081), .Z(n26970) );
    VMW_AO22 U1383 ( .A(matrixInput[2004]), .B(n25096), .C(matrixInput[1996]), 
        .D(n25081), .Z(n25260) );
    VMW_AO22 U1402 ( .A(matrixInput[1987]), .B(n25096), .C(matrixInput[1979]), 
        .D(n25081), .Z(n25277) );
    VMW_AO22 U1425 ( .A(matrixInput[1966]), .B(n25096), .C(matrixInput[1958]), 
        .D(n25081), .Z(n25298) );
    VMW_AO22 U1857 ( .A(matrixInput[1577]), .B(n25096), .C(matrixInput[1569]), 
        .D(n25081), .Z(n25687) );
    VMW_AO22 U2223 ( .A(matrixInput[1247]), .B(n25096), .C(matrixInput[1239]), 
        .D(n25081), .Z(n26017) );
    VMW_AO22 U2432 ( .A(matrixInput[1058]), .B(n25096), .C(matrixInput[1050]), 
        .D(n25081), .Z(n26206) );
    VMW_FD \matrixInput_reg[1151]  ( .D(n26105), .CP(Clk), .Q(matrixInput
        [1151]) );
    VMW_FD \matrixInput_reg[746]  ( .D(n26510), .CP(Clk), .Q(matrixInput[746])
         );
    VMW_FD \matrixInput_reg[1148]  ( .D(n26108), .CP(Clk), .Q(matrixInput
        [1148]) );
    VMW_AO22 U2204 ( .A(matrixInput[1264]), .B(n25096), .C(matrixInput[1256]), 
        .D(n25081), .Z(n26000) );
    VMW_OAI21 U2585 ( .A(n25156), .B(n25157), .C(n25093), .Z(n25162) );
    VMW_FD \matrixInput_reg[1476]  ( .D(n25780), .CP(Clk), .Q(matrixInput
        [1476]) );
    VMW_FD \matrixInput_reg[278]  ( .D(n26978), .CP(Clk), .Q(matrixInput[278])
         );
    VMW_FD \matrixInput_reg[261]  ( .D(n26995), .CP(Clk), .Q(matrixInput[261])
         );
    VMW_FD \matrixInput_reg[1775]  ( .D(n25481), .CP(Clk), .Q(matrixInput
        [1775]) );
    VMW_AO22 U2394 ( .A(matrixInput[1093]), .B(n25096), .C(matrixInput[1085]), 
        .D(n25081), .Z(n26171) );
    VMW_AO22 U2415 ( .A(matrixInput[1074]), .B(n25096), .C(matrixInput[1066]), 
        .D(n25081), .Z(n26190) );
    VMW_FD \matrixInput_reg[252]  ( .D(n27004), .CP(Clk), .Q(matrixInput[252])
         );
    VMW_FD \matrixInput_reg[162]  ( .D(n27094), .CP(Clk), .Q(matrixInput[162])
         );
    VMW_AO22 U1104 ( .A(matrixInput[410]), .B(n25096), .C(matrixInput[402]), 
        .D(n25081), .Z(n26854) );
    VMW_AO22 U1715 ( .A(matrixInput[1705]), .B(n25096), .C(matrixInput[1697]), 
        .D(n25081), .Z(n25559) );
    VMW_AO22 U1685 ( .A(matrixInput[1731]), .B(n25096), .C(matrixInput[1723]), 
        .D(n25081), .Z(n25533) );
    VMW_FD \matrixInput_reg[1445]  ( .D(n25811), .CP(Clk), .Q(matrixInput
        [1445]) );
    VMW_AO22 U1839 ( .A(matrixInput[1593]), .B(n25096), .C(matrixInput[1585]), 
        .D(n25081), .Z(n25671) );
    VMW_AO22 U2134 ( .A(matrixInput[1327]), .B(n25096), .C(matrixInput[1319]), 
        .D(n25081), .Z(n25937) );
    VMW_FD \matrixInput_reg[1746]  ( .D(n25510), .CP(Clk), .Q(matrixInput
        [1746]) );
    VMW_FD \matrixInput_reg[151]  ( .D(n27105), .CP(Clk), .Q(matrixInput[151])
         );
    VMW_FD \matrixInput_reg[148]  ( .D(n27108), .CP(Clk), .Q(matrixInput[148])
         );
    VMW_FD \matrixInput_reg[959]  ( .D(n26297), .CP(Clk), .Q(matrixInput[959])
         );
    VMW_FD \matrixInput_reg[940]  ( .D(n26316), .CP(Clk), .Q(matrixInput[940])
         );
    VMW_FD \vectorInput_reg[39]  ( .D(n27345), .CP(Clk), .Q(vectorInput[39])
         );
    VMW_FD \vectorInput_reg[20]  ( .D(n27364), .CP(Clk), .Q(vectorInput[20])
         );
    VMW_FD \vectorInput_reg[13]  ( .D(n27371), .CP(Clk), .Q(vectorInput[13])
         );
    VMW_AO22 U404 ( .A(vectorInput[25]), .B(n25095), .C(vectorInput[17]), .D(
        n25080), .Z(n27367) );
    VMW_AO22 U423 ( .A(vectorInput[123]), .B(n25095), .C(vectorInput[115]), 
        .D(n25080), .Z(n27269) );
    VMW_AO22 U594 ( .A(matrixInput[870]), .B(n25096), .C(matrixInput[862]), 
        .D(n25081), .Z(n26394) );
    VMW_AO22 U876 ( .A(matrixInput[616]), .B(n25096), .C(matrixInput[608]), 
        .D(n25081), .Z(n26648) );
    VMW_FD \matrixInput_reg[973]  ( .D(n26283), .CP(Clk), .Q(matrixInput[973])
         );
    VMW_AO22 U538 ( .A(matrixInput[920]), .B(n25096), .C(matrixInput[912]), 
        .D(n25081), .Z(n26344) );
    VMW_AO22 U683 ( .A(matrixInput[790]), .B(n25096), .C(matrixInput[782]), 
        .D(n25081), .Z(n26474) );
    VMW_AO22 U851 ( .A(matrixInput[638]), .B(n25096), .C(matrixInput[630]), 
        .D(n25081), .Z(n26626) );
    VMW_FD \matrixInput_reg[1959]  ( .D(n25297), .CP(Clk), .Q(matrixInput
        [1959]) );
    VMW_FD \matrixInput_reg[1940]  ( .D(n25316), .CP(Clk), .Q(matrixInput
        [1940]) );
    VMW_FD \matrixInput_reg[89]  ( .D(n27167), .CP(Clk), .Q(matrixInput[89])
         );
    VMW_FD \matrixInput_reg[90]  ( .D(n27166), .CP(Clk), .Q(matrixInput[90])
         );
    VMW_FD \matrixInput_reg[1973]  ( .D(n25283), .CP(Clk), .Q(matrixInput
        [1973]) );
    VMW_AO22 U713 ( .A(matrixInput[763]), .B(n25096), .C(matrixInput[755]), 
        .D(n25081), .Z(n26501) );
    VMW_AO22 U1071 ( .A(matrixInput[440]), .B(n25096), .C(matrixInput[432]), 
        .D(n25081), .Z(n26824) );
    VMW_AO22 U1341 ( .A(matrixInput[2040]), .B(n25096), .C(matrixInput[2032]), 
        .D(n25081), .Z(n25224) );
    VMW_AO22 U1550 ( .A(matrixInput[1853]), .B(n25096), .C(matrixInput[1845]), 
        .D(n25081), .Z(n25411) );
    VMW_AO22 U1922 ( .A(matrixInput[158]), .B(n25096), .C(matrixInput[150]), 
        .D(n25081), .Z(n27106) );
    VMW_AO22 U2371 ( .A(matrixInput[1113]), .B(n25096), .C(matrixInput[1105]), 
        .D(n25081), .Z(n26151) );
    VMW_AND3 U2560 ( .A(n25182), .B(n25183), .C(n25184), .Z(n25058) );
    VMW_FD \matrixInput_reg[1183]  ( .D(n26073), .CP(Clk), .Q(matrixInput
        [1183]) );
    VMW_FD \matrixInput_reg[1507]  ( .D(n25749), .CP(Clk), .Q(matrixInput
        [1507]) );
    VMW_FD \matrixInput_reg[794]  ( .D(n26462), .CP(Clk), .Q(matrixInput[794])
         );
    VMW_FD \matrixInput_reg[310]  ( .D(n26946), .CP(Clk), .Q(matrixInput[310])
         );
    VMW_FD \matrixInput_reg[309]  ( .D(n26947), .CP(Clk), .Q(matrixInput[309])
         );
    VMW_FD \matrixInput_reg[1604]  ( .D(n25652), .CP(Clk), .Q(matrixInput
        [1604]) );
    VMW_FD \matrixInput_reg[1299]  ( .D(n25957), .CP(Clk), .Q(matrixInput
        [1299]) );
    VMW_FD \matrixInput_reg[1280]  ( .D(n25976), .CP(Clk), .Q(matrixInput
        [1280]) );
    VMW_AO22 U1660 ( .A(matrixInput[1754]), .B(n25096), .C(matrixInput[1746]), 
        .D(n25081), .Z(n25510) );
    VMW_AO22 U2041 ( .A(matrixInput[1410]), .B(n25096), .C(matrixInput[1402]), 
        .D(n25081), .Z(n25854) );
    VMW_FD \matrixInput_reg[1534]  ( .D(n25722), .CP(Clk), .Q(matrixInput
        [1534]) );
    VMW_FD \matrixInput_reg[497]  ( .D(n26759), .CP(Clk), .Q(matrixInput[497])
         );
    VMW_FD \matrixInput_reg[323]  ( .D(n26933), .CP(Clk), .Q(matrixInput[323])
         );
    VMW_FD \matrixInput_reg[1794]  ( .D(n25462), .CP(Clk), .Q(matrixInput
        [1794]) );
    VMW_FD \matrixInput_reg[1637]  ( .D(n25619), .CP(Clk), .Q(matrixInput
        [1637]) );
    VMW_FD \matrixInput_reg[507]  ( .D(n26749), .CP(Clk), .Q(matrixInput[507])
         );
    VMW_FD \matrixInput_reg[183]  ( .D(n27073), .CP(Clk), .Q(matrixInput[183])
         );
    VMW_AO22 U2066 ( .A(matrixInput[1388]), .B(n25096), .C(matrixInput[1380]), 
        .D(n25081), .Z(n25876) );
    VMW_AO22 U382 ( .A(vectorInput[45]), .B(n25095), .C(vectorInput[37]), .D(
        n25080), .Z(n27347) );
    VMW_AO22 U403 ( .A(vectorInput[26]), .B(n25095), .C(vectorInput[18]), .D(
        n25080), .Z(n27366) );
    VMW_AO22 U424 ( .A(vectorInput[122]), .B(n25095), .C(vectorInput[114]), 
        .D(n25080), .Z(n27270) );
    VMW_AO22 U608 ( .A(matrixInput[92]), .B(n25096), .C(matrixInput[84]), .D(
        n25081), .Z(n27172) );
    VMW_AO22 U1056 ( .A(matrixInput[454]), .B(n25096), .C(matrixInput[446]), 
        .D(n25081), .Z(n26810) );
    VMW_FD \matrixInput_reg[1310]  ( .D(n25946), .CP(Clk), .Q(matrixInput
        [1310]) );
    VMW_FD \matrixInput_reg[1309]  ( .D(n25947), .CP(Clk), .Q(matrixInput
        [1309]) );
    VMW_AO22 U1647 ( .A(matrixInput[1766]), .B(n25096), .C(matrixInput[1758]), 
        .D(n25081), .Z(n25498) );
    VMW_FD \matrixInput_reg[604]  ( .D(n26652), .CP(Clk), .Q(matrixInput[604])
         );
    VMW_AO22 U2547 ( .A(cOutput[81]), .B(n25087), .C(cOutput[65]), .D(n25084), 
        .Z(n25167) );
    VMW_FD \matrixInput_reg[1497]  ( .D(n25759), .CP(Clk), .Q(matrixInput
        [1497]) );
    VMW_FD \matrixInput_reg[1013]  ( .D(n26243), .CP(Clk), .Q(matrixInput
        [1013]) );
    VMW_FD \matrixInput_reg[1323]  ( .D(n25933), .CP(Clk), .Q(matrixInput
        [1323]) );
    VMW_FD \matrixInput_reg[299]  ( .D(n26957), .CP(Clk), .Q(matrixInput[299])
         );
    VMW_FD \matrixInput_reg[280]  ( .D(n26976), .CP(Clk), .Q(matrixInput[280])
         );
    VMW_AO22 U684 ( .A(matrixInput[789]), .B(n25096), .C(matrixInput[781]), 
        .D(n25081), .Z(n26475) );
    VMW_AO22 U714 ( .A(matrixInput[762]), .B(n25096), .C(matrixInput[754]), 
        .D(n25081), .Z(n26502) );
    VMW_AO22 U798 ( .A(matrixInput[687]), .B(n25096), .C(matrixInput[679]), 
        .D(n25081), .Z(n26577) );
    VMW_FD \matrixInput_reg[534]  ( .D(n26722), .CP(Clk), .Q(matrixInput[534])
         );
    VMW_AO22 U1366 ( .A(matrixInput[208]), .B(n25096), .C(matrixInput[200]), 
        .D(n25081), .Z(n27056) );
    VMW_AO22 U1895 ( .A(matrixInput[1542]), .B(n25096), .C(matrixInput[1534]), 
        .D(n25081), .Z(n25722) );
    VMW_AO22 U2356 ( .A(matrixInput[1127]), .B(n25096), .C(matrixInput[1119]), 
        .D(n25081), .Z(n26137) );
    VMW_AO22 U1905 ( .A(matrixInput[1533]), .B(n25096), .C(matrixInput[1525]), 
        .D(n25081), .Z(n25731) );
    VMW_FD \matrixInput_reg[1039]  ( .D(n26217), .CP(Clk), .Q(matrixInput
        [1039]) );
    VMW_FD \matrixInput_reg[1020]  ( .D(n26236), .CP(Clk), .Q(matrixInput
        [1020]) );
    VMW_AO22 U1577 ( .A(matrixInput[1828]), .B(n25096), .C(matrixInput[1820]), 
        .D(n25081), .Z(n25436) );
    VMW_FD \matrixInput_reg[637]  ( .D(n26619), .CP(Clk), .Q(matrixInput[637])
         );
    VMW_AO22 U856 ( .A(matrixInput[634]), .B(n25096), .C(matrixInput[626]), 
        .D(n25081), .Z(n26630) );
    VMW_AO22 U1819 ( .A(matrixInput[1610]), .B(n25096), .C(matrixInput[1602]), 
        .D(n25081), .Z(n25654) );
    VMW_AO22 U1989 ( .A(matrixInput[152]), .B(n25096), .C(matrixInput[144]), 
        .D(n25081), .Z(n27112) );
    VMW_FD \matrixInput_reg[942]  ( .D(n26314), .CP(Clk), .Q(matrixInput[942])
         );
    VMW_FD \vectorInput_reg[22]  ( .D(n27362), .CP(Clk), .Q(vectorInput[22])
         );
    VMW_FD \matrixInput_reg[971]  ( .D(n26285), .CP(Clk), .Q(matrixInput[971])
         );
    VMW_FD \matrixInput_reg[968]  ( .D(n26288), .CP(Clk), .Q(matrixInput[968])
         );
    VMW_AO22 U593 ( .A(matrixInput[871]), .B(n25096), .C(matrixInput[863]), 
        .D(n25081), .Z(n26393) );
    VMW_AO22 U871 ( .A(matrixInput[620]), .B(n25096), .C(matrixInput[612]), 
        .D(n25081), .Z(n26644) );
    VMW_FD \vectorInput_reg[11]  ( .D(n27373), .CP(Clk), .Q(vectorInput[11])
         );
    VMW_FD \matrixInput_reg[1942]  ( .D(n25314), .CP(Clk), .Q(matrixInput
        [1942]) );
    VMW_FD \matrixInput_reg[92]  ( .D(n27164), .CP(Clk), .Q(matrixInput[92])
         );
    VMW_AO22 U518 ( .A(matrixInput[938]), .B(n25096), .C(matrixInput[930]), 
        .D(n25081), .Z(n26326) );
    VMW_AO22 U733 ( .A(matrixInput[745]), .B(n25096), .C(matrixInput[737]), 
        .D(n25081), .Z(n26519) );
    VMW_AO22 U1051 ( .A(matrixInput[458]), .B(n25096), .C(matrixInput[450]), 
        .D(n25081), .Z(n26806) );
    VMW_AO22 U1361 ( .A(matrixInput[2022]), .B(n25096), .C(matrixInput[2014]), 
        .D(n25081), .Z(n25242) );
    VMW_AO22 U1570 ( .A(matrixInput[1835]), .B(n25096), .C(matrixInput[1827]), 
        .D(n25081), .Z(n25429) );
    VMW_FD \matrixInput_reg[1971]  ( .D(n25285), .CP(Clk), .Q(matrixInput
        [1971]) );
    VMW_FD \matrixInput_reg[1968]  ( .D(n25288), .CP(Clk), .Q(matrixInput
        [1968]) );
    VMW_FD \matrixInput_reg[1282]  ( .D(n25974), .CP(Clk), .Q(matrixInput
        [1282]) );
    VMW_FD \matrixInput_reg[495]  ( .D(n26761), .CP(Clk), .Q(matrixInput[495])
         );
    VMW_AO22 U1640 ( .A(matrixInput[1772]), .B(n25096), .C(matrixInput[1764]), 
        .D(n25081), .Z(n25492) );
    VMW_AO22 U1892 ( .A(matrixInput[1545]), .B(n25096), .C(matrixInput[1537]), 
        .D(n25081), .Z(n25719) );
    VMW_AO22 U1902 ( .A(matrixInput[1536]), .B(n25096), .C(matrixInput[1528]), 
        .D(n25081), .Z(n25728) );
    VMW_FD \matrixInput_reg[1606]  ( .D(n25650), .CP(Clk), .Q(matrixInput
        [1606]) );
    VMW_AO22 U2351 ( .A(matrixInput[1131]), .B(n25096), .C(matrixInput[1123]), 
        .D(n25081), .Z(n26133) );
    VMW_FD \matrixInput_reg[1505]  ( .D(n25751), .CP(Clk), .Q(matrixInput
        [1505]) );
    VMW_FD \matrixInput_reg[796]  ( .D(n26460), .CP(Clk), .Q(matrixInput[796])
         );
    VMW_FD \matrixInput_reg[312]  ( .D(n26944), .CP(Clk), .Q(matrixInput[312])
         );
    VMW_AO22 U2540 ( .A(cOutput[114]), .B(n25087), .C(cOutput[98]), .D(n25084), 
        .Z(n25158) );
    VMW_FD \matrixInput_reg[1198]  ( .D(n26058), .CP(Clk), .Q(matrixInput
        [1198]) );
    VMW_FD \matrixInput_reg[1635]  ( .D(n25621), .CP(Clk), .Q(matrixInput
        [1635]) );
    VMW_FD \matrixInput_reg[1181]  ( .D(n26075), .CP(Clk), .Q(matrixInput
        [1181]) );
    VMW_AO22 U1076 ( .A(matrixInput[436]), .B(n25096), .C(matrixInput[428]), 
        .D(n25081), .Z(n26828) );
    VMW_AO22 U2061 ( .A(matrixInput[1393]), .B(n25096), .C(matrixInput[1385]), 
        .D(n25081), .Z(n25871) );
    VMW_FD \matrixInput_reg[1536]  ( .D(n25720), .CP(Clk), .Q(matrixInput
        [1536]) );
    VMW_FD \matrixInput_reg[338]  ( .D(n26918), .CP(Clk), .Q(matrixInput[338])
         );
    VMW_FD \matrixInput_reg[321]  ( .D(n26935), .CP(Clk), .Q(matrixInput[321])
         );
    VMW_FD \matrixInput_reg[1495]  ( .D(n25761), .CP(Clk), .Q(matrixInput
        [1495]) );
    VMW_FD \matrixInput_reg[282]  ( .D(n26974), .CP(Clk), .Q(matrixInput[282])
         );
    VMW_FD \matrixInput_reg[1011]  ( .D(n26245), .CP(Clk), .Q(matrixInput
        [1011]) );
    VMW_FD \matrixInput_reg[1008]  ( .D(n26248), .CP(Clk), .Q(matrixInput
        [1008]) );
    VMW_AO22 U1667 ( .A(matrixInput[181]), .B(n25096), .C(matrixInput[173]), 
        .D(n25081), .Z(n27083) );
    VMW_FD \matrixInput_reg[1312]  ( .D(n25944), .CP(Clk), .Q(matrixInput
        [1312]) );
    VMW_FD \matrixInput_reg[606]  ( .D(n26650), .CP(Clk), .Q(matrixInput[606])
         );
    VMW_NOR2 U309 ( .A(Addr[3]), .B(Addr[2]), .Z(n25090) );
    VMW_AO22 U488 ( .A(matrixInput[966]), .B(n25096), .C(matrixInput[958]), 
        .D(n25081), .Z(n26298) );
    VMW_FD \matrixInput_reg[505]  ( .D(n26751), .CP(Clk), .Q(matrixInput[505])
         );
    VMW_AO22 U2046 ( .A(matrixInput[1407]), .B(n25096), .C(matrixInput[1399]), 
        .D(n25081), .Z(n25857) );
    VMW_AO22 U340 ( .A(vectorInput[83]), .B(n25095), .C(vectorInput[75]), .D(
        n25080), .Z(n27309) );
    VMW_AO22 U367 ( .A(vectorInput[58]), .B(n25095), .C(vectorInput[50]), .D(
        n25080), .Z(n27334) );
    VMW_AO22 U628 ( .A(matrixInput[839]), .B(n25096), .C(matrixInput[831]), 
        .D(n25081), .Z(n26425) );
    VMW_AO22 U1346 ( .A(matrixInput[2036]), .B(n25096), .C(matrixInput[2028]), 
        .D(n25081), .Z(n25228) );
    VMW_FD \matrixInput_reg[1796]  ( .D(n25460), .CP(Clk), .Q(matrixInput
        [1796]) );
    VMW_FD \matrixInput_reg[198]  ( .D(n27058), .CP(Clk), .Q(matrixInput[198])
         );
    VMW_FD \matrixInput_reg[181]  ( .D(n27075), .CP(Clk), .Q(matrixInput[181])
         );
    VMW_AO22 U1557 ( .A(matrixInput[1847]), .B(n25096), .C(matrixInput[1839]), 
        .D(n25081), .Z(n25417) );
    VMW_FD \matrixInput_reg[635]  ( .D(n26621), .CP(Clk), .Q(matrixInput[635])
         );
    VMW_AO22 U1925 ( .A(matrixInput[1515]), .B(n25096), .C(matrixInput[1507]), 
        .D(n25081), .Z(n25749) );
    VMW_FD \matrixInput_reg[1022]  ( .D(n26234), .CP(Clk), .Q(matrixInput
        [1022]) );
    VMW_OAI21 U2567 ( .A(n25108), .B(n25109), .C(n25090), .Z(n25117) );
    VMW_FD \matrixInput_reg[536]  ( .D(n26720), .CP(Clk), .Q(matrixInput[536])
         );
    VMW_AO22 U894 ( .A(matrixInput[600]), .B(n25096), .C(matrixInput[592]), 
        .D(n25081), .Z(n26664) );
    VMW_AO22 U1018 ( .A(matrixInput[488]), .B(n25096), .C(matrixInput[480]), 
        .D(n25081), .Z(n26776) );
    VMW_AO22 U1188 ( .A(matrixInput[335]), .B(n25096), .C(matrixInput[327]), 
        .D(n25081), .Z(n26929) );
    VMW_AO22 U1609 ( .A(matrixInput[1800]), .B(n25096), .C(matrixInput[1792]), 
        .D(n25081), .Z(n25464) );
    VMW_AO22 U2376 ( .A(matrixInput[1108]), .B(n25096), .C(matrixInput[1100]), 
        .D(n25081), .Z(n26156) );
    VMW_FD \matrixInput_reg[1338]  ( .D(n25918), .CP(Clk), .Q(matrixInput
        [1338]) );
    VMW_FD \matrixInput_reg[1321]  ( .D(n25935), .CP(Clk), .Q(matrixInput
        [1321]) );
    VMW_AO22 U1799 ( .A(matrixInput[1628]), .B(n25096), .C(matrixInput[1620]), 
        .D(n25081), .Z(n25636) );
    VMW_FD \matrixInput_reg[1833]  ( .D(n25423), .CP(Clk), .Q(matrixInput
        [1833]) );
    VMW_AO22 U904 ( .A(matrixInput[591]), .B(n25096), .C(matrixInput[583]), 
        .D(n25081), .Z(n26673) );
    VMW_AO22 U2028 ( .A(matrixInput[1422]), .B(n25096), .C(matrixInput[1414]), 
        .D(n25081), .Z(n25842) );
    VMW_AO22 U551 ( .A(matrixInput[908]), .B(n25096), .C(matrixInput[900]), 
        .D(n25081), .Z(n26356) );
    VMW_AO22 U576 ( .A(matrixInput[887]), .B(n25096), .C(matrixInput[879]), 
        .D(n25081), .Z(n26377) );
    VMW_BUFIZ U2639 ( .A(n25208), .E(RD), .Z(\DataOut[8]1 ) );
    VMW_AO22 U646 ( .A(matrixInput[823]), .B(n25096), .C(matrixInput[815]), 
        .D(n25081), .Z(n26441) );
    VMW_AO22 U1328 ( .A(DataIn[4]), .B(n25096), .C(matrixInput[2044]), .D(
        n25081), .Z(n25212) );
    VMW_AO22 U1539 ( .A(matrixInput[1863]), .B(n25096), .C(matrixInput[1855]), 
        .D(n25081), .Z(n25401) );
    VMW_FD \matrixInput_reg[1819]  ( .D(n25437), .CP(Clk), .Q(matrixInput
        [1819]) );
    VMW_FD \matrixInput_reg[1800]  ( .D(n25456), .CP(Clk), .Q(matrixInput
        [1800]) );
    VMW_AO22 U2288 ( .A(matrixInput[1188]), .B(n25096), .C(matrixInput[1180]), 
        .D(n25081), .Z(n26076) );
    VMW_AO22 U2318 ( .A(matrixInput[1161]), .B(n25096), .C(matrixInput[1153]), 
        .D(n25081), .Z(n26103) );
    VMW_AO22 U2499 ( .A(cOutput[30]), .B(n25089), .C(cOutput[14]), .D(n25088), 
        .Z(n25109) );
    VMW_FD \matrixInput_reg[989]  ( .D(n26267), .CP(Clk), .Q(matrixInput[989])
         );
    VMW_AO22 U2509 ( .A(cOutput[53]), .B(n25087), .C(cOutput[37]), .D(n25084), 
        .Z(n25121) );
    VMW_FD \matrixInput_reg[990]  ( .D(n26266), .CP(Clk), .Q(matrixInput[990])
         );
    VMW_AO22 U661 ( .A(matrixInput[809]), .B(n25096), .C(matrixInput[801]), 
        .D(n25081), .Z(n26455) );
    VMW_FD \matrixInput_reg[833]  ( .D(n26423), .CP(Clk), .Q(matrixInput[833])
         );
    VMW_AO22 U923 ( .A(matrixInput[574]), .B(n25096), .C(matrixInput[566]), 
        .D(n25081), .Z(n26690) );
    VMW_FD \matrixInput_reg[819]  ( .D(n26437), .CP(Clk), .Q(matrixInput[819])
         );
    VMW_FD \matrixInput_reg[73]  ( .D(n27183), .CP(Clk), .Q(matrixInput[73])
         );
    VMW_FD \matrixInput_reg[800]  ( .D(n26456), .CP(Clk), .Q(matrixInput[800])
         );
    VMW_FD \matrixInput_reg[1990]  ( .D(n25266), .CP(Clk), .Q(matrixInput
        [1990]) );
    VMW_FD \matrixInput_reg[1989]  ( .D(n25267), .CP(Clk), .Q(matrixInput
        [1989]) );
    VMW_FD \matrixInput_reg[40]  ( .D(n27216), .CP(Clk), .Q(matrixInput[40])
         );
    VMW_FD \matrixInput_reg[59]  ( .D(n27197), .CP(Clk), .Q(matrixInput[59])
         );
    VMW_AO22 U451 ( .A(matrixInput[999]), .B(n25096), .C(matrixInput[991]), 
        .D(n25081), .Z(n26265) );
    VMW_AO22 U823 ( .A(matrixInput[664]), .B(n25096), .C(matrixInput[656]), 
        .D(n25081), .Z(n26600) );
    VMW_AO22 U838 ( .A(matrixInput[650]), .B(n25096), .C(matrixInput[642]), 
        .D(n25081), .Z(n26614) );
    VMW_AO22 U1093 ( .A(matrixInput[420]), .B(n25096), .C(matrixInput[412]), 
        .D(n25081), .Z(n26844) );
    VMW_AO22 U1103 ( .A(matrixInput[411]), .B(n25096), .C(matrixInput[403]), 
        .D(n25081), .Z(n26853) );
    VMW_AO22 U1682 ( .A(matrixInput[1734]), .B(n25096), .C(matrixInput[1726]), 
        .D(n25081), .Z(n25530) );
    VMW_AO22 U2133 ( .A(matrixInput[139]), .B(n25096), .C(matrixInput[131]), 
        .D(n25081), .Z(n27125) );
    VMW_FD \matrixInput_reg[1263]  ( .D(n25993), .CP(Clk), .Q(matrixInput
        [1263]) );
    VMW_FD \matrixInput_reg[1179]  ( .D(n26077), .CP(Clk), .Q(matrixInput
        [1179]) );
    VMW_FD \matrixInput_reg[1160]  ( .D(n26096), .CP(Clk), .Q(matrixInput
        [1160]) );
    VMW_FD \matrixInput_reg[777]  ( .D(n26479), .CP(Clk), .Q(matrixInput[777])
         );
    VMW_FD \matrixInput_reg[474]  ( .D(n26782), .CP(Clk), .Q(matrixInput[474])
         );
    VMW_AO22 U1712 ( .A(matrixInput[177]), .B(n25096), .C(matrixInput[169]), 
        .D(n25081), .Z(n27087) );
    VMW_AO22 U1214 ( .A(matrixInput[311]), .B(n25096), .C(matrixInput[303]), 
        .D(n25081), .Z(n26953) );
    VMW_AO22 U1233 ( .A(matrixInput[295]), .B(n25096), .C(matrixInput[287]), 
        .D(n25081), .Z(n26969) );
    VMW_AO22 U2203 ( .A(matrixInput[1265]), .B(n25096), .C(matrixInput[1257]), 
        .D(n25081), .Z(n25999) );
    VMW_AO22 U2393 ( .A(matrixInput[1094]), .B(n25096), .C(matrixInput[1086]), 
        .D(n25081), .Z(n26170) );
    VMW_FD \matrixInput_reg[1153]  ( .D(n26103), .CP(Clk), .Q(matrixInput
        [1153]) );
    VMW_FD \matrixInput_reg[744]  ( .D(n26512), .CP(Clk), .Q(matrixInput[744])
         );
    VMW_AO22 U2412 ( .A(matrixInput[1077]), .B(n25096), .C(matrixInput[1069]), 
        .D(n25081), .Z(n26187) );
    VMW_OAI21 U2582 ( .A(n25147), .B(n25148), .C(n25094), .Z(n25066) );
    VMW_AO22 U1384 ( .A(matrixInput[2003]), .B(n25096), .C(matrixInput[1995]), 
        .D(n25081), .Z(n25261) );
    VMW_AO22 U1422 ( .A(matrixInput[1968]), .B(n25096), .C(matrixInput[1960]), 
        .D(n25081), .Z(n25296) );
    VMW_AO22 U1850 ( .A(matrixInput[1583]), .B(n25096), .C(matrixInput[1575]), 
        .D(n25081), .Z(n25681) );
    VMW_FD \matrixInput_reg[1249]  ( .D(n26007), .CP(Clk), .Q(matrixInput
        [1249]) );
    VMW_AO22 U2224 ( .A(matrixInput[1246]), .B(n25096), .C(matrixInput[1238]), 
        .D(n25081), .Z(n26018) );
    VMW_FD \matrixInput_reg[1777]  ( .D(n25479), .CP(Clk), .Q(matrixInput
        [1777]) );
    VMW_FD \matrixInput_reg[1250]  ( .D(n26006), .CP(Clk), .Q(matrixInput
        [1250]) );
    VMW_FD \matrixInput_reg[447]  ( .D(n26809), .CP(Clk), .Q(matrixInput[447])
         );
    VMW_FD \matrixInput_reg[179]  ( .D(n27077), .CP(Clk), .Q(matrixInput[179])
         );
    VMW_FD \matrixInput_reg[160]  ( .D(n27096), .CP(Clk), .Q(matrixInput[160])
         );
    VMW_AO22 U2435 ( .A(matrixInput[1056]), .B(n25096), .C(matrixInput[1048]), 
        .D(n25081), .Z(n26208) );
    VMW_FD \matrixInput_reg[263]  ( .D(n26993), .CP(Clk), .Q(matrixInput[263])
         );
    VMW_AO22 U1405 ( .A(matrixInput[1984]), .B(n25096), .C(matrixInput[1976]), 
        .D(n25081), .Z(n25280) );
    VMW_AO22 U1595 ( .A(matrixInput[1812]), .B(n25096), .C(matrixInput[1804]), 
        .D(n25081), .Z(n25452) );
    VMW_FD \matrixInput_reg[1474]  ( .D(n25782), .CP(Clk), .Q(matrixInput
        [1474]) );
    VMW_AO22 U1877 ( .A(matrixInput[1558]), .B(n25096), .C(matrixInput[1550]), 
        .D(n25081), .Z(n25706) );
    VMW_AO22 U2084 ( .A(matrixInput[1372]), .B(n25096), .C(matrixInput[1364]), 
        .D(n25081), .Z(n25892) );
    VMW_AO22 U2114 ( .A(matrixInput[1345]), .B(n25096), .C(matrixInput[1337]), 
        .D(n25081), .Z(n25919) );
    VMW_FD \matrixInput_reg[1744]  ( .D(n25512), .CP(Clk), .Q(matrixInput
        [1744]) );
    VMW_FD \matrixInput_reg[153]  ( .D(n27103), .CP(Clk), .Q(matrixInput[153])
         );
    VMW_AO22 U1124 ( .A(matrixInput[393]), .B(n25096), .C(matrixInput[385]), 
        .D(n25081), .Z(n26871) );
    VMW_AO22 U1735 ( .A(matrixInput[1687]), .B(n25096), .C(matrixInput[1679]), 
        .D(n25081), .Z(n25577) );
    VMW_FD \matrixInput_reg[1999]  ( .D(n25257), .CP(Clk), .Q(matrixInput
        [1999]) );
    VMW_FD \matrixInput_reg[1980]  ( .D(n25276), .CP(Clk), .Q(matrixInput
        [1980]) );
    VMW_FD \matrixInput_reg[1447]  ( .D(n25809), .CP(Clk), .Q(matrixInput
        [1447]) );
    VMW_FD \matrixInput_reg[810]  ( .D(n26446), .CP(Clk), .Q(matrixInput[810])
         );
    VMW_FD \matrixInput_reg[250]  ( .D(n27006), .CP(Clk), .Q(matrixInput[250])
         );
    VMW_FD \matrixInput_reg[249]  ( .D(n27007), .CP(Clk), .Q(matrixInput[249])
         );
    VMW_FD \matrixInput_reg[809]  ( .D(n26447), .CP(Clk), .Q(matrixInput[809])
         );
    VMW_FD \matrixInput_reg[49]  ( .D(n27207), .CP(Clk), .Q(matrixInput[49])
         );
    VMW_FD \matrixInput_reg[50]  ( .D(n27206), .CP(Clk), .Q(matrixInput[50])
         );
    VMW_AO22 U476 ( .A(matrixInput[977]), .B(n25096), .C(matrixInput[969]), 
        .D(n25081), .Z(n26287) );
    VMW_AO22 U746 ( .A(matrixInput[733]), .B(n25096), .C(matrixInput[725]), 
        .D(n25081), .Z(n26531) );
    VMW_AO22 U761 ( .A(matrixInput[719]), .B(n25096), .C(matrixInput[711]), 
        .D(n25081), .Z(n26545) );
    VMW_FD \matrixInput_reg[823]  ( .D(n26433), .CP(Clk), .Q(matrixInput[823])
         );
    VMW_AO22 U1228 ( .A(matrixInput[299]), .B(n25096), .C(matrixInput[291]), 
        .D(n25081), .Z(n26965) );
    VMW_FD \matrixInput_reg[1810]  ( .D(n25446), .CP(Clk), .Q(matrixInput
        [1810]) );
    VMW_FD \matrixInput_reg[63]  ( .D(n27193), .CP(Clk), .Q(matrixInput[63])
         );
    VMW_FD \matrixInput_reg[1809]  ( .D(n25447), .CP(Clk), .Q(matrixInput
        [1809]) );
    VMW_AO22 U1439 ( .A(matrixInput[1953]), .B(n25096), .C(matrixInput[1945]), 
        .D(n25081), .Z(n25311) );
    VMW_AO22 U2388 ( .A(matrixInput[1098]), .B(n25096), .C(matrixInput[1090]), 
        .D(n25081), .Z(n26166) );
    VMW_AO22 U2409 ( .A(matrixInput[1079]), .B(n25096), .C(matrixInput[1071]), 
        .D(n25081), .Z(n26185) );
    VMW_FD \matrixInput_reg[980]  ( .D(n26276), .CP(Clk), .Q(matrixInput[980])
         );
    VMW_AO22 U804 ( .A(matrixInput[681]), .B(n25096), .C(matrixInput[673]), 
        .D(n25081), .Z(n26583) );
    VMW_AO22 U1088 ( .A(matrixInput[425]), .B(n25096), .C(matrixInput[417]), 
        .D(n25081), .Z(n26839) );
    VMW_AO22 U1118 ( .A(matrixInput[398]), .B(n25096), .C(matrixInput[390]), 
        .D(n25081), .Z(n26866) );
    VMW_AO22 U1699 ( .A(matrixInput[1718]), .B(n25096), .C(matrixInput[1710]), 
        .D(n25081), .Z(n25546) );
    VMW_AO22 U2218 ( .A(matrixInput[1251]), .B(n25096), .C(matrixInput[1243]), 
        .D(n25081), .Z(n26013) );
    VMW_INV U2599 ( .A(Addr[0]), .Z(n25085) );
    VMW_FD \matrixInput_reg[999]  ( .D(n26257), .CP(Clk), .Q(matrixInput[999])
         );
    VMW_AO22 U1709 ( .A(matrixInput[1709]), .B(n25096), .C(matrixInput[1701]), 
        .D(n25081), .Z(n25555) );
    VMW_FD \matrixInput_reg[1823]  ( .D(n25433), .CP(Clk), .Q(matrixInput
        [1823]) );
    VMW_AO22 U994 ( .A(matrixInput[509]), .B(n25096), .C(matrixInput[501]), 
        .D(n25081), .Z(n26755) );
    VMW_AO22 U2128 ( .A(matrixInput[1332]), .B(n25096), .C(matrixInput[1324]), 
        .D(n25081), .Z(n25932) );
    VMW_PULLDOWN U268 ( .Z(n25186) );
    VMW_PULLDOWN U273 ( .Z(n25191) );
    VMW_PULLDOWN U274 ( .Z(n25192) );
    VMW_PULLDOWN U275 ( .Z(n25193) );
    VMW_PULLDOWN U282 ( .Z(n25200) );
    VMW_AO22 U503 ( .A(matrixInput[952]), .B(n25096), .C(matrixInput[944]), 
        .D(n25081), .Z(n26312) );
    VMW_AO22 U633 ( .A(matrixInput[835]), .B(n25096), .C(matrixInput[827]), 
        .D(n25081), .Z(n26429) );
    VMW_AO22 U938 ( .A(matrixInput[560]), .B(n25096), .C(matrixInput[552]), 
        .D(n25081), .Z(n26704) );
    VMW_AO22 U2014 ( .A(matrixInput[1435]), .B(n25096), .C(matrixInput[1427]), 
        .D(n25081), .Z(n25829) );
    VMW_AO22 U2184 ( .A(matrixInput[1282]), .B(n25096), .C(matrixInput[1274]), 
        .D(n25081), .Z(n25982) );
    VMW_INV U2605 ( .A(\holder[6] ), .Z(n25074) );
    VMW_FD \matrixInput_reg[143]  ( .D(n27113), .CP(Clk), .Q(matrixInput[143])
         );
    VMW_FD \matrixInput_reg[1754]  ( .D(n25502), .CP(Clk), .Q(matrixInput
        [1754]) );
    VMW_AO22 U1003 ( .A(matrixInput[502]), .B(n25096), .C(matrixInput[494]), 
        .D(n25081), .Z(n26762) );
    VMW_AO22 U1024 ( .A(matrixInput[483]), .B(n25096), .C(matrixInput[475]), 
        .D(n25081), .Z(n26781) );
    VMW_FD \matrixInput_reg[259]  ( .D(n26997), .CP(Clk), .Q(matrixInput[259])
         );
    VMW_FD \matrixInput_reg[240]  ( .D(n27016), .CP(Clk), .Q(matrixInput[240])
         );
    VMW_AO22 U1193 ( .A(matrixInput[330]), .B(n25096), .C(matrixInput[322]), 
        .D(n25081), .Z(n26934) );
    VMW_AO22 U1284 ( .A(matrixInput[248]), .B(n25096), .C(matrixInput[240]), 
        .D(n25081), .Z(n27016) );
    VMW_AO22 U1314 ( .A(matrixInput[221]), .B(n25096), .C(matrixInput[213]), 
        .D(n25081), .Z(n27043) );
    VMW_AO22 U1635 ( .A(matrixInput[1777]), .B(n25096), .C(matrixInput[1769]), 
        .D(n25081), .Z(n25487) );
    VMW_FD \matrixInput_reg[1457]  ( .D(n25799), .CP(Clk), .Q(matrixInput
        [1457]) );
    VMW_AO22 U2324 ( .A(matrixInput[1156]), .B(n25096), .C(matrixInput[1148]), 
        .D(n25081), .Z(n26108) );
    VMW_AO22 U2535 ( .A(cOutput[26]), .B(n25089), .C(cOutput[10]), .D(n25088), 
        .Z(n25153) );
    VMW_FD \matrixInput_reg[1767]  ( .D(n25489), .CP(Clk), .Q(matrixInput
        [1767]) );
    VMW_FD \matrixInput_reg[170]  ( .D(n27086), .CP(Clk), .Q(matrixInput[170])
         );
    VMW_FD \matrixInput_reg[169]  ( .D(n27087), .CP(Clk), .Q(matrixInput[169])
         );
    VMW_AO22 U1495 ( .A(matrixInput[1903]), .B(n25096), .C(matrixInput[1895]), 
        .D(n25081), .Z(n25361) );
    VMW_FD \matrixInput_reg[1464]  ( .D(n25792), .CP(Clk), .Q(matrixInput
        [1464]) );
    VMW_AO22 U1333 ( .A(matrixInput[211]), .B(n25096), .C(matrixInput[203]), 
        .D(n25081), .Z(n27053) );
    VMW_AO22 U1505 ( .A(matrixInput[1894]), .B(n25096), .C(matrixInput[1886]), 
        .D(n25081), .Z(n25370) );
    VMW_AO22 U1522 ( .A(matrixInput[1878]), .B(n25096), .C(matrixInput[1870]), 
        .D(n25081), .Z(n25386) );
    VMW_AO22 U1977 ( .A(matrixInput[1468]), .B(n25096), .C(matrixInput[1460]), 
        .D(n25081), .Z(n25796) );
    VMW_FD \matrixInput_reg[273]  ( .D(n26983), .CP(Clk), .Q(matrixInput[273])
         );
    VMW_AO22 U2293 ( .A(matrixInput[1184]), .B(n25096), .C(matrixInput[1176]), 
        .D(n25081), .Z(n26080) );
    VMW_AO22 U2303 ( .A(matrixInput[1175]), .B(n25096), .C(matrixInput[1167]), 
        .D(n25081), .Z(n26089) );
    VMW_FD \matrixInput_reg[1143]  ( .D(n26113), .CP(Clk), .Q(matrixInput
        [1143]) );
    VMW_FD \matrixInput_reg[754]  ( .D(n26502), .CP(Clk), .Q(matrixInput[754])
         );
    VMW_AO22 U2482 ( .A(matrixInput[1013]), .B(n25096), .C(matrixInput[1005]), 
        .D(n25081), .Z(n26251) );
    VMW_AO22 U2512 ( .A(cOutput[93]), .B(n25089), .C(cOutput[77]), .D(n25088), 
        .Z(n25124) );
    VMW_AO22 U1612 ( .A(matrixInput[186]), .B(n25096), .C(matrixInput[178]), 
        .D(n25081), .Z(n27078) );
    VMW_AO22 U1950 ( .A(matrixInput[1493]), .B(n25096), .C(matrixInput[1485]), 
        .D(n25081), .Z(n25771) );
    VMW_FD \matrixInput_reg[1240]  ( .D(n26016), .CP(Clk), .Q(matrixInput
        [1240]) );
    VMW_FD \matrixInput_reg[457]  ( .D(n26799), .CP(Clk), .Q(matrixInput[457])
         );
    VMW_AO22 U2033 ( .A(matrixInput[148]), .B(n25096), .C(matrixInput[140]), 
        .D(n25081), .Z(n27116) );
    VMW_FD \matrixInput_reg[1259]  ( .D(n25997), .CP(Clk), .Q(matrixInput
        [1259]) );
    VMW_BUFIZ U2622 ( .A(n25196), .E(RD), .Z(\DataOut[28]1 ) );
    VMW_FD \matrixInput_reg[1273]  ( .D(n25983), .CP(Clk), .Q(matrixInput
        [1273]) );
    VMW_FD \matrixInput_reg[1170]  ( .D(n26086), .CP(Clk), .Q(matrixInput
        [1170]) );
    VMW_FD \matrixInput_reg[1169]  ( .D(n26087), .CP(Clk), .Q(matrixInput
        [1169]) );
    VMW_FD \matrixInput_reg[767]  ( .D(n26489), .CP(Clk), .Q(matrixInput[767])
         );
    VMW_FD \matrixInput_reg[464]  ( .D(n26792), .CP(Clk), .Q(matrixInput[464])
         );
    VMW_AO22 U1782 ( .A(matrixInput[1644]), .B(n25096), .C(matrixInput[1636]), 
        .D(n25081), .Z(n25620) );
    VMW_FD \matrixInput_reg[1978]  ( .D(n25278), .CP(Clk), .Q(matrixInput
        [1978]) );
    VMW_FD \matrixInput_reg[1961]  ( .D(n25295), .CP(Clk), .Q(matrixInput
        [1961]) );
    VMW_AO22 U971 ( .A(matrixInput[530]), .B(n25096), .C(matrixInput[522]), 
        .D(n25081), .Z(n26734) );
    VMW_PULLDOWN U290 ( .Z(n25208) );
    VMW_OAI211 U300 ( .A(n25055), .B(n25074), .C(n25075), .D(n25076), .Z(
        n27386) );
    VMW_AND2 U312 ( .A(Addr[3]), .B(Addr[2]), .Z(n25094) );
    VMW_AO22 U493 ( .A(matrixInput[961]), .B(n25096), .C(matrixInput[953]), 
        .D(n25081), .Z(n26303) );
    VMW_AO22 U335 ( .A(vectorInput[15]), .B(n25095), .C(vectorInput[7]), .D(
        n25080), .Z(n27377) );
    VMW_AO22 U956 ( .A(matrixInput[544]), .B(n25096), .C(matrixInput[536]), 
        .D(n25081), .Z(n26720) );
    VMW_FD \matrixInput_reg[1952]  ( .D(n25304), .CP(Clk), .Q(matrixInput
        [1952]) );
    VMW_FD \matrixInput_reg[82]  ( .D(n27174), .CP(Clk), .Q(matrixInput[82])
         );
    VMW_FD \matrixInput_reg[978]  ( .D(n26278), .CP(Clk), .Q(matrixInput[978])
         );
    VMW_FD \matrixInput_reg[961]  ( .D(n26295), .CP(Clk), .Q(matrixInput[961])
         );
    VMW_AO22 U399 ( .A(vectorInput[29]), .B(n25095), .C(vectorInput[21]), .D(
        n25080), .Z(n27363) );
    VMW_AO22 U418 ( .A(vectorInput[19]), .B(n25095), .C(vectorInput[11]), .D(
        n25080), .Z(n27373) );
    VMW_AO22 U524 ( .A(matrixInput[933]), .B(n25096), .C(matrixInput[925]), 
        .D(n25081), .Z(n26331) );
    VMW_AO22 U588 ( .A(matrixInput[876]), .B(n25096), .C(matrixInput[868]), 
        .D(n25081), .Z(n26388) );
    VMW_AO22 U614 ( .A(matrixInput[852]), .B(n25096), .C(matrixInput[844]), 
        .D(n25081), .Z(n26412) );
    VMW_AO22 U784 ( .A(matrixInput[699]), .B(n25096), .C(matrixInput[691]), 
        .D(n25081), .Z(n26565) );
    VMW_FD \vectorInput_reg[18]  ( .D(n27366), .CP(Clk), .Q(vectorInput[18])
         );
    VMW_AO22 U728 ( .A(matrixInput[749]), .B(n25096), .C(matrixInput[741]), 
        .D(n25081), .Z(n26515) );
    VMW_AO22 U1246 ( .A(matrixInput[283]), .B(n25096), .C(matrixInput[275]), 
        .D(n25081), .Z(n26981) );
    VMW_AO22 U1457 ( .A(matrixInput[1937]), .B(n25096), .C(matrixInput[1929]), 
        .D(n25081), .Z(n25327) );
    VMW_AO22 U1889 ( .A(matrixInput[161]), .B(n25096), .C(matrixInput[153]), 
        .D(n25081), .Z(n27103) );
    VMW_AO22 U1919 ( .A(matrixInput[1520]), .B(n25096), .C(matrixInput[1512]), 
        .D(n25081), .Z(n25744) );
    VMW_FD \matrixInput_reg[952]  ( .D(n26304), .CP(Clk), .Q(matrixInput[952])
         );
    VMW_FD \matrixInput_reg[1032]  ( .D(n26224), .CP(Clk), .Q(matrixInput
        [1032]) );
    VMW_FD \vectorInput_reg[32]  ( .D(n27352), .CP(Clk), .Q(vectorInput[32])
         );
    VMW_FD \matrixInput_reg[625]  ( .D(n26631), .CP(Clk), .Q(matrixInput[625])
         );
    VMW_AO22 U1825 ( .A(matrixInput[1606]), .B(n25096), .C(matrixInput[1598]), 
        .D(n25081), .Z(n25658) );
    VMW_AO22 U2276 ( .A(matrixInput[1199]), .B(n25096), .C(matrixInput[1191]), 
        .D(n25081), .Z(n26065) );
    VMW_FD \matrixInput_reg[1331]  ( .D(n25925), .CP(Clk), .Q(matrixInput
        [1331]) );
    VMW_FD \matrixInput_reg[1328]  ( .D(n25928), .CP(Clk), .Q(matrixInput
        [1328]) );
    VMW_FD \holder_reg[4]  ( .D(n27388), .CP(Clk), .Q(\holder[4] ) );
    VMW_AO22 U2467 ( .A(matrixInput[1027]), .B(n25096), .C(matrixInput[1019]), 
        .D(n25081), .Z(n26237) );
    VMW_FD \matrixInput_reg[526]  ( .D(n26730), .CP(Clk), .Q(matrixInput[526])
         );
    VMW_AO22 U1176 ( .A(matrixInput[346]), .B(n25096), .C(matrixInput[338]), 
        .D(n25081), .Z(n26918) );
    VMW_AO22 U1767 ( .A(matrixInput[172]), .B(n25096), .C(matrixInput[164]), 
        .D(n25081), .Z(n27092) );
    VMW_FD \matrixInput_reg[1485]  ( .D(n25771), .CP(Clk), .Q(matrixInput
        [1485]) );
    VMW_FD \matrixInput_reg[292]  ( .D(n26964), .CP(Clk), .Q(matrixInput[292])
         );
    VMW_FD \matrixInput_reg[616]  ( .D(n26640), .CP(Clk), .Q(matrixInput[616])
         );
    VMW_FD \matrixInput_reg[1018]  ( .D(n26238), .CP(Clk), .Q(matrixInput
        [1018]) );
    VMW_FD \matrixInput_reg[1001]  ( .D(n26255), .CP(Clk), .Q(matrixInput
        [1001]) );
    VMW_AO22 U2146 ( .A(matrixInput[1316]), .B(n25096), .C(matrixInput[1308]), 
        .D(n25081), .Z(n25948) );
    VMW_FD \matrixInput_reg[515]  ( .D(n26741), .CP(Clk), .Q(matrixInput[515])
         );
    VMW_AO22 U481 ( .A(matrixInput[972]), .B(n25096), .C(matrixInput[964]), 
        .D(n25081), .Z(n26292) );
    VMW_AO22 U621 ( .A(matrixInput[846]), .B(n25096), .C(matrixInput[838]), 
        .D(n25081), .Z(n26418) );
    VMW_AO22 U878 ( .A(matrixInput[614]), .B(n25096), .C(matrixInput[606]), 
        .D(n25081), .Z(n26650) );
    VMW_AO22 U1151 ( .A(matrixInput[368]), .B(n25096), .C(matrixInput[360]), 
        .D(n25081), .Z(n26896) );
    VMW_FD \matrixInput_reg[1786]  ( .D(n25470), .CP(Clk), .Q(matrixInput
        [1786]) );
    VMW_FD \matrixInput_reg[1302]  ( .D(n25954), .CP(Clk), .Q(matrixInput
        [1302]) );
    VMW_FD \matrixInput_reg[1625]  ( .D(n25631), .CP(Clk), .Q(matrixInput
        [1625]) );
    VMW_FD \matrixInput_reg[191]  ( .D(n27065), .CP(Clk), .Q(matrixInput[191])
         );
    VMW_FD \matrixInput_reg[188]  ( .D(n27068), .CP(Clk), .Q(matrixInput[188])
         );
    VMW_AO22 U1164 ( .A(matrixInput[357]), .B(n25096), .C(matrixInput[349]), 
        .D(n25081), .Z(n26907) );
    VMW_AO22 U1254 ( .A(matrixInput[276]), .B(n25096), .C(matrixInput[268]), 
        .D(n25081), .Z(n26988) );
    VMW_AO22 U1261 ( .A(matrixInput[269]), .B(n25096), .C(matrixInput[261]), 
        .D(n25081), .Z(n26995) );
    VMW_AO22 U1740 ( .A(matrixInput[1682]), .B(n25096), .C(matrixInput[1674]), 
        .D(n25081), .Z(n25582) );
    VMW_AO22 U2161 ( .A(matrixInput[1303]), .B(n25096), .C(matrixInput[1295]), 
        .D(n25081), .Z(n25961) );
    VMW_FD \matrixInput_reg[2042]  ( .D(n25214), .CP(Clk), .Q(matrixInput
        [2042]) );
    VMW_FD \matrixInput_reg[1526]  ( .D(n25730), .CP(Clk), .Q(matrixInput
        [1526]) );
    VMW_FD \matrixInput_reg[331]  ( .D(n26925), .CP(Clk), .Q(matrixInput[331])
         );
    VMW_FD \matrixInput_reg[328]  ( .D(n26928), .CP(Clk), .Q(matrixInput[328])
         );
    VMW_AO22 U1470 ( .A(matrixInput[1925]), .B(n25096), .C(matrixInput[1917]), 
        .D(n25081), .Z(n25339) );
    VMW_AO22 U1802 ( .A(matrixInput[1626]), .B(n25096), .C(matrixInput[1618]), 
        .D(n25081), .Z(n25638) );
    VMW_AO22 U1992 ( .A(matrixInput[1455]), .B(n25096), .C(matrixInput[1447]), 
        .D(n25081), .Z(n25809) );
    VMW_FD \matrixInput_reg[1292]  ( .D(n25964), .CP(Clk), .Q(matrixInput
        [1292]) );
    VMW_FD \matrixInput_reg[485]  ( .D(n26771), .CP(Clk), .Q(matrixInput[485])
         );
    VMW_AO22 U1837 ( .A(matrixInput[1595]), .B(n25096), .C(matrixInput[1587]), 
        .D(n25081), .Z(n25669) );
    VMW_AO22 U2251 ( .A(matrixInput[1221]), .B(n25096), .C(matrixInput[1213]), 
        .D(n25081), .Z(n26043) );
    VMW_AO22 U2440 ( .A(matrixInput[1051]), .B(n25096), .C(matrixInput[1043]), 
        .D(n25081), .Z(n26213) );
    VMW_FD \matrixInput_reg[1616]  ( .D(n25640), .CP(Clk), .Q(matrixInput
        [1616]) );
    VMW_FD \matrixInput_reg[1515]  ( .D(n25741), .CP(Clk), .Q(matrixInput
        [1515]) );
    VMW_FD \matrixInput_reg[302]  ( .D(n26954), .CP(Clk), .Q(matrixInput[302])
         );
    VMW_FD \matrixInput_reg[1191]  ( .D(n26065), .CP(Clk), .Q(matrixInput
        [1191]) );
    VMW_FD \matrixInput_reg[1188]  ( .D(n26068), .CP(Clk), .Q(matrixInput
        [1188]) );
    VMW_FD \matrixInput_reg[786]  ( .D(n26470), .CP(Clk), .Q(matrixInput[786])
         );
    VMW_AO22 U1445 ( .A(matrixInput[201]), .B(n25096), .C(matrixInput[193]), 
        .D(n25081), .Z(n27063) );
    VMW_FD \matrixInput_reg[1470]  ( .D(n25786), .CP(Clk), .Q(matrixInput
        [1470]) );
    VMW_FD \matrixInput_reg[1469]  ( .D(n25787), .CP(Clk), .Q(matrixInput
        [1469]) );
    VMW_AO22 U2264 ( .A(matrixInput[1209]), .B(n25096), .C(matrixInput[1201]), 
        .D(n25081), .Z(n26055) );
    VMW_AO22 U2475 ( .A(matrixInput[1019]), .B(n25096), .C(matrixInput[1011]), 
        .D(n25081), .Z(n26245) );
    VMW_FD \matrixInput_reg[267]  ( .D(n26989), .CP(Clk), .Q(matrixInput[267])
         );
    VMW_FD \matrixInput_reg[1773]  ( .D(n25483), .CP(Clk), .Q(matrixInput
        [1773]) );
    VMW_FD \matrixInput_reg[254]  ( .D(n27002), .CP(Clk), .Q(matrixInput[254])
         );
    VMW_FD \matrixInput_reg[164]  ( .D(n27092), .CP(Clk), .Q(matrixInput[164])
         );
    VMW_AO22 U1775 ( .A(matrixInput[1650]), .B(n25096), .C(matrixInput[1642]), 
        .D(n25081), .Z(n25614) );
    VMW_FD \matrixInput_reg[1443]  ( .D(n25813), .CP(Clk), .Q(matrixInput
        [1443]) );
    VMW_AO22 U1143 ( .A(matrixInput[376]), .B(n25096), .C(matrixInput[368]), 
        .D(n25081), .Z(n26888) );
    VMW_AO22 U1752 ( .A(matrixInput[1671]), .B(n25096), .C(matrixInput[1663]), 
        .D(n25081), .Z(n25593) );
    VMW_AO22 U2154 ( .A(matrixInput[1308]), .B(n25096), .C(matrixInput[1300]), 
        .D(n25081), .Z(n25956) );
    VMW_FD \matrixInput_reg[1759]  ( .D(n25497), .CP(Clk), .Q(matrixInput
        [1759]) );
    VMW_FD \matrixInput_reg[157]  ( .D(n27099), .CP(Clk), .Q(matrixInput[157])
         );
    VMW_FD \matrixInput_reg[1740]  ( .D(n25516), .CP(Clk), .Q(matrixInput
        [1740]) );
    VMW_AO22 U1273 ( .A(matrixInput[258]), .B(n25096), .C(matrixInput[250]), 
        .D(n25081), .Z(n27006) );
    VMW_AO22 U1462 ( .A(matrixInput[1932]), .B(n25096), .C(matrixInput[1924]), 
        .D(n25081), .Z(n25332) );
    VMW_AO22 U1810 ( .A(matrixInput[1618]), .B(n25096), .C(matrixInput[1610]), 
        .D(n25081), .Z(n25646) );
    VMW_AO22 U2173 ( .A(matrixInput[1292]), .B(n25096), .C(matrixInput[1284]), 
        .D(n25081), .Z(n25972) );
    VMW_FD \matrixInput_reg[1267]  ( .D(n25989), .CP(Clk), .Q(matrixInput
        [1267]) );
    VMW_FD \matrixInput_reg[1164]  ( .D(n26092), .CP(Clk), .Q(matrixInput
        [1164]) );
    VMW_FD \matrixInput_reg[470]  ( .D(n26786), .CP(Clk), .Q(matrixInput[470])
         );
    VMW_FD \matrixInput_reg[469]  ( .D(n26787), .CP(Clk), .Q(matrixInput[469])
         );
    VMW_FD \matrixInput_reg[773]  ( .D(n26483), .CP(Clk), .Q(matrixInput[773])
         );
    VMW_FD \matrixInput_reg[1254]  ( .D(n26002), .CP(Clk), .Q(matrixInput
        [1254]) );
    VMW_FD \matrixInput_reg[443]  ( .D(n26813), .CP(Clk), .Q(matrixInput[443])
         );
    VMW_AO22 U1980 ( .A(matrixInput[1466]), .B(n25096), .C(matrixInput[1458]), 
        .D(n25081), .Z(n25798) );
    VMW_AO22 U2243 ( .A(matrixInput[1228]), .B(n25096), .C(matrixInput[1220]), 
        .D(n25081), .Z(n26036) );
    VMW_AO22 U2452 ( .A(matrixInput[1040]), .B(n25096), .C(matrixInput[1032]), 
        .D(n25081), .Z(n26224) );
    VMW_FD \matrixInput_reg[1157]  ( .D(n26099), .CP(Clk), .Q(matrixInput
        [1157]) );
    VMW_FD \matrixInput_reg[759]  ( .D(n26497), .CP(Clk), .Q(matrixInput[759])
         );
    VMW_FD \matrixInput_reg[740]  ( .D(n26516), .CP(Clk), .Q(matrixInput[740])
         );
    VMW_FD \matrixInput_reg[77]  ( .D(n27179), .CP(Clk), .Q(matrixInput[77])
         );
    VMW_FD \matrixInput_reg[837]  ( .D(n26419), .CP(Clk), .Q(matrixInput[837])
         );
    VMW_AO22 U511 ( .A(matrixInput[945]), .B(n25096), .C(matrixInput[937]), 
        .D(n25081), .Z(n26319) );
    VMW_AO22 U327 ( .A(vectorInput[95]), .B(n25095), .C(vectorInput[87]), .D(
        n25080), .Z(n27297) );
    VMW_AO22 U536 ( .A(matrixInput[922]), .B(n25096), .C(matrixInput[914]), 
        .D(n25081), .Z(n26342) );
    VMW_AO22 U963 ( .A(matrixInput[60]), .B(n25096), .C(matrixInput[52]), .D(
        n25081), .Z(n27204) );
    VMW_FD \matrixInput_reg[1994]  ( .D(n25262), .CP(Clk), .Q(matrixInput
        [1994]) );
    VMW_FD \matrixInput_reg[44]  ( .D(n27212), .CP(Clk), .Q(matrixInput[44])
         );
    VMW_FD \matrixInput_reg[804]  ( .D(n26452), .CP(Clk), .Q(matrixInput[804])
         );
    VMW_AO22 U2068 ( .A(matrixInput[1387]), .B(n25096), .C(matrixInput[1379]), 
        .D(n25081), .Z(n25877) );
    VMW_AO22 U349 ( .A(vectorInput[75]), .B(n25095), .C(vectorInput[67]), .D(
        n25080), .Z(n27317) );
    VMW_AO22 U606 ( .A(matrixInput[859]), .B(n25096), .C(matrixInput[851]), 
        .D(n25081), .Z(n26405) );
    VMW_AO22 U944 ( .A(matrixInput[555]), .B(n25096), .C(matrixInput[547]), 
        .D(n25081), .Z(n26709) );
    VMW_AO22 U1058 ( .A(matrixInput[452]), .B(n25096), .C(matrixInput[444]), 
        .D(n25081), .Z(n26812) );
    VMW_FD \matrixInput_reg[1837]  ( .D(n25419), .CP(Clk), .Q(matrixInput
        [1837]) );
    VMW_AO22 U1649 ( .A(matrixInput[1764]), .B(n25096), .C(matrixInput[1756]), 
        .D(n25081), .Z(n25500) );
    VMW_AO22 U2549 ( .A(cOutput[113]), .B(n25087), .C(cOutput[97]), .D(n25084), 
        .Z(n25169) );
    VMW_FD \matrixInput_reg[994]  ( .D(n26262), .CP(Clk), .Q(matrixInput[994])
         );
    VMW_AO22 U796 ( .A(matrixInput[688]), .B(n25096), .C(matrixInput[680]), 
        .D(n25081), .Z(n26576) );
    VMW_AO22 U2358 ( .A(matrixInput[1125]), .B(n25096), .C(matrixInput[1117]), 
        .D(n25081), .Z(n26139) );
    VMW_AO22 U1368 ( .A(matrixInput[2016]), .B(n25096), .C(matrixInput[2008]), 
        .D(n25081), .Z(n25248) );
    VMW_AO22 U1579 ( .A(matrixInput[1827]), .B(n25096), .C(matrixInput[1819]), 
        .D(n25081), .Z(n25437) );
    VMW_AO22 U2006 ( .A(matrixInput[1442]), .B(n25096), .C(matrixInput[1434]), 
        .D(n25081), .Z(n25822) );
    VMW_FD \matrixInput_reg[1804]  ( .D(n25452), .CP(Clk), .Q(matrixInput
        [1804]) );
    VMW_FD \matrixInput_reg[1792]  ( .D(n25464), .CP(Clk), .Q(matrixInput
        [1792]) );
    VMW_FD \matrixInput_reg[185]  ( .D(n27071), .CP(Clk), .Q(matrixInput[185])
         );
    VMW_AO22 U443 ( .A(matrixInput[1007]), .B(n25096), .C(matrixInput[999]), 
        .D(n25081), .Z(n26257) );
    VMW_AO22 U558 ( .A(matrixInput[903]), .B(n25096), .C(matrixInput[895]), 
        .D(n25081), .Z(n26361) );
    VMW_BUFIZ U2617 ( .A(n25192), .E(RD), .Z(\DataOut[16]1 ) );
    VMW_FD \matrixInput_reg[518]  ( .D(n26738), .CP(Clk), .Q(matrixInput[518])
         );
    VMW_AO22 U668 ( .A(matrixInput[804]), .B(n25096), .C(matrixInput[796]), 
        .D(n25081), .Z(n26460) );
    VMW_AO22 U1036 ( .A(matrixInput[472]), .B(n25096), .C(matrixInput[464]), 
        .D(n25081), .Z(n26792) );
    VMW_AO22 U1627 ( .A(matrixInput[1784]), .B(n25096), .C(matrixInput[1776]), 
        .D(n25081), .Z(n25480) );
    VMW_AO22 U2196 ( .A(matrixInput[1271]), .B(n25096), .C(matrixInput[1263]), 
        .D(n25081), .Z(n25993) );
    VMW_FD \matrixInput_reg[1316]  ( .D(n25940), .CP(Clk), .Q(matrixInput
        [1316]) );
    VMW_FD \matrixInput_reg[501]  ( .D(n26755), .CP(Clk), .Q(matrixInput[501])
         );
    VMW_FD \matrixInput_reg[602]  ( .D(n26654), .CP(Clk), .Q(matrixInput[602])
         );
    VMW_AO22 U2336 ( .A(matrixInput[1145]), .B(n25096), .C(matrixInput[1137]), 
        .D(n25081), .Z(n26119) );
    VMW_FD \matrixInput_reg[1491]  ( .D(n25765), .CP(Clk), .Q(matrixInput
        [1491]) );
    VMW_FD \matrixInput_reg[1488]  ( .D(n25768), .CP(Clk), .Q(matrixInput
        [1488]) );
    VMW_FD \matrixInput_reg[1015]  ( .D(n26241), .CP(Clk), .Q(matrixInput
        [1015]) );
    VMW_FD \matrixInput_reg[1325]  ( .D(n25931), .CP(Clk), .Q(matrixInput
        [1325]) );
    VMW_FD \matrixInput_reg[286]  ( .D(n26970), .CP(Clk), .Q(matrixInput[286])
         );
    VMW_AO22 U2527 ( .A(cOutput[51]), .B(n25087), .C(cOutput[35]), .D(n25084), 
        .Z(n25143) );
    VMW_FD \matrixInput_reg[532]  ( .D(n26724), .CP(Clk), .Q(matrixInput[532])
         );
    VMW_AO22 U1011 ( .A(matrixInput[495]), .B(n25096), .C(matrixInput[487]), 
        .D(n25081), .Z(n26769) );
    VMW_AO22 U1296 ( .A(matrixInput[30]), .B(n25096), .C(matrixInput[22]), .D(
        n25081), .Z(n27234) );
    VMW_AO22 U1965 ( .A(matrixInput[1479]), .B(n25096), .C(matrixInput[1471]), 
        .D(n25081), .Z(n25785) );
    VMW_FD \matrixInput_reg[1026]  ( .D(n26230), .CP(Clk), .Q(matrixInput
        [1026]) );
    VMW_FD \matrixInput_reg[631]  ( .D(n26625), .CP(Clk), .Q(matrixInput[631])
         );
    VMW_AO22 U1306 ( .A(matrixInput[228]), .B(n25096), .C(matrixInput[220]), 
        .D(n25081), .Z(n27036) );
    VMW_AO22 U1517 ( .A(matrixInput[1883]), .B(n25096), .C(matrixInput[1875]), 
        .D(n25081), .Z(n25381) );
    VMW_FD \matrixInput_reg[628]  ( .D(n26628), .CP(Clk), .Q(matrixInput[628])
         );
    VMW_AO22 U1321 ( .A(matrixInput[215]), .B(n25096), .C(matrixInput[207]), 
        .D(n25081), .Z(n27049) );
    VMW_AO22 U1487 ( .A(matrixInput[1909]), .B(n25096), .C(matrixInput[1901]), 
        .D(n25081), .Z(n25355) );
    VMW_AO22 U1942 ( .A(matrixInput[1500]), .B(n25096), .C(matrixInput[1492]), 
        .D(n25081), .Z(n25764) );
    VMW_AO22 U2281 ( .A(matrixInput[1195]), .B(n25096), .C(matrixInput[1187]), 
        .D(n25081), .Z(n26069) );
    VMW_AO22 U2311 ( .A(matrixInput[123]), .B(n25096), .C(matrixInput[115]), 
        .D(n25081), .Z(n27141) );
    VMW_AO22 U2500 ( .A(cOutput[54]), .B(n25087), .C(cOutput[38]), .D(n25084), 
        .Z(n25110) );
    VMW_FD \matrixInput_reg[1185]  ( .D(n26071), .CP(Clk), .Q(matrixInput
        [1185]) );
    VMW_AO22 U2490 ( .A(cOutput[31]), .B(n25089), .C(cOutput[15]), .D(n25088), 
        .Z(n25098) );
    VMW_FD \matrixInput_reg[1518]  ( .D(n25738), .CP(Clk), .Q(matrixInput
        [1518]) );
    VMW_FD \matrixInput_reg[792]  ( .D(n26464), .CP(Clk), .Q(matrixInput[792])
         );
    VMW_FD \matrixInput_reg[316]  ( .D(n26940), .CP(Clk), .Q(matrixInput[316])
         );
    VMW_FD \matrixInput_reg[1501]  ( .D(n25755), .CP(Clk), .Q(matrixInput
        [1501]) );
    VMW_FD \matrixInput_reg[1602]  ( .D(n25654), .CP(Clk), .Q(matrixInput
        [1602]) );
    VMW_AO22 U1530 ( .A(matrixInput[1871]), .B(n25096), .C(matrixInput[1863]), 
        .D(n25081), .Z(n25393) );
    VMW_AO22 U1790 ( .A(matrixInput[1637]), .B(n25096), .C(matrixInput[1629]), 
        .D(n25081), .Z(n25627) );
    VMW_AO22 U2021 ( .A(matrixInput[1428]), .B(n25096), .C(matrixInput[1420]), 
        .D(n25081), .Z(n25836) );
    VMW_BUFIZ U2630 ( .A(n25203), .E(RD), .Z(\DataOut[17]1 ) );
    VMW_FD \matrixInput_reg[1532]  ( .D(n25724), .CP(Clk), .Q(matrixInput
        [1532]) );
    VMW_FD \matrixInput_reg[1286]  ( .D(n25970), .CP(Clk), .Q(matrixInput
        [1286]) );
    VMW_FD \matrixInput_reg[491]  ( .D(n26765), .CP(Clk), .Q(matrixInput[491])
         );
    VMW_FD \matrixInput_reg[488]  ( .D(n26768), .CP(Clk), .Q(matrixInput[488])
         );
    VMW_FD \matrixInput_reg[325]  ( .D(n26931), .CP(Clk), .Q(matrixInput[325])
         );
    VMW_AO22 U1181 ( .A(matrixInput[341]), .B(n25096), .C(matrixInput[333]), 
        .D(n25081), .Z(n26923) );
    VMW_AO22 U1600 ( .A(matrixInput[25]), .B(n25096), .C(matrixInput[17]), .D(
        n25081), .Z(n27239) );
    VMW_FD \matrixInput_reg[1631]  ( .D(n25625), .CP(Clk), .Q(matrixInput
        [1631]) );
    VMW_FD \matrixInput_reg[1628]  ( .D(n25628), .CP(Clk), .Q(matrixInput
        [1628]) );
    VMW_AO22 U754 ( .A(matrixInput[726]), .B(n25096), .C(matrixInput[718]), 
        .D(n25081), .Z(n26538) );
    VMW_AO22 U773 ( .A(matrixInput[708]), .B(n25096), .C(matrixInput[700]), 
        .D(n25081), .Z(n26556) );
    VMW_AO22 U831 ( .A(matrixInput[657]), .B(n25096), .C(matrixInput[649]), 
        .D(n25081), .Z(n26607) );
    VMW_FD \matrixInput_reg[1946]  ( .D(n25310), .CP(Clk), .Q(matrixInput
        [1946]) );
    VMW_FD \matrixInput_reg[96]  ( .D(n27160), .CP(Clk), .Q(matrixInput[96])
         );
    VMW_FD \matrixInput_reg[1975]  ( .D(n25281), .CP(Clk), .Q(matrixInput
        [1975]) );
    VMW_AO22 U1859 ( .A(matrixInput[1575]), .B(n25096), .C(matrixInput[1567]), 
        .D(n25081), .Z(n25689) );
    VMW_FD \matrixInput_reg[946]  ( .D(n26310), .CP(Clk), .Q(matrixInput[946])
         );
    VMW_FD \vectorInput_reg[26]  ( .D(n27358), .CP(Clk), .Q(vectorInput[26])
         );
    VMW_FD \vectorInput_reg[15]  ( .D(n27369), .CP(Clk), .Q(vectorInput[15])
         );
    VMW_PULLDOWN U283 ( .Z(n25201) );
    VMW_AO22 U313 ( .A(vectorInput[17]), .B(n25095), .C(vectorInput[9]), .D(
        n25080), .Z(n27375) );
    VMW_AO22 U352 ( .A(vectorInput[72]), .B(n25095), .C(vectorInput[64]), .D(
        n25080), .Z(n27320) );
    VMW_AO22 U375 ( .A(vectorInput[51]), .B(n25095), .C(vectorInput[43]), .D(
        n25080), .Z(n27341) );
    VMW_AO22 U458 ( .A(matrixInput[993]), .B(n25096), .C(matrixInput[985]), 
        .D(n25081), .Z(n26271) );
    VMW_AO22 U464 ( .A(matrixInput[105]), .B(n25096), .C(matrixInput[97]), .D(
        n25081), .Z(n27159) );
    VMW_AO22 U768 ( .A(matrixInput[713]), .B(n25096), .C(matrixInput[705]), 
        .D(n25081), .Z(n26551) );
    VMW_AO22 U816 ( .A(matrixInput[670]), .B(n25096), .C(matrixInput[662]), 
        .D(n25081), .Z(n26594) );
    VMW_AO22 U986 ( .A(matrixInput[517]), .B(n25096), .C(matrixInput[509]), 
        .D(n25081), .Z(n26747) );
    VMW_AO22 U1081 ( .A(matrixInput[431]), .B(n25096), .C(matrixInput[423]), 
        .D(n25081), .Z(n26833) );
    VMW_AO22 U1700 ( .A(matrixInput[178]), .B(n25096), .C(matrixInput[170]), 
        .D(n25081), .Z(n27086) );
    VMW_AO22 U2121 ( .A(matrixInput[1338]), .B(n25096), .C(matrixInput[1330]), 
        .D(n25081), .Z(n25926) );
    VMW_FD \matrixInput_reg[1522]  ( .D(n25734), .CP(Clk), .Q(matrixInput
        [1522]) );
    VMW_FD \matrixInput_reg[975]  ( .D(n26281), .CP(Clk), .Q(matrixInput[975])
         );
    VMW_FD \matrixInput_reg[335]  ( .D(n26921), .CP(Clk), .Q(matrixInput[335])
         );
    VMW_FD \matrixInput_reg[2046]  ( .D(n25210), .CP(Clk), .Q(matrixInput
        [2046]) );
    VMW_AO22 U1111 ( .A(matrixInput[405]), .B(n25096), .C(matrixInput[397]), 
        .D(n25081), .Z(n26859) );
    VMW_AO22 U1690 ( .A(matrixInput[1727]), .B(n25096), .C(matrixInput[1719]), 
        .D(n25081), .Z(n25537) );
    VMW_AO22 U1221 ( .A(matrixInput[306]), .B(n25096), .C(matrixInput[298]), 
        .D(n25081), .Z(n26958) );
    VMW_AO22 U1430 ( .A(matrixInput[1961]), .B(n25096), .C(matrixInput[1953]), 
        .D(n25081), .Z(n25303) );
    VMW_AO22 U1842 ( .A(matrixInput[1590]), .B(n25096), .C(matrixInput[1582]), 
        .D(n25081), .Z(n25674) );
    VMW_AO22 U2211 ( .A(matrixInput[132]), .B(n25096), .C(matrixInput[124]), 
        .D(n25081), .Z(n27132) );
    VMW_FD \matrixInput_reg[1638]  ( .D(n25618), .CP(Clk), .Q(matrixInput
        [1638]) );
    VMW_FD \matrixInput_reg[1621]  ( .D(n25635), .CP(Clk), .Q(matrixInput
        [1621]) );
    VMW_FD \matrixInput_reg[782]  ( .D(n26474), .CP(Clk), .Q(matrixInput[782])
         );
    VMW_AO22 U2381 ( .A(matrixInput[1105]), .B(n25096), .C(matrixInput[1097]), 
        .D(n25081), .Z(n26159) );
    VMW_OAI21 U2590 ( .A(n25169), .B(n25170), .C(n25094), .Z(n25060) );
    VMW_AO22 U2400 ( .A(matrixInput[115]), .B(n25096), .C(matrixInput[107]), 
        .D(n25081), .Z(n27149) );
    VMW_FD \matrixInput_reg[1612]  ( .D(n25644), .CP(Clk), .Q(matrixInput
        [1612]) );
    VMW_FD \matrixInput_reg[1511]  ( .D(n25745), .CP(Clk), .Q(matrixInput
        [1511]) );
    VMW_FD \matrixInput_reg[1195]  ( .D(n26061), .CP(Clk), .Q(matrixInput
        [1195]) );
    VMW_FD \matrixInput_reg[1508]  ( .D(n25748), .CP(Clk), .Q(matrixInput
        [1508]) );
    VMW_FD \matrixInput_reg[306]  ( .D(n26950), .CP(Clk), .Q(matrixInput[306])
         );
    VMW_FD \matrixInput_reg[1296]  ( .D(n25960), .CP(Clk), .Q(matrixInput
        [1296]) );
    VMW_FD \matrixInput_reg[498]  ( .D(n26758), .CP(Clk), .Q(matrixInput[498])
         );
    VMW_FD \matrixInput_reg[481]  ( .D(n26775), .CP(Clk), .Q(matrixInput[481])
         );
    VMW_AO22 U2427 ( .A(matrixInput[1063]), .B(n25096), .C(matrixInput[1055]), 
        .D(n25081), .Z(n26201) );
    VMW_FD \matrixInput_reg[522]  ( .D(n26734), .CP(Clk), .Q(matrixInput[522])
         );
    VMW_AO22 U1206 ( .A(matrixInput[318]), .B(n25096), .C(matrixInput[310]), 
        .D(n25081), .Z(n26946) );
    VMW_AO22 U1865 ( .A(matrixInput[1569]), .B(n25096), .C(matrixInput[1561]), 
        .D(n25081), .Z(n25695) );
    VMW_AO22 U2236 ( .A(matrixInput[1235]), .B(n25096), .C(matrixInput[1227]), 
        .D(n25081), .Z(n26029) );
    VMW_FD \matrixInput_reg[1335]  ( .D(n25921), .CP(Clk), .Q(matrixInput
        [1335]) );
    VMW_FD \holder_reg[0]  ( .D(n27392), .CP(Clk), .Q(\holder[0] ) );
    VMW_FD \matrixInput_reg[638]  ( .D(n26618), .CP(Clk), .Q(matrixInput[638])
         );
    VMW_AO22 U1396 ( .A(matrixInput[1992]), .B(n25096), .C(matrixInput[1984]), 
        .D(n25081), .Z(n25272) );
    VMW_AO22 U1587 ( .A(matrixInput[1819]), .B(n25096), .C(matrixInput[1811]), 
        .D(n25081), .Z(n25445) );
    VMW_FD \matrixInput_reg[621]  ( .D(n26635), .CP(Clk), .Q(matrixInput[621])
         );
    VMW_AO22 U1417 ( .A(matrixInput[1973]), .B(n25096), .C(matrixInput[1965]), 
        .D(n25081), .Z(n25291) );
    VMW_FD \matrixInput_reg[1782]  ( .D(n25474), .CP(Clk), .Q(matrixInput
        [1782]) );
    VMW_FD \matrixInput_reg[1036]  ( .D(n26220), .CP(Clk), .Q(matrixInput
        [1036]) );
    VMW_FD \matrixInput_reg[195]  ( .D(n27061), .CP(Clk), .Q(matrixInput[195])
         );
    VMW_FD \matrixInput_reg[1306]  ( .D(n25950), .CP(Clk), .Q(matrixInput
        [1306]) );
    VMW_AO22 U564 ( .A(matrixInput[96]), .B(n25096), .C(matrixInput[88]), .D(
        n25081), .Z(n27168) );
    VMW_AO22 U1136 ( .A(matrixInput[382]), .B(n25096), .C(matrixInput[374]), 
        .D(n25081), .Z(n26882) );
    VMW_AO22 U2096 ( .A(matrixInput[1361]), .B(n25096), .C(matrixInput[1353]), 
        .D(n25081), .Z(n25903) );
    VMW_AO22 U2106 ( .A(matrixInput[1352]), .B(n25096), .C(matrixInput[1344]), 
        .D(n25081), .Z(n25912) );
    VMW_FD \matrixInput_reg[511]  ( .D(n26745), .CP(Clk), .Q(matrixInput[511])
         );
    VMW_FD \matrixInput_reg[1005]  ( .D(n26251), .CP(Clk), .Q(matrixInput
        [1005]) );
    VMW_FD \matrixInput_reg[508]  ( .D(n26748), .CP(Clk), .Q(matrixInput[508])
         );
    VMW_AO22 U1727 ( .A(matrixInput[1694]), .B(n25096), .C(matrixInput[1686]), 
        .D(n25081), .Z(n25570) );
    VMW_FD \matrixInput_reg[1498]  ( .D(n25758), .CP(Clk), .Q(matrixInput
        [1498]) );
    VMW_FD \matrixInput_reg[1481]  ( .D(n25775), .CP(Clk), .Q(matrixInput
        [1481]) );
    VMW_FD \matrixInput_reg[612]  ( .D(n26644), .CP(Clk), .Q(matrixInput[612])
         );
    VMW_FD \matrixInput_reg[296]  ( .D(n26960), .CP(Clk), .Q(matrixInput[296])
         );
    VMW_AO22 U654 ( .A(matrixInput[816]), .B(n25096), .C(matrixInput[808]), 
        .D(n25081), .Z(n26448) );
    VMW_AO22 U886 ( .A(matrixInput[67]), .B(n25096), .C(matrixInput[59]), .D(
        n25081), .Z(n27197) );
    VMW_AO22 U916 ( .A(matrixInput[580]), .B(n25096), .C(matrixInput[572]), 
        .D(n25081), .Z(n26684) );
    VMW_FD \matrixInput_reg[965]  ( .D(n26291), .CP(Clk), .Q(matrixInput[965])
         );
    VMW_AO22 U1959 ( .A(matrixInput[1485]), .B(n25096), .C(matrixInput[1477]), 
        .D(n25081), .Z(n25779) );
    VMW_FD \vectorInput_reg[36]  ( .D(n27348), .CP(Clk), .Q(vectorInput[36])
         );
    VMW_FD \matrixInput_reg[956]  ( .D(n26300), .CP(Clk), .Q(matrixInput[956])
         );
    VMW_AO22 U673 ( .A(matrixInput[799]), .B(n25096), .C(matrixInput[791]), 
        .D(n25081), .Z(n26465) );
    VMW_FD \matrixInput_reg[1965]  ( .D(n25291), .CP(Clk), .Q(matrixInput
        [1965]) );
    VMW_FD \matrixInput_reg[1956]  ( .D(n25300), .CP(Clk), .Q(matrixInput
        [1956]) );
    VMW_FD \matrixInput_reg[86]  ( .D(n27170), .CP(Clk), .Q(matrixInput[86])
         );
    VMW_AO22 U390 ( .A(vectorInput[10]), .B(n25095), .C(vectorInput[2]), .D(
        n25080), .Z(n27382) );
    VMW_AO22 U411 ( .A(DataIn[6]), .B(n25095), .C(vectorInput[126]), .D(n25080
        ), .Z(n27258) );
    VMW_AO22 U436 ( .A(vectorInput[111]), .B(n25095), .C(vectorInput[103]), 
        .D(n25080), .Z(n27281) );
    VMW_AO22 U543 ( .A(matrixInput[916]), .B(n25096), .C(matrixInput[908]), 
        .D(n25081), .Z(n26348) );
    VMW_AO22 U696 ( .A(matrixInput[778]), .B(n25096), .C(matrixInput[770]), 
        .D(n25081), .Z(n26486) );
    VMW_AO22 U931 ( .A(matrixInput[567]), .B(n25096), .C(matrixInput[559]), 
        .D(n25081), .Z(n26697) );
    VMW_AO22 U978 ( .A(matrixInput[524]), .B(n25096), .C(matrixInput[516]), 
        .D(n25081), .Z(n26740) );
    VMW_AO22 U1043 ( .A(matrixInput[466]), .B(n25096), .C(matrixInput[458]), 
        .D(n25081), .Z(n26798) );
    VMW_AO22 U1373 ( .A(matrixInput[2011]), .B(n25096), .C(matrixInput[2003]), 
        .D(n25081), .Z(n25253) );
    VMW_AO22 U1880 ( .A(matrixInput[1556]), .B(n25096), .C(matrixInput[1548]), 
        .D(n25081), .Z(n25708) );
    VMW_AO22 U1910 ( .A(matrixInput[1528]), .B(n25096), .C(matrixInput[1520]), 
        .D(n25081), .Z(n25736) );
    VMW_FD \matrixInput_reg[1244]  ( .D(n26012), .CP(Clk), .Q(matrixInput
        [1244]) );
    VMW_FD \matrixInput_reg[453]  ( .D(n26803), .CP(Clk), .Q(matrixInput[453])
         );
    VMW_AO22 U1562 ( .A(matrixInput[1842]), .B(n25096), .C(matrixInput[1834]), 
        .D(n25081), .Z(n25422) );
    VMW_AO22 U2343 ( .A(matrixInput[1138]), .B(n25096), .C(matrixInput[1130]), 
        .D(n25081), .Z(n26126) );
    VMW_AO22 U2552 ( .A(cOutput[16]), .B(n25087), .C(cOutput[0]), .D(n25084), 
        .Z(n25174) );
    VMW_FD \matrixInput_reg[1147]  ( .D(n26109), .CP(Clk), .Q(matrixInput
        [1147]) );
    VMW_FD \matrixInput_reg[750]  ( .D(n26506), .CP(Clk), .Q(matrixInput[750])
         );
    VMW_FD \matrixInput_reg[749]  ( .D(n26507), .CP(Clk), .Q(matrixInput[749])
         );
    VMW_AO22 U1064 ( .A(matrixInput[447]), .B(n25096), .C(matrixInput[439]), 
        .D(n25081), .Z(n26817) );
    VMW_AO22 U1652 ( .A(matrixInput[1761]), .B(n25096), .C(matrixInput[1753]), 
        .D(n25081), .Z(n25503) );
    VMW_AO22 U1675 ( .A(matrixInput[1740]), .B(n25096), .C(matrixInput[1732]), 
        .D(n25081), .Z(n25524) );
    VMW_AO22 U2073 ( .A(matrixInput[1382]), .B(n25096), .C(matrixInput[1374]), 
        .D(n25081), .Z(n25882) );
    VMW_FD \matrixInput_reg[1277]  ( .D(n25979), .CP(Clk), .Q(matrixInput
        [1277]) );
    VMW_FD \matrixInput_reg[479]  ( .D(n26777), .CP(Clk), .Q(matrixInput[479])
         );
    VMW_FD \matrixInput_reg[460]  ( .D(n26796), .CP(Clk), .Q(matrixInput[460])
         );
    VMW_FD \matrixInput_reg[1174]  ( .D(n26082), .CP(Clk), .Q(matrixInput
        [1174]) );
    VMW_FD \matrixInput_reg[763]  ( .D(n26493), .CP(Clk), .Q(matrixInput[763])
         );
    VMW_FD \matrixInput_reg[1453]  ( .D(n25803), .CP(Clk), .Q(matrixInput
        [1453]) );
    VMW_FD \matrixInput_reg[244]  ( .D(n27012), .CP(Clk), .Q(matrixInput[244])
         );
    VMW_AO22 U1354 ( .A(matrixInput[2028]), .B(n25096), .C(matrixInput[2020]), 
        .D(n25081), .Z(n25236) );
    VMW_AO22 U1545 ( .A(matrixInput[192]), .B(n25096), .C(matrixInput[184]), 
        .D(n25081), .Z(n27072) );
    VMW_AO22 U1937 ( .A(matrixInput[1505]), .B(n25096), .C(matrixInput[1497]), 
        .D(n25081), .Z(n25759) );
    VMW_AO22 U2054 ( .A(matrixInput[1399]), .B(n25096), .C(matrixInput[1391]), 
        .D(n25081), .Z(n25865) );
    VMW_FD \matrixInput_reg[1750]  ( .D(n25506), .CP(Clk), .Q(matrixInput
        [1750]) );
    VMW_FD \matrixInput_reg[1749]  ( .D(n25507), .CP(Clk), .Q(matrixInput
        [1749]) );
    VMW_FD \matrixInput_reg[147]  ( .D(n27109), .CP(Clk), .Q(matrixInput[147])
         );
    VMW_FD \matrixInput_reg[1479]  ( .D(n25777), .CP(Clk), .Q(matrixInput
        [1479]) );
    VMW_FD \matrixInput_reg[277]  ( .D(n26979), .CP(Clk), .Q(matrixInput[277])
         );
    VMW_AO22 U2258 ( .A(matrixInput[1215]), .B(n25096), .C(matrixInput[1207]), 
        .D(n25081), .Z(n26049) );
    VMW_AO22 U2364 ( .A(matrixInput[1119]), .B(n25096), .C(matrixInput[1111]), 
        .D(n25081), .Z(n26145) );
    VMW_FD \matrixInput_reg[1763]  ( .D(n25493), .CP(Clk), .Q(matrixInput
        [1763]) );
    VMW_FD \matrixInput_reg[1460]  ( .D(n25796), .CP(Clk), .Q(matrixInput
        [1460]) );
    VMW_FD \matrixInput_reg[174]  ( .D(n27082), .CP(Clk), .Q(matrixInput[174])
         );
    VMW_OAI21 U2575 ( .A(n25130), .B(n25131), .C(n25090), .Z(n25139) );
    VMW_AO22 U706 ( .A(matrixInput[769]), .B(n25096), .C(matrixInput[761]), 
        .D(n25081), .Z(n26495) );
    VMW_AO22 U2449 ( .A(matrixInput[1043]), .B(n25096), .C(matrixInput[1035]), 
        .D(n25081), .Z(n26221) );
    VMW_FD \matrixInput_reg[984]  ( .D(n26272), .CP(Clk), .Q(matrixInput[984])
         );
    VMW_AO22 U1268 ( .A(matrixInput[263]), .B(n25096), .C(matrixInput[255]), 
        .D(n25081), .Z(n27001) );
    VMW_AO22 U1479 ( .A(matrixInput[1917]), .B(n25096), .C(matrixInput[1909]), 
        .D(n25081), .Z(n25347) );
    VMW_AO22 U2168 ( .A(matrixInput[1297]), .B(n25096), .C(matrixInput[1289]), 
        .D(n25081), .Z(n25967) );
    VMW_FD \matrixInput_reg[1814]  ( .D(n25442), .CP(Clk), .Q(matrixInput
        [1814]) );
    VMW_AO22 U844 ( .A(matrixInput[645]), .B(n25096), .C(matrixInput[637]), 
        .D(n25081), .Z(n26619) );
    VMW_AO22 U1158 ( .A(matrixInput[362]), .B(n25096), .C(matrixInput[354]), 
        .D(n25081), .Z(n26902) );
    VMW_AO22 U1749 ( .A(matrixInput[1674]), .B(n25096), .C(matrixInput[1666]), 
        .D(n25081), .Z(n25590) );
    VMW_FD \matrixInput_reg[1827]  ( .D(n25429), .CP(Clk), .Q(matrixInput
        [1827]) );
    VMW_AO22 U581 ( .A(matrixInput[882]), .B(n25096), .C(matrixInput[874]), 
        .D(n25081), .Z(n26382) );
    VMW_AO22 U632 ( .A(matrixInput[836]), .B(n25096), .C(matrixInput[828]), 
        .D(n25081), .Z(n26428) );
    VMW_AO22 U721 ( .A(matrixInput[756]), .B(n25096), .C(matrixInput[748]), 
        .D(n25081), .Z(n26508) );
    VMW_AO22 U863 ( .A(matrixInput[69]), .B(n25096), .C(matrixInput[61]), .D(
        n25081), .Z(n27195) );
    VMW_FD \matrixInput_reg[1984]  ( .D(n25272), .CP(Clk), .Q(matrixInput
        [1984]) );
    VMW_FD \matrixInput_reg[54]  ( .D(n27202), .CP(Clk), .Q(matrixInput[54])
         );
    VMW_FD \matrixInput_reg[814]  ( .D(n26442), .CP(Clk), .Q(matrixInput[814])
         );
    VMW_FD \matrixInput_reg[67]  ( .D(n27189), .CP(Clk), .Q(matrixInput[67])
         );
    VMW_FD \matrixInput_reg[1919]  ( .D(n25337), .CP(Clk), .Q(matrixInput
        [1919]) );
    VMW_FD \matrixInput_reg[890]  ( .D(n26366), .CP(Clk), .Q(matrixInput[890])
         );
    VMW_FD \matrixInput_reg[889]  ( .D(n26367), .CP(Clk), .Q(matrixInput[889])
         );
    VMW_FD \matrixInput_reg[827]  ( .D(n26429), .CP(Clk), .Q(matrixInput[827])
         );
    VMW_FD \matrixInput_reg[1900]  ( .D(n25356), .CP(Clk), .Q(matrixInput
        [1900]) );
    VMW_AO22 U970 ( .A(matrixInput[531]), .B(n25096), .C(matrixInput[523]), 
        .D(n25081), .Z(n26733) );
    VMW_AO22 U492 ( .A(matrixInput[962]), .B(n25096), .C(matrixInput[954]), 
        .D(n25081), .Z(n26302) );
    VMW_OAI211 U298 ( .A(n25055), .B(n25068), .C(n25069), .D(n25070), .Z(
        n27388) );
    VMW_AND2 U308 ( .A(n25086), .B(Addr[0]), .Z(n25089) );
    VMW_AO22 U334 ( .A(vectorInput[88]), .B(n25095), .C(vectorInput[80]), .D(
        n25080), .Z(n27304) );
    VMW_AO22 U502 ( .A(matrixInput[953]), .B(n25096), .C(matrixInput[945]), 
        .D(n25081), .Z(n26311) );
    VMW_AO22 U525 ( .A(matrixInput[932]), .B(n25096), .C(matrixInput[924]), 
        .D(n25081), .Z(n26332) );
    VMW_AO22 U957 ( .A(matrixInput[543]), .B(n25096), .C(matrixInput[535]), 
        .D(n25081), .Z(n26721) );
    VMW_FD \matrixInput_reg[1933]  ( .D(n25323), .CP(Clk), .Q(matrixInput
        [1933]) );
    VMW_FD \matrixInput_reg[9]  ( .D(n27247), .CP(Clk), .Q(matrixInput[9]) );
    VMW_FD \matrixInput_reg[1890]  ( .D(n25366), .CP(Clk), .Q(matrixInput
        [1890]) );
    VMW_FD \matrixInput_reg[1889]  ( .D(n25367), .CP(Clk), .Q(matrixInput
        [1889]) );
    VMW_FD \vectorInput_reg[79]  ( .D(n27305), .CP(Clk), .Q(vectorInput[79])
         );
    VMW_FD \vectorInput_reg[60]  ( .D(n27324), .CP(Clk), .Q(vectorInput[60])
         );
    VMW_FD \matrixInput_reg[919]  ( .D(n26337), .CP(Clk), .Q(matrixInput[919])
         );
    VMW_FD \matrixInput_reg[900]  ( .D(n26356), .CP(Clk), .Q(matrixInput[900])
         );
    VMW_AO22 U341 ( .A(vectorInput[82]), .B(n25095), .C(vectorInput[74]), .D(
        n25080), .Z(n27310) );
    VMW_AO22 U366 ( .A(vectorInput[59]), .B(n25095), .C(vectorInput[51]), .D(
        n25080), .Z(n27333) );
    VMW_AO22 U398 ( .A(vectorInput[30]), .B(n25095), .C(vectorInput[22]), .D(
        n25080), .Z(n27362) );
    VMW_AO22 U615 ( .A(matrixInput[851]), .B(n25096), .C(matrixInput[843]), 
        .D(n25081), .Z(n26413) );
    VMW_AO22 U1888 ( .A(matrixInput[1548]), .B(n25096), .C(matrixInput[1540]), 
        .D(n25081), .Z(n25716) );
    VMW_AO22 U1918 ( .A(matrixInput[1521]), .B(n25096), .C(matrixInput[1513]), 
        .D(n25081), .Z(n25743) );
    VMW_FD \vectorInput_reg[53]  ( .D(n27331), .CP(Clk), .Q(vectorInput[53])
         );
    VMW_AO22 U729 ( .A(matrixInput[748]), .B(n25096), .C(matrixInput[740]), 
        .D(n25081), .Z(n26516) );
    VMW_AO22 U785 ( .A(matrixInput[698]), .B(n25096), .C(matrixInput[690]), 
        .D(n25081), .Z(n26566) );
    VMW_FD \matrixInput_reg[1350]  ( .D(n25906), .CP(Clk), .Q(matrixInput
        [1350]) );
    VMW_FD \matrixInput_reg[1349]  ( .D(n25907), .CP(Clk), .Q(matrixInput
        [1349]) );
    VMW_FD \matrixInput_reg[933]  ( .D(n26323), .CP(Clk), .Q(matrixInput[933])
         );
    VMW_AO22 U1247 ( .A(matrixInput[282]), .B(n25096), .C(matrixInput[274]), 
        .D(n25081), .Z(n26982) );
    VMW_AO22 U2277 ( .A(matrixInput[1198]), .B(n25096), .C(matrixInput[1190]), 
        .D(n25081), .Z(n26066) );
    VMW_AO22 U2466 ( .A(matrixInput[109]), .B(n25096), .C(matrixInput[101]), 
        .D(n25081), .Z(n27155) );
    VMW_FD \matrixInput_reg[547]  ( .D(n26709), .CP(Clk), .Q(matrixInput[547])
         );
    VMW_FD \matrixInput_reg[1053]  ( .D(n26203), .CP(Clk), .Q(matrixInput
        [1053]) );
    VMW_FD \matrixInput_reg[644]  ( .D(n26612), .CP(Clk), .Q(matrixInput[644])
         );
    VMW_AO22 U1456 ( .A(matrixInput[200]), .B(n25096), .C(matrixInput[192]), 
        .D(n25081), .Z(n27064) );
    VMW_AO22 U1824 ( .A(matrixInput[1607]), .B(n25096), .C(matrixInput[1599]), 
        .D(n25081), .Z(n25657) );
    VMW_AO22 U419 ( .A(vectorInput[127]), .B(n25095), .C(vectorInput[119]), 
        .D(n25080), .Z(n27265) );
    VMW_AO22 U450 ( .A(matrixInput[1000]), .B(n25096), .C(matrixInput[992]), 
        .D(n25081), .Z(n26264) );
    VMW_AO22 U589 ( .A(matrixInput[875]), .B(n25096), .C(matrixInput[867]), 
        .D(n25081), .Z(n26389) );
    VMW_AO22 U2147 ( .A(matrixInput[1315]), .B(n25096), .C(matrixInput[1307]), 
        .D(n25081), .Z(n25949) );
    VMW_AO22 U822 ( .A(matrixInput[665]), .B(n25096), .C(matrixInput[657]), 
        .D(n25081), .Z(n26599) );
    VMW_AO22 U1150 ( .A(matrixInput[369]), .B(n25096), .C(matrixInput[361]), 
        .D(n25081), .Z(n26895) );
    VMW_AO22 U1177 ( .A(matrixInput[345]), .B(n25096), .C(matrixInput[337]), 
        .D(n25081), .Z(n26919) );
    VMW_FD \matrixInput_reg[1363]  ( .D(n25893), .CP(Clk), .Q(matrixInput
        [1363]) );
    VMW_FD \matrixInput_reg[574]  ( .D(n26682), .CP(Clk), .Q(matrixInput[574])
         );
    VMW_AO22 U1741 ( .A(matrixInput[1681]), .B(n25096), .C(matrixInput[1673]), 
        .D(n25081), .Z(n25583) );
    VMW_AO22 U1766 ( .A(matrixInput[1658]), .B(n25096), .C(matrixInput[1650]), 
        .D(n25081), .Z(n25606) );
    VMW_FD \matrixInput_reg[677]  ( .D(n26579), .CP(Clk), .Q(matrixInput[677])
         );
    VMW_AO22 U2160 ( .A(matrixInput[1304]), .B(n25096), .C(matrixInput[1296]), 
        .D(n25081), .Z(n25960) );
    VMW_FD \matrixInput_reg[2023]  ( .D(n25233), .CP(Clk), .Q(matrixInput
        [2023]) );
    VMW_FD \matrixInput_reg[1079]  ( .D(n26177), .CP(Clk), .Q(matrixInput
        [1079]) );
    VMW_FD \matrixInput_reg[1060]  ( .D(n26196), .CP(Clk), .Q(matrixInput
        [1060]) );
    VMW_FD \matrixInput_reg[1644]  ( .D(n25612), .CP(Clk), .Q(matrixInput
        [1644]) );
    VMW_FD \matrixInput_reg[1547]  ( .D(n25709), .CP(Clk), .Q(matrixInput
        [1547]) );
    VMW_FD \matrixInput_reg[350]  ( .D(n26906), .CP(Clk), .Q(matrixInput[350])
         );
    VMW_FD \matrixInput_reg[349]  ( .D(n26907), .CP(Clk), .Q(matrixInput[349])
         );
    VMW_AO22 U1260 ( .A(matrixInput[270]), .B(n25096), .C(matrixInput[262]), 
        .D(n25081), .Z(n26994) );
    VMW_AO22 U1471 ( .A(matrixInput[1924]), .B(n25096), .C(matrixInput[1916]), 
        .D(n25081), .Z(n25340) );
    VMW_AO22 U2250 ( .A(matrixInput[1222]), .B(n25096), .C(matrixInput[1214]), 
        .D(n25081), .Z(n26042) );
    VMW_FD \matrixInput_reg[1574]  ( .D(n25682), .CP(Clk), .Q(matrixInput
        [1574]) );
    VMW_FD \matrixInput_reg[363]  ( .D(n26893), .CP(Clk), .Q(matrixInput[363])
         );
    VMW_AO22 U2441 ( .A(matrixInput[1050]), .B(n25096), .C(matrixInput[1042]), 
        .D(n25081), .Z(n26214) );
    VMW_FD \matrixInput_reg[2010]  ( .D(n25246), .CP(Clk), .Q(matrixInput
        [2010]) );
    VMW_FD \matrixInput_reg[2009]  ( .D(n25247), .CP(Clk), .Q(matrixInput
        [2009]) );
    VMW_AO22 U1803 ( .A(matrixInput[1625]), .B(n25096), .C(matrixInput[1617]), 
        .D(n25081), .Z(n25639) );
    VMW_AO22 U1993 ( .A(matrixInput[1454]), .B(n25096), .C(matrixInput[1446]), 
        .D(n25081), .Z(n25810) );
    VMW_FD \matrixInput_reg[1677]  ( .D(n25579), .CP(Clk), .Q(matrixInput
        [1677]) );
    VMW_FD \matrixInput_reg[31]  ( .D(n27225), .CP(Clk), .Q(matrixInput[31])
         );
    VMW_FD \matrixInput_reg[28]  ( .D(n27228), .CP(Clk), .Q(matrixInput[28])
         );
    VMW_AO22 U477 ( .A(matrixInput[976]), .B(n25096), .C(matrixInput[968]), 
        .D(n25081), .Z(n26288) );
    VMW_AO22 U747 ( .A(matrixInput[732]), .B(n25096), .C(matrixInput[724]), 
        .D(n25081), .Z(n26532) );
    VMW_AO22 U760 ( .A(matrixInput[720]), .B(n25096), .C(matrixInput[712]), 
        .D(n25081), .Z(n26544) );
    VMW_FD \matrixInput_reg[871]  ( .D(n26385), .CP(Clk), .Q(matrixInput[871])
         );
    VMW_FD \matrixInput_reg[868]  ( .D(n26388), .CP(Clk), .Q(matrixInput[868])
         );
    VMW_AO22 U2219 ( .A(matrixInput[1250]), .B(n25096), .C(matrixInput[1242]), 
        .D(n25081), .Z(n26014) );
    VMW_INV U2598 ( .A(Addr[3]), .Z(n25092) );
    VMW_FD \matrixInput_reg[842]  ( .D(n26414), .CP(Clk), .Q(matrixInput[842])
         );
    VMW_AO22 U805 ( .A(matrixInput[680]), .B(n25096), .C(matrixInput[672]), 
        .D(n25081), .Z(n26584) );
    VMW_AO22 U995 ( .A(matrixInput[508]), .B(n25096), .C(matrixInput[500]), 
        .D(n25081), .Z(n26756) );
    VMW_AO22 U1229 ( .A(matrixInput[298]), .B(n25096), .C(matrixInput[290]), 
        .D(n25081), .Z(n26966) );
    VMW_AO22 U1438 ( .A(matrixInput[1954]), .B(n25096), .C(matrixInput[1946]), 
        .D(n25081), .Z(n25310) );
    VMW_AO22 U2389 ( .A(matrixInput[116]), .B(n25096), .C(matrixInput[108]), 
        .D(n25081), .Z(n27148) );
    VMW_AO22 U2408 ( .A(matrixInput[1080]), .B(n25096), .C(matrixInput[1072]), 
        .D(n25081), .Z(n26184) );
    VMW_FD \matrixInput_reg[1871]  ( .D(n25385), .CP(Clk), .Q(matrixInput
        [1871]) );
    VMW_FD \matrixInput_reg[1868]  ( .D(n25388), .CP(Clk), .Q(matrixInput
        [1868]) );
    VMW_FD \vectorInput_reg[98]  ( .D(n27286), .CP(Clk), .Q(vectorInput[98])
         );
    VMW_FD \vectorInput_reg[81]  ( .D(n27303), .CP(Clk), .Q(vectorInput[81])
         );
    VMW_AO22 U2129 ( .A(matrixInput[1331]), .B(n25096), .C(matrixInput[1323]), 
        .D(n25081), .Z(n25933) );
    VMW_FD \vectorInput_reg[102]  ( .D(n27282), .CP(Clk), .Q(vectorInput[102])
         );
    VMW_AO22 U577 ( .A(matrixInput[886]), .B(n25096), .C(matrixInput[878]), 
        .D(n25081), .Z(n26378) );
    VMW_AO22 U895 ( .A(matrixInput[599]), .B(n25096), .C(matrixInput[591]), 
        .D(n25081), .Z(n26665) );
    VMW_AO22 U905 ( .A(matrixInput[590]), .B(n25096), .C(matrixInput[582]), 
        .D(n25081), .Z(n26674) );
    VMW_AO22 U939 ( .A(matrixInput[559]), .B(n25096), .C(matrixInput[551]), 
        .D(n25081), .Z(n26705) );
    VMW_AO22 U1025 ( .A(matrixInput[482]), .B(n25096), .C(matrixInput[474]), 
        .D(n25081), .Z(n26782) );
    VMW_AO22 U1089 ( .A(matrixInput[424]), .B(n25096), .C(matrixInput[416]), 
        .D(n25081), .Z(n26840) );
    VMW_AO22 U1119 ( .A(matrixInput[46]), .B(n25096), .C(matrixInput[38]), .D(
        n25081), .Z(n27218) );
    VMW_AO22 U1708 ( .A(matrixInput[1710]), .B(n25096), .C(matrixInput[1702]), 
        .D(n25081), .Z(n25554) );
    VMW_AO22 U1634 ( .A(matrixInput[184]), .B(n25096), .C(matrixInput[176]), 
        .D(n25081), .Z(n27080) );
    VMW_AO22 U1698 ( .A(matrixInput[1719]), .B(n25096), .C(matrixInput[1711]), 
        .D(n25081), .Z(n25545) );
    VMW_FD \matrixInput_reg[1842]  ( .D(n25414), .CP(Clk), .Q(matrixInput
        [1842]) );
    VMW_FD \matrixInput_reg[1436]  ( .D(n25820), .CP(Clk), .Q(matrixInput
        [1436]) );
    VMW_FD \matrixInput_reg[238]  ( .D(n27018), .CP(Clk), .Q(matrixInput[238])
         );
    VMW_FD \matrixInput_reg[221]  ( .D(n27035), .CP(Clk), .Q(matrixInput[221])
         );
    VMW_AO22 U2015 ( .A(matrixInput[1434]), .B(n25096), .C(matrixInput[1426]), 
        .D(n25081), .Z(n25830) );
    VMW_FD \matrixInput_reg[122]  ( .D(n27134), .CP(Clk), .Q(matrixInput[122])
         );
    VMW_AO22 U2185 ( .A(matrixInput[1281]), .B(n25096), .C(matrixInput[1273]), 
        .D(n25081), .Z(n25983) );
    VMW_INV U2604 ( .A(\holder[2] ), .Z(n25062) );
    VMW_FD \matrixInput_reg[1735]  ( .D(n25521), .CP(Clk), .Q(matrixInput
        [1735]) );
    VMW_AO22 U1002 ( .A(matrixInput[503]), .B(n25096), .C(matrixInput[495]), 
        .D(n25081), .Z(n26761) );
    VMW_AO22 U1285 ( .A(matrixInput[31]), .B(n25096), .C(matrixInput[23]), .D(
        n25081), .Z(n27233) );
    VMW_AO22 U1504 ( .A(matrixInput[1895]), .B(n25096), .C(matrixInput[1887]), 
        .D(n25081), .Z(n25369) );
    VMW_FD \matrixInput_reg[1405]  ( .D(n25851), .CP(Clk), .Q(matrixInput
        [1405]) );
    VMW_AO22 U1315 ( .A(matrixInput[220]), .B(n25096), .C(matrixInput[212]), 
        .D(n25081), .Z(n27044) );
    VMW_AO22 U1494 ( .A(matrixInput[1904]), .B(n25096), .C(matrixInput[1896]), 
        .D(n25081), .Z(n25360) );
    VMW_AO22 U1332 ( .A(DataIn[0]), .B(n25096), .C(matrixInput[2040]), .D(
        n25081), .Z(n25216) );
    VMW_AO22 U1976 ( .A(matrixInput[1469]), .B(n25096), .C(matrixInput[1461]), 
        .D(n25081), .Z(n25795) );
    VMW_FD \matrixInput_reg[212]  ( .D(n27044), .CP(Clk), .Q(matrixInput[212])
         );
    VMW_AO22 U2325 ( .A(matrixInput[1155]), .B(n25096), .C(matrixInput[1147]), 
        .D(n25081), .Z(n26109) );
    VMW_FD \matrixInput_reg[1382]  ( .D(n25874), .CP(Clk), .Q(matrixInput
        [1382]) );
    VMW_FD \matrixInput_reg[1098]  ( .D(n26158), .CP(Clk), .Q(matrixInput
        [1098]) );
    VMW_FD \matrixInput_reg[696]  ( .D(n26560), .CP(Clk), .Q(matrixInput[696])
         );
    VMW_FD \matrixInput_reg[1081]  ( .D(n26175), .CP(Clk), .Q(matrixInput
        [1081]) );
    VMW_FD \matrixInput_reg[595]  ( .D(n26661), .CP(Clk), .Q(matrixInput[595])
         );
    VMW_AO22 U2534 ( .A(cOutput[18]), .B(n25087), .C(cOutput[2]), .D(n25084), 
        .Z(n25152) );
    VMW_FD \matrixInput_reg[1706]  ( .D(n25550), .CP(Clk), .Q(matrixInput
        [1706]) );
    VMW_FD \matrixInput_reg[111]  ( .D(n27145), .CP(Clk), .Q(matrixInput[111])
         );
    VMW_FD \matrixInput_reg[108]  ( .D(n27148), .CP(Clk), .Q(matrixInput[108])
         );
    VMW_AO22 U1523 ( .A(matrixInput[194]), .B(n25096), .C(matrixInput[186]), 
        .D(n25081), .Z(n27070) );
    VMW_AO22 U1951 ( .A(matrixInput[1492]), .B(n25096), .C(matrixInput[1484]), 
        .D(n25081), .Z(n25772) );
    VMW_FD \matrixInput_reg[1221]  ( .D(n26035), .CP(Clk), .Q(matrixInput
        [1221]) );
    VMW_FD \matrixInput_reg[436]  ( .D(n26820), .CP(Clk), .Q(matrixInput[436])
         );
    VMW_AO22 U2292 ( .A(matrixInput[1185]), .B(n25096), .C(matrixInput[1177]), 
        .D(n25081), .Z(n26079) );
    VMW_AO22 U2513 ( .A(cOutput[117]), .B(n25087), .C(cOutput[101]), .D(n25084
        ), .Z(n25125) );
    VMW_FD \matrixInput_reg[1238]  ( .D(n26018), .CP(Clk), .Q(matrixInput
        [1238]) );
    VMW_FD \matrixInput_reg[1122]  ( .D(n26134), .CP(Clk), .Q(matrixInput
        [1122]) );
    VMW_FD \matrixInput_reg[735]  ( .D(n26521), .CP(Clk), .Q(matrixInput[735])
         );
    VMW_AO22 U2302 ( .A(matrixInput[1176]), .B(n25096), .C(matrixInput[1168]), 
        .D(n25081), .Z(n26088) );
    VMW_AO22 U2483 ( .A(matrixInput[1012]), .B(n25096), .C(matrixInput[1004]), 
        .D(n25081), .Z(n26252) );
    VMW_FD \matrixInput_reg[1212]  ( .D(n26044), .CP(Clk), .Q(matrixInput
        [1212]) );
    VMW_FD \matrixInput_reg[405]  ( .D(n26851), .CP(Clk), .Q(matrixInput[405])
         );
    VMW_AO22 U1192 ( .A(matrixInput[331]), .B(n25096), .C(matrixInput[323]), 
        .D(n25081), .Z(n26933) );
    VMW_AO22 U1783 ( .A(matrixInput[1643]), .B(n25096), .C(matrixInput[1635]), 
        .D(n25081), .Z(n25621) );
    VMW_AO22 U1613 ( .A(matrixInput[1797]), .B(n25096), .C(matrixInput[1789]), 
        .D(n25081), .Z(n25467) );
    VMW_AO22 U2032 ( .A(matrixInput[1418]), .B(n25096), .C(matrixInput[1410]), 
        .D(n25081), .Z(n25846) );
    VMW_BUFIZ U2623 ( .A(\holder[2] ), .E(RD), .Z(\DataOut[2]1 ) );
    VMW_FD \matrixInput_reg[1696]  ( .D(n25560), .CP(Clk), .Q(matrixInput
        [1696]) );
    VMW_FD \matrixInput_reg[382]  ( .D(n26874), .CP(Clk), .Q(matrixInput[382])
         );
    VMW_FD \matrixInput_reg[1595]  ( .D(n25661), .CP(Clk), .Q(matrixInput
        [1595]) );
    VMW_FD \matrixInput_reg[1111]  ( .D(n26145), .CP(Clk), .Q(matrixInput
        [1111]) );
    VMW_FD \matrixInput_reg[1108]  ( .D(n26148), .CP(Clk), .Q(matrixInput
        [1108]) );
    VMW_FD \matrixInput_reg[706]  ( .D(n26550), .CP(Clk), .Q(matrixInput[706])
         );
    VMW_BUFIZ U2638 ( .A(\holder[1] ), .E(RD), .Z(\DataOut[1]1 ) );
    VMW_AO22 U647 ( .A(matrixInput[822]), .B(n25096), .C(matrixInput[814]), 
        .D(n25081), .Z(n26442) );
    VMW_AO22 U1019 ( .A(matrixInput[55]), .B(n25096), .C(matrixInput[47]), .D(
        n25081), .Z(n27209) );
    VMW_AO22 U2029 ( .A(matrixInput[1421]), .B(n25096), .C(matrixInput[1413]), 
        .D(n25081), .Z(n25843) );
    VMW_FD \vectorInput_reg[112]  ( .D(n27272), .CP(Clk), .Q(vectorInput[112])
         );
    VMW_AO22 U1189 ( .A(matrixInput[334]), .B(n25096), .C(matrixInput[326]), 
        .D(n25081), .Z(n26930) );
    VMW_AO22 U1798 ( .A(matrixInput[1629]), .B(n25096), .C(matrixInput[1621]), 
        .D(n25081), .Z(n25635) );
    VMW_AO22 U1608 ( .A(matrixInput[1801]), .B(n25096), .C(matrixInput[1793]), 
        .D(n25081), .Z(n25463) );
    VMW_FD \matrixInput_reg[1852]  ( .D(n25404), .CP(Clk), .Q(matrixInput
        [1852]) );
    VMW_AO22 U660 ( .A(matrixInput[810]), .B(n25096), .C(matrixInput[802]), 
        .D(n25081), .Z(n26454) );
    VMW_AO22 U1329 ( .A(DataIn[3]), .B(n25096), .C(matrixInput[2043]), .D(
        n25081), .Z(n25213) );
    VMW_AO22 U2289 ( .A(matrixInput[125]), .B(n25096), .C(matrixInput[117]), 
        .D(n25081), .Z(n27139) );
    VMW_AO22 U2508 ( .A(cOutput[29]), .B(n25089), .C(cOutput[13]), .D(n25088), 
        .Z(n25120) );
    VMW_AO22 U2319 ( .A(matrixInput[1160]), .B(n25096), .C(matrixInput[1152]), 
        .D(n25081), .Z(n26104) );
    VMW_AO22 U2498 ( .A(cOutput[22]), .B(n25087), .C(cOutput[6]), .D(n25084), 
        .Z(n25108) );
    VMW_FD \vectorInput_reg[121]  ( .D(n27263), .CP(Clk), .Q(vectorInput[121])
         );
    VMW_FD \matrixInput_reg[1878]  ( .D(n25378), .CP(Clk), .Q(matrixInput
        [1878]) );
    VMW_FD \matrixInput_reg[1861]  ( .D(n25395), .CP(Clk), .Q(matrixInput
        [1861]) );
    VMW_AO22 U1538 ( .A(matrixInput[1864]), .B(n25096), .C(matrixInput[1856]), 
        .D(n25081), .Z(n25400) );
    VMW_FD \vectorInput_reg[91]  ( .D(n27293), .CP(Clk), .Q(vectorInput[91])
         );
    VMW_FD \vectorInput_reg[88]  ( .D(n27296), .CP(Clk), .Q(vectorInput[88])
         );
    VMW_AO22 U922 ( .A(matrixInput[575]), .B(n25096), .C(matrixInput[567]), 
        .D(n25081), .Z(n26689) );
    VMW_FD \matrixInput_reg[852]  ( .D(n26404), .CP(Clk), .Q(matrixInput[852])
         );
    VMW_FD \matrixInput_reg[12]  ( .D(n27244), .CP(Clk), .Q(matrixInput[12])
         );
    VMW_FD \matrixInput_reg[38]  ( .D(n27218), .CP(Clk), .Q(matrixInput[38])
         );
    VMW_FD \matrixInput_reg[21]  ( .D(n27235), .CP(Clk), .Q(matrixInput[21])
         );
    VMW_AO22 U383 ( .A(vectorInput[44]), .B(n25095), .C(vectorInput[36]), .D(
        n25080), .Z(n27348) );
    VMW_AO22 U425 ( .A(vectorInput[121]), .B(n25095), .C(vectorInput[113]), 
        .D(n25080), .Z(n27271) );
    VMW_AO22 U550 ( .A(matrixInput[909]), .B(n25096), .C(matrixInput[901]), 
        .D(n25081), .Z(n26355) );
    VMW_AO22 U685 ( .A(matrixInput[788]), .B(n25096), .C(matrixInput[780]), 
        .D(n25081), .Z(n26476) );
    VMW_AO22 U839 ( .A(matrixInput[649]), .B(n25096), .C(matrixInput[641]), 
        .D(n25081), .Z(n26615) );
    VMW_AO22 U1092 ( .A(matrixInput[421]), .B(n25096), .C(matrixInput[413]), 
        .D(n25081), .Z(n26843) );
    VMW_FD \matrixInput_reg[1686]  ( .D(n25570), .CP(Clk), .Q(matrixInput
        [1686]) );
    VMW_FD \matrixInput_reg[1202]  ( .D(n26054), .CP(Clk), .Q(matrixInput
        [1202]) );
    VMW_FD \matrixInput_reg[878]  ( .D(n26378), .CP(Clk), .Q(matrixInput[878])
         );
    VMW_FD \matrixInput_reg[861]  ( .D(n26395), .CP(Clk), .Q(matrixInput[861])
         );
    VMW_FD \matrixInput_reg[415]  ( .D(n26841), .CP(Clk), .Q(matrixInput[415])
         );
    VMW_AO22 U1102 ( .A(matrixInput[412]), .B(n25096), .C(matrixInput[404]), 
        .D(n25081), .Z(n26852) );
    VMW_AO22 U1713 ( .A(matrixInput[1707]), .B(n25096), .C(matrixInput[1699]), 
        .D(n25081), .Z(n25557) );
    VMW_AO22 U1125 ( .A(matrixInput[392]), .B(n25096), .C(matrixInput[384]), 
        .D(n25081), .Z(n26872) );
    VMW_AO22 U1215 ( .A(matrixInput[310]), .B(n25096), .C(matrixInput[302]), 
        .D(n25081), .Z(n26954) );
    VMW_AO22 U1232 ( .A(matrixInput[296]), .B(n25096), .C(matrixInput[288]), 
        .D(n25081), .Z(n26968) );
    VMW_AO22 U1423 ( .A(matrixInput[203]), .B(n25096), .C(matrixInput[195]), 
        .D(n25081), .Z(n27061) );
    VMW_AO22 U1683 ( .A(matrixInput[1733]), .B(n25096), .C(matrixInput[1725]), 
        .D(n25081), .Z(n25531) );
    VMW_AO22 U2132 ( .A(matrixInput[1328]), .B(n25096), .C(matrixInput[1320]), 
        .D(n25081), .Z(n25936) );
    VMW_FD \matrixInput_reg[1585]  ( .D(n25671), .CP(Clk), .Q(matrixInput
        [1585]) );
    VMW_FD \matrixInput_reg[1118]  ( .D(n26138), .CP(Clk), .Q(matrixInput
        [1118]) );
    VMW_FD \matrixInput_reg[1101]  ( .D(n26155), .CP(Clk), .Q(matrixInput
        [1101]) );
    VMW_FD \matrixInput_reg[716]  ( .D(n26540), .CP(Clk), .Q(matrixInput[716])
         );
    VMW_FD \matrixInput_reg[392]  ( .D(n26864), .CP(Clk), .Q(matrixInput[392])
         );
    VMW_AO22 U1594 ( .A(matrixInput[1813]), .B(n25096), .C(matrixInput[1805]), 
        .D(n25081), .Z(n25451) );
    VMW_AO22 U1851 ( .A(matrixInput[1582]), .B(n25096), .C(matrixInput[1574]), 
        .D(n25081), .Z(n25682) );
    VMW_AO22 U2202 ( .A(matrixInput[1266]), .B(n25096), .C(matrixInput[1258]), 
        .D(n25081), .Z(n25998) );
    VMW_OAI21 U2583 ( .A(n25152), .B(n25153), .C(n25090), .Z(n25161) );
    VMW_FD \matrixInput_reg[1231]  ( .D(n26025), .CP(Clk), .Q(matrixInput
        [1231]) );
    VMW_FD \matrixInput_reg[1228]  ( .D(n26028), .CP(Clk), .Q(matrixInput
        [1228]) );
    VMW_FD \matrixInput_reg[1132]  ( .D(n26124), .CP(Clk), .Q(matrixInput
        [1132]) );
    VMW_FD \matrixInput_reg[426]  ( .D(n26830), .CP(Clk), .Q(matrixInput[426])
         );
    VMW_FD \matrixInput_reg[725]  ( .D(n26531), .CP(Clk), .Q(matrixInput[725])
         );
    VMW_FD \vectorInput_reg[6]  ( .D(n27378), .CP(Clk), .Q(vectorInput[6]) );
    VMW_AO22 U2392 ( .A(matrixInput[1095]), .B(n25096), .C(matrixInput[1087]), 
        .D(n25081), .Z(n26169) );
    VMW_AO22 U2413 ( .A(matrixInput[1076]), .B(n25096), .C(matrixInput[1068]), 
        .D(n25081), .Z(n26188) );
    VMW_FD \matrixInput_reg[202]  ( .D(n27054), .CP(Clk), .Q(matrixInput[202])
         );
    VMW_AO22 U1385 ( .A(matrixInput[2002]), .B(n25096), .C(matrixInput[1994]), 
        .D(n25081), .Z(n25262) );
    VMW_AO22 U1404 ( .A(matrixInput[1985]), .B(n25096), .C(matrixInput[1977]), 
        .D(n25081), .Z(n25279) );
    VMW_FD \matrixInput_reg[1415]  ( .D(n25841), .CP(Clk), .Q(matrixInput
        [1415]) );
    VMW_AO22 U1876 ( .A(matrixInput[1559]), .B(n25096), .C(matrixInput[1551]), 
        .D(n25081), .Z(n25705) );
    VMW_FD \matrixInput_reg[1091]  ( .D(n26165), .CP(Clk), .Q(matrixInput
        [1091]) );
    VMW_FD \matrixInput_reg[1088]  ( .D(n26168), .CP(Clk), .Q(matrixInput
        [1088]) );
    VMW_FD \matrixInput_reg[686]  ( .D(n26570), .CP(Clk), .Q(matrixInput[686])
         );
    VMW_AO22 U2225 ( .A(matrixInput[1245]), .B(n25096), .C(matrixInput[1237]), 
        .D(n25081), .Z(n26019) );
    VMW_AO22 U2434 ( .A(matrixInput[1057]), .B(n25096), .C(matrixInput[1049]), 
        .D(n25081), .Z(n26207) );
    VMW_FD \matrixInput_reg[1392]  ( .D(n25864), .CP(Clk), .Q(matrixInput
        [1392]) );
    VMW_FD \matrixInput_reg[585]  ( .D(n26671), .CP(Clk), .Q(matrixInput[585])
         );
    VMW_FD \matrixInput_reg[118]  ( .D(n27138), .CP(Clk), .Q(matrixInput[118])
         );
    VMW_FD \matrixInput_reg[101]  ( .D(n27155), .CP(Clk), .Q(matrixInput[101])
         );
    VMW_FD \matrixInput_reg[1716]  ( .D(n25540), .CP(Clk), .Q(matrixInput
        [1716]) );
    VMW_AO22 U1734 ( .A(matrixInput[175]), .B(n25096), .C(matrixInput[167]), 
        .D(n25081), .Z(n27089) );
    VMW_FD \matrixInput_reg[1426]  ( .D(n25830), .CP(Clk), .Q(matrixInput
        [1426]) );
    VMW_AO22 U2085 ( .A(matrixInput[1371]), .B(n25096), .C(matrixInput[1363]), 
        .D(n25081), .Z(n25893) );
    VMW_FD \matrixInput_reg[231]  ( .D(n27025), .CP(Clk), .Q(matrixInput[231])
         );
    VMW_FD \matrixInput_reg[228]  ( .D(n27028), .CP(Clk), .Q(matrixInput[228])
         );
    VMW_AO22 U2115 ( .A(matrixInput[1344]), .B(n25096), .C(matrixInput[1336]), 
        .D(n25081), .Z(n25920) );
    VMW_FD \matrixInput_reg[1725]  ( .D(n25531), .CP(Clk), .Q(matrixInput
        [1725]) );
    VMW_FD \matrixInput_reg[132]  ( .D(n27124), .CP(Clk), .Q(matrixInput[132])
         );
    VMW_AO22 U1818 ( .A(matrixInput[1611]), .B(n25096), .C(matrixInput[1603]), 
        .D(n25081), .Z(n25653) );
    VMW_FD \vectorInput_reg[43]  ( .D(n27341), .CP(Clk), .Q(vectorInput[43])
         );
    VMW_AO22 U1988 ( .A(matrixInput[1458]), .B(n25096), .C(matrixInput[1450]), 
        .D(n25081), .Z(n25806) );
    VMW_AO22 U715 ( .A(matrixInput[761]), .B(n25096), .C(matrixInput[753]), 
        .D(n25081), .Z(n26503) );
    VMW_AO22 U857 ( .A(matrixInput[633]), .B(n25096), .C(matrixInput[625]), 
        .D(n25081), .Z(n26631) );
    VMW_FD \matrixInput_reg[1899]  ( .D(n25357), .CP(Clk), .Q(matrixInput
        [1899]) );
    VMW_FD \matrixInput_reg[1880]  ( .D(n25376), .CP(Clk), .Q(matrixInput
        [1880]) );
    VMW_FD \matrixInput_reg[923]  ( .D(n26333), .CP(Clk), .Q(matrixInput[923])
         );
    VMW_FD \matrixInput_reg[910]  ( .D(n26346), .CP(Clk), .Q(matrixInput[910])
         );
    VMW_FD \vectorInput_reg[70]  ( .D(n27314), .CP(Clk), .Q(vectorInput[70])
         );
    VMW_FD \vectorInput_reg[69]  ( .D(n27315), .CP(Clk), .Q(vectorInput[69])
         );
    VMW_FD \matrixInput_reg[909]  ( .D(n26347), .CP(Clk), .Q(matrixInput[909])
         );
    VMW_AO22 U870 ( .A(matrixInput[621]), .B(n25096), .C(matrixInput[613]), 
        .D(n25081), .Z(n26643) );
    VMW_FD \matrixInput_reg[1923]  ( .D(n25333), .CP(Clk), .Q(matrixInput
        [1923]) );
    VMW_FD \matrixInput_reg[0]  ( .D(n27256), .CP(Clk), .Q(matrixInput[0]) );
    VMW_AO22 U402 ( .A(vectorInput[27]), .B(n25095), .C(vectorInput[19]), .D(
        n25080), .Z(n27365) );
    VMW_AO22 U592 ( .A(matrixInput[872]), .B(n25096), .C(matrixInput[864]), 
        .D(n25081), .Z(n26392) );
    VMW_AO22 U732 ( .A(matrixInput[746]), .B(n25096), .C(matrixInput[738]), 
        .D(n25081), .Z(n26518) );
    VMW_FD \matrixInput_reg[899]  ( .D(n26357), .CP(Clk), .Q(matrixInput[899])
         );
    VMW_FD \matrixInput_reg[880]  ( .D(n26376), .CP(Clk), .Q(matrixInput[880])
         );
    VMW_AO22 U1050 ( .A(matrixInput[459]), .B(n25096), .C(matrixInput[451]), 
        .D(n25081), .Z(n26805) );
    VMW_AO22 U1360 ( .A(matrixInput[2023]), .B(n25096), .C(matrixInput[2015]), 
        .D(n25081), .Z(n25241) );
    VMW_AO22 U2350 ( .A(matrixInput[1132]), .B(n25096), .C(matrixInput[1124]), 
        .D(n25081), .Z(n26132) );
    VMW_AO22 U2541 ( .A(cOutput[122]), .B(n25089), .C(cOutput[106]), .D(n25088
        ), .Z(n25159) );
    VMW_FD \matrixInput_reg[2019]  ( .D(n25237), .CP(Clk), .Q(matrixInput
        [2019]) );
    VMW_FD \matrixInput_reg[2000]  ( .D(n25256), .CP(Clk), .Q(matrixInput
        [2000]) );
    VMW_FD \matrixInput_reg[1910]  ( .D(n25346), .CP(Clk), .Q(matrixInput
        [1910]) );
    VMW_FD \matrixInput_reg[1909]  ( .D(n25347), .CP(Clk), .Q(matrixInput
        [1909]) );
    VMW_FD \matrixInput_reg[1564]  ( .D(n25692), .CP(Clk), .Q(matrixInput
        [1564]) );
    VMW_FD \matrixInput_reg[373]  ( .D(n26883), .CP(Clk), .Q(matrixInput[373])
         );
    VMW_AO22 U1571 ( .A(matrixInput[1834]), .B(n25096), .C(matrixInput[1826]), 
        .D(n25081), .Z(n25430) );
    VMW_AO22 U1893 ( .A(matrixInput[1544]), .B(n25096), .C(matrixInput[1536]), 
        .D(n25081), .Z(n25720) );
    VMW_FD \matrixInput_reg[1667]  ( .D(n25589), .CP(Clk), .Q(matrixInput
        [1667]) );
    VMW_AO22 U1903 ( .A(matrixInput[1535]), .B(n25096), .C(matrixInput[1527]), 
        .D(n25081), .Z(n25729) );
    VMW_AO22 U2060 ( .A(matrixInput[1394]), .B(n25096), .C(matrixInput[1386]), 
        .D(n25081), .Z(n25870) );
    VMW_FD \matrixInput_reg[2033]  ( .D(n25223), .CP(Clk), .Q(matrixInput
        [2033]) );
    VMW_FD \matrixInput_reg[1654]  ( .D(n25602), .CP(Clk), .Q(matrixInput
        [1654]) );
    VMW_FD \matrixInput_reg[1557]  ( .D(n25699), .CP(Clk), .Q(matrixInput
        [1557]) );
    VMW_FD \matrixInput_reg[359]  ( .D(n26897), .CP(Clk), .Q(matrixInput[359])
         );
    VMW_FD \matrixInput_reg[340]  ( .D(n26916), .CP(Clk), .Q(matrixInput[340])
         );
    VMW_AO22 U1641 ( .A(matrixInput[1771]), .B(n25096), .C(matrixInput[1763]), 
        .D(n25081), .Z(n25493) );
    VMW_FD \matrixInput_reg[1373]  ( .D(n25883), .CP(Clk), .Q(matrixInput
        [1373]) );
    VMW_AO22 U489 ( .A(matrixInput[965]), .B(n25096), .C(matrixInput[957]), 
        .D(n25081), .Z(n26299) );
    VMW_AO22 U2047 ( .A(matrixInput[1406]), .B(n25096), .C(matrixInput[1398]), 
        .D(n25081), .Z(n25858) );
    VMW_FD \matrixInput_reg[564]  ( .D(n26692), .CP(Clk), .Q(matrixInput[564])
         );
    VMW_AO22 U348 ( .A(vectorInput[76]), .B(n25095), .C(vectorInput[68]), .D(
        n25080), .Z(n27316) );
    VMW_AO22 U353 ( .A(vectorInput[71]), .B(n25095), .C(vectorInput[63]), .D(
        n25080), .Z(n27321) );
    VMW_AO22 U374 ( .A(vectorInput[52]), .B(n25095), .C(vectorInput[44]), .D(
        n25080), .Z(n27340) );
    VMW_AO22 U391 ( .A(vectorInput[37]), .B(n25095), .C(vectorInput[29]), .D(
        n25080), .Z(n27355) );
    VMW_AO22 U437 ( .A(vectorInput[110]), .B(n25095), .C(vectorInput[102]), 
        .D(n25080), .Z(n27282) );
    VMW_AO22 U519 ( .A(matrixInput[100]), .B(n25096), .C(matrixInput[92]), .D(
        n25081), .Z(n27164) );
    VMW_AO22 U629 ( .A(matrixInput[838]), .B(n25096), .C(matrixInput[830]), 
        .D(n25081), .Z(n26426) );
    VMW_AO22 U1077 ( .A(matrixInput[435]), .B(n25096), .C(matrixInput[427]), 
        .D(n25081), .Z(n26829) );
    VMW_AO22 U1666 ( .A(matrixInput[1748]), .B(n25096), .C(matrixInput[1740]), 
        .D(n25081), .Z(n25516) );
    VMW_FD \matrixInput_reg[1070]  ( .D(n26186), .CP(Clk), .Q(matrixInput
        [1070]) );
    VMW_FD \matrixInput_reg[1069]  ( .D(n26187), .CP(Clk), .Q(matrixInput
        [1069]) );
    VMW_AO22 U2377 ( .A(matrixInput[18]), .B(n25096), .C(matrixInput[10]), .D(
        n25081), .Z(n27246) );
    VMW_FD \matrixInput_reg[667]  ( .D(n26589), .CP(Clk), .Q(matrixInput[667])
         );
    VMW_FD \matrixInput_reg[557]  ( .D(n26699), .CP(Clk), .Q(matrixInput[557])
         );
    VMW_AO22 U697 ( .A(matrixInput[84]), .B(n25096), .C(matrixInput[76]), .D(
        n25081), .Z(n27180) );
    VMW_AO22 U707 ( .A(matrixInput[768]), .B(n25096), .C(matrixInput[760]), 
        .D(n25081), .Z(n26496) );
    VMW_AO22 U979 ( .A(matrixInput[523]), .B(n25096), .C(matrixInput[515]), 
        .D(n25081), .Z(n26741) );
    VMW_AO22 U1042 ( .A(matrixInput[467]), .B(n25096), .C(matrixInput[459]), 
        .D(n25081), .Z(n26797) );
    VMW_AO22 U1347 ( .A(matrixInput[2035]), .B(n25096), .C(matrixInput[2027]), 
        .D(n25081), .Z(n25229) );
    VMW_AO22 U1556 ( .A(matrixInput[191]), .B(n25096), .C(matrixInput[183]), 
        .D(n25081), .Z(n27073) );
    VMW_OAI21 U2566 ( .A(n25103), .B(n25104), .C(n25094), .Z(n25078) );
    VMW_FD \matrixInput_reg[1359]  ( .D(n25897), .CP(Clk), .Q(matrixInput
        [1359]) );
    VMW_FD \matrixInput_reg[1340]  ( .D(n25916), .CP(Clk), .Q(matrixInput
        [1340]) );
    VMW_FD \matrixInput_reg[654]  ( .D(n26602), .CP(Clk), .Q(matrixInput[654])
         );
    VMW_AO22 U1372 ( .A(matrixInput[2012]), .B(n25096), .C(matrixInput[2004]), 
        .D(n25081), .Z(n25252) );
    VMW_AO22 U1563 ( .A(matrixInput[1841]), .B(n25096), .C(matrixInput[1833]), 
        .D(n25081), .Z(n25423) );
    VMW_AO22 U1881 ( .A(matrixInput[1555]), .B(n25096), .C(matrixInput[1547]), 
        .D(n25081), .Z(n25709) );
    VMW_AO22 U1911 ( .A(matrixInput[159]), .B(n25096), .C(matrixInput[151]), 
        .D(n25081), .Z(n27105) );
    VMW_AO22 U1924 ( .A(matrixInput[1516]), .B(n25096), .C(matrixInput[1508]), 
        .D(n25081), .Z(n25748) );
    VMW_FD \matrixInput_reg[1043]  ( .D(n26213), .CP(Clk), .Q(matrixInput
        [1043]) );
    VMW_AO22 U2342 ( .A(matrixInput[1139]), .B(n25096), .C(matrixInput[1131]), 
        .D(n25081), .Z(n26125) );
    VMW_AO22 U2553 ( .A(cOutput[24]), .B(n25089), .C(cOutput[8]), .D(n25088), 
        .Z(n25175) );
    VMW_FD \matrixInput_reg[1126]  ( .D(n26130), .CP(Clk), .Q(matrixInput
        [1126]) );
    VMW_FD \matrixInput_reg[731]  ( .D(n26525), .CP(Clk), .Q(matrixInput[731])
         );
    VMW_FD \matrixInput_reg[728]  ( .D(n26528), .CP(Clk), .Q(matrixInput[728])
         );
    VMW_FD \matrixInput_reg[1225]  ( .D(n26031), .CP(Clk), .Q(matrixInput
        [1225]) );
    VMW_FD \matrixInput_reg[432]  ( .D(n26824), .CP(Clk), .Q(matrixInput[432])
         );
    VMW_AO22 U1653 ( .A(matrixInput[1760]), .B(n25096), .C(matrixInput[1752]), 
        .D(n25081), .Z(n25504) );
    VMW_AO22 U2072 ( .A(matrixInput[1383]), .B(n25096), .C(matrixInput[1375]), 
        .D(n25081), .Z(n25881) );
    VMW_FD \matrixInput_reg[1591]  ( .D(n25665), .CP(Clk), .Q(matrixInput
        [1591]) );
    VMW_FD \matrixInput_reg[1588]  ( .D(n25668), .CP(Clk), .Q(matrixInput
        [1588]) );
    VMW_FD \matrixInput_reg[1115]  ( .D(n26141), .CP(Clk), .Q(matrixInput
        [1115]) );
    VMW_FD \matrixInput_reg[702]  ( .D(n26554), .CP(Clk), .Q(matrixInput[702])
         );
    VMW_FD \matrixInput_reg[1692]  ( .D(n25564), .CP(Clk), .Q(matrixInput
        [1692]) );
    VMW_FD \matrixInput_reg[386]  ( .D(n26870), .CP(Clk), .Q(matrixInput[386])
         );
    VMW_FD \matrixInput_reg[1216]  ( .D(n26040), .CP(Clk), .Q(matrixInput
        [1216]) );
    VMW_FD \matrixInput_reg[418]  ( .D(n26838), .CP(Clk), .Q(matrixInput[418])
         );
    VMW_FD \matrixInput_reg[401]  ( .D(n26855), .CP(Clk), .Q(matrixInput[401])
         );
    VMW_AO22 U1065 ( .A(matrixInput[446]), .B(n25096), .C(matrixInput[438]), 
        .D(n25081), .Z(n26818) );
    VMW_AO22 U2055 ( .A(matrixInput[1398]), .B(n25096), .C(matrixInput[1390]), 
        .D(n25081), .Z(n25866) );
    VMW_FD \matrixInput_reg[1731]  ( .D(n25525), .CP(Clk), .Q(matrixInput
        [1731]) );
    VMW_FD \matrixInput_reg[1728]  ( .D(n25528), .CP(Clk), .Q(matrixInput
        [1728]) );
    VMW_FD \matrixInput_reg[126]  ( .D(n27130), .CP(Clk), .Q(matrixInput[126])
         );
    VMW_AO22 U1269 ( .A(matrixInput[262]), .B(n25096), .C(matrixInput[254]), 
        .D(n25081), .Z(n27002) );
    VMW_AO22 U1355 ( .A(matrixInput[209]), .B(n25096), .C(matrixInput[201]), 
        .D(n25081), .Z(n27055) );
    VMW_AO22 U1674 ( .A(matrixInput[1741]), .B(n25096), .C(matrixInput[1733]), 
        .D(n25081), .Z(n25523) );
    VMW_FD \matrixInput_reg[1432]  ( .D(n25824), .CP(Clk), .Q(matrixInput
        [1432]) );
    VMW_AO22 U1936 ( .A(matrixInput[1506]), .B(n25096), .C(matrixInput[1498]), 
        .D(n25081), .Z(n25758) );
    VMW_AO22 U2365 ( .A(matrixInput[1118]), .B(n25096), .C(matrixInput[1110]), 
        .D(n25081), .Z(n26146) );
    VMW_OAI21 U2574 ( .A(n25125), .B(n25126), .C(n25094), .Z(n25072) );
    VMW_FD \matrixInput_reg[225]  ( .D(n27031), .CP(Clk), .Q(matrixInput[225])
         );
    VMW_FD \matrixInput_reg[115]  ( .D(n27141), .CP(Clk), .Q(matrixInput[115])
         );
    VMW_FD \matrixInput_reg[1702]  ( .D(n25554), .CP(Clk), .Q(matrixInput
        [1702]) );
    VMW_FD \matrixInput_reg[1386]  ( .D(n25870), .CP(Clk), .Q(matrixInput
        [1386]) );
    VMW_FD \matrixInput_reg[1085]  ( .D(n26171), .CP(Clk), .Q(matrixInput
        [1085]) );
    VMW_FD \matrixInput_reg[591]  ( .D(n26665), .CP(Clk), .Q(matrixInput[591])
         );
    VMW_FD \matrixInput_reg[588]  ( .D(n26668), .CP(Clk), .Q(matrixInput[588])
         );
    VMW_FD \matrixInput_reg[692]  ( .D(n26564), .CP(Clk), .Q(matrixInput[692])
         );
    VMW_FD \matrixInput_reg[1418]  ( .D(n25838), .CP(Clk), .Q(matrixInput
        [1418]) );
    VMW_FD \matrixInput_reg[216]  ( .D(n27040), .CP(Clk), .Q(matrixInput[216])
         );
    VMW_AO22 U1544 ( .A(matrixInput[1858]), .B(n25096), .C(matrixInput[1850]), 
        .D(n25081), .Z(n25406) );
    VMW_FD \matrixInput_reg[1401]  ( .D(n25855), .CP(Clk), .Q(matrixInput
        [1401]) );
    VMW_AO22 U1478 ( .A(matrixInput[198]), .B(n25096), .C(matrixInput[190]), 
        .D(n25081), .Z(n27066) );
    VMW_FD \matrixInput_reg[1875]  ( .D(n25381), .CP(Clk), .Q(matrixInput
        [1875]) );
    VMW_FD \vectorInput_reg[85]  ( .D(n27299), .CP(Clk), .Q(vectorInput[85])
         );
    VMW_AO22 U2448 ( .A(matrixInput[1044]), .B(n25096), .C(matrixInput[1036]), 
        .D(n25081), .Z(n26220) );
    VMW_AO22 U1159 ( .A(matrixInput[361]), .B(n25096), .C(matrixInput[353]), 
        .D(n25081), .Z(n26903) );
    VMW_AO22 U2259 ( .A(matrixInput[1214]), .B(n25096), .C(matrixInput[1206]), 
        .D(n25081), .Z(n26050) );
    VMW_FD \matrixInput_reg[1846]  ( .D(n25410), .CP(Clk), .Q(matrixInput
        [1846]) );
    VMW_AO22 U1748 ( .A(matrixInput[1675]), .B(n25096), .C(matrixInput[1667]), 
        .D(n25081), .Z(n25589) );
    VMW_AO22 U580 ( .A(matrixInput[883]), .B(n25096), .C(matrixInput[875]), 
        .D(n25081), .Z(n26381) );
    VMW_AO22 U845 ( .A(matrixInput[644]), .B(n25096), .C(matrixInput[636]), 
        .D(n25081), .Z(n26620) );
    VMW_AO22 U2169 ( .A(matrixInput[1296]), .B(n25096), .C(matrixInput[1288]), 
        .D(n25081), .Z(n25968) );
    VMW_FD \vectorInput_reg[106]  ( .D(n27278), .CP(Clk), .Q(vectorInput[106])
         );
    VMW_FD \matrixInput_reg[875]  ( .D(n26381), .CP(Clk), .Q(matrixInput[875])
         );
    VMW_AO22 U410 ( .A(DataIn[7]), .B(n25095), .C(vectorInput[127]), .D(n25080
        ), .Z(n27257) );
    VMW_AO22 U459 ( .A(matrixInput[992]), .B(n25096), .C(matrixInput[984]), 
        .D(n25081), .Z(n26272) );
    VMW_AO22 U720 ( .A(matrixInput[757]), .B(n25096), .C(matrixInput[749]), 
        .D(n25081), .Z(n26507) );
    VMW_AO22 U862 ( .A(matrixInput[628]), .B(n25096), .C(matrixInput[620]), 
        .D(n25081), .Z(n26636) );
    VMW_FD \matrixInput_reg[846]  ( .D(n26410), .CP(Clk), .Q(matrixInput[846])
         );
    VMW_FD \matrixInput_reg[35]  ( .D(n27221), .CP(Clk), .Q(matrixInput[35])
         );
    VMW_AO22 U769 ( .A(matrixInput[712]), .B(n25096), .C(matrixInput[704]), 
        .D(n25081), .Z(n26552) );
    VMW_AO22 U1080 ( .A(matrixInput[432]), .B(n25096), .C(matrixInput[424]), 
        .D(n25081), .Z(n26832) );
    VMW_AO22 U1110 ( .A(matrixInput[406]), .B(n25096), .C(matrixInput[398]), 
        .D(n25081), .Z(n26858) );
    VMW_AO22 U1691 ( .A(matrixInput[1726]), .B(n25096), .C(matrixInput[1718]), 
        .D(n25081), .Z(n25538) );
    VMW_AO22 U1207 ( .A(matrixInput[38]), .B(n25096), .C(matrixInput[30]), .D(
        n25081), .Z(n27226) );
    VMW_AO22 U1220 ( .A(matrixInput[307]), .B(n25096), .C(matrixInput[299]), 
        .D(n25081), .Z(n26957) );
    VMW_AO22 U1701 ( .A(matrixInput[1717]), .B(n25096), .C(matrixInput[1709]), 
        .D(n25081), .Z(n25547) );
    VMW_AO22 U1843 ( .A(matrixInput[1589]), .B(n25096), .C(matrixInput[1581]), 
        .D(n25081), .Z(n25675) );
    VMW_AO22 U2120 ( .A(matrixInput[1339]), .B(n25096), .C(matrixInput[1331]), 
        .D(n25081), .Z(n25925) );
    VMW_FD \matrixInput_reg[1659]  ( .D(n25597), .CP(Clk), .Q(matrixInput
        [1659]) );
    VMW_FD \matrixInput_reg[1640]  ( .D(n25616), .CP(Clk), .Q(matrixInput
        [1640]) );
    VMW_FD \matrixInput_reg[1543]  ( .D(n25713), .CP(Clk), .Q(matrixInput
        [1543]) );
    VMW_FD \matrixInput_reg[354]  ( .D(n26902), .CP(Clk), .Q(matrixInput[354])
         );
    VMW_FD \matrixInput_reg[2027]  ( .D(n25229), .CP(Clk), .Q(matrixInput
        [2027]) );
    VMW_FD \matrixInput_reg[1673]  ( .D(n25583), .CP(Clk), .Q(matrixInput
        [1673]) );
    VMW_AO22 U1397 ( .A(matrixInput[1991]), .B(n25096), .C(matrixInput[1983]), 
        .D(n25081), .Z(n25273) );
    VMW_AO22 U1416 ( .A(matrixInput[1974]), .B(n25096), .C(matrixInput[1966]), 
        .D(n25081), .Z(n25290) );
    VMW_AO22 U1431 ( .A(matrixInput[1960]), .B(n25096), .C(matrixInput[1952]), 
        .D(n25081), .Z(n25304) );
    VMW_AO22 U1864 ( .A(matrixInput[1570]), .B(n25096), .C(matrixInput[1562]), 
        .D(n25081), .Z(n25694) );
    VMW_AO22 U2210 ( .A(matrixInput[1258]), .B(n25096), .C(matrixInput[1250]), 
        .D(n25081), .Z(n26006) );
    VMW_AO22 U2380 ( .A(matrixInput[1106]), .B(n25096), .C(matrixInput[1098]), 
        .D(n25081), .Z(n26158) );
    VMW_AO22 U2401 ( .A(matrixInput[1087]), .B(n25096), .C(matrixInput[1079]), 
        .D(n25081), .Z(n26177) );
    VMW_FD \matrixInput_reg[2014]  ( .D(n25242), .CP(Clk), .Q(matrixInput
        [2014]) );
    VMW_OAI21 U2591 ( .A(n25174), .B(n25175), .C(n25090), .Z(n25183) );
    VMW_FD \matrixInput_reg[1570]  ( .D(n25686), .CP(Clk), .Q(matrixInput
        [1570]) );
    VMW_FD \matrixInput_reg[1569]  ( .D(n25687), .CP(Clk), .Q(matrixInput
        [1569]) );
    VMW_FD \matrixInput_reg[367]  ( .D(n26889), .CP(Clk), .Q(matrixInput[367])
         );
    VMW_FD \matrixInput_reg[659]  ( .D(n26597), .CP(Clk), .Q(matrixInput[659])
         );
    VMW_AO22 U1586 ( .A(matrixInput[1820]), .B(n25096), .C(matrixInput[1812]), 
        .D(n25081), .Z(n25444) );
    VMW_FD \matrixInput_reg[640]  ( .D(n26616), .CP(Clk), .Q(matrixInput[640])
         );
    VMW_AO22 U2237 ( .A(matrixInput[1234]), .B(n25096), .C(matrixInput[1226]), 
        .D(n25081), .Z(n26030) );
    VMW_FD \matrixInput_reg[1057]  ( .D(n26199), .CP(Clk), .Q(matrixInput
        [1057]) );
    VMW_FD \matrixInput_reg[543]  ( .D(n26713), .CP(Clk), .Q(matrixInput[543])
         );
    VMW_AO22 U1137 ( .A(matrixInput[381]), .B(n25096), .C(matrixInput[373]), 
        .D(n25081), .Z(n26883) );
    VMW_AO22 U1726 ( .A(matrixInput[1695]), .B(n25096), .C(matrixInput[1687]), 
        .D(n25081), .Z(n25569) );
    VMW_AO22 U2426 ( .A(matrixInput[1064]), .B(n25096), .C(matrixInput[1056]), 
        .D(n25081), .Z(n26200) );
    VMW_FD \matrixInput_reg[1354]  ( .D(n25902), .CP(Clk), .Q(matrixInput
        [1354]) );
    VMW_FD \matrixInput_reg[1064]  ( .D(n26192), .CP(Clk), .Q(matrixInput
        [1064]) );
    VMW_AO22 U2097 ( .A(matrixInput[1360]), .B(n25096), .C(matrixInput[1352]), 
        .D(n25081), .Z(n25904) );
    VMW_AO22 U2107 ( .A(matrixInput[1351]), .B(n25096), .C(matrixInput[1343]), 
        .D(n25081), .Z(n25913) );
    VMW_FD \matrixInput_reg[1367]  ( .D(n25889), .CP(Clk), .Q(matrixInput
        [1367]) );
    VMW_FD \matrixInput_reg[673]  ( .D(n26583), .CP(Clk), .Q(matrixInput[673])
         );
    VMW_FD \matrixInput_reg[570]  ( .D(n26686), .CP(Clk), .Q(matrixInput[570])
         );
    VMW_FD \matrixInput_reg[569]  ( .D(n26687), .CP(Clk), .Q(matrixInput[569])
         );
    VMW_AO22 U542 ( .A(matrixInput[917]), .B(n25096), .C(matrixInput[909]), 
        .D(n25081), .Z(n26347) );
    VMW_AO22 U565 ( .A(matrixInput[897]), .B(n25096), .C(matrixInput[889]), 
        .D(n25081), .Z(n26367) );
    VMW_AO22 U655 ( .A(matrixInput[815]), .B(n25096), .C(matrixInput[807]), 
        .D(n25081), .Z(n26449) );
    VMW_AO22 U887 ( .A(matrixInput[607]), .B(n25096), .C(matrixInput[599]), 
        .D(n25081), .Z(n26657) );
    VMW_AO22 U917 ( .A(matrixInput[579]), .B(n25096), .C(matrixInput[571]), 
        .D(n25081), .Z(n26685) );
    VMW_FD \matrixInput_reg[904]  ( .D(n26352), .CP(Clk), .Q(matrixInput[904])
         );
    VMW_FD \matrixInput_reg[1894]  ( .D(n25362), .CP(Clk), .Q(matrixInput
        [1894]) );
    VMW_FD \vectorInput_reg[64]  ( .D(n27320), .CP(Clk), .Q(vectorInput[64])
         );
    VMW_FD \matrixInput_reg[937]  ( .D(n26319), .CP(Clk), .Q(matrixInput[937])
         );
    VMW_AO22 U672 ( .A(matrixInput[800]), .B(n25096), .C(matrixInput[792]), 
        .D(n25081), .Z(n26464) );
    VMW_AO22 U1958 ( .A(matrixInput[1486]), .B(n25096), .C(matrixInput[1478]), 
        .D(n25081), .Z(n25778) );
    VMW_FD \vectorInput_reg[57]  ( .D(n27327), .CP(Clk), .Q(vectorInput[57])
         );
    VMW_FD \matrixInput_reg[1937]  ( .D(n25319), .CP(Clk), .Q(matrixInput
        [1937]) );
    VMW_FD \matrixInput_reg[1904]  ( .D(n25352), .CP(Clk), .Q(matrixInput
        [1904]) );
    VMW_FD \matrixInput_reg[894]  ( .D(n26362), .CP(Clk), .Q(matrixInput[894])
         );
    VMW_AO22 U559 ( .A(matrixInput[902]), .B(n25096), .C(matrixInput[894]), 
        .D(n25081), .Z(n26362) );
    VMW_AO22 U930 ( .A(matrixInput[63]), .B(n25096), .C(matrixInput[55]), .D(
        n25081), .Z(n27201) );
    VMW_AO22 U1037 ( .A(matrixInput[471]), .B(n25096), .C(matrixInput[463]), 
        .D(n25081), .Z(n26793) );
    VMW_AO22 U1626 ( .A(matrixInput[1785]), .B(n25096), .C(matrixInput[1777]), 
        .D(n25081), .Z(n25479) );
    VMW_FD \matrixInput_reg[663]  ( .D(n26593), .CP(Clk), .Q(matrixInput[663])
         );
    VMW_AO22 U2197 ( .A(matrixInput[1270]), .B(n25096), .C(matrixInput[1262]), 
        .D(n25081), .Z(n25994) );
    VMW_FD \matrixInput_reg[1074]  ( .D(n26182), .CP(Clk), .Q(matrixInput
        [1074]) );
    VMW_FD \matrixInput_reg[579]  ( .D(n26677), .CP(Clk), .Q(matrixInput[579])
         );
    VMW_BUFIZ U2616 ( .A(n25191), .E(RD), .Z(\DataOut[25]1 ) );
    VMW_AO22 U442 ( .A(matrixInput[107]), .B(n25096), .C(matrixInput[99]), .D(
        n25081), .Z(n27157) );
    VMW_AO22 U669 ( .A(matrixInput[803]), .B(n25096), .C(matrixInput[795]), 
        .D(n25081), .Z(n26461) );
    VMW_AO22 U1297 ( .A(matrixInput[237]), .B(n25096), .C(matrixInput[229]), 
        .D(n25081), .Z(n27027) );
    VMW_AO22 U1307 ( .A(matrixInput[29]), .B(n25096), .C(matrixInput[21]), .D(
        n25081), .Z(n27235) );
    VMW_AO22 U1486 ( .A(matrixInput[1910]), .B(n25096), .C(matrixInput[1902]), 
        .D(n25081), .Z(n25354) );
    VMW_AO22 U1964 ( .A(matrixInput[1480]), .B(n25096), .C(matrixInput[1472]), 
        .D(n25081), .Z(n25784) );
    VMW_AO22 U2007 ( .A(matrixInput[1441]), .B(n25096), .C(matrixInput[1433]), 
        .D(n25081), .Z(n25823) );
    VMW_FD \matrixInput_reg[1377]  ( .D(n25879), .CP(Clk), .Q(matrixInput
        [1377]) );
    VMW_FD \matrixInput_reg[560]  ( .D(n26696), .CP(Clk), .Q(matrixInput[560])
         );
    VMW_FD \matrixInput_reg[1047]  ( .D(n26209), .CP(Clk), .Q(matrixInput
        [1047]) );
    VMW_FD \matrixInput_reg[650]  ( .D(n26606), .CP(Clk), .Q(matrixInput[650])
         );
    VMW_AO22 U1516 ( .A(matrixInput[1884]), .B(n25096), .C(matrixInput[1876]), 
        .D(n25081), .Z(n25380) );
    VMW_FD \matrixInput_reg[649]  ( .D(n26607), .CP(Clk), .Q(matrixInput[649])
         );
    VMW_FD \matrixInput_reg[1344]  ( .D(n25912), .CP(Clk), .Q(matrixInput
        [1344]) );
    VMW_AO22 U1010 ( .A(matrixInput[496]), .B(n25096), .C(matrixInput[488]), 
        .D(n25081), .Z(n26768) );
    VMW_AO22 U1180 ( .A(matrixInput[342]), .B(n25096), .C(matrixInput[334]), 
        .D(n25081), .Z(n26922) );
    VMW_AO22 U1320 ( .A(matrixInput[216]), .B(n25096), .C(matrixInput[208]), 
        .D(n25081), .Z(n27048) );
    VMW_AO22 U1531 ( .A(matrixInput[1870]), .B(n25096), .C(matrixInput[1862]), 
        .D(n25081), .Z(n25394) );
    VMW_AO22 U1943 ( .A(matrixInput[1499]), .B(n25096), .C(matrixInput[1491]), 
        .D(n25081), .Z(n25765) );
    VMW_AO22 U2337 ( .A(matrixInput[1144]), .B(n25096), .C(matrixInput[1136]), 
        .D(n25081), .Z(n26120) );
    VMW_AO22 U2526 ( .A(cOutput[27]), .B(n25089), .C(cOutput[11]), .D(n25088), 
        .Z(n25142) );
    VMW_FD \matrixInput_reg[553]  ( .D(n26703), .CP(Clk), .Q(matrixInput[553])
         );
    VMW_FD \matrixInput_reg[1663]  ( .D(n25593), .CP(Clk), .Q(matrixInput
        [1663]) );
    VMW_AO22 U2280 ( .A(matrixInput[1196]), .B(n25096), .C(matrixInput[1188]), 
        .D(n25081), .Z(n26068) );
    VMW_AO22 U2310 ( .A(matrixInput[1168]), .B(n25096), .C(matrixInput[1160]), 
        .D(n25081), .Z(n26096) );
    VMW_AO22 U2491 ( .A(cOutput[55]), .B(n25087), .C(cOutput[39]), .D(n25084), 
        .Z(n25099) );
    VMW_AO22 U2501 ( .A(cOutput[62]), .B(n25089), .C(cOutput[46]), .D(n25088), 
        .Z(n25111) );
    VMW_FD \matrixInput_reg[2004]  ( .D(n25252), .CP(Clk), .Q(matrixInput
        [2004]) );
    VMW_FD \matrixInput_reg[1579]  ( .D(n25677), .CP(Clk), .Q(matrixInput
        [1579]) );
    VMW_FD \matrixInput_reg[377]  ( .D(n26879), .CP(Clk), .Q(matrixInput[377])
         );
    VMW_FD \matrixInput_reg[1560]  ( .D(n25696), .CP(Clk), .Q(matrixInput
        [1560]) );
    VMW_AO22 U1601 ( .A(matrixInput[187]), .B(n25096), .C(matrixInput[179]), 
        .D(n25081), .Z(n27077) );
    VMW_AO22 U1791 ( .A(matrixInput[1636]), .B(n25096), .C(matrixInput[1628]), 
        .D(n25081), .Z(n25628) );
    VMW_AO22 U2020 ( .A(matrixInput[1429]), .B(n25096), .C(matrixInput[1421]), 
        .D(n25081), .Z(n25835) );
    VMW_FD \matrixInput_reg[2037]  ( .D(n25219), .CP(Clk), .Q(matrixInput
        [2037]) );
    VMW_FD \matrixInput_reg[1650]  ( .D(n25606), .CP(Clk), .Q(matrixInput
        [1650]) );
    VMW_FD \matrixInput_reg[1649]  ( .D(n25607), .CP(Clk), .Q(matrixInput
        [1649]) );
    VMW_FD \matrixInput_reg[1553]  ( .D(n25703), .CP(Clk), .Q(matrixInput
        [1553]) );
    VMW_FD \matrixInput_reg[344]  ( .D(n26912), .CP(Clk), .Q(matrixInput[344])
         );
    VMW_BUFIZ U2631 ( .A(\holder[3] ), .E(RD), .Z(\DataOut[3]1 ) );
    VMW_AO22 U465 ( .A(matrixInput[987]), .B(n25096), .C(matrixInput[979]), 
        .D(n25081), .Z(n26277) );
    VMW_AO22 U755 ( .A(matrixInput[725]), .B(n25096), .C(matrixInput[717]), 
        .D(n25081), .Z(n26539) );
    VMW_AO22 U772 ( .A(matrixInput[709]), .B(n25096), .C(matrixInput[701]), 
        .D(n25081), .Z(n26555) );
    VMW_AO22 U830 ( .A(matrixInput[72]), .B(n25096), .C(matrixInput[64]), .D(
        n25081), .Z(n27192) );
    VMW_FD \matrixInput_reg[1927]  ( .D(n25329), .CP(Clk), .Q(matrixInput
        [1927]) );
    VMW_FD \matrixInput_reg[4]  ( .D(n27252), .CP(Clk), .Q(matrixInput[4]) );
    VMW_FD \matrixInput_reg[1914]  ( .D(n25342), .CP(Clk), .Q(matrixInput
        [1914]) );
    VMW_FD \matrixInput_reg[927]  ( .D(n26329), .CP(Clk), .Q(matrixInput[927])
         );
    VMW_FD \matrixInput_reg[884]  ( .D(n26372), .CP(Clk), .Q(matrixInput[884])
         );
    VMW_AO22 U1858 ( .A(matrixInput[1576]), .B(n25096), .C(matrixInput[1568]), 
        .D(n25081), .Z(n25688) );
    VMW_FD \vectorInput_reg[47]  ( .D(n27337), .CP(Clk), .Q(vectorInput[47])
         );
    VMW_PULLDOWN U291 ( .Z(n27393) );
    VMW_AO22 U620 ( .A(matrixInput[847]), .B(n25096), .C(matrixInput[839]), 
        .D(n25081), .Z(n26417) );
    VMW_AO22 U817 ( .A(matrixInput[669]), .B(n25096), .C(matrixInput[661]), 
        .D(n25081), .Z(n26595) );
    VMW_AO22 U879 ( .A(matrixInput[613]), .B(n25096), .C(matrixInput[605]), 
        .D(n25081), .Z(n26651) );
    VMW_AO22 U987 ( .A(matrixInput[516]), .B(n25096), .C(matrixInput[508]), 
        .D(n25081), .Z(n26748) );
    VMW_FD \matrixInput_reg[914]  ( .D(n26342), .CP(Clk), .Q(matrixInput[914])
         );
    VMW_AO22 U1255 ( .A(matrixInput[275]), .B(n25096), .C(matrixInput[267]), 
        .D(n25081), .Z(n26989) );
    VMW_AO22 U1444 ( .A(matrixInput[1948]), .B(n25096), .C(matrixInput[1940]), 
        .D(n25081), .Z(n25316) );
    VMW_AO22 U1836 ( .A(matrixInput[1596]), .B(n25096), .C(matrixInput[1588]), 
        .D(n25081), .Z(n25668) );
    VMW_AO22 U2265 ( .A(matrixInput[1208]), .B(n25096), .C(matrixInput[1200]), 
        .D(n25081), .Z(n26056) );
    VMW_FD \matrixInput_reg[1884]  ( .D(n25372), .CP(Clk), .Q(matrixInput
        [1884]) );
    VMW_FD \vectorInput_reg[74]  ( .D(n27310), .CP(Clk), .Q(vectorInput[74])
         );
    VMW_AO22 U2474 ( .A(matrixInput[1020]), .B(n25096), .C(matrixInput[1012]), 
        .D(n25081), .Z(n26244) );
    VMW_FD \matrixInput_reg[1712]  ( .D(n25544), .CP(Clk), .Q(matrixInput
        [1712]) );
    VMW_FD \matrixInput_reg[1396]  ( .D(n25860), .CP(Clk), .Q(matrixInput
        [1396]) );
    VMW_FD \matrixInput_reg[598]  ( .D(n26658), .CP(Clk), .Q(matrixInput[598])
         );
    VMW_FD \matrixInput_reg[581]  ( .D(n26675), .CP(Clk), .Q(matrixInput[581])
         );
    VMW_FD \matrixInput_reg[105]  ( .D(n27151), .CP(Clk), .Q(matrixInput[105])
         );
    VMW_FD \matrixInput_reg[1411]  ( .D(n25845), .CP(Clk), .Q(matrixInput
        [1411]) );
    VMW_FD \matrixInput_reg[1095]  ( .D(n26161), .CP(Clk), .Q(matrixInput
        [1095]) );
    VMW_FD \matrixInput_reg[682]  ( .D(n26574), .CP(Clk), .Q(matrixInput[682])
         );
    VMW_FD \matrixInput_reg[1408]  ( .D(n25848), .CP(Clk), .Q(matrixInput
        [1408]) );
    VMW_FD \matrixInput_reg[206]  ( .D(n27050), .CP(Clk), .Q(matrixInput[206])
         );
    VMW_AO22 U1142 ( .A(matrixInput[377]), .B(n25096), .C(matrixInput[369]), 
        .D(n25081), .Z(n26887) );
    VMW_AO22 U1165 ( .A(matrixInput[356]), .B(n25096), .C(matrixInput[348]), 
        .D(n25081), .Z(n26908) );
    VMW_AO22 U1774 ( .A(matrixInput[1651]), .B(n25096), .C(matrixInput[1643]), 
        .D(n25081), .Z(n25613) );
    VMW_AO22 U2155 ( .A(matrixInput[20]), .B(n25096), .C(matrixInput[12]), .D(
        n25081), .Z(n27244) );
    VMW_FD \matrixInput_reg[136]  ( .D(n27120), .CP(Clk), .Q(matrixInput[136])
         );
    VMW_FD \matrixInput_reg[1738]  ( .D(n25518), .CP(Clk), .Q(matrixInput
        [1738]) );
    VMW_FD \matrixInput_reg[1721]  ( .D(n25535), .CP(Clk), .Q(matrixInput
        [1721]) );
    VMW_FD \matrixInput_reg[1422]  ( .D(n25834), .CP(Clk), .Q(matrixInput
        [1422]) );
    VMW_FD \matrixInput_reg[235]  ( .D(n27021), .CP(Clk), .Q(matrixInput[235])
         );
    VMW_AO22 U2172 ( .A(matrixInput[1293]), .B(n25096), .C(matrixInput[1285]), 
        .D(n25081), .Z(n25971) );
    VMW_FD \matrixInput_reg[1105]  ( .D(n26151), .CP(Clk), .Q(matrixInput
        [1105]) );
    VMW_FD \matrixInput_reg[712]  ( .D(n26544), .CP(Clk), .Q(matrixInput[712])
         );
    VMW_FD \matrixInput_reg[396]  ( .D(n26860), .CP(Clk), .Q(matrixInput[396])
         );
    VMW_FD \matrixInput_reg[1598]  ( .D(n25658), .CP(Clk), .Q(matrixInput
        [1598]) );
    VMW_FD \matrixInput_reg[1581]  ( .D(n25675), .CP(Clk), .Q(matrixInput
        [1581]) );
    VMW_AO22 U1272 ( .A(matrixInput[259]), .B(n25096), .C(matrixInput[251]), 
        .D(n25081), .Z(n27005) );
    VMW_AO22 U1753 ( .A(matrixInput[1670]), .B(n25096), .C(matrixInput[1662]), 
        .D(n25081), .Z(n25594) );
    VMW_AO22 U1811 ( .A(matrixInput[168]), .B(n25096), .C(matrixInput[160]), 
        .D(n25081), .Z(n27096) );
    VMW_AO22 U1981 ( .A(matrixInput[1465]), .B(n25096), .C(matrixInput[1457]), 
        .D(n25081), .Z(n25799) );
    VMW_AO22 U2242 ( .A(matrixInput[1229]), .B(n25096), .C(matrixInput[1221]), 
        .D(n25081), .Z(n26035) );
    VMW_AO22 U2453 ( .A(matrixInput[1039]), .B(n25096), .C(matrixInput[1031]), 
        .D(n25081), .Z(n26225) );
    VMW_FD \matrixInput_reg[1682]  ( .D(n25574), .CP(Clk), .Q(matrixInput
        [1682]) );
    VMW_FD \matrixInput_reg[1206]  ( .D(n26050), .CP(Clk), .Q(matrixInput
        [1206]) );
    VMW_FD \matrixInput_reg[411]  ( .D(n26845), .CP(Clk), .Q(matrixInput[411])
         );
    VMW_FD \matrixInput_reg[408]  ( .D(n26848), .CP(Clk), .Q(matrixInput[408])
         );
    VMW_FD \matrixInput_reg[1136]  ( .D(n26120), .CP(Clk), .Q(matrixInput
        [1136]) );
    VMW_FD \matrixInput_reg[738]  ( .D(n26518), .CP(Clk), .Q(matrixInput[738])
         );
    VMW_FD \matrixInput_reg[721]  ( .D(n26535), .CP(Clk), .Q(matrixInput[721])
         );
    VMW_FD \vectorInput_reg[2]  ( .D(n27382), .CP(Clk), .Q(vectorInput[2]) );
    VMW_FD \matrixInput_reg[422]  ( .D(n26834), .CP(Clk), .Q(matrixInput[422])
         );
    VMW_FD \matrixInput_reg[1235]  ( .D(n26021), .CP(Clk), .Q(matrixInput
        [1235]) );
    VMW_AO22 U1463 ( .A(matrixInput[1931]), .B(n25096), .C(matrixInput[1923]), 
        .D(n25081), .Z(n25333) );
    VMW_FD \matrixInput_reg[856]  ( .D(n26400), .CP(Clk), .Q(matrixInput[856])
         );
    VMW_FD \matrixInput_reg[16]  ( .D(n27240), .CP(Clk), .Q(matrixInput[16])
         );
    VMW_FD \matrixInput_reg[865]  ( .D(n26391), .CP(Clk), .Q(matrixInput[865])
         );
    VMW_OAI211 U296 ( .A(n25055), .B(n25062), .C(n25063), .D(n25064), .Z(
        n27390) );
    VMW_OAI211 U301 ( .A(n25055), .B(n25077), .C(n25078), .D(n25079), .Z(
        n27385) );
    VMW_AO22 U510 ( .A(matrixInput[946]), .B(n25096), .C(matrixInput[938]), 
        .D(n25081), .Z(n26318) );
    VMW_AND2 U306 ( .A(n25086), .B(n25085), .Z(n25087) );
    VMW_AO22 U321 ( .A(vectorInput[100]), .B(n25095), .C(vectorInput[92]), .D(
        n25080), .Z(n27292) );
    VMW_AO22 U326 ( .A(vectorInput[96]), .B(n25095), .C(vectorInput[88]), .D(
        n25080), .Z(n27296) );
    VMW_AO22 U480 ( .A(matrixInput[973]), .B(n25096), .C(matrixInput[965]), 
        .D(n25081), .Z(n26291) );
    VMW_AO22 U962 ( .A(matrixInput[538]), .B(n25096), .C(matrixInput[530]), 
        .D(n25081), .Z(n26726) );
    VMW_FD \matrixInput_reg[25]  ( .D(n27231), .CP(Clk), .Q(matrixInput[25])
         );
    VMW_AO22 U1059 ( .A(matrixInput[451]), .B(n25096), .C(matrixInput[443]), 
        .D(n25081), .Z(n26813) );
    VMW_AO22 U1648 ( .A(matrixInput[1765]), .B(n25096), .C(matrixInput[1757]), 
        .D(n25081), .Z(n25499) );
    VMW_FD \matrixInput_reg[1856]  ( .D(n25400), .CP(Clk), .Q(matrixInput
        [1856]) );
    VMW_AO22 U530 ( .A(matrixInput[99]), .B(n25096), .C(matrixInput[91]), .D(
        n25081), .Z(n27165) );
    VMW_AO22 U537 ( .A(matrixInput[921]), .B(n25096), .C(matrixInput[913]), 
        .D(n25081), .Z(n26343) );
    VMW_AO22 U2069 ( .A(matrixInput[1386]), .B(n25096), .C(matrixInput[1378]), 
        .D(n25081), .Z(n25878) );
    VMW_FD \vectorInput_reg[116]  ( .D(n27268), .CP(Clk), .Q(vectorInput[116])
         );
    VMW_AO22 U600 ( .A(matrixInput[865]), .B(n25096), .C(matrixInput[857]), 
        .D(n25081), .Z(n26399) );
    VMW_AO22 U607 ( .A(matrixInput[858]), .B(n25096), .C(matrixInput[850]), 
        .D(n25081), .Z(n26406) );
    VMW_AO22 U797 ( .A(matrixInput[75]), .B(n25096), .C(matrixInput[67]), .D(
        n25081), .Z(n27189) );
    VMW_AO22 U945 ( .A(matrixInput[554]), .B(n25096), .C(matrixInput[546]), 
        .D(n25081), .Z(n26710) );
    VMW_AO22 U1369 ( .A(matrixInput[2015]), .B(n25096), .C(matrixInput[2007]), 
        .D(n25081), .Z(n25249) );
    VMW_AO22 U1578 ( .A(matrixInput[189]), .B(n25096), .C(matrixInput[181]), 
        .D(n25081), .Z(n27075) );
    VMW_FD \vectorInput_reg[95]  ( .D(n27289), .CP(Clk), .Q(vectorInput[95])
         );
    VMW_FD \matrixInput_reg[1865]  ( .D(n25391), .CP(Clk), .Q(matrixInput
        [1865]) );
    VMW_AO22 U2359 ( .A(matrixInput[1124]), .B(n25096), .C(matrixInput[1116]), 
        .D(n25081), .Z(n26140) );
    VMW_FD \vectorInput_reg[125]  ( .D(n27259), .CP(Clk), .Q(vectorInput[125])
         );
    VMW_AO22 U859 ( .A(matrixInput[631]), .B(n25096), .C(matrixInput[623]), 
        .D(n25081), .Z(n26633) );
    VMW_AO22 U1145 ( .A(matrixInput[374]), .B(n25096), .C(matrixInput[366]), 
        .D(n25081), .Z(n26890) );
    VMW_AO22 U1275 ( .A(matrixInput[257]), .B(n25096), .C(matrixInput[249]), 
        .D(n25081), .Z(n27007) );
    VMW_AO22 U1464 ( .A(matrixInput[1930]), .B(n25096), .C(matrixInput[1922]), 
        .D(n25081), .Z(n25334) );
    VMW_AO22 U2548 ( .A(cOutput[89]), .B(n25089), .C(cOutput[73]), .D(n25088), 
        .Z(n25168) );
    VMW_FD \matrixInput_reg[1413]  ( .D(n25843), .CP(Clk), .Q(matrixInput
        [1413]) );
    VMW_FD \matrixInput_reg[204]  ( .D(n27052), .CP(Clk), .Q(matrixInput[204])
         );
    VMW_AO22 U1754 ( .A(matrixInput[1669]), .B(n25096), .C(matrixInput[1661]), 
        .D(n25081), .Z(n25595) );
    VMW_AO22 U1816 ( .A(matrixInput[1613]), .B(n25096), .C(matrixInput[1605]), 
        .D(n25081), .Z(n25651) );
    VMW_FD \matrixInput_reg[1097]  ( .D(n26159), .CP(Clk), .Q(matrixInput
        [1097]) );
    VMW_AO22 U1986 ( .A(matrixInput[1460]), .B(n25096), .C(matrixInput[1452]), 
        .D(n25081), .Z(n25804) );
    VMW_FD \matrixInput_reg[699]  ( .D(n26557), .CP(Clk), .Q(matrixInput[699])
         );
    VMW_AO22 U2245 ( .A(matrixInput[1227]), .B(n25096), .C(matrixInput[1219]), 
        .D(n25081), .Z(n26037) );
    VMW_FD \matrixInput_reg[1394]  ( .D(n25862), .CP(Clk), .Q(matrixInput
        [1394]) );
    VMW_FD \matrixInput_reg[680]  ( .D(n26576), .CP(Clk), .Q(matrixInput[680])
         );
    VMW_FD \matrixInput_reg[583]  ( .D(n26673), .CP(Clk), .Q(matrixInput[583])
         );
    VMW_FD \matrixInput_reg[107]  ( .D(n27149), .CP(Clk), .Q(matrixInput[107])
         );
    VMW_AO22 U2454 ( .A(matrixInput[1038]), .B(n25096), .C(matrixInput[1030]), 
        .D(n25081), .Z(n26226) );
    VMW_FD \matrixInput_reg[1709]  ( .D(n25547), .CP(Clk), .Q(matrixInput
        [1709]) );
    VMW_FD \matrixInput_reg[1710]  ( .D(n25546), .CP(Clk), .Q(matrixInput
        [1710]) );
    VMW_FD \matrixInput_reg[1420]  ( .D(n25836), .CP(Clk), .Q(matrixInput
        [1420]) );
    VMW_FD \matrixInput_reg[1439]  ( .D(n25817), .CP(Clk), .Q(matrixInput
        [1439]) );
    VMW_AO22 U2175 ( .A(matrixInput[1290]), .B(n25096), .C(matrixInput[1282]), 
        .D(n25081), .Z(n25974) );
    VMW_FD \matrixInput_reg[237]  ( .D(n27019), .CP(Clk), .Q(matrixInput[237])
         );
    VMW_FD \matrixInput_reg[1723]  ( .D(n25533), .CP(Clk), .Q(matrixInput
        [1723]) );
    VMW_FD \matrixInput_reg[134]  ( .D(n27122), .CP(Clk), .Q(matrixInput[134])
         );
    VMW_AO22 U1162 ( .A(matrixInput[358]), .B(n25096), .C(matrixInput[350]), 
        .D(n25081), .Z(n26906) );
    VMW_FD \matrixInput_reg[1699]  ( .D(n25557), .CP(Clk), .Q(matrixInput
        [1699]) );
    VMW_FD \matrixInput_reg[1204]  ( .D(n26052), .CP(Clk), .Q(matrixInput
        [1204]) );
    VMW_FD \matrixInput_reg[413]  ( .D(n26843), .CP(Clk), .Q(matrixInput[413])
         );
    VMW_FD \matrixInput_reg[1680]  ( .D(n25576), .CP(Clk), .Q(matrixInput
        [1680]) );
    VMW_AO22 U1252 ( .A(matrixInput[34]), .B(n25096), .C(matrixInput[26]), .D(
        n25081), .Z(n27230) );
    VMW_AO22 U1773 ( .A(matrixInput[1652]), .B(n25096), .C(matrixInput[1644]), 
        .D(n25081), .Z(n25612) );
    VMW_AO22 U2152 ( .A(matrixInput[1310]), .B(n25096), .C(matrixInput[1302]), 
        .D(n25081), .Z(n25954) );
    VMW_FD \matrixInput_reg[1583]  ( .D(n25673), .CP(Clk), .Q(matrixInput
        [1583]) );
    VMW_FD \matrixInput_reg[394]  ( .D(n26862), .CP(Clk), .Q(matrixInput[394])
         );
    VMW_FD \matrixInput_reg[1107]  ( .D(n26149), .CP(Clk), .Q(matrixInput
        [1107]) );
    VMW_FD \matrixInput_reg[710]  ( .D(n26546), .CP(Clk), .Q(matrixInput[710])
         );
    VMW_FD \matrixInput_reg[709]  ( .D(n26547), .CP(Clk), .Q(matrixInput[709])
         );
    VMW_AO22 U1443 ( .A(matrixInput[1949]), .B(n25096), .C(matrixInput[1941]), 
        .D(n25081), .Z(n25315) );
    VMW_AO22 U1831 ( .A(matrixInput[1600]), .B(n25096), .C(matrixInput[1592]), 
        .D(n25081), .Z(n25664) );
    VMW_FD \matrixInput_reg[1237]  ( .D(n26019), .CP(Clk), .Q(matrixInput
        [1237]) );
    VMW_AO22 U2262 ( .A(matrixInput[1211]), .B(n25096), .C(matrixInput[1203]), 
        .D(n25081), .Z(n26053) );
    VMW_AO22 U2473 ( .A(matrixInput[1021]), .B(n25096), .C(matrixInput[1013]), 
        .D(n25081), .Z(n26243) );
    VMW_FD \matrixInput_reg[1134]  ( .D(n26122), .CP(Clk), .Q(matrixInput
        [1134]) );
    VMW_FD \matrixInput_reg[439]  ( .D(n26817), .CP(Clk), .Q(matrixInput[439])
         );
    VMW_FD \matrixInput_reg[420]  ( .D(n26836), .CP(Clk), .Q(matrixInput[420])
         );
    VMW_FD \matrixInput_reg[723]  ( .D(n26533), .CP(Clk), .Q(matrixInput[723])
         );
    VMW_FD \vectorInput_reg[0]  ( .D(n27384), .CP(Clk), .Q(vectorInput[0]) );
    VMW_AO22 U790 ( .A(matrixInput[694]), .B(n25096), .C(matrixInput[686]), 
        .D(n25081), .Z(n26570) );
    VMW_AO22 U942 ( .A(matrixInput[557]), .B(n25096), .C(matrixInput[549]), 
        .D(n25081), .Z(n26707) );
    VMW_FD \matrixInput_reg[854]  ( .D(n26402), .CP(Clk), .Q(matrixInput[854])
         );
    VMW_FD \matrixInput_reg[14]  ( .D(n27242), .CP(Clk), .Q(matrixInput[14])
         );
    VMW_FD \matrixInput_reg[27]  ( .D(n27229), .CP(Clk), .Q(matrixInput[27])
         );
    VMW_AO22 U487 ( .A(matrixInput[967]), .B(n25096), .C(matrixInput[959]), 
        .D(n25081), .Z(n26297) );
    VMW_AO22 U965 ( .A(matrixInput[536]), .B(n25096), .C(matrixInput[528]), 
        .D(n25081), .Z(n26728) );
    VMW_FD \matrixInput_reg[867]  ( .D(n26389), .CP(Clk), .Q(matrixInput[867])
         );
    VMW_FD \vectorInput_reg[114]  ( .D(n27270), .CP(Clk), .Q(vectorInput[114])
         );
    VMW_AO22 U517 ( .A(matrixInput[939]), .B(n25096), .C(matrixInput[931]), 
        .D(n25081), .Z(n26325) );
    VMW_AO22 U2049 ( .A(matrixInput[1404]), .B(n25096), .C(matrixInput[1396]), 
        .D(n25081), .Z(n25860) );
    VMW_AO22 U368 ( .A(vectorInput[12]), .B(n25095), .C(vectorInput[4]), .D(
        n25080), .Z(n27380) );
    VMW_AO22 U579 ( .A(matrixInput[884]), .B(n25096), .C(matrixInput[876]), 
        .D(n25081), .Z(n26380) );
    VMW_AO22 U627 ( .A(matrixInput[840]), .B(n25096), .C(matrixInput[832]), 
        .D(n25081), .Z(n26424) );
    VMW_AO22 U1079 ( .A(matrixInput[433]), .B(n25096), .C(matrixInput[425]), 
        .D(n25081), .Z(n26831) );
    VMW_AO22 U1668 ( .A(matrixInput[1747]), .B(n25096), .C(matrixInput[1739]), 
        .D(n25081), .Z(n25517) );
    VMW_AO22 U2379 ( .A(matrixInput[1107]), .B(n25096), .C(matrixInput[1099]), 
        .D(n25081), .Z(n26157) );
    VMW_FD \matrixInput_reg[1854]  ( .D(n25402), .CP(Clk), .Q(matrixInput
        [1854]) );
    VMW_FD \vectorInput_reg[127]  ( .D(n27257), .CP(Clk), .Q(vectorInput[127])
         );
    VMW_AO22 U1349 ( .A(matrixInput[2033]), .B(n25096), .C(matrixInput[2025]), 
        .D(n25081), .Z(n25231) );
    VMW_AO22 U1558 ( .A(matrixInput[1846]), .B(n25096), .C(matrixInput[1838]), 
        .D(n25081), .Z(n25418) );
    VMW_OAI21 U2568 ( .A(n25110), .B(n25111), .C(n25091), .Z(n25116) );
    VMW_FD \matrixInput_reg[1867]  ( .D(n25389), .CP(Clk), .Q(matrixInput
        [1867]) );
    VMW_FD \matrixInput_reg[1375]  ( .D(n25881), .CP(Clk), .Q(matrixInput
        [1375]) );
    VMW_FD \vectorInput_reg[97]  ( .D(n27287), .CP(Clk), .Q(vectorInput[97])
         );
    VMW_BUFIZ U2636 ( .A(n25206), .E(RD), .Z(\DataOut[18]1 ) );
    VMW_FD \matrixInput_reg[562]  ( .D(n26694), .CP(Clk), .Q(matrixInput[562])
         );
    VMW_AO22 U649 ( .A(matrixInput[820]), .B(n25096), .C(matrixInput[812]), 
        .D(n25081), .Z(n26444) );
    VMW_AO22 U1017 ( .A(matrixInput[489]), .B(n25096), .C(matrixInput[481]), 
        .D(n25081), .Z(n26775) );
    VMW_AO22 U1796 ( .A(matrixInput[1631]), .B(n25096), .C(matrixInput[1623]), 
        .D(n25081), .Z(n25633) );
    VMW_AO22 U2027 ( .A(matrixInput[1423]), .B(n25096), .C(matrixInput[1415]), 
        .D(n25081), .Z(n25841) );
    VMW_FD \matrixInput_reg[1076]  ( .D(n26180), .CP(Clk), .Q(matrixInput
        [1076]) );
    VMW_FD \matrixInput_reg[661]  ( .D(n26595), .CP(Clk), .Q(matrixInput[661])
         );
    VMW_AO22 U1187 ( .A(matrixInput[336]), .B(n25096), .C(matrixInput[328]), 
        .D(n25081), .Z(n26928) );
    VMW_AO22 U1606 ( .A(matrixInput[1803]), .B(n25096), .C(matrixInput[1795]), 
        .D(n25081), .Z(n25461) );
    VMW_FD \matrixInput_reg[678]  ( .D(n26578), .CP(Clk), .Q(matrixInput[678])
         );
    VMW_AO22 U2287 ( .A(matrixInput[1189]), .B(n25096), .C(matrixInput[1181]), 
        .D(n25081), .Z(n26075) );
    VMW_FD \matrixInput_reg[548]  ( .D(n26708), .CP(Clk), .Q(matrixInput[548])
         );
    VMW_AO22 U810 ( .A(matrixInput[676]), .B(n25096), .C(matrixInput[668]), 
        .D(n25081), .Z(n26588) );
    VMW_AO22 U980 ( .A(matrixInput[522]), .B(n25096), .C(matrixInput[514]), 
        .D(n25081), .Z(n26742) );
    VMW_AO22 U1030 ( .A(matrixInput[54]), .B(n25096), .C(matrixInput[46]), .D(
        n25081), .Z(n27210) );
    VMW_AO22 U1290 ( .A(matrixInput[243]), .B(n25096), .C(matrixInput[235]), 
        .D(n25081), .Z(n27021) );
    VMW_AO22 U1327 ( .A(DataIn[5]), .B(n25096), .C(matrixInput[2045]), .D(
        n25081), .Z(n25211) );
    VMW_AO22 U2317 ( .A(matrixInput[1162]), .B(n25096), .C(matrixInput[1154]), 
        .D(n25081), .Z(n26102) );
    VMW_AND3 U2506 ( .A(n25116), .B(n25117), .C(n25118), .Z(n25076) );
    VMW_AO22 U2496 ( .A(cOutput[127]), .B(n25089), .C(cOutput[111]), .D(n25088
        ), .Z(n25104) );
    VMW_FD \matrixInput_reg[551]  ( .D(n26705), .CP(Clk), .Q(matrixInput[551])
         );
    VMW_FD \matrixInput_reg[1346]  ( .D(n25910), .CP(Clk), .Q(matrixInput
        [1346]) );
    VMW_AO22 U1536 ( .A(matrixInput[1866]), .B(n25096), .C(matrixInput[1858]), 
        .D(n25081), .Z(n25398) );
    VMW_FD \matrixInput_reg[652]  ( .D(n26604), .CP(Clk), .Q(matrixInput[652])
         );
    VMW_AO22 U1944 ( .A(matrixInput[1498]), .B(n25096), .C(matrixInput[1490]), 
        .D(n25081), .Z(n25766) );
    VMW_FD \matrixInput_reg[1045]  ( .D(n26211), .CP(Clk), .Q(matrixInput
        [1045]) );
    VMW_AO22 U2330 ( .A(matrixInput[1150]), .B(n25096), .C(matrixInput[1142]), 
        .D(n25081), .Z(n26114) );
    VMW_FD \matrixInput_reg[2006]  ( .D(n25250), .CP(Clk), .Q(matrixInput
        [2006]) );
    VMW_FD \matrixInput_reg[1562]  ( .D(n25694), .CP(Clk), .Q(matrixInput
        [1562]) );
    VMW_FD \matrixInput_reg[375]  ( .D(n26881), .CP(Clk), .Q(matrixInput[375])
         );
    VMW_AO22 U2521 ( .A(cOutput[92]), .B(n25089), .C(cOutput[76]), .D(n25088), 
        .Z(n25135) );
    VMW_AO22 U1300 ( .A(matrixInput[234]), .B(n25096), .C(matrixInput[226]), 
        .D(n25081), .Z(n27030) );
    VMW_AO22 U1511 ( .A(matrixInput[1888]), .B(n25096), .C(matrixInput[1880]), 
        .D(n25081), .Z(n25376) );
    VMW_AO22 U1481 ( .A(matrixInput[1915]), .B(n25096), .C(matrixInput[1907]), 
        .D(n25081), .Z(n25349) );
    VMW_AO22 U1621 ( .A(matrixInput[1789]), .B(n25096), .C(matrixInput[1781]), 
        .D(n25081), .Z(n25475) );
    VMW_AO22 U1963 ( .A(matrixInput[1481]), .B(n25096), .C(matrixInput[1473]), 
        .D(n25081), .Z(n25783) );
    VMW_FD \matrixInput_reg[1678]  ( .D(n25578), .CP(Clk), .Q(matrixInput
        [1678]) );
    VMW_FD \matrixInput_reg[1661]  ( .D(n25595), .CP(Clk), .Q(matrixInput
        [1661]) );
    VMW_AO22 U2000 ( .A(matrixInput[151]), .B(n25096), .C(matrixInput[143]), 
        .D(n25081), .Z(n27113) );
    VMW_AO22 U2190 ( .A(matrixInput[1277]), .B(n25096), .C(matrixInput[1269]), 
        .D(n25081), .Z(n25987) );
    VMW_BUFIZ U2611 ( .A(n25188), .E(RD), .Z(\DataOut[10]1 ) );
    VMW_FD \matrixInput_reg[2035]  ( .D(n25221), .CP(Clk), .Q(matrixInput
        [2035]) );
    VMW_FD \matrixInput_reg[1652]  ( .D(n25604), .CP(Clk), .Q(matrixInput
        [1652]) );
    VMW_FD \matrixInput_reg[1551]  ( .D(n25705), .CP(Clk), .Q(matrixInput
        [1551]) );
    VMW_FD \matrixInput_reg[1548]  ( .D(n25708), .CP(Clk), .Q(matrixInput
        [1548]) );
    VMW_FD \matrixInput_reg[346]  ( .D(n26910), .CP(Clk), .Q(matrixInput[346])
         );
    VMW_FD \matrixInput_reg[1925]  ( .D(n25331), .CP(Clk), .Q(matrixInput
        [1925]) );
    VMW_FD \matrixInput_reg[6]  ( .D(n27250), .CP(Clk), .Q(matrixInput[6]) );
    VMW_AO22 U445 ( .A(matrixInput[1005]), .B(n25096), .C(matrixInput[997]), 
        .D(n25081), .Z(n26259) );
    VMW_AO22 U462 ( .A(matrixInput[989]), .B(n25096), .C(matrixInput[981]), 
        .D(n25081), .Z(n26275) );
    VMW_AO22 U752 ( .A(matrixInput[79]), .B(n25096), .C(matrixInput[71]), .D(
        n25081), .Z(n27185) );
    VMW_FD \matrixInput_reg[886]  ( .D(n26370), .CP(Clk), .Q(matrixInput[886])
         );
    VMW_AO22 U775 ( .A(matrixInput[77]), .B(n25096), .C(matrixInput[69]), .D(
        n25081), .Z(n27187) );
    VMW_AO22 U1878 ( .A(matrixInput[162]), .B(n25096), .C(matrixInput[154]), 
        .D(n25081), .Z(n27102) );
    VMW_FD \matrixInput_reg[1916]  ( .D(n25340), .CP(Clk), .Q(matrixInput
        [1916]) );
    VMW_FD \vectorInput_reg[45]  ( .D(n27339), .CP(Clk), .Q(vectorInput[45])
         );
    VMW_AO22 U837 ( .A(matrixInput[651]), .B(n25096), .C(matrixInput[643]), 
        .D(n25081), .Z(n26613) );
    VMW_FD \matrixInput_reg[1886]  ( .D(n25370), .CP(Clk), .Q(matrixInput
        [1886]) );
    VMW_FD \matrixInput_reg[925]  ( .D(n26331), .CP(Clk), .Q(matrixInput[925])
         );
    VMW_FD \vectorInput_reg[76]  ( .D(n27308), .CP(Clk), .Q(vectorInput[76])
         );
    VMW_FD \matrixInput_reg[916]  ( .D(n26340), .CP(Clk), .Q(matrixInput[916])
         );
    VMW_AO22 U749 ( .A(matrixInput[730]), .B(n25096), .C(matrixInput[722]), 
        .D(n25081), .Z(n26534) );
    VMW_AO22 U1130 ( .A(matrixInput[45]), .B(n25096), .C(matrixInput[37]), .D(
        n25081), .Z(n27219) );
    VMW_AO22 U2090 ( .A(matrixInput[1367]), .B(n25096), .C(matrixInput[1359]), 
        .D(n25081), .Z(n25897) );
    VMW_FD \matrixInput_reg[2025]  ( .D(n25231), .CP(Clk), .Q(matrixInput
        [2025]) );
    VMW_AO22 U2100 ( .A(matrixInput[142]), .B(n25096), .C(matrixInput[134]), 
        .D(n25081), .Z(n27122) );
    VMW_FD \matrixInput_reg[1642]  ( .D(n25614), .CP(Clk), .Q(matrixInput
        [1642]) );
    VMW_FD \matrixInput_reg[1558]  ( .D(n25698), .CP(Clk), .Q(matrixInput
        [1558]) );
    VMW_FD \matrixInput_reg[1541]  ( .D(n25715), .CP(Clk), .Q(matrixInput
        [1541]) );
    VMW_FD \matrixInput_reg[356]  ( .D(n26900), .CP(Clk), .Q(matrixInput[356])
         );
    VMW_AO22 U1200 ( .A(matrixInput[324]), .B(n25096), .C(matrixInput[316]), 
        .D(n25081), .Z(n26940) );
    VMW_AO22 U1721 ( .A(matrixInput[1699]), .B(n25096), .C(matrixInput[1691]), 
        .D(n25081), .Z(n25565) );
    VMW_AO22 U2230 ( .A(matrixInput[1240]), .B(n25096), .C(matrixInput[1232]), 
        .D(n25081), .Z(n26024) );
    VMW_AO22 U2421 ( .A(matrixInput[1068]), .B(n25096), .C(matrixInput[1060]), 
        .D(n25081), .Z(n26196) );
    VMW_FD \matrixInput_reg[1572]  ( .D(n25684), .CP(Clk), .Q(matrixInput
        [1572]) );
    VMW_FD \matrixInput_reg[365]  ( .D(n26891), .CP(Clk), .Q(matrixInput[365])
         );
    VMW_FD \matrixInput_reg[2016]  ( .D(n25240), .CP(Clk), .Q(matrixInput
        [2016]) );
    VMW_AO22 U1390 ( .A(matrixInput[206]), .B(n25096), .C(matrixInput[198]), 
        .D(n25081), .Z(n27058) );
    VMW_AO22 U1581 ( .A(matrixInput[1825]), .B(n25096), .C(matrixInput[1817]), 
        .D(n25081), .Z(n25439) );
    VMW_AO22 U1411 ( .A(matrixInput[1978]), .B(n25096), .C(matrixInput[1970]), 
        .D(n25081), .Z(n25286) );
    VMW_AO22 U1863 ( .A(matrixInput[1571]), .B(n25096), .C(matrixInput[1563]), 
        .D(n25081), .Z(n25693) );
    VMW_AO22 U2217 ( .A(matrixInput[1252]), .B(n25096), .C(matrixInput[1244]), 
        .D(n25081), .Z(n26012) );
    VMW_FD \matrixInput_reg[1671]  ( .D(n25585), .CP(Clk), .Q(matrixInput
        [1671]) );
    VMW_FD \matrixInput_reg[1668]  ( .D(n25588), .CP(Clk), .Q(matrixInput
        [1668]) );
    VMW_FD \matrixInput_reg[1356]  ( .D(n25900), .CP(Clk), .Q(matrixInput
        [1356]) );
    VMW_AO22 U2387 ( .A(matrixInput[1099]), .B(n25096), .C(matrixInput[1091]), 
        .D(n25081), .Z(n26165) );
    VMW_INV U2596 ( .A(n25081), .Z(n25096) );
    VMW_FD \matrixInput_reg[541]  ( .D(n26715), .CP(Clk), .Q(matrixInput[541])
         );
    VMW_AO22 U1227 ( .A(matrixInput[300]), .B(n25096), .C(matrixInput[292]), 
        .D(n25081), .Z(n26964) );
    VMW_AO22 U1436 ( .A(matrixInput[1956]), .B(n25096), .C(matrixInput[1948]), 
        .D(n25081), .Z(n25308) );
    VMW_AO22 U2406 ( .A(matrixInput[1082]), .B(n25096), .C(matrixInput[1074]), 
        .D(n25081), .Z(n26182) );
    VMW_FD \matrixInput_reg[558]  ( .D(n26698), .CP(Clk), .Q(matrixInput[558])
         );
    VMW_FD \matrixInput_reg[1055]  ( .D(n26201), .CP(Clk), .Q(matrixInput
        [1055]) );
    VMW_AO22 U1844 ( .A(matrixInput[1588]), .B(n25096), .C(matrixInput[1580]), 
        .D(n25081), .Z(n25676) );
    VMW_FD \matrixInput_reg[642]  ( .D(n26614), .CP(Clk), .Q(matrixInput[642])
         );
    VMW_FD \matrixInput_reg[572]  ( .D(n26684), .CP(Clk), .Q(matrixInput[572])
         );
    VMW_PULLDOWN U284 ( .Z(n25202) );
    VMW_AO22 U328 ( .A(vectorInput[94]), .B(n25095), .C(vectorInput[86]), .D(
        n25080), .Z(n27298) );
    VMW_AO22 U354 ( .A(vectorInput[70]), .B(n25095), .C(vectorInput[62]), .D(
        n25080), .Z(n27322) );
    VMW_AO22 U479 ( .A(matrixInput[974]), .B(n25096), .C(matrixInput[966]), 
        .D(n25081), .Z(n26290) );
    VMW_AO22 U2127 ( .A(matrixInput[1333]), .B(n25096), .C(matrixInput[1325]), 
        .D(n25081), .Z(n25931) );
    VMW_AO22 U937 ( .A(matrixInput[561]), .B(n25096), .C(matrixInput[553]), 
        .D(n25081), .Z(n26703) );
    VMW_AO22 U1087 ( .A(matrixInput[426]), .B(n25096), .C(matrixInput[418]), 
        .D(n25081), .Z(n26838) );
    VMW_AO22 U1706 ( .A(matrixInput[1712]), .B(n25096), .C(matrixInput[1704]), 
        .D(n25081), .Z(n25552) );
    VMW_FD \matrixInput_reg[1365]  ( .D(n25891), .CP(Clk), .Q(matrixInput
        [1365]) );
    VMW_FD \matrixInput_reg[668]  ( .D(n26588), .CP(Clk), .Q(matrixInput[668])
         );
    VMW_AO22 U1117 ( .A(matrixInput[399]), .B(n25096), .C(matrixInput[391]), 
        .D(n25081), .Z(n26865) );
    VMW_AO22 U1696 ( .A(matrixInput[1721]), .B(n25096), .C(matrixInput[1713]), 
        .D(n25081), .Z(n25543) );
    VMW_FD \matrixInput_reg[671]  ( .D(n26585), .CP(Clk), .Q(matrixInput[671])
         );
    VMW_FD \matrixInput_reg[1896]  ( .D(n25360), .CP(Clk), .Q(matrixInput
        [1896]) );
    VMW_FD \matrixInput_reg[1066]  ( .D(n26190), .CP(Clk), .Q(matrixInput
        [1066]) );
    VMW_FD \matrixInput_reg[906]  ( .D(n26350), .CP(Clk), .Q(matrixInput[906])
         );
    VMW_FD \vectorInput_reg[66]  ( .D(n27318), .CP(Clk), .Q(vectorInput[66])
         );
    VMW_AO22 U373 ( .A(vectorInput[53]), .B(n25095), .C(vectorInput[45]), .D(
        n25080), .Z(n27339) );
    VMW_AO22 U545 ( .A(matrixInput[914]), .B(n25096), .C(matrixInput[906]), 
        .D(n25081), .Z(n26350) );
    VMW_AO22 U562 ( .A(matrixInput[899]), .B(n25096), .C(matrixInput[891]), 
        .D(n25081), .Z(n26365) );
    VMW_AO22 U652 ( .A(matrixInput[88]), .B(n25096), .C(matrixInput[80]), .D(
        n25081), .Z(n27176) );
    VMW_AO22 U675 ( .A(matrixInput[86]), .B(n25096), .C(matrixInput[78]), .D(
        n25081), .Z(n27178) );
    VMW_AO22 U1978 ( .A(matrixInput[153]), .B(n25096), .C(matrixInput[145]), 
        .D(n25081), .Z(n27111) );
    VMW_FD \vectorInput_reg[55]  ( .D(n27329), .CP(Clk), .Q(vectorInput[55])
         );
    VMW_FD \matrixInput_reg[1906]  ( .D(n25350), .CP(Clk), .Q(matrixInput
        [1906]) );
    VMW_FD \matrixInput_reg[935]  ( .D(n26321), .CP(Clk), .Q(matrixInput[935])
         );
    VMW_FD \matrixInput_reg[896]  ( .D(n26360), .CP(Clk), .Q(matrixInput[896])
         );
    VMW_AO22 U880 ( .A(matrixInput[612]), .B(n25096), .C(matrixInput[604]), 
        .D(n25081), .Z(n26652) );
    VMW_AO22 U910 ( .A(matrixInput[586]), .B(n25096), .C(matrixInput[578]), 
        .D(n25081), .Z(n26678) );
    VMW_AO22 U384 ( .A(vectorInput[43]), .B(n25095), .C(vectorInput[35]), .D(
        n25080), .Z(n27349) );
    VMW_AO22 U396 ( .A(vectorInput[32]), .B(n25095), .C(vectorInput[24]), .D(
        n25080), .Z(n27360) );
    VMW_AO22 U417 ( .A(DataIn[0]), .B(n25095), .C(vectorInput[120]), .D(n25080
        ), .Z(n27264) );
    VMW_AO22 U727 ( .A(matrixInput[750]), .B(n25096), .C(matrixInput[742]), 
        .D(n25081), .Z(n26514) );
    VMW_AO22 U959 ( .A(matrixInput[541]), .B(n25096), .C(matrixInput[533]), 
        .D(n25081), .Z(n26723) );
    VMW_AO22 U1045 ( .A(matrixInput[464]), .B(n25096), .C(matrixInput[456]), 
        .D(n25081), .Z(n26800) );
    VMW_AO22 U1062 ( .A(matrixInput[448]), .B(n25096), .C(matrixInput[440]), 
        .D(n25081), .Z(n26816) );
    VMW_AO22 U1352 ( .A(matrixInput[2030]), .B(n25096), .C(matrixInput[2022]), 
        .D(n25081), .Z(n25234) );
    VMW_AO22 U1543 ( .A(matrixInput[1859]), .B(n25096), .C(matrixInput[1851]), 
        .D(n25081), .Z(n25405) );
    VMW_FD \matrixInput_reg[1935]  ( .D(n25321), .CP(Clk), .Q(matrixInput
        [1935]) );
    VMW_AO22 U1673 ( .A(matrixInput[1742]), .B(n25096), .C(matrixInput[1734]), 
        .D(n25081), .Z(n25522) );
    VMW_AO22 U1931 ( .A(matrixInput[1509]), .B(n25096), .C(matrixInput[1501]), 
        .D(n25081), .Z(n25755) );
    VMW_FD \matrixInput_reg[430]  ( .D(n26826), .CP(Clk), .Q(matrixInput[430])
         );
    VMW_FD \matrixInput_reg[429]  ( .D(n26827), .CP(Clk), .Q(matrixInput[429])
         );
    VMW_AO22 U2362 ( .A(matrixInput[1121]), .B(n25096), .C(matrixInput[1113]), 
        .D(n25081), .Z(n26143) );
    VMW_FD \matrixInput_reg[1227]  ( .D(n26029), .CP(Clk), .Q(matrixInput
        [1227]) );
    VMW_FD \matrixInput_reg[1124]  ( .D(n26132), .CP(Clk), .Q(matrixInput
        [1124]) );
    VMW_FD \matrixInput_reg[733]  ( .D(n26523), .CP(Clk), .Q(matrixInput[733])
         );
    VMW_FD \vectorInput_reg[9]  ( .D(n27375), .CP(Clk), .Q(vectorInput[9]) );
    VMW_OAI21 U2573 ( .A(n25123), .B(n25124), .C(n25093), .Z(n25129) );
    VMW_FD \matrixInput_reg[1214]  ( .D(n26042), .CP(Clk), .Q(matrixInput
        [1214]) );
    VMW_FD \matrixInput_reg[403]  ( .D(n26853), .CP(Clk), .Q(matrixInput[403])
         );
    VMW_AO22 U2052 ( .A(matrixInput[1401]), .B(n25096), .C(matrixInput[1393]), 
        .D(n25081), .Z(n25863) );
    VMW_FD \matrixInput_reg[1690]  ( .D(n25566), .CP(Clk), .Q(matrixInput
        [1690]) );
    VMW_FD \matrixInput_reg[1689]  ( .D(n25567), .CP(Clk), .Q(matrixInput
        [1689]) );
    VMW_FD \matrixInput_reg[1593]  ( .D(n25663), .CP(Clk), .Q(matrixInput
        [1593]) );
    VMW_FD \matrixInput_reg[384]  ( .D(n26872), .CP(Clk), .Q(matrixInput[384])
         );
    VMW_FD \matrixInput_reg[1429]  ( .D(n25827), .CP(Clk), .Q(matrixInput
        [1429]) );
    VMW_FD \matrixInput_reg[1117]  ( .D(n26139), .CP(Clk), .Q(matrixInput
        [1117]) );
    VMW_FD \matrixInput_reg[719]  ( .D(n26537), .CP(Clk), .Q(matrixInput[719])
         );
    VMW_FD \matrixInput_reg[700]  ( .D(n26556), .CP(Clk), .Q(matrixInput[700])
         );
    VMW_FD \matrixInput_reg[227]  ( .D(n27029), .CP(Clk), .Q(matrixInput[227])
         );
    VMW_AO22 U1654 ( .A(matrixInput[1759]), .B(n25096), .C(matrixInput[1751]), 
        .D(n25081), .Z(n25505) );
    VMW_FD \matrixInput_reg[1430]  ( .D(n25826), .CP(Clk), .Q(matrixInput
        [1430]) );
    VMW_AO22 U2075 ( .A(matrixInput[1380]), .B(n25096), .C(matrixInput[1372]), 
        .D(n25081), .Z(n25884) );
    VMW_FD \matrixInput_reg[1733]  ( .D(n25523), .CP(Clk), .Q(matrixInput
        [1733]) );
    VMW_FD \matrixInput_reg[124]  ( .D(n27132), .CP(Clk), .Q(matrixInput[124])
         );
    VMW_AO22 U1375 ( .A(matrixInput[2009]), .B(n25096), .C(matrixInput[2001]), 
        .D(n25081), .Z(n25255) );
    VMW_AO22 U1564 ( .A(matrixInput[1840]), .B(n25096), .C(matrixInput[1832]), 
        .D(n25081), .Z(n25424) );
    VMW_FD \matrixInput_reg[1403]  ( .D(n25853), .CP(Clk), .Q(matrixInput
        [1403]) );
    VMW_AO22 U1886 ( .A(matrixInput[1550]), .B(n25096), .C(matrixInput[1542]), 
        .D(n25081), .Z(n25714) );
    VMW_FD \matrixInput_reg[214]  ( .D(n27042), .CP(Clk), .Q(matrixInput[214])
         );
    VMW_AO22 U1916 ( .A(matrixInput[1523]), .B(n25096), .C(matrixInput[1515]), 
        .D(n25081), .Z(n25741) );
    VMW_FD \matrixInput_reg[690]  ( .D(n26566), .CP(Clk), .Q(matrixInput[690])
         );
    VMW_AO22 U2345 ( .A(matrixInput[1137]), .B(n25096), .C(matrixInput[1129]), 
        .D(n25081), .Z(n26127) );
    VMW_AO22 U2554 ( .A(cOutput[48]), .B(n25087), .C(cOutput[32]), .D(n25084), 
        .Z(n25176) );
    VMW_FD \matrixInput_reg[1384]  ( .D(n25872), .CP(Clk), .Q(matrixInput
        [1384]) );
    VMW_FD \matrixInput_reg[1087]  ( .D(n26169), .CP(Clk), .Q(matrixInput
        [1087]) );
    VMW_FD \matrixInput_reg[689]  ( .D(n26567), .CP(Clk), .Q(matrixInput[689])
         );
    VMW_FD \matrixInput_reg[593]  ( .D(n26663), .CP(Clk), .Q(matrixInput[593])
         );
    VMW_FD \matrixInput_reg[1700]  ( .D(n25556), .CP(Clk), .Q(matrixInput
        [1700]) );
    VMW_FD \matrixInput_reg[1719]  ( .D(n25537), .CP(Clk), .Q(matrixInput
        [1719]) );
    VMW_FD \matrixInput_reg[117]  ( .D(n27139), .CP(Clk), .Q(matrixInput[117])
         );
    VMW_AO22 U865 ( .A(matrixInput[626]), .B(n25096), .C(matrixInput[618]), 
        .D(n25081), .Z(n26638) );
    VMW_AO22 U1249 ( .A(matrixInput[280]), .B(n25096), .C(matrixInput[272]), 
        .D(n25081), .Z(n26984) );
    VMW_AO22 U2279 ( .A(matrixInput[1197]), .B(n25096), .C(matrixInput[1189]), 
        .D(n25081), .Z(n26067) );
    VMW_AO22 U2468 ( .A(matrixInput[1026]), .B(n25096), .C(matrixInput[1018]), 
        .D(n25081), .Z(n26238) );
    VMW_FD \matrixInput_reg[1877]  ( .D(n25379), .CP(Clk), .Q(matrixInput
        [1877]) );
    VMW_FD \vectorInput_reg[87]  ( .D(n27297), .CP(Clk), .Q(vectorInput[87])
         );
    VMW_AO22 U1458 ( .A(matrixInput[1936]), .B(n25096), .C(matrixInput[1928]), 
        .D(n25081), .Z(n25328) );
    VMW_AO22 U405 ( .A(vectorInput[24]), .B(n25095), .C(vectorInput[16]), .D(
        n25080), .Z(n27368) );
    VMW_AO22 U430 ( .A(vectorInput[117]), .B(n25095), .C(vectorInput[109]), 
        .D(n25080), .Z(n27275) );
    VMW_AO22 U587 ( .A(matrixInput[877]), .B(n25096), .C(matrixInput[869]), 
        .D(n25081), .Z(n26387) );
    VMW_AO22 U842 ( .A(matrixInput[647]), .B(n25096), .C(matrixInput[639]), 
        .D(n25081), .Z(n26617) );
    VMW_AO22 U1179 ( .A(matrixInput[343]), .B(n25096), .C(matrixInput[335]), 
        .D(n25081), .Z(n26921) );
    VMW_AO22 U2149 ( .A(matrixInput[1313]), .B(n25096), .C(matrixInput[1305]), 
        .D(n25081), .Z(n25951) );
    VMW_FD \vectorInput_reg[104]  ( .D(n27280), .CP(Clk), .Q(vectorInput[104])
         );
    VMW_AO22 U1768 ( .A(matrixInput[1657]), .B(n25096), .C(matrixInput[1649]), 
        .D(n25081), .Z(n25607) );
    VMW_FD \matrixInput_reg[1844]  ( .D(n25412), .CP(Clk), .Q(matrixInput
        [1844]) );
    VMW_FD \matrixInput_reg[37]  ( .D(n27219), .CP(Clk), .Q(matrixInput[37])
         );
    VMW_AO22 U595 ( .A(matrixInput[869]), .B(n25096), .C(matrixInput[861]), 
        .D(n25081), .Z(n26395) );
    VMW_AO22 U690 ( .A(matrixInput[784]), .B(n25096), .C(matrixInput[776]), 
        .D(n25081), .Z(n26480) );
    VMW_FD \matrixInput_reg[877]  ( .D(n26379), .CP(Clk), .Q(matrixInput[877])
         );
    VMW_AO22 U700 ( .A(matrixInput[775]), .B(n25096), .C(matrixInput[767]), 
        .D(n25081), .Z(n26489) );
    VMW_AO22 U735 ( .A(matrixInput[743]), .B(n25096), .C(matrixInput[735]), 
        .D(n25081), .Z(n26521) );
    VMW_FD \matrixInput_reg[938]  ( .D(n26318), .CP(Clk), .Q(matrixInput[938])
         );
    VMW_FD \matrixInput_reg[921]  ( .D(n26335), .CP(Clk), .Q(matrixInput[921])
         );
    VMW_FD \matrixInput_reg[844]  ( .D(n26412), .CP(Clk), .Q(matrixInput[844])
         );
    VMW_AO22 U1838 ( .A(matrixInput[1594]), .B(n25096), .C(matrixInput[1586]), 
        .D(n25081), .Z(n25670) );
    VMW_FD \vectorInput_reg[58]  ( .D(n27326), .CP(Clk), .Q(vectorInput[58])
         );
    VMW_FD \vectorInput_reg[41]  ( .D(n27343), .CP(Clk), .Q(vectorInput[41])
         );
    VMW_AO22 U422 ( .A(vectorInput[124]), .B(n25095), .C(vectorInput[116]), 
        .D(n25080), .Z(n27268) );
    VMW_AO22 U877 ( .A(matrixInput[615]), .B(n25096), .C(matrixInput[607]), 
        .D(n25081), .Z(n26649) );
    VMW_FD \matrixInput_reg[912]  ( .D(n26344), .CP(Clk), .Q(matrixInput[912])
         );
    VMW_FD \matrixInput_reg[1882]  ( .D(n25374), .CP(Clk), .Q(matrixInput
        [1882]) );
    VMW_FD \vectorInput_reg[72]  ( .D(n27312), .CP(Clk), .Q(vectorInput[72])
         );
    VMW_AO22 U682 ( .A(matrixInput[791]), .B(n25096), .C(matrixInput[783]), 
        .D(n25081), .Z(n26473) );
    VMW_AO22 U712 ( .A(matrixInput[764]), .B(n25096), .C(matrixInput[756]), 
        .D(n25081), .Z(n26500) );
    VMW_AO22 U850 ( .A(matrixInput[639]), .B(n25096), .C(matrixInput[631]), 
        .D(n25081), .Z(n26625) );
    VMW_FD \matrixInput_reg[1938]  ( .D(n25318), .CP(Clk), .Q(matrixInput
        [1938]) );
    VMW_FD \matrixInput_reg[1921]  ( .D(n25335), .CP(Clk), .Q(matrixInput
        [1921]) );
    VMW_FD \matrixInput_reg[2]  ( .D(n27254), .CP(Clk), .Q(matrixInput[2]) );
    VMW_FD \matrixInput_reg[1912]  ( .D(n25344), .CP(Clk), .Q(matrixInput
        [1912]) );
    VMW_AO22 U1057 ( .A(matrixInput[453]), .B(n25096), .C(matrixInput[445]), 
        .D(n25081), .Z(n26811) );
    VMW_AO22 U1070 ( .A(matrixInput[441]), .B(n25096), .C(matrixInput[433]), 
        .D(n25081), .Z(n26823) );
    VMW_AO22 U1340 ( .A(matrixInput[2041]), .B(n25096), .C(matrixInput[2033]), 
        .D(n25081), .Z(n25223) );
    VMW_AO22 U1923 ( .A(matrixInput[1517]), .B(n25096), .C(matrixInput[1509]), 
        .D(n25081), .Z(n25747) );
    VMW_FD \matrixInput_reg[882]  ( .D(n26374), .CP(Clk), .Q(matrixInput[882])
         );
    VMW_FD \matrixInput_reg[1665]  ( .D(n25591), .CP(Clk), .Q(matrixInput
        [1665]) );
    VMW_AO22 U1551 ( .A(matrixInput[1852]), .B(n25096), .C(matrixInput[1844]), 
        .D(n25081), .Z(n25412) );
    VMW_AO22 U2370 ( .A(matrixInput[1114]), .B(n25096), .C(matrixInput[1106]), 
        .D(n25081), .Z(n26150) );
    VMW_NAND3 U2561 ( .A(n25085), .B(n25083), .C(WR), .Z(n25081) );
    VMW_FD \matrixInput_reg[2002]  ( .D(n25254), .CP(Clk), .Q(matrixInput
        [2002]) );
    VMW_FD \matrixInput_reg[1566]  ( .D(n25690), .CP(Clk), .Q(matrixInput
        [1566]) );
    VMW_FD \matrixInput_reg[371]  ( .D(n26885), .CP(Clk), .Q(matrixInput[371])
         );
    VMW_FD \matrixInput_reg[368]  ( .D(n26888), .CP(Clk), .Q(matrixInput[368])
         );
    VMW_AO22 U1646 ( .A(matrixInput[1767]), .B(n25096), .C(matrixInput[1759]), 
        .D(n25081), .Z(n25497) );
    VMW_AO22 U1661 ( .A(matrixInput[1753]), .B(n25096), .C(matrixInput[1745]), 
        .D(n25081), .Z(n25511) );
    VMW_AO22 U2040 ( .A(matrixInput[1411]), .B(n25096), .C(matrixInput[1403]), 
        .D(n25081), .Z(n25853) );
    VMW_FD \matrixInput_reg[2031]  ( .D(n25225), .CP(Clk), .Q(matrixInput
        [2031]) );
    VMW_FD \matrixInput_reg[1656]  ( .D(n25600), .CP(Clk), .Q(matrixInput
        [1656]) );
    VMW_FD \matrixInput_reg[1555]  ( .D(n25701), .CP(Clk), .Q(matrixInput
        [1555]) );
    VMW_FD \matrixInput_reg[342]  ( .D(n26914), .CP(Clk), .Q(matrixInput[342])
         );
    VMW_FD \matrixInput_reg[2028]  ( .D(n25228), .CP(Clk), .Q(matrixInput
        [2028]) );
    VMW_FD \matrixInput_reg[665]  ( .D(n26591), .CP(Clk), .Q(matrixInput[665])
         );
    VMW_FD \matrixInput_reg[1072]  ( .D(n26184), .CP(Clk), .Q(matrixInput
        [1072]) );
    VMW_FD \matrixInput_reg[566]  ( .D(n26690), .CP(Clk), .Q(matrixInput[566])
         );
    VMW_AO22 U333 ( .A(vectorInput[89]), .B(n25095), .C(vectorInput[81]), .D(
        n25080), .Z(n27303) );
    VMW_AO22 U346 ( .A(vectorInput[14]), .B(n25095), .C(vectorInput[6]), .D(
        n25080), .Z(n27378) );
    VMW_AO22 U539 ( .A(matrixInput[919]), .B(n25096), .C(matrixInput[911]), 
        .D(n25081), .Z(n26345) );
    VMW_AO22 U2067 ( .A(matrixInput[145]), .B(n25096), .C(matrixInput[137]), 
        .D(n25081), .Z(n27119) );
    VMW_AO22 U557 ( .A(matrixInput[904]), .B(n25096), .C(matrixInput[896]), 
        .D(n25081), .Z(n26360) );
    VMW_AO22 U609 ( .A(matrixInput[857]), .B(n25096), .C(matrixInput[849]), 
        .D(n25081), .Z(n26407) );
    VMW_AO22 U799 ( .A(matrixInput[686]), .B(n25096), .C(matrixInput[678]), 
        .D(n25081), .Z(n26578) );
    VMW_AO22 U1367 ( .A(matrixInput[2017]), .B(n25096), .C(matrixInput[2009]), 
        .D(n25081), .Z(n25247) );
    VMW_AO22 U1576 ( .A(matrixInput[1829]), .B(n25096), .C(matrixInput[1821]), 
        .D(n25081), .Z(n25435) );
    VMW_AO22 U1894 ( .A(matrixInput[1543]), .B(n25096), .C(matrixInput[1535]), 
        .D(n25081), .Z(n25721) );
    VMW_AO22 U1904 ( .A(matrixInput[1534]), .B(n25096), .C(matrixInput[1526]), 
        .D(n25081), .Z(n25730) );
    VMW_FD \matrixInput_reg[1371]  ( .D(n25885), .CP(Clk), .Q(matrixInput
        [1371]) );
    VMW_FD \matrixInput_reg[1368]  ( .D(n25888), .CP(Clk), .Q(matrixInput
        [1368]) );
    VMW_FD \matrixInput_reg[1058]  ( .D(n26198), .CP(Clk), .Q(matrixInput
        [1058]) );
    VMW_FD \matrixInput_reg[1041]  ( .D(n26215), .CP(Clk), .Q(matrixInput
        [1041]) );
    VMW_AO22 U2357 ( .A(matrixInput[1126]), .B(n25096), .C(matrixInput[1118]), 
        .D(n25081), .Z(n26138) );
    VMW_FD \matrixInput_reg[1342]  ( .D(n25914), .CP(Clk), .Q(matrixInput
        [1342]) );
    VMW_FD \matrixInput_reg[656]  ( .D(n26600), .CP(Clk), .Q(matrixInput[656])
         );
    VMW_FD \matrixInput_reg[555]  ( .D(n26701), .CP(Clk), .Q(matrixInput[555])
         );
    VMW_AO22 U1039 ( .A(matrixInput[469]), .B(n25096), .C(matrixInput[461]), 
        .D(n25081), .Z(n26795) );
    VMW_AO22 U2546 ( .A(cOutput[57]), .B(n25089), .C(cOutput[41]), .D(n25088), 
        .Z(n25166) );
    VMW_FD \matrixInput_reg[1850]  ( .D(n25406), .CP(Clk), .Q(matrixInput
        [1850]) );
    VMW_FD \matrixInput_reg[1849]  ( .D(n25407), .CP(Clk), .Q(matrixInput
        [1849]) );
    VMW_AO22 U1628 ( .A(matrixInput[1783]), .B(n25096), .C(matrixInput[1775]), 
        .D(n25081), .Z(n25481) );
    VMW_AO22 U2199 ( .A(matrixInput[1268]), .B(n25096), .C(matrixInput[1260]), 
        .D(n25081), .Z(n25996) );
    VMW_BUFIZ U2618 ( .A(n25193), .E(RD), .Z(\DataOut[31] ) );
    VMW_FD \vectorInput_reg[109]  ( .D(n27275), .CP(Clk), .Q(vectorInput[109])
         );
    VMW_FD \vectorInput_reg[110]  ( .D(n27274), .CP(Clk), .Q(vectorInput[110])
         );
    VMW_AO22 U361 ( .A(vectorInput[64]), .B(n25095), .C(vectorInput[56]), .D(
        n25080), .Z(n27328) );
    VMW_AO22 U640 ( .A(matrixInput[828]), .B(n25096), .C(matrixInput[820]), 
        .D(n25081), .Z(n26436) );
    VMW_AO22 U667 ( .A(matrixInput[805]), .B(n25096), .C(matrixInput[797]), 
        .D(n25081), .Z(n26459) );
    VMW_AO22 U925 ( .A(matrixInput[572]), .B(n25096), .C(matrixInput[564]), 
        .D(n25081), .Z(n26692) );
    VMW_AO22 U2009 ( .A(matrixInput[1439]), .B(n25096), .C(matrixInput[1431]), 
        .D(n25081), .Z(n25825) );
    VMW_AO22 U1299 ( .A(matrixInput[235]), .B(n25096), .C(matrixInput[227]), 
        .D(n25081), .Z(n27029) );
    VMW_AO22 U1309 ( .A(matrixInput[226]), .B(n25096), .C(matrixInput[218]), 
        .D(n25081), .Z(n27038) );
    VMW_FD \vectorInput_reg[93]  ( .D(n27291), .CP(Clk), .Q(vectorInput[93])
         );
    VMW_AO22 U1488 ( .A(matrixInput[1908]), .B(n25096), .C(matrixInput[1900]), 
        .D(n25081), .Z(n25356) );
    VMW_AO22 U1518 ( .A(matrixInput[1882]), .B(n25096), .C(matrixInput[1874]), 
        .D(n25081), .Z(n25382) );
    VMW_FD \matrixInput_reg[1863]  ( .D(n25393), .CP(Clk), .Q(matrixInput
        [1863]) );
    VMW_AO22 U2339 ( .A(matrixInput[1142]), .B(n25096), .C(matrixInput[1134]), 
        .D(n25081), .Z(n26122) );
    VMW_AO22 U2528 ( .A(cOutput[59]), .B(n25089), .C(cOutput[43]), .D(n25088), 
        .Z(n25144) );
    VMW_FD \matrixInput_reg[850]  ( .D(n26406), .CP(Clk), .Q(matrixInput[850])
         );
    VMW_FD \matrixInput_reg[849]  ( .D(n26407), .CP(Clk), .Q(matrixInput[849])
         );
    VMW_FD \vectorInput_reg[123]  ( .D(n27261), .CP(Clk), .Q(vectorInput[123])
         );
    VMW_FD \matrixInput_reg[10]  ( .D(n27246), .CP(Clk), .Q(matrixInput[10])
         );
    VMW_FD \matrixInput_reg[863]  ( .D(n26393), .CP(Clk), .Q(matrixInput[863])
         );
    VMW_AO22 U457 ( .A(matrixInput[994]), .B(n25096), .C(matrixInput[986]), 
        .D(n25081), .Z(n26270) );
    VMW_AO22 U470 ( .A(matrixInput[982]), .B(n25096), .C(matrixInput[974]), 
        .D(n25081), .Z(n26282) );
    VMW_AO22 U570 ( .A(matrixInput[892]), .B(n25096), .C(matrixInput[884]), 
        .D(n25081), .Z(n26372) );
    VMW_AO22 U819 ( .A(matrixInput[73]), .B(n25096), .C(matrixInput[65]), .D(
        n25081), .Z(n27191) );
    VMW_AO22 U892 ( .A(matrixInput[602]), .B(n25096), .C(matrixInput[594]), 
        .D(n25081), .Z(n26662) );
    VMW_FD \matrixInput_reg[23]  ( .D(n27233), .CP(Clk), .Q(matrixInput[23])
         );
    VMW_AO22 U902 ( .A(matrixInput[593]), .B(n25096), .C(matrixInput[585]), 
        .D(n25081), .Z(n26671) );
    VMW_AO22 U1122 ( .A(matrixInput[395]), .B(n25096), .C(matrixInput[387]), 
        .D(n25081), .Z(n26869) );
    VMW_AO22 U1733 ( .A(matrixInput[1688]), .B(n25096), .C(matrixInput[1680]), 
        .D(n25081), .Z(n25576) );
    VMW_AO22 U2082 ( .A(matrixInput[1374]), .B(n25096), .C(matrixInput[1366]), 
        .D(n25081), .Z(n25890) );
    VMW_AO22 U2112 ( .A(matrixInput[1347]), .B(n25096), .C(matrixInput[1339]), 
        .D(n25081), .Z(n25917) );
    VMW_FD \matrixInput_reg[1103]  ( .D(n26153), .CP(Clk), .Q(matrixInput
        [1103]) );
    VMW_FD \matrixInput_reg[714]  ( .D(n26542), .CP(Clk), .Q(matrixInput[714])
         );
    VMW_FD \matrixInput_reg[389]  ( .D(n26867), .CP(Clk), .Q(matrixInput[389])
         );
    VMW_FD \matrixInput_reg[390]  ( .D(n26866), .CP(Clk), .Q(matrixInput[390])
         );
    VMW_FD \matrixInput_reg[1587]  ( .D(n25669), .CP(Clk), .Q(matrixInput
        [1587]) );
    VMW_AO22 U1212 ( .A(matrixInput[313]), .B(n25096), .C(matrixInput[305]), 
        .D(n25081), .Z(n26951) );
    VMW_AO22 U1382 ( .A(matrixInput[2005]), .B(n25096), .C(matrixInput[1997]), 
        .D(n25081), .Z(n25259) );
    VMW_AO22 U1871 ( .A(matrixInput[1564]), .B(n25096), .C(matrixInput[1556]), 
        .D(n25081), .Z(n25700) );
    VMW_AO22 U2222 ( .A(matrixInput[131]), .B(n25096), .C(matrixInput[123]), 
        .D(n25081), .Z(n27133) );
    VMW_FD \matrixInput_reg[1684]  ( .D(n25572), .CP(Clk), .Q(matrixInput
        [1684]) );
    VMW_FD \matrixInput_reg[1219]  ( .D(n26037), .CP(Clk), .Q(matrixInput
        [1219]) );
    VMW_FD \matrixInput_reg[1200]  ( .D(n26056), .CP(Clk), .Q(matrixInput
        [1200]) );
    VMW_FD \matrixInput_reg[417]  ( .D(n26839), .CP(Clk), .Q(matrixInput[417])
         );
    VMW_AO22 U2433 ( .A(matrixInput[112]), .B(n25096), .C(matrixInput[104]), 
        .D(n25081), .Z(n27152) );
    VMW_FD \matrixInput_reg[1130]  ( .D(n26126), .CP(Clk), .Q(matrixInput
        [1130]) );
    VMW_FD \matrixInput_reg[727]  ( .D(n26529), .CP(Clk), .Q(matrixInput[727])
         );
    VMW_FD \vectorInput_reg[4]  ( .D(n27380), .CP(Clk), .Q(vectorInput[4]) );
    VMW_FD \matrixInput_reg[1129]  ( .D(n26127), .CP(Clk), .Q(matrixInput
        [1129]) );
    VMW_FD \matrixInput_reg[424]  ( .D(n26832), .CP(Clk), .Q(matrixInput[424])
         );
    VMW_FD \matrixInput_reg[1233]  ( .D(n26023), .CP(Clk), .Q(matrixInput
        [1233]) );
    VMW_AO22 U1403 ( .A(matrixInput[1986]), .B(n25096), .C(matrixInput[1978]), 
        .D(n25081), .Z(n25278) );
    VMW_AO22 U1235 ( .A(matrixInput[293]), .B(n25096), .C(matrixInput[285]), 
        .D(n25081), .Z(n26971) );
    VMW_AO22 U1593 ( .A(matrixInput[1814]), .B(n25096), .C(matrixInput[1806]), 
        .D(n25081), .Z(n25450) );
    VMW_AO22 U1856 ( .A(matrixInput[164]), .B(n25096), .C(matrixInput[156]), 
        .D(n25081), .Z(n27100) );
    VMW_AO22 U2205 ( .A(matrixInput[1263]), .B(n25096), .C(matrixInput[1255]), 
        .D(n25081), .Z(n26001) );
    VMW_AO22 U2395 ( .A(matrixInput[1092]), .B(n25096), .C(matrixInput[1084]), 
        .D(n25081), .Z(n26172) );
    VMW_AO22 U2414 ( .A(matrixInput[1075]), .B(n25096), .C(matrixInput[1067]), 
        .D(n25081), .Z(n26189) );
    VMW_FD \matrixInput_reg[1714]  ( .D(n25542), .CP(Clk), .Q(matrixInput
        [1714]) );
    VMW_OAI21 U2584 ( .A(n25154), .B(n25155), .C(n25091), .Z(n25160) );
    VMW_FD \matrixInput_reg[1390]  ( .D(n25866), .CP(Clk), .Q(matrixInput
        [1390]) );
    VMW_FD \matrixInput_reg[1389]  ( .D(n25867), .CP(Clk), .Q(matrixInput
        [1389]) );
    VMW_FD \matrixInput_reg[587]  ( .D(n26669), .CP(Clk), .Q(matrixInput[587])
         );
    VMW_FD \matrixInput_reg[103]  ( .D(n27153), .CP(Clk), .Q(matrixInput[103])
         );
    VMW_FD \matrixInput_reg[684]  ( .D(n26572), .CP(Clk), .Q(matrixInput[684])
         );
    VMW_FD \matrixInput_reg[1093]  ( .D(n26163), .CP(Clk), .Q(matrixInput
        [1093]) );
    VMW_AO22 U1424 ( .A(matrixInput[1967]), .B(n25096), .C(matrixInput[1959]), 
        .D(n25081), .Z(n25297) );
    VMW_FD \matrixInput_reg[1417]  ( .D(n25839), .CP(Clk), .Q(matrixInput
        [1417]) );
    VMW_FD \matrixInput_reg[219]  ( .D(n27037), .CP(Clk), .Q(matrixInput[219])
         );
    VMW_FD \matrixInput_reg[200]  ( .D(n27056), .CP(Clk), .Q(matrixInput[200])
         );
    VMW_AO22 U989 ( .A(matrixInput[514]), .B(n25096), .C(matrixInput[506]), 
        .D(n25081), .Z(n26750) );
    VMW_AO22 U1095 ( .A(matrixInput[418]), .B(n25096), .C(matrixInput[410]), 
        .D(n25081), .Z(n26846) );
    VMW_AO22 U1105 ( .A(matrixInput[409]), .B(n25096), .C(matrixInput[401]), 
        .D(n25081), .Z(n26855) );
    VMW_AO22 U1684 ( .A(matrixInput[1732]), .B(n25096), .C(matrixInput[1724]), 
        .D(n25081), .Z(n25532) );
    VMW_AO22 U2135 ( .A(matrixInput[1326]), .B(n25096), .C(matrixInput[1318]), 
        .D(n25081), .Z(n25938) );
    VMW_FD \matrixInput_reg[1727]  ( .D(n25529), .CP(Clk), .Q(matrixInput
        [1727]) );
    VMW_FD \matrixInput_reg[130]  ( .D(n27126), .CP(Clk), .Q(matrixInput[130])
         );
    VMW_FD \matrixInput_reg[129]  ( .D(n27127), .CP(Clk), .Q(matrixInput[129])
         );
    VMW_FD \matrixInput_reg[233]  ( .D(n27023), .CP(Clk), .Q(matrixInput[233])
         );
    VMW_AO22 U1714 ( .A(matrixInput[1706]), .B(n25096), .C(matrixInput[1698]), 
        .D(n25081), .Z(n25558) );
    VMW_FD \matrixInput_reg[1424]  ( .D(n25832), .CP(Clk), .Q(matrixInput
        [1424]) );
    VMW_FD \matrixInput_reg[873]  ( .D(n26383), .CP(Clk), .Q(matrixInput[873])
         );
    VMW_AO22 U740 ( .A(matrixInput[738]), .B(n25096), .C(matrixInput[730]), 
        .D(n25081), .Z(n26526) );
    VMW_AO22 U802 ( .A(matrixInput[683]), .B(n25096), .C(matrixInput[675]), 
        .D(n25081), .Z(n26581) );
    VMW_AO22 U992 ( .A(matrixInput[511]), .B(n25096), .C(matrixInput[503]), 
        .D(n25081), .Z(n26753) );
    VMW_FD \matrixInput_reg[859]  ( .D(n26397), .CP(Clk), .Q(matrixInput[859])
         );
    VMW_FD \matrixInput_reg[840]  ( .D(n26416), .CP(Clk), .Q(matrixInput[840])
         );
    VMW_FD \matrixInput_reg[33]  ( .D(n27223), .CP(Clk), .Q(matrixInput[33])
         );
    VMW_FD \matrixInput_reg[19]  ( .D(n27237), .CP(Clk), .Q(matrixInput[19])
         );
    VMW_AO22 U767 ( .A(matrixInput[714]), .B(n25096), .C(matrixInput[706]), 
        .D(n25081), .Z(n26550) );
    VMW_AO22 U1209 ( .A(matrixInput[316]), .B(n25096), .C(matrixInput[308]), 
        .D(n25081), .Z(n26948) );
    VMW_AO22 U1399 ( .A(matrixInput[1989]), .B(n25096), .C(matrixInput[1981]), 
        .D(n25081), .Z(n25275) );
    VMW_AO22 U1418 ( .A(matrixInput[1972]), .B(n25096), .C(matrixInput[1964]), 
        .D(n25081), .Z(n25292) );
    VMW_AO22 U1588 ( .A(matrixInput[1818]), .B(n25096), .C(matrixInput[1810]), 
        .D(n25081), .Z(n25446) );
    VMW_AO22 U2239 ( .A(matrixInput[1232]), .B(n25096), .C(matrixInput[1224]), 
        .D(n25081), .Z(n26032) );
    VMW_FD \matrixInput_reg[1873]  ( .D(n25383), .CP(Clk), .Q(matrixInput
        [1873]) );
    VMW_FD \vectorInput_reg[83]  ( .D(n27301), .CP(Clk), .Q(vectorInput[83])
         );
    VMW_AO22 U1139 ( .A(matrixInput[379]), .B(n25096), .C(matrixInput[371]), 
        .D(n25081), .Z(n26885) );
    VMW_AO22 U1728 ( .A(matrixInput[1693]), .B(n25096), .C(matrixInput[1685]), 
        .D(n25081), .Z(n25571) );
    VMW_AO22 U2428 ( .A(matrixInput[1062]), .B(n25096), .C(matrixInput[1054]), 
        .D(n25081), .Z(n26202) );
    VMW_FD \matrixInput_reg[1859]  ( .D(n25397), .CP(Clk), .Q(matrixInput
        [1859]) );
    VMW_FD \matrixInput_reg[1840]  ( .D(n25416), .CP(Clk), .Q(matrixInput
        [1840]) );
    VMW_AO22 U2109 ( .A(matrixInput[1349]), .B(n25096), .C(matrixInput[1341]), 
        .D(n25081), .Z(n25915) );
    VMW_FD \vectorInput_reg[100]  ( .D(n27284), .CP(Clk), .Q(vectorInput[100])
         );
    VMW_AO22 U612 ( .A(matrixInput[854]), .B(n25096), .C(matrixInput[846]), 
        .D(n25081), .Z(n26410) );
    VMW_AO22 U782 ( .A(matrixInput[701]), .B(n25096), .C(matrixInput[693]), 
        .D(n25081), .Z(n26563) );
    VMW_AO22 U825 ( .A(matrixInput[662]), .B(n25096), .C(matrixInput[654]), 
        .D(n25081), .Z(n26602) );
    VMW_AO22 U2099 ( .A(matrixInput[1358]), .B(n25096), .C(matrixInput[1350]), 
        .D(n25081), .Z(n25906) );
    VMW_FD \vectorInput_reg[119]  ( .D(n27265), .CP(Clk), .Q(vectorInput[119])
         );
    VMW_AO22 U889 ( .A(matrixInput[605]), .B(n25096), .C(matrixInput[597]), 
        .D(n25081), .Z(n26659) );
    VMW_AO22 U919 ( .A(matrixInput[64]), .B(n25096), .C(matrixInput[56]), .D(
        n25081), .Z(n27200) );
    VMW_AO22 U1005 ( .A(matrixInput[500]), .B(n25096), .C(matrixInput[492]), 
        .D(n25081), .Z(n26764) );
    VMW_AO22 U1195 ( .A(matrixInput[328]), .B(n25096), .C(matrixInput[320]), 
        .D(n25081), .Z(n26936) );
    VMW_AO22 U1614 ( .A(matrixInput[1796]), .B(n25096), .C(matrixInput[1788]), 
        .D(n25081), .Z(n25468) );
    VMW_AO22 U2035 ( .A(matrixInput[1416]), .B(n25096), .C(matrixInput[1408]), 
        .D(n25081), .Z(n25848) );
    VMW_BUFIZ U2624 ( .A(n25197), .E(RD), .Z(\DataOut[13]1 ) );
    VMW_FD \matrixInput_reg[1737]  ( .D(n25519), .CP(Clk), .Q(matrixInput
        [1737]) );
    VMW_FD \matrixInput_reg[1434]  ( .D(n25822), .CP(Clk), .Q(matrixInput
        [1434]) );
    VMW_FD \matrixInput_reg[139]  ( .D(n27117), .CP(Clk), .Q(matrixInput[139])
         );
    VMW_FD \matrixInput_reg[120]  ( .D(n27136), .CP(Clk), .Q(matrixInput[120])
         );
    VMW_AO22 U1784 ( .A(matrixInput[1642]), .B(n25096), .C(matrixInput[1634]), 
        .D(n25081), .Z(n25622) );
    VMW_AO22 U1022 ( .A(matrixInput[485]), .B(n25096), .C(matrixInput[477]), 
        .D(n25081), .Z(n26779) );
    VMW_AO22 U1282 ( .A(matrixInput[250]), .B(n25096), .C(matrixInput[242]), 
        .D(n25081), .Z(n27014) );
    VMW_AO22 U1312 ( .A(matrixInput[223]), .B(n25096), .C(matrixInput[215]), 
        .D(n25081), .Z(n27041) );
    VMW_AO22 U1335 ( .A(matrixInput[2046]), .B(n25096), .C(matrixInput[2038]), 
        .D(n25081), .Z(n25218) );
    VMW_AO22 U1524 ( .A(matrixInput[1877]), .B(n25096), .C(matrixInput[1869]), 
        .D(n25081), .Z(n25387) );
    VMW_AO22 U1956 ( .A(matrixInput[155]), .B(n25096), .C(matrixInput[147]), 
        .D(n25081), .Z(n27109) );
    VMW_AO22 U2295 ( .A(matrixInput[1182]), .B(n25096), .C(matrixInput[1174]), 
        .D(n25081), .Z(n26082) );
    VMW_AO22 U2305 ( .A(matrixInput[1173]), .B(n25096), .C(matrixInput[1165]), 
        .D(n25081), .Z(n26091) );
    VMW_FD \matrixInput_reg[223]  ( .D(n27033), .CP(Clk), .Q(matrixInput[223])
         );
    VMW_FD \matrixInput_reg[113]  ( .D(n27143), .CP(Clk), .Q(matrixInput[113])
         );
    VMW_AO22 U2484 ( .A(matrixInput[1011]), .B(n25096), .C(matrixInput[1003]), 
        .D(n25081), .Z(n26253) );
    VMW_AO22 U2514 ( .A(cOutput[125]), .B(n25089), .C(cOutput[109]), .D(n25088
        ), .Z(n25126) );
    VMW_FD \matrixInput_reg[1704]  ( .D(n25552), .CP(Clk), .Q(matrixInput
        [1704]) );
    VMW_FD \matrixInput_reg[1399]  ( .D(n25857), .CP(Clk), .Q(matrixInput
        [1399]) );
    VMW_FD \matrixInput_reg[1380]  ( .D(n25876), .CP(Clk), .Q(matrixInput
        [1380]) );
    VMW_FD \matrixInput_reg[1083]  ( .D(n26173), .CP(Clk), .Q(matrixInput
        [1083]) );
    VMW_FD \matrixInput_reg[597]  ( .D(n26659), .CP(Clk), .Q(matrixInput[597])
         );
    VMW_FD \matrixInput_reg[1407]  ( .D(n25849), .CP(Clk), .Q(matrixInput
        [1407]) );
    VMW_FD \matrixInput_reg[694]  ( .D(n26562), .CP(Clk), .Q(matrixInput[694])
         );
    VMW_FD \matrixInput_reg[210]  ( .D(n27046), .CP(Clk), .Q(matrixInput[210])
         );
    VMW_FD \matrixInput_reg[209]  ( .D(n27047), .CP(Clk), .Q(matrixInput[209])
         );
    VMW_AO22 U1971 ( .A(matrixInput[1474]), .B(n25096), .C(matrixInput[1466]), 
        .D(n25081), .Z(n25790) );
    VMW_AO22 U2322 ( .A(matrixInput[122]), .B(n25096), .C(matrixInput[114]), 
        .D(n25081), .Z(n27142) );
    VMW_AND3 U2533 ( .A(n25149), .B(n25150), .C(n25151), .Z(n25067) );
    VMW_FD \matrixInput_reg[1223]  ( .D(n26033), .CP(Clk), .Q(matrixInput
        [1223]) );
    VMW_FD \matrixInput_reg[1139]  ( .D(n26117), .CP(Clk), .Q(matrixInput
        [1139]) );
    VMW_FD \matrixInput_reg[1120]  ( .D(n26136), .CP(Clk), .Q(matrixInput
        [1120]) );
    VMW_FD \matrixInput_reg[737]  ( .D(n26519), .CP(Clk), .Q(matrixInput[737])
         );
    VMW_FD \matrixInput_reg[434]  ( .D(n26822), .CP(Clk), .Q(matrixInput[434])
         );
    VMW_AO22 U1493 ( .A(matrixInput[1905]), .B(n25096), .C(matrixInput[1897]), 
        .D(n25081), .Z(n25359) );
    VMW_AO22 U1503 ( .A(matrixInput[1896]), .B(n25096), .C(matrixInput[1888]), 
        .D(n25081), .Z(n25368) );
    VMW_AO22 U2012 ( .A(matrixInput[1437]), .B(n25096), .C(matrixInput[1429]), 
        .D(n25081), .Z(n25827) );
    VMW_AO22 U2182 ( .A(matrixInput[1284]), .B(n25096), .C(matrixInput[1276]), 
        .D(n25081), .Z(n25980) );
    VMW_INV U2603 ( .A(\holder[3] ), .Z(n25065) );
    VMW_FD \matrixInput_reg[1597]  ( .D(n25659), .CP(Clk), .Q(matrixInput
        [1597]) );
    VMW_FD \matrixInput_reg[1113]  ( .D(n26143), .CP(Clk), .Q(matrixInput
        [1113]) );
    VMW_FD \matrixInput_reg[704]  ( .D(n26552), .CP(Clk), .Q(matrixInput[704])
         );
    VMW_FD \matrixInput_reg[380]  ( .D(n26876), .CP(Clk), .Q(matrixInput[380])
         );
    VMW_FD \matrixInput_reg[1694]  ( .D(n25562), .CP(Clk), .Q(matrixInput
        [1694]) );
    VMW_FD \matrixInput_reg[399]  ( .D(n26857), .CP(Clk), .Q(matrixInput[399])
         );
    VMW_AO22 U1633 ( .A(matrixInput[1778]), .B(n25096), .C(matrixInput[1770]), 
        .D(n25081), .Z(n25486) );
    VMW_FD \matrixInput_reg[1210]  ( .D(n26046), .CP(Clk), .Q(matrixInput
        [1210]) );
    VMW_FD \matrixInput_reg[407]  ( .D(n26849), .CP(Clk), .Q(matrixInput[407])
         );
    VMW_FD \matrixInput_reg[1209]  ( .D(n26047), .CP(Clk), .Q(matrixInput
        [1209]) );
    VMW_FD \matrixInput_reg[1931]  ( .D(n25325), .CP(Clk), .Q(matrixInput
        [1931]) );
    VMW_FD \matrixInput_reg[1928]  ( .D(n25328), .CP(Clk), .Q(matrixInput
        [1928]) );
    VMW_FD \matrixInput_reg[1902]  ( .D(n25354), .CP(Clk), .Q(matrixInput
        [1902]) );
    VMW_FD \matrixInput_reg[892]  ( .D(n26364), .CP(Clk), .Q(matrixInput[892])
         );
    VMW_AO22 U505 ( .A(matrixInput[950]), .B(n25096), .C(matrixInput[942]), 
        .D(n25081), .Z(n26314) );
    VMW_AO22 U522 ( .A(matrixInput[935]), .B(n25096), .C(matrixInput[927]), 
        .D(n25081), .Z(n26329) );
    VMW_AO22 U950 ( .A(matrixInput[549]), .B(n25096), .C(matrixInput[541]), 
        .D(n25081), .Z(n26715) );
    VMW_AO22 U314 ( .A(vectorInput[107]), .B(n25095), .C(vectorInput[99]), .D(
        n25080), .Z(n27285) );
    VMW_AO22 U495 ( .A(matrixInput[959]), .B(n25096), .C(matrixInput[951]), 
        .D(n25081), .Z(n26305) );
    VMW_AO22 U439 ( .A(vectorInput[108]), .B(n25095), .C(vectorInput[100]), 
        .D(n25080), .Z(n27284) );
    VMW_AO22 U635 ( .A(matrixInput[833]), .B(n25096), .C(matrixInput[825]), 
        .D(n25081), .Z(n26431) );
    VMW_AO22 U977 ( .A(matrixInput[525]), .B(n25096), .C(matrixInput[517]), 
        .D(n25081), .Z(n26739) );
    VMW_FD \matrixInput_reg[1892]  ( .D(n25364), .CP(Clk), .Q(matrixInput
        [1892]) );
    VMW_FD \matrixInput_reg[902]  ( .D(n26354), .CP(Clk), .Q(matrixInput[902])
         );
    VMW_FD \vectorInput_reg[62]  ( .D(n27322), .CP(Clk), .Q(vectorInput[62])
         );
    VMW_FD \matrixInput_reg[931]  ( .D(n26325), .CP(Clk), .Q(matrixInput[931])
         );
    VMW_FD \matrixInput_reg[928]  ( .D(n26328), .CP(Clk), .Q(matrixInput[928])
         );
    VMW_AO22 U699 ( .A(matrixInput[776]), .B(n25096), .C(matrixInput[768]), 
        .D(n25081), .Z(n26488) );
    VMW_AO22 U709 ( .A(matrixInput[767]), .B(n25096), .C(matrixInput[759]), 
        .D(n25081), .Z(n26497) );
    VMW_AO22 U1267 ( .A(matrixInput[264]), .B(n25096), .C(matrixInput[256]), 
        .D(n25081), .Z(n27000) );
    VMW_AO22 U1804 ( .A(matrixInput[1624]), .B(n25096), .C(matrixInput[1616]), 
        .D(n25081), .Z(n25640) );
    VMW_AO22 U1938 ( .A(matrixInput[1504]), .B(n25096), .C(matrixInput[1496]), 
        .D(n25081), .Z(n25760) );
    VMW_FD \vectorInput_reg[51]  ( .D(n27333), .CP(Clk), .Q(vectorInput[51])
         );
    VMW_FD \vectorInput_reg[48]  ( .D(n27336), .CP(Clk), .Q(vectorInput[48])
         );
    VMW_AO22 U1994 ( .A(matrixInput[1453]), .B(n25096), .C(matrixInput[1445]), 
        .D(n25081), .Z(n25811) );
    VMW_AO22 U1476 ( .A(matrixInput[1919]), .B(n25096), .C(matrixInput[1911]), 
        .D(n25081), .Z(n25345) );
    VMW_FD \matrixInput_reg[646]  ( .D(n26610), .CP(Clk), .Q(matrixInput[646])
         );
    VMW_FD \matrixInput_reg[1051]  ( .D(n26205), .CP(Clk), .Q(matrixInput
        [1051]) );
    VMW_FD \matrixInput_reg[1048]  ( .D(n26208), .CP(Clk), .Q(matrixInput
        [1048]) );
    VMW_AO22 U2257 ( .A(matrixInput[1216]), .B(n25096), .C(matrixInput[1208]), 
        .D(n25081), .Z(n26048) );
    VMW_AO22 U2446 ( .A(matrixInput[1046]), .B(n25096), .C(matrixInput[1038]), 
        .D(n25081), .Z(n26218) );
    VMW_AO22 U1157 ( .A(matrixInput[363]), .B(n25096), .C(matrixInput[355]), 
        .D(n25081), .Z(n26901) );
    VMW_FD \matrixInput_reg[1352]  ( .D(n25904), .CP(Clk), .Q(matrixInput
        [1352]) );
    VMW_FD \matrixInput_reg[545]  ( .D(n26711), .CP(Clk), .Q(matrixInput[545])
         );
    VMW_FD \matrixInput_reg[1062]  ( .D(n26194), .CP(Clk), .Q(matrixInput
        [1062]) );
    VMW_FD \matrixInput_reg[675]  ( .D(n26581), .CP(Clk), .Q(matrixInput[675])
         );
    VMW_AO22 U1746 ( .A(matrixInput[1677]), .B(n25096), .C(matrixInput[1669]), 
        .D(n25081), .Z(n25587) );
    VMW_FD \matrixInput_reg[1378]  ( .D(n25878), .CP(Clk), .Q(matrixInput
        [1378]) );
    VMW_FD \matrixInput_reg[1361]  ( .D(n25895), .CP(Clk), .Q(matrixInput
        [1361]) );
    VMW_AO22 U1170 ( .A(matrixInput[351]), .B(n25096), .C(matrixInput[343]), 
        .D(n25081), .Z(n26913) );
    VMW_AO22 U1761 ( .A(matrixInput[1663]), .B(n25096), .C(matrixInput[1655]), 
        .D(n25081), .Z(n25601) );
    VMW_AO22 U2167 ( .A(matrixInput[136]), .B(n25096), .C(matrixInput[128]), 
        .D(n25081), .Z(n27128) );
    VMW_FD \matrixInput_reg[576]  ( .D(n26680), .CP(Clk), .Q(matrixInput[576])
         );
    VMW_AO22 U1240 ( .A(matrixInput[288]), .B(n25096), .C(matrixInput[280]), 
        .D(n25081), .Z(n26976) );
    VMW_AO22 U1451 ( .A(matrixInput[1942]), .B(n25096), .C(matrixInput[1934]), 
        .D(n25081), .Z(n25322) );
    VMW_AO22 U1823 ( .A(matrixInput[167]), .B(n25096), .C(matrixInput[159]), 
        .D(n25081), .Z(n27097) );
    VMW_AO22 U2140 ( .A(matrixInput[1321]), .B(n25096), .C(matrixInput[1313]), 
        .D(n25081), .Z(n25943) );
    VMW_FD \matrixInput_reg[1646]  ( .D(n25610), .CP(Clk), .Q(matrixInput
        [1646]) );
    VMW_FD \matrixInput_reg[1545]  ( .D(n25711), .CP(Clk), .Q(matrixInput
        [1545]) );
    VMW_FD \matrixInput_reg[352]  ( .D(n26904), .CP(Clk), .Q(matrixInput[352])
         );
    VMW_FD \matrixInput_reg[2038]  ( .D(n25218), .CP(Clk), .Q(matrixInput
        [2038]) );
    VMW_FD \matrixInput_reg[2021]  ( .D(n25235), .CP(Clk), .Q(matrixInput
        [2021]) );
    VMW_FD \matrixInput_reg[1675]  ( .D(n25581), .CP(Clk), .Q(matrixInput
        [1675]) );
    VMW_AO22 U2270 ( .A(matrixInput[1205]), .B(n25096), .C(matrixInput[1197]), 
        .D(n25081), .Z(n26059) );
    VMW_FD \matrixInput_reg[2012]  ( .D(n25244), .CP(Clk), .Q(matrixInput
        [2012]) );
    VMW_AO22 U2461 ( .A(matrixInput[1032]), .B(n25096), .C(matrixInput[1024]), 
        .D(n25081), .Z(n26232) );
    VMW_FD \matrixInput_reg[1576]  ( .D(n25680), .CP(Clk), .Q(matrixInput
        [1576]) );
    VMW_FD \matrixInput_reg[378]  ( .D(n26878), .CP(Clk), .Q(matrixInput[378])
         );
    VMW_FD \matrixInput_reg[361]  ( .D(n26895), .CP(Clk), .Q(matrixInput[361])
         );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_14 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n1, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_13 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n2, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n2) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n2), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_12 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n3, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n3) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_15 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_15 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n31, n32, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , \CARRYB[2][1] , 
        \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \ab[3][3] , 
        \A1[2] , n33, n34, n35, \A2[3] , \ab[2][0] , \ab[6][0] , \ab[2][2] , 
        \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , 
        \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[4][2] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[1][1] , \ab[0][7] , 
        \CARRYB[1][5] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , n36, \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , \A2[4] , 
        \A2[2] , \A2[6] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n31) );
    VMW_PULLDOWN U5 ( .Z(n33) );
    VMW_PULLDOWN U6 ( .Z(n34) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n32), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n35) );
    VMW_PULLDOWN U8 ( .Z(n36) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n33), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n34), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n31), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_15 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n36), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n32) );
    VMW_FADD S0_1 ( .CI(n35), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_11 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n4, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n4) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n4), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_14 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_14 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n37, n38, n40, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n41, \A2[3] , \ab[6][0] , \ab[2][2] , 
        \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , 
        \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[0][7] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , 
        \ab[4][3] , \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , n39, n42, 
        \SUMB[1][3] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , \CARRYB[2][2] , 
        \A2[2] , \A2[6] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , 
        \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , 
        \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n37) );
    VMW_PULLDOWN U5 ( .Z(n39) );
    VMW_PULLDOWN U6 ( .Z(n40) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n38), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n41) );
    VMW_PULLDOWN U8 ( .Z(n42) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n39), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n40), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n37), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_14 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n42), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n38) );
    VMW_FADD S0_1 ( .CI(n41), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_13 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_13 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n43, n44, n46, n47, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n48, lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[0][6] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[0][7] , \CARRYB[1][5] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \CARRYB[1][1] , \SUMB[3][3] , \ab[1][4] , \CARRYB[4][0] , 
        n45, \A2[2] , \A2[6] , \ab[1][6] , \SUMB[3][1] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n43) );
    VMW_PULLDOWN U5 ( .Z(n45) );
    VMW_PULLDOWN U6 ( .Z(n46) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n44), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n47) );
    VMW_PULLDOWN U8 ( .Z(n48) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n45), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n46), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n43), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_13 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n48), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n44) );
    VMW_FADD S0_1 ( .CI(n47), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_12 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_12 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n49, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , n50, n51, n52, 
        \SUMB[1][2] , \CARRYB[2][3] , n53, \ab[1][3] , \A1[4] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , n54, lsb_0, \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , 
        \CARRYB[1][0] , \SUMB[2][1] , \ab[0][7] , \ab[1][5] , \SUMB[3][2] , 
        \CARRYB[1][5] , \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , 
        \SUMB[2][5] , \ab[0][2] , \ab[1][1] , \ab[4][1] , \ab[0][3] , 
        \SUMB[2][4] , \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , 
        \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , 
        \CARRYB[4][2] , \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , 
        \SUMB[2][2] , \ab[4][3] , \ab[5][0] , \A2[6] , \SUMB[1][3] , 
        \ab[0][1] , \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \A2[4] , \A2[2] , \ab[6][1] , 
        \ab[2][3] , \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , 
        \ab[7][0] , \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , 
        \CARRYB[2][0] , \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n49) );
    VMW_PULLDOWN U5 ( .Z(n51) );
    VMW_PULLDOWN U6 ( .Z(n52) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n50), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n53) );
    VMW_PULLDOWN U8 ( .Z(n54) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n51), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n52), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n49), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_12 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n54), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n50) );
    VMW_FADD S0_1 ( .CI(n53), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_10 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n5, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n5) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n5), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_11 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_11 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n55, n56, n60, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , n57, n58, \ab[0][7] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \SUMB[2][2] , n59, \ab[1][2] , 
        \ab[0][1] , \ab[4][3] , \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , 
        \A2[2] , \A2[6] , \SUMB[1][3] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n55) );
    VMW_PULLDOWN U5 ( .Z(n57) );
    VMW_PULLDOWN U6 ( .Z(n58) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n56), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n59) );
    VMW_PULLDOWN U8 ( .Z(n60) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n57), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n58), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n55), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_11 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n60), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n56) );
    VMW_FADD S0_1 ( .CI(n59), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_10 ( A, B, CI, 
    SUM, CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_10 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n61, n66, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , \CARRYB[1][0] , 
        \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , 
        \SUMB[2][5] , \ab[0][2] , n62, n63, \ab[0][7] , \CARRYB[1][5] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \CARRYB[1][1] , n64, \ab[1][4] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , n65, \ab[1][6] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A2[2] , \A2[6] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n61) );
    VMW_PULLDOWN U5 ( .Z(n63) );
    VMW_PULLDOWN U6 ( .Z(n64) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n62), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n65) );
    VMW_PULLDOWN U8 ( .Z(n66) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n63), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n64), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n61), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_10 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n66), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n62) );
    VMW_FADD S0_1 ( .CI(n65), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_9 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n6, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n6) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n6), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_9 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_9 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n67, n69, n72, \A1[13] , \A2[5] , \CARRYB[2][1] , \SUMB[5][2] , 
        \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \A2[1] , \SUMB[1][4] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n68, lsb_0, \A2[3] , \ab[6][0] , 
        \ab[2][2] , \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , n70, n71, \ab[0][6] , 
        \ab[1][5] , \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \SUMB[2][4] , \A2[2] , \A2[6] , \ab[0][7] , 
        \ab[0][3] , \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , 
        \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , 
        \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , \CARRYB[5][1] , 
        \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n67) );
    VMW_PULLDOWN U5 ( .Z(n69) );
    VMW_PULLDOWN U6 ( .Z(n70) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n68), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n71) );
    VMW_PULLDOWN U8 ( .Z(n72) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n69), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n70), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n67), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_9 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n72), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n68) );
    VMW_FADD S0_1 ( .CI(n71), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_8 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n7, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n7) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n7), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_8 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_8 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n73, n74, n75, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , 
        \CARRYB[2][3] , \ab[1][3] , \A1[4] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , lsb_0, \ab[0][6] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \CARRYB[1][0] , 
        \SUMB[2][1] , n76, n78, \ab[1][5] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \ab[0][7] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , 
        \ab[4][3] , \ab[5][0] , n77, \A2[6] , \SUMB[1][3] , \SUMB[4][2] , 
        \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \A2[4] , \A2[2] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n73) );
    VMW_PULLDOWN U5 ( .Z(n75) );
    VMW_PULLDOWN U6 ( .Z(n76) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n74), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n77) );
    VMW_PULLDOWN U8 ( .Z(n78) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n75), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n76), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n73), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_8 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n78), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n74) );
    VMW_FADD S0_1 ( .CI(n77), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_7 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_7 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n79, n80, n81, n82, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , n83, \A2[3] , 
        \A1[0] , \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , 
        \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[5][1] , 
        \SUMB[3][4] , n84, lsb_0, \ab[4][2] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[0][7] , \CARRYB[1][5] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , \CARRYB[4][2] , \ab[0][5] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , 
        \ab[4][3] , \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , \SUMB[5][1] , 
        \CARRYB[6][0] , \A2[4] , \A2[2] , \A2[6] , \SUMB[1][3] , \ab[3][4] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \SUMB[1][5] , \A1[1] , 
        \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , \ab[3][2] , 
        \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , \CARRYB[3][3] , \ab[2][5] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n79) );
    VMW_PULLDOWN U5 ( .Z(n81) );
    VMW_PULLDOWN U6 ( .Z(n82) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n80), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n83) );
    VMW_PULLDOWN U8 ( .Z(n84) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n81), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n82), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n79), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_7 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n84), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n80) );
    VMW_FADD S0_1 ( .CI(n83), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_7 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n8, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n8) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n8), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_6 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_6 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n85, \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , \CARRYB[2][1] , 
        \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \ab[3][3] , 
        \ab[2][0] , \A1[2] , n86, n90, \A2[3] , \ab[6][0] , \ab[2][2] , 
        \A1[0] , \SUMB[1][6] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , lsb_0, 
        \ab[1][3] , \SUMB[1][2] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , \ab[0][7] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \CARRYB[1][1] , n87, n88, \ab[1][6] , \ab[1][4] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , n89, \A2[2] , 
        \A2[6] , \SUMB[1][3] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \A1[1] , \A2[4] , 
        \SUMB[1][5] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , 
        \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n85) );
    VMW_PULLDOWN U5 ( .Z(n87) );
    VMW_PULLDOWN U6 ( .Z(n88) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n86), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n89) );
    VMW_PULLDOWN U8 ( .Z(n90) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n87), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n88), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n85), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_6 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n90), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n86) );
    VMW_FADD S0_1 ( .CI(n89), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_5 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_5 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n91, lsb_0, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , n92, n93, n94, n96, \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , 
        \CARRYB[1][0] , \SUMB[2][1] , \ab[1][5] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[0][7] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[5][0] , 
        \A2[6] , \SUMB[1][3] , \ab[0][1] , \ab[4][3] , \SUMB[4][2] , 
        \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[2][3] , n95, \A2[2] , \ab[6][1] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n91) );
    VMW_PULLDOWN U5 ( .Z(n93) );
    VMW_PULLDOWN U6 ( .Z(n94) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n92), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n95) );
    VMW_PULLDOWN U8 ( .Z(n96) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n93), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n94), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] ), 
        .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n91), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_5 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n96), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n92) );
    VMW_FADD S0_1 ( .CI(n95), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] ), 
        .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_4 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_4 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n97, \A1[13] , \A2[5] , n98, n99, n100, \CARRYB[2][1] , \SUMB[5][2] , 
        \CARRYB[3][2] , \A2[1] , \SUMB[1][4] , \ab[2][4] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A2[3] , 
        \A1[0] , \SUMB[1][6] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , n101, lsb_0, \ab[1][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , 
        \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , n102, \A2[2] , \A2[6] , 
        \ab[0][7] , \ab[0][6] , \ab[1][5] , \CARRYB[1][0] , \SUMB[2][1] , 
        \SUMB[3][2] , \CARRYB[1][5] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[1][1] , \ab[4][1] , 
        \ab[0][3] , \SUMB[2][4] , \ab[1][0] , \ab[5][2] , \ab[1][6] , 
        \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , 
        \ab[0][5] , \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , 
        \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , 
        \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \A2[4] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n97) );
    VMW_PULLDOWN U5 ( .Z(n99) );
    VMW_PULLDOWN U6 ( .Z(n100) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n98), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] ), 
        .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n101) );
    VMW_PULLDOWN U8 ( .Z(n102) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n99), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] ), 
        .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n100), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] 
        ), .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n97), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] ), 
        .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_4 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n102), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n98) );
    VMW_FADD S0_1 ( .CI(n101), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] 
        ), .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_6 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n9, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n9) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n9), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_3 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_3 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n103, n106, n107, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , lsb_0, 
        \ab[1][3] , \SUMB[1][2] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , 
        \ab[5][1] , \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , \SUMB[2][3] , 
        \CARRYB[5][0] , \SUMB[6][1] , n108, \ab[0][6] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , \ab[4][0] , 
        \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \CARRYB[1][5] , \ab[1][1] , 
        \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , \ab[5][2] , n104, 
        \ab[0][7] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , 
        \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \SUMB[2][2] , n105, \A2[2] , \A2[6] , 
        \SUMB[1][3] , \ab[1][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \A1[1] , \A2[4] , 
        \SUMB[1][5] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \ab[2][1] , 
        \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , \ab[2][5] , 
        \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n103) );
    VMW_PULLDOWN U5 ( .Z(n105) );
    VMW_PULLDOWN U6 ( .Z(n106) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n104), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] 
        ), .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n107) );
    VMW_PULLDOWN U8 ( .Z(n108) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n105), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] 
        ), .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n106), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] 
        ), .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n103), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] 
        ), .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_3 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n108), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n104) );
    VMW_FADD S0_1 ( .CI(n107), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] 
        ), .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_2 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_2 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n109, n112, \A1[13] , \A2[5] , \CARRYB[2][1] , \SUMB[5][2] , 
        \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , \A2[1] , \SUMB[1][4] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , n110, n111, n113, n114, \A2[3] , 
        \ab[6][0] , \ab[2][2] , \A1[0] , \SUMB[1][6] , \SUMB[1][2] , 
        \ab[3][1] , \CARRYB[3][0] , \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , 
        lsb_0, \ab[1][3] , \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][6] , 
        \ab[0][4] , \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , 
        \ab[1][5] , \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][4] , 
        \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , \ab[1][1] , 
        \CARRYB[1][5] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \A2[4] , \A2[2] , \A2[6] , \ab[0][7] , \ab[1][6] , 
        \ab[1][4] , \CARRYB[1][1] , \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , 
        \ab[0][5] , \CARRYB[4][2] , \SUMB[1][3] , \CARRYB[1][3] , 
        \CARRYB[5][1] , \ab[1][2] , \SUMB[2][2] , \ab[0][1] , \ab[4][3] , 
        \ab[5][0] , \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , 
        \CARRYB[3][3] , \ab[2][5] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n109) );
    VMW_PULLDOWN U5 ( .Z(n111) );
    VMW_PULLDOWN U6 ( .Z(n112) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n110), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] 
        ), .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n113) );
    VMW_PULLDOWN U8 ( .Z(n114) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n111), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] 
        ), .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n112), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] 
        ), .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n109), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] 
        ), .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_2 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n114), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n110) );
    VMW_FADD S0_1 ( .CI(n113), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] 
        ), .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_5 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n10, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n10) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n10), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_4 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n11, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n11) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n11), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_1 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_1 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n115, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , n116, n118, n120, \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , lsb_0, \ab[1][3] , \SUMB[1][2] , \A1[4] , \CARRYB[2][3] , 
        \ab[4][2] , \ab[5][1] , \SUMB[3][4] , \ab[0][6] , \ab[0][4] , 
        \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , \SUMB[6][1] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \SUMB[2][4] , \ab[0][7] , \ab[0][3] , 
        \ab[1][0] , \ab[5][2] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \SUMB[2][2] , n117, \ab[1][2] , 
        \ab[0][1] , \ab[4][3] , \ab[5][0] , \CARRYB[3][1] , n119, \A2[2] , 
        \A2[6] , \SUMB[1][3] , \SUMB[4][2] , \ab[3][4] , \SUMB[5][1] , 
        \CARRYB[6][0] , \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , 
        \SUMB[1][5] , \A1[1] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \A2[4] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n115) );
    VMW_PULLDOWN U5 ( .Z(n117) );
    VMW_PULLDOWN U6 ( .Z(n118) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n116), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] 
        ), .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n119) );
    VMW_PULLDOWN U8 ( .Z(n120) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n117), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] 
        ), .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n118), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] 
        ), .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n115), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] 
        ), .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_1 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n120), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n116) );
    VMW_FADD S0_1 ( .CI(n119), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] 
        ), .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_0 ( A, B, CI, SUM, 
    CO );
input  [13:0] A;
input  [13:0] B;
output [13:0] SUM;
input  CI;
output CO;
    wire \A[4] , \A[0] , \A[2] , \A[3] , \A[5] , \A[1] ;
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    assign SUM[5] = \A[5] ;
    assign SUM[4] = \A[4] ;
    assign SUM[3] = \A[3] ;
    assign SUM[2] = \A[2] ;
    assign SUM[1] = \A[1] ;
    assign SUM[0] = \A[0] ;
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_0 ( A, B, TC, 
    PRODUCT );
input  [7:0] A;
input  [7:0] B;
output [15:0] PRODUCT;
input  TC;
    wire n121, lsb_0, \A2[3] , \A2[1] , \A1[13] , \A2[5] , \SUMB[1][4] , 
        \CARRYB[2][1] , \SUMB[5][2] , \ab[2][4] , \CARRYB[3][2] , \SUMB[4][1] , 
        \ab[3][3] , \ab[2][0] , \A1[2] , \ab[6][0] , \ab[2][2] , \A1[0] , 
        \SUMB[1][6] , \ab[1][3] , \SUMB[1][2] , \ab[3][1] , \CARRYB[3][0] , 
        \SUMB[4][3] , \A1[4] , \CARRYB[2][3] , \ab[4][2] , \ab[5][1] , 
        \SUMB[3][4] , \ab[0][4] , \CARRYB[1][2] , \SUMB[2][3] , \CARRYB[5][0] , 
        \SUMB[6][1] , n122, n123, n124, n126, \ab[0][6] , \ab[1][5] , 
        \CARRYB[1][0] , \SUMB[2][1] , \SUMB[3][2] , \CARRYB[1][5] , 
        \CARRYB[1][4] , \ab[4][0] , \CARRYB[4][1] , \SUMB[2][5] , \ab[0][2] , 
        \ab[1][1] , \ab[4][1] , \ab[0][3] , \SUMB[2][4] , \ab[1][0] , 
        \ab[5][2] , \ab[0][7] , \ab[1][6] , \ab[1][4] , \CARRYB[1][1] , 
        \SUMB[3][3] , \SUMB[3][1] , \CARRYB[4][0] , \ab[0][5] , \CARRYB[4][2] , 
        \CARRYB[1][3] , \CARRYB[5][1] , \SUMB[2][2] , \A2[2] , \A2[6] , 
        \SUMB[1][3] , \ab[1][2] , \ab[0][1] , \ab[4][3] , \ab[5][0] , 
        \SUMB[4][2] , \CARRYB[3][1] , \ab[3][4] , \SUMB[5][1] , \CARRYB[6][0] , 
        \CARRYB[2][2] , \A1[5] , \ab[6][1] , \ab[2][3] , \A1[1] , n125, 
        \SUMB[1][5] , \ab[3][0] , \CARRYB[2][4] , \ab[7][0] , \A2[4] , 
        \ab[2][1] , \ab[3][2] , \A1[3] , \SUMB[1][1] , \CARRYB[2][0] , 
        \ab[2][5] , \CARRYB[3][3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 ;
    VMW_PULLDOWN U3 ( .Z(n121) );
    VMW_PULLDOWN U5 ( .Z(n123) );
    VMW_PULLDOWN U6 ( .Z(n124) );
    VMW_PULLDOWN U14 ( .Z(\A2[1] ) );
    VMW_FADD S0_4 ( .CI(n122), .A(\ab[0][5] ), .B(\ab[1][4] ), .S(\SUMB[1][4] 
        ), .CO(\CARRYB[1][4] ) );
    VMW_FADD S2_2_2 ( .CI(\SUMB[1][3] ), .A(\ab[2][2] ), .B(\CARRYB[1][2] ), 
        .S(\SUMB[2][2] ), .CO(\CARRYB[2][2] ) );
    VMW_AND2 U21 ( .A(A[1]), .B(B[3]), .Z(\ab[1][3] ) );
    VMW_FADD S2_3_2 ( .CI(\SUMB[2][3] ), .A(\ab[3][2] ), .B(\CARRYB[2][2] ), 
        .S(\SUMB[3][2] ), .CO(\CARRYB[3][2] ) );
    VMW_FADD S2_5_1 ( .CI(\SUMB[4][2] ), .A(\ab[5][1] ), .B(\CARRYB[4][1] ), 
        .S(\SUMB[5][1] ), .CO(\CARRYB[5][1] ) );
    VMW_AND2 U28 ( .A(A[0]), .B(B[5]), .Z(\ab[0][5] ) );
    VMW_AND2 U33 ( .A(B[0]), .B(A[7]), .Z(\ab[7][0] ) );
    VMW_PULLDOWN U7 ( .Z(n125) );
    VMW_PULLDOWN U8 ( .Z(n126) );
    VMW_PULLDOWN U13 ( .Z(\A2[3] ) );
    VMW_AND2 U34 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
    VMW_AND2 U41 ( .A(A[5]), .B(B[1]), .Z(\ab[5][1] ) );
    VMW_AND2 U46 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
    VMW_FADD S2_4_1 ( .CI(\SUMB[3][2] ), .A(\ab[4][1] ), .B(\CARRYB[3][1] ), 
        .S(\SUMB[4][1] ), .CO(\CARRYB[4][1] ) );
    VMW_FADD S1_6_0 ( .CI(\SUMB[5][1] ), .A(\ab[6][0] ), .B(\CARRYB[5][0] ), 
        .S(\A1[4] ), .CO(\CARRYB[6][0] ) );
    VMW_AND2 U26 ( .A(A[2]), .B(B[1]), .Z(\ab[2][1] ) );
    VMW_AND2 U48 ( .A(A[2]), .B(B[3]), .Z(\ab[2][3] ) );
    VMW_PULLDOWN U9 ( .Z(\A2[4] ) );
    VMW_PULLDOWN U12 ( .Z(lsb_0) );
    VMW_FADD S0_3 ( .CI(n123), .A(\ab[0][4] ), .B(\ab[1][3] ), .S(\SUMB[1][3] 
        ), .CO(\CARRYB[1][3] ) );
    VMW_AND2 U35 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
    VMW_AND2 U53 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    VMW_FADD S2_2_5 ( .CI(\SUMB[1][6] ), .A(\ab[2][5] ), .B(\CARRYB[1][5] ), 
        .S(\SUMB[2][5] ) );
    VMW_FADD S0_2 ( .CI(n124), .A(\ab[0][3] ), .B(\ab[1][2] ), .S(\SUMB[1][2] 
        ), .CO(\CARRYB[1][2] ) );
    VMW_AND2 U40 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
    VMW_AND2 U52 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    VMW_FADD S2_2_4 ( .CI(\SUMB[1][5] ), .A(\ab[2][4] ), .B(\CARRYB[1][4] ), 
        .S(\SUMB[2][4] ), .CO(\CARRYB[2][4] ) );
    VMW_AND2 U27 ( .A(A[0]), .B(B[2]), .Z(\ab[0][2] ) );
    VMW_FADD S0_5 ( .CI(n121), .A(\ab[0][6] ), .B(\ab[1][5] ), .S(\SUMB[1][5] 
        ), .CO(\CARRYB[1][5] ) );
    VMW_AND2 U20 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    VMW_AND2 U49 ( .A(A[3]), .B(B[3]), .Z(\ab[3][3] ) );
    VMW_FADD S2_3_4 ( .CI(\SUMB[2][5] ), .A(\ab[3][4] ), .B(\CARRYB[2][4] ), 
        .S(\SUMB[3][4] ) );
    VMW_FADD S2_3_3 ( .CI(\SUMB[2][4] ), .A(\ab[3][3] ), .B(\CARRYB[2][3] ), 
        .S(\SUMB[3][3] ), .CO(\CARRYB[3][3] ) );
    VMW_AND2 U29 ( .A(A[1]), .B(B[5]), .Z(\ab[1][5] ) );
    VMW_AND2 U47 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
    VMW_FADD S2_2_3 ( .CI(\SUMB[1][4] ), .A(\ab[2][3] ), .B(\CARRYB[1][3] ), 
        .S(\SUMB[2][3] ), .CO(\CARRYB[2][3] ) );
    VMW_FADD S1_3_0 ( .CI(\SUMB[2][1] ), .A(\ab[3][0] ), .B(\CARRYB[2][0] ), 
        .S(\A1[1] ), .CO(\CARRYB[3][0] ) );
    VMW_PULLDOWN U15 ( .Z(\A1[13] ) );
    VMW_XOR2 U17 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
    VMW_AND2 U22 ( .A(A[1]), .B(B[4]), .Z(\ab[1][4] ) );
    VMW_AND2 U32 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    VMW_AND2 U39 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_14_0 FS ( .A({\A1[13] , 
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({UNCONNECTED_8, UNCONNECTED_9, 
        UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, UNCONNECTED_13, 
        UNCONNECTED_14, \A2[6] , \A2[5] , \A2[4] , \A2[3] , \A2[2] , \A2[1] , 
        lsb_0}), .CI(lsb_0), .SUM({UNCONNECTED_15, UNCONNECTED_16, 
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, PRODUCT[7], PRODUCT[6], PRODUCT[5], 
        PRODUCT[4], PRODUCT[3], PRODUCT[2]}) );
    VMW_FADD S1_2_0 ( .CI(\SUMB[1][1] ), .A(\ab[2][0] ), .B(\CARRYB[1][0] ), 
        .S(\A1[0] ), .CO(\CARRYB[2][0] ) );
    VMW_FADD S2_2_1 ( .CI(\SUMB[1][2] ), .A(\ab[2][1] ), .B(\CARRYB[1][1] ), 
        .S(\SUMB[2][1] ), .CO(\CARRYB[2][1] ) );
    VMW_AND2 U30 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
    VMW_FADD S2_3_1 ( .CI(\SUMB[2][2] ), .A(\ab[3][1] ), .B(\CARRYB[2][1] ), 
        .S(\SUMB[3][1] ), .CO(\CARRYB[3][1] ) );
    VMW_FADD S2_5_2 ( .CI(\SUMB[4][3] ), .A(\ab[5][2] ), .B(\CARRYB[4][2] ), 
        .S(\SUMB[5][2] ) );
    VMW_PULLDOWN U10 ( .Z(\A2[2] ) );
    VMW_AND2 U42 ( .A(A[5]), .B(B[2]), .Z(\ab[5][2] ) );
    VMW_AND2 U45 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    VMW_FADD S2_4_2 ( .CI(\SUMB[3][3] ), .A(\ab[4][2] ), .B(\CARRYB[3][2] ), 
        .S(\SUMB[4][2] ), .CO(\CARRYB[4][2] ) );
    VMW_PULLDOWN U11 ( .Z(\A2[6] ) );
    VMW_FADD S0_0 ( .CI(n126), .A(\ab[0][1] ), .B(\ab[1][0] ), .S(PRODUCT[1]), 
        .CO(\CARRYB[1][0] ) );
    VMW_AND2 U19 ( .A(A[0]), .B(B[3]), .Z(\ab[0][3] ) );
    VMW_AND2 U25 ( .A(A[0]), .B(B[7]), .Z(\ab[0][7] ) );
    VMW_AND2 U37 ( .A(B[5]), .B(A[2]), .Z(\ab[2][5] ) );
    VMW_AND2 U50 ( .A(B[4]), .B(A[3]), .Z(\ab[3][4] ) );
    VMW_AND2 U36 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    VMW_PULLDOWN U4 ( .Z(n122) );
    VMW_FADD S0_1 ( .CI(n125), .A(\ab[0][2] ), .B(\ab[1][1] ), .S(\SUMB[1][1] 
        ), .CO(\CARRYB[1][1] ) );
    VMW_AND2 U18 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
    VMW_AND2 U43 ( .A(A[0]), .B(B[6]), .Z(\ab[0][6] ) );
    VMW_AND2 U51 ( .A(A[2]), .B(B[4]), .Z(\ab[2][4] ) );
    VMW_AND2 U23 ( .A(A[0]), .B(B[4]), .Z(\ab[0][4] ) );
    VMW_AND2 U24 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    VMW_FADD S1_4_0 ( .CI(\SUMB[3][1] ), .A(\ab[4][0] ), .B(\CARRYB[3][0] ), 
        .S(\A1[2] ), .CO(\CARRYB[4][0] ) );
    VMW_FADD S2_6_1 ( .CI(\SUMB[5][2] ), .A(\ab[6][1] ), .B(\CARRYB[5][1] ), 
        .S(\SUMB[6][1] ) );
    VMW_AND2 U38 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
    VMW_FADD S4_0 ( .CI(\SUMB[6][1] ), .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .S(
        \A1[5] ) );
    VMW_AND2 U44 ( .A(B[6]), .B(A[1]), .Z(\ab[1][6] ) );
    VMW_FADD S2_4_3 ( .CI(\SUMB[3][4] ), .A(\ab[4][3] ), .B(\CARRYB[3][3] ), 
        .S(\SUMB[4][3] ) );
    VMW_FADD S1_5_0 ( .CI(\SUMB[4][1] ), .A(\ab[5][0] ), .B(\CARRYB[4][0] ), 
        .S(\A1[3] ), .CO(\CARRYB[5][0] ) );
    VMW_PULLDOWN U16 ( .Z(\A2[5] ) );
    VMW_AND2 U31 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_3 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n12, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n12) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n12), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_2 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n13, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n13) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n13), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_1 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n14, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n14) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n14), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_0 ( A, B, CI, SUM, 
    CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n15, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n15) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n15), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module VectorDotProduct_pVectorSize16_pWordSize8 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, vectorAInput, vectorBInput, cOutput );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [127:0] vectorAInput;
output [7:0] cOutput;
input  [127:0] vectorBInput;
input  Clk, Reset, RD, WR;
    wire n1539, n1532, n1548, \result60[1] , \n642[8] , \result1264[2] , 
        \result1086[6] , \result1175[4] , \result463[5] , n1554, n1534, n1541, 
        n1553, \n998[2] , \n1176[4] , \n553[7] , \n464[7] , \result552[2] , 
        \n642[1] , \result997[1] , \n909[5] , \result60[5] , \result285[2] , 
        \n820[4] , \result463[1] , \result1175[0] , \n909[8] , \result1264[6] , 
        \result1353[6] , \result1086[2] , \n642[5] , \result285[6] , 
        \result552[6] , \result997[5] , \n909[1] , \n998[6] , \n553[3] , 
        \n464[3] , n1561, n1546, n1533, \result552[4] , \result908[4] , 
        \n909[3] , \n553[1] , \n464[1] , \n642[7] , \result908[6] , \n998[4] , 
        \result997[7] , \result285[4] , \n995[8] , \result1353[4] , 
        \result1086[0] , \result60[7] , \n642[3] , \result997[3] , \n820[6] , 
        \n1176[2] , \result463[3] , \result1175[2] , \n553[8] , \n1262[4] , 
        \n464[8] , \result285[0] , n1547, \result60[3] , \result552[0] , 
        \result908[2] , \n464[5] , \n553[5] , \result1175[6] , \n909[7] , 
        \n820[2] , \result463[7] , \n1176[6] , \result641[1] , \result1264[0] , 
        \result1353[0] , \result1086[4] , \n286[2] , \n731[8] , \result819[3] , 
        \n197[4] , n1560, \result196[1] , \n106[3] , \result374[5] , 
        \n1442[6] , \n731[1] , \result730[4] , n1537, n1549, n1552, n1555, 
        \result641[5] , \result196[5] , \n1265[7] , \n1087[3] , \n106[7] , 
        \n375[4] , \result374[1] , \result819[7] , \n1354[4] , \n286[6] , 
        \n1265[3] , \n906[8] , \n1087[7] , \n731[5] , \n1442[2] , 
        \result730[0] , \n731[7] , \n1265[1] , \n1087[5] , \result641[7] , 
        \result730[2] , \n1354[6] , \n286[4] , \n1265[8] , n1559, n1540, n1535, 
        \result196[7] , \n106[5] , \result374[3] , \n375[6] , \n197[2] , 
        \result819[5] , \n1442[4] , \result730[6] , \n731[3] , \n1265[5] , 
        \n1351[6] , \result196[3] , \n1087[1] , \n106[8] , \n375[2] , 
        \n197[6] , \n106[1] , \result374[7] , n1542, n1550, \result641[3] , 
        \n1087[8] , \n286[8] , \n1442[5] , \result730[7] , \n1354[2] , 
        \n731[2] , \n1265[4] , \n375[3] , \n197[7] , \result819[0] , 
        \result641[2] , \result196[2] , \result374[6] , \n1354[3] , \n286[1] , 
        \n731[6] , \result641[6] , \n1442[1] , \n1087[4] , \result730[3] , 
        \n286[5] , \n1354[7] , \n1442[8] , n1545, n1562, \result641[4] , 
        \result196[6] , \result196[4] , \n106[4] , \result374[2] , \n375[7] , 
        \result819[4] , \n197[3] , \n106[6] , \result374[0] , \result819[6] , 
        \n375[5] , \n197[1] , \n286[7] , \n1354[5] , \n731[4] , \n1442[3] , 
        \n1265[2] , \n1087[6] , \result730[1] , \n197[8] , n1543, n1558, n1544, 
        n1557, \result641[0] , \n1354[1] , \n286[3] , \n375[1] , \n197[5] , 
        \result819[2] , \n642[2] , \result997[2] , \result196[0] , \n106[2] , 
        \result374[4] , \n375[8] , \n1442[7] , \result730[5] , \n1265[6] , 
        \n1087[2] , \n1354[8] , \result285[1] , \n553[4] , \n464[4] , n1538, 
        n1556, \result60[2] , \result552[1] , \result908[3] , \n998[1] , 
        \n909[6] , \n998[8] , \result1175[7] , \n820[3] , \n1176[7] , 
        \result463[6] , \result552[5] , \result1264[1] , \result1353[1] , 
        \result1086[5] , \n642[6] , \result908[7] , \n998[5] , \n909[2] , 
        \result60[6] , \result997[6] , \result285[5] , \result1353[5] , 
        \result1264[5] , \result1086[1] , n1551, \n820[7] , \result463[2] , 
        \result1175[3] , \n1176[3] , \n820[5] , \result463[0] , \n1176[1] , 
        \result1175[1] , \result1264[7] , \result1353[7] , \result1086[3] , 
        n1536, \result60[4] , \n642[4] , \result285[7] , \result60[0] , 
        \result552[7] , \result997[4] , \n1176[8] , \result908[5] , \n998[7] , 
        \n553[2] , \n464[2] , \result1353[3] , \result1264[3] , 
        \result1175[5] , \result1086[7] , \n1176[5] , \n820[1] , 
        \result463[4] , \n464[6] , \n553[6] , \result552[3] , \result908[1] , 
        \n998[3] , \n820[8] , \n909[4] , \n817[7] , \result285[3] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 , UNCONNECTED_23 , UNCONNECTED_24 , 
	UNCONNECTED_25 , UNCONNECTED_26 , UNCONNECTED_27 , UNCONNECTED_28 , 
	UNCONNECTED_29 , UNCONNECTED_30 , UNCONNECTED_31 , UNCONNECTED_32 , 
	UNCONNECTED_33 , UNCONNECTED_34 , UNCONNECTED_35 , UNCONNECTED_36 , 
	UNCONNECTED_37 , UNCONNECTED_38 , UNCONNECTED_39 , UNCONNECTED_40 , 
	UNCONNECTED_41 , UNCONNECTED_42 , UNCONNECTED_43 , UNCONNECTED_44 , 
	UNCONNECTED_45 , UNCONNECTED_46 , UNCONNECTED_47 , UNCONNECTED_48 , 
	UNCONNECTED_49 , UNCONNECTED_50 , UNCONNECTED_51 , UNCONNECTED_52 , 
	UNCONNECTED_53 , UNCONNECTED_54 , UNCONNECTED_55 , UNCONNECTED_56 , 
	UNCONNECTED_57 , UNCONNECTED_58 , UNCONNECTED_59 , UNCONNECTED_60 , 
	UNCONNECTED_61 , UNCONNECTED_62 , UNCONNECTED_63 , UNCONNECTED_64 , 
	UNCONNECTED_65 , UNCONNECTED_66 , UNCONNECTED_67 , UNCONNECTED_68 , 
	UNCONNECTED_69 , UNCONNECTED_70 , UNCONNECTED_71 , UNCONNECTED_72 , 
	UNCONNECTED_73 , UNCONNECTED_74 , UNCONNECTED_75 , UNCONNECTED_76 , 
	UNCONNECTED_77 , UNCONNECTED_78 , UNCONNECTED_79 , UNCONNECTED_80 , 
	UNCONNECTED_81 , UNCONNECTED_82 , UNCONNECTED_83 , UNCONNECTED_84 , 
	UNCONNECTED_85 , UNCONNECTED_86 , UNCONNECTED_87 , UNCONNECTED_88 , 
	UNCONNECTED_89 , UNCONNECTED_90 , UNCONNECTED_91 , UNCONNECTED_92 , 
	UNCONNECTED_93 , UNCONNECTED_94 , UNCONNECTED_95 , UNCONNECTED_96 , 
	UNCONNECTED_97 , UNCONNECTED_98 , UNCONNECTED_99 , UNCONNECTED_100 , 
	UNCONNECTED_101 , UNCONNECTED_102 , UNCONNECTED_103 , UNCONNECTED_104 , 
	UNCONNECTED_105 , UNCONNECTED_106 , UNCONNECTED_107 , UNCONNECTED_108 , 
	UNCONNECTED_109 , UNCONNECTED_110 , UNCONNECTED_111 , UNCONNECTED_112 , 
	UNCONNECTED_113 , UNCONNECTED_114 , UNCONNECTED_115 , UNCONNECTED_116 , 
	UNCONNECTED_117 , UNCONNECTED_118 , UNCONNECTED_119 , UNCONNECTED_120 , 
	UNCONNECTED_121 , UNCONNECTED_122 , UNCONNECTED_123 , UNCONNECTED_124 , 
	UNCONNECTED_125 , UNCONNECTED_126 , UNCONNECTED_127 , UNCONNECTED_128 ;
    VMW_PULLDOWN U36 ( .Z(n1539) );
    VMW_PULLDOWN U37 ( .Z(n1532) );
    VMW_PULLDOWN U39 ( .Z(n1554) );
    VMW_PULLDOWN U40 ( .Z(n1537) );
    VMW_PULLDOWN U41 ( .Z(n1534) );
    VMW_PULLDOWN U46 ( .Z(n1561) );
    VMW_PULLDOWN U54 ( .Z(n1562) );
    VMW_PULLDOWN U61 ( .Z(n1547) );
    VMW_FD \cOutput_reg[6]  ( .D(\result60[6] ), .CP(Clk), .Q(cOutput[6]) );
    VMW_FD \cOutput_reg[2]  ( .D(\result60[2] ), .CP(Clk), .Q(cOutput[2]) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_8 add_48_11 ( .A({
        \result997[7] , \result997[6] , \result997[5] , \result997[4] , 
        \result997[3] , \result997[2] , \result997[1] , \n995[8] }), .B({
        \n1087[1] , \n1087[2] , \n1087[3] , \n1087[4] , \n1087[5] , \n1087[6] , 
        \n1087[7] , \n1087[8] }), .CI(n1549), .SUM({\result1086[7] , 
        \result1086[6] , \result1086[5] , \result1086[4] , \result1086[3] , 
        \result1086[2] , \result1086[1] , \result1086[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_5 mul_48_6 ( .A(
        vectorAInput[55:48]), .B(vectorBInput[55:48]), .TC(n1544), .PRODUCT({
        UNCONNECTED_1, UNCONNECTED_2, UNCONNECTED_3, UNCONNECTED_4, 
        UNCONNECTED_5, UNCONNECTED_6, UNCONNECTED_7, UNCONNECTED_8, \n642[1] , 
        \n642[2] , \n642[3] , \n642[4] , \n642[5] , \n642[6] , \n642[7] , 
        \n642[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_1 add_48_8 ( .A({
        \result730[7] , \result730[6] , \result730[5] , \result730[4] , 
        \result730[3] , \result730[2] , \result730[1] , \result730[0] }), .B({
        \n820[1] , \n820[2] , \n820[3] , \n820[4] , \n820[5] , \n820[6] , 
        \n820[7] , \n820[8] }), .CI(n1533), .SUM({\result819[7] , 
        \result819[6] , \result819[5] , \result819[4] , \result819[3] , 
        \result819[2] , \n817[7] , \result819[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_6 add_48_1 ( .A({
        \n106[1] , \n106[2] , \n106[3] , \n106[4] , \n106[5] , \n106[6] , 
        \n106[7] , \n106[8] }), .B({\n197[1] , \n197[2] , \n197[3] , \n197[4] , 
        \n197[5] , \n197[6] , \n197[7] , \n197[8] }), .CI(n1542), .SUM({
        \result196[7] , \result196[6] , \result196[5] , \result196[4] , 
        \result196[3] , \result196[2] , \result196[1] , \result196[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_14 add_48_6 ( .A({
        \result552[7] , \result552[6] , \result552[5] , \result552[4] , 
        \result552[3] , \result552[2] , \result552[1] , \result552[0] }), .B({
        \n642[1] , \n642[2] , \n642[3] , \n642[4] , \n642[5] , \n642[6] , 
        \n642[7] , \n642[8] }), .CI(n1562), .SUM({\result641[7] , 
        \result641[6] , \result641[5] , \result641[4] , \result641[3] , 
        \result641[2] , \result641[1] , \result641[0] }) );
    VMW_PULLDOWN U48 ( .Z(n1546) );
    VMW_PULLDOWN U66 ( .Z(n1557) );
    VMW_FD \cOutput_reg[4]  ( .D(\result60[4] ), .CP(Clk), .Q(cOutput[4]) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_9 mul_48_1 ( .A(
        vectorAInput[15:8]), .B(vectorBInput[15:8]), .TC(n1550), .PRODUCT({
        UNCONNECTED_9, UNCONNECTED_10, UNCONNECTED_11, UNCONNECTED_12, 
        UNCONNECTED_13, UNCONNECTED_14, UNCONNECTED_15, UNCONNECTED_16, 
        \n197[1] , \n197[2] , \n197[3] , \n197[4] , \n197[5] , \n197[6] , 
        \n197[7] , \n197[8] }) );
    VMW_PULLDOWN U53 ( .Z(n1541) );
    VMW_FD \cOutput_reg[0]  ( .D(\result60[0] ), .CP(Clk), .Q(cOutput[0]) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_12 mul_48_8 ( .A(
        vectorAInput[71:64]), .B(vectorBInput[71:64]), .TC(n1555), .PRODUCT({
        UNCONNECTED_17, UNCONNECTED_18, UNCONNECTED_19, UNCONNECTED_20, 
        UNCONNECTED_21, UNCONNECTED_22, UNCONNECTED_23, UNCONNECTED_24, 
        \n820[1] , \n820[2] , \n820[3] , \n820[4] , \n820[5] , \n820[6] , 
        \n820[7] , \n820[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_11 add_48_7 ( .A({
        \result641[7] , \result641[6] , \result641[5] , \result641[4] , 
        \result641[3] , \result641[2] , \result641[1] , \result641[0] }), .B({
        \n731[1] , \n731[2] , \n731[3] , \n731[4] , \n731[5] , \n731[6] , 
        \n731[7] , \n731[8] }), .CI(n1558), .SUM({\result730[7] , 
        \result730[6] , \result730[5] , \result730[4] , \result730[3] , 
        \result730[2] , \result730[1] , \result730[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_4 mul_48_11 ( .A(
        vectorAInput[95:88]), .B(vectorBInput[95:88]), .TC(n1543), .PRODUCT({
        UNCONNECTED_25, UNCONNECTED_26, UNCONNECTED_27, UNCONNECTED_28, 
        UNCONNECTED_29, UNCONNECTED_30, UNCONNECTED_31, UNCONNECTED_32, 
        \n1087[1] , \n1087[2] , \n1087[3] , \n1087[4] , \n1087[5] , \n1087[6] , 
        \n1087[7] , \n1087[8] }) );
    VMW_PULLDOWN U47 ( .Z(n1540) );
    VMW_PULLDOWN U49 ( .Z(n1552) );
    VMW_PULLDOWN U52 ( .Z(n1558) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_10 mul_48_9 ( .A(
        vectorAInput[79:72]), .B(vectorBInput[79:72]), .TC(n1552), .PRODUCT({
        UNCONNECTED_33, UNCONNECTED_34, UNCONNECTED_35, UNCONNECTED_36, 
        UNCONNECTED_37, UNCONNECTED_38, UNCONNECTED_39, UNCONNECTED_40, 
        \n909[1] , \n909[2] , \n909[3] , \n909[4] , \n909[5] , \n909[6] , 
        \n909[7] , \n909[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_14 mul_48 ( .A(
        vectorAInput[7:0]), .B(vectorBInput[7:0]), .TC(n1557), .PRODUCT({
        UNCONNECTED_41, UNCONNECTED_42, UNCONNECTED_43, UNCONNECTED_44, 
        UNCONNECTED_45, UNCONNECTED_46, UNCONNECTED_47, UNCONNECTED_48, 
        \n106[1] , \n106[2] , \n106[3] , \n106[4] , \n106[5] , \n106[6] , 
        \n106[7] , \n106[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_2 mul_48_10 ( .A(
        vectorAInput[87:80]), .B(vectorBInput[87:80]), .TC(n1540), .PRODUCT({
        UNCONNECTED_49, UNCONNECTED_50, UNCONNECTED_51, UNCONNECTED_52, 
        UNCONNECTED_53, UNCONNECTED_54, UNCONNECTED_55, UNCONNECTED_56, 
        \n998[1] , \n998[2] , \n998[3] , \n998[4] , \n998[5] , \n998[6] , 
        \n998[7] , \n998[8] }) );
    VMW_PULLDOWN U55 ( .Z(n1544) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_13 add_48_10 ( .A({
        \result908[7] , \result908[6] , \result908[5] , \result908[4] , 
        \result908[3] , \result908[2] , \result908[1] , \n906[8] }), .B({
        \n998[1] , \n998[2] , \n998[3] , \n998[4] , \n998[5] , \n998[6] , 
        \n998[7] , \n998[8] }), .CI(n1561), .SUM({\result997[7] , 
        \result997[6] , \result997[5] , \result997[4] , \result997[3] , 
        \result997[2] , \result997[1] , \n995[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_7 add_48_9 ( .A({
        \result819[7] , \result819[6] , \result819[5] , \result819[4] , 
        \result819[3] , \result819[2] , \n817[7] , \result819[0] }), .B({
        \n909[1] , \n909[2] , \n909[3] , \n909[4] , \n909[5] , \n909[6] , 
        \n909[7] , \n909[8] }), .CI(n1546), .SUM({\result908[7] , 
        \result908[6] , \result908[5] , \result908[4] , \result908[3] , 
        \result908[2] , \result908[1] , \n906[8] }) );
    VMW_PULLDOWN U60 ( .Z(n1551) );
    VMW_PULLDOWN U57 ( .Z(n1556) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_15 mul_48_15 ( .A(
        vectorAInput[127:120]), .B(vectorBInput[127:120]), .TC(n1559), 
        .PRODUCT({UNCONNECTED_57, UNCONNECTED_58, UNCONNECTED_59, 
        UNCONNECTED_60, UNCONNECTED_61, UNCONNECTED_62, UNCONNECTED_63, 
        UNCONNECTED_64, \n1442[1] , \n1442[2] , \n1442[3] , \n1442[4] , 
        \n1442[5] , \n1442[6] , \n1442[7] , \n1442[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_3 mul_48_7 ( .A(
        vectorAInput[63:56]), .B(vectorBInput[63:56]), .TC(n1541), .PRODUCT({
        UNCONNECTED_65, UNCONNECTED_66, UNCONNECTED_67, UNCONNECTED_68, 
        UNCONNECTED_69, UNCONNECTED_70, UNCONNECTED_71, UNCONNECTED_72, 
        \n731[1] , \n731[2] , \n731[3] , \n731[4] , \n731[5] , \n731[6] , 
        \n731[7] , \n731[8] }) );
    VMW_PULLDOWN U42 ( .Z(n1545) );
    VMW_PULLDOWN U45 ( .Z(n1559) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_13 mul_48_5 ( .A(
        vectorAInput[47:40]), .B(vectorBInput[47:40]), .TC(n1556), .PRODUCT({
        UNCONNECTED_73, UNCONNECTED_74, UNCONNECTED_75, UNCONNECTED_76, 
        UNCONNECTED_77, UNCONNECTED_78, UNCONNECTED_79, UNCONNECTED_80, 
        \n553[1] , \n553[2] , \n553[3] , \n553[4] , \n553[5] , \n553[6] , 
        \n553[7] , \n553[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_2 add_48_12 ( .A({
        \result1086[7] , \result1086[6] , \result1086[5] , \result1086[4] , 
        \result1086[3] , \result1086[2] , \result1086[1] , \result1086[0] }), 
        .B({\n1176[1] , \n1176[2] , \n1176[3] , \n1176[4] , \n1176[5] , 
        \n1176[6] , \n1176[7] , \n1176[8] }), .CI(n1534), .SUM({
        \result1175[7] , \result1175[6] , \result1175[5] , \result1175[4] , 
        \result1175[3] , \result1175[2] , \result1175[1] , \result1175[0] })
         );
    VMW_PULLDOWN U62 ( .Z(n1560) );
    VMW_PULLDOWN U65 ( .Z(n1550) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_12 add_48_2 ( .A({
        \result196[7] , \result196[6] , \result196[5] , \result196[4] , 
        \result196[3] , \result196[2] , \result196[1] , \result196[0] }), .B({
        \n286[1] , \n286[2] , \n286[3] , \n286[4] , \n286[5] , \n286[6] , 
        \n286[7] , \n286[8] }), .CI(n1560), .SUM({\result285[7] , 
        \result285[6] , \result285[5] , \result285[4] , \result285[3] , 
        \result285[2] , \result285[1] , \result285[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_4 add_48_5 ( .A({
        \result463[7] , \result463[6] , \result463[5] , \result463[4] , 
        \result463[3] , \result463[2] , \result463[1] , \result463[0] }), .B({
        \n553[1] , \n553[2] , \n553[3] , \n553[4] , \n553[5] , \n553[6] , 
        \n553[7] , \n553[8] }), .CI(n1538), .SUM({\result552[7] , 
        \result552[6] , \result552[5] , \result552[4] , \result552[3] , 
        \result552[2] , \result552[1] , \result552[0] }) );
    VMW_PULLDOWN U50 ( .Z(n1533) );
    VMW_PULLDOWN U59 ( .Z(n1553) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_6 mul_48_12 ( .A(
        vectorAInput[103:96]), .B(vectorBInput[103:96]), .TC(n1545), .PRODUCT(
        {UNCONNECTED_81, UNCONNECTED_82, UNCONNECTED_83, UNCONNECTED_84, 
        UNCONNECTED_85, UNCONNECTED_86, UNCONNECTED_87, UNCONNECTED_88, 
        \n1176[1] , \n1176[2] , \n1176[3] , \n1176[4] , \n1176[5] , \n1176[6] , 
        \n1176[7] , \n1176[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_5 add_48_15 ( .A({
        \result1353[7] , \result1353[6] , \result1353[5] , \result1353[4] , 
        \result1353[3] , \n1351[6] , \result1353[1] , \result1353[0] }), .B({
        \n1442[1] , \n1442[2] , \n1442[3] , \n1442[4] , \n1442[5] , \n1442[6] , 
        \n1442[7] , \n1442[8] }), .CI(n1539), .SUM({\result60[7] , 
        \result60[6] , \result60[5] , \result60[4] , \result60[3] , 
        \result60[2] , \result60[1] , \result60[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_0 mul_48_2 ( .A(
        vectorAInput[23:16]), .B(vectorBInput[23:16]), .TC(n1536), .PRODUCT({
        UNCONNECTED_89, UNCONNECTED_90, UNCONNECTED_91, UNCONNECTED_92, 
        UNCONNECTED_93, UNCONNECTED_94, UNCONNECTED_95, UNCONNECTED_96, 
        \n286[1] , \n286[2] , \n286[3] , \n286[4] , \n286[5] , \n286[6] , 
        \n286[7] , \n286[8] }) );
    VMW_PULLDOWN U58 ( .Z(n1535) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_7 mul_48_3 ( .A(
        vectorAInput[31:24]), .B(vectorBInput[31:24]), .TC(n1547), .PRODUCT({
        UNCONNECTED_97, UNCONNECTED_98, UNCONNECTED_99, UNCONNECTED_100, 
        UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, UNCONNECTED_104, 
        \n375[1] , \n375[2] , \n375[3] , \n375[4] , \n375[5] , \n375[6] , 
        \n375[7] , \n375[8] }) );
    VMW_PULLDOWN U38 ( .Z(n1548) );
    VMW_PULLDOWN U43 ( .Z(n1549) );
    VMW_PULLDOWN U64 ( .Z(n1542) );
    VMW_FD \cOutput_reg[1]  ( .D(\result60[1] ), .CP(Clk), .Q(cOutput[1]) );
    VMW_PULLDOWN U51 ( .Z(n1555) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_1 mul_48_13 ( .A(
        vectorAInput[111:104]), .B(vectorBInput[111:104]), .TC(n1537), 
        .PRODUCT({UNCONNECTED_105, UNCONNECTED_106, UNCONNECTED_107, 
        UNCONNECTED_108, UNCONNECTED_109, UNCONNECTED_110, UNCONNECTED_111, 
        UNCONNECTED_112, \n1265[1] , \n1265[2] , \n1265[3] , \n1265[4] , 
        \n1265[5] , \n1265[6] , \n1265[7] , \n1265[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_3 add_48_4 ( .A({
        \result374[7] , \result374[6] , \result374[5] , \result374[4] , 
        \result374[3] , \result374[2] , \result374[1] , \result374[0] }), .B({
        \n464[1] , \n464[2] , \n464[3] , \n464[4] , \n464[5] , \n464[6] , 
        \n464[7] , \n464[8] }), .CI(n1535), .SUM({\result463[7] , 
        \result463[6] , \result463[5] , \result463[4] , \result463[3] , 
        \result463[2] , \result463[1] , \result463[0] }) );
    VMW_FD \cOutput_reg[7]  ( .D(\result60[7] ), .CP(Clk), .Q(cOutput[7]) );
    VMW_FD \cOutput_reg[5]  ( .D(\result60[5] ), .CP(Clk), .Q(cOutput[5]) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_0 add_48_14 ( .A({
        \result1264[7] , \result1264[6] , \result1264[5] , \n1262[4] , 
        \result1264[3] , \result1264[2] , \result1264[1] , \result1264[0] }), 
        .B({\n1354[1] , \n1354[2] , \n1354[3] , \n1354[4] , \n1354[5] , 
        \n1354[6] , \n1354[7] , \n1354[8] }), .CI(n1532), .SUM({
        \result1353[7] , \result1353[6] , \result1353[5] , \result1353[4] , 
        \result1353[3] , \n1351[6] , \result1353[1] , \result1353[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_10 add_48_13 ( .A({
        \result1175[7] , \result1175[6] , \result1175[5] , \result1175[4] , 
        \result1175[3] , \result1175[2] , \result1175[1] , \result1175[0] }), 
        .B({\n1265[1] , \n1265[2] , \n1265[3] , \n1265[4] , \n1265[5] , 
        \n1265[6] , \n1265[7] , \n1265[8] }), .CI(n1554), .SUM({
        \result1264[7] , \result1264[6] , \result1264[5] , \n1262[4] , 
        \result1264[3] , \result1264[2] , \result1264[1] , \result1264[0] })
         );
    VMW_PULLDOWN U44 ( .Z(n1543) );
    VMW_PULLDOWN U56 ( .Z(n1538) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_8 mul_48_14 ( .A(
        vectorAInput[119:112]), .B(vectorBInput[119:112]), .TC(n1548), 
        .PRODUCT({UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
        UNCONNECTED_116, UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119, 
        UNCONNECTED_120, \n1354[1] , \n1354[2] , \n1354[3] , \n1354[4] , 
        \n1354[5] , \n1354[6] , \n1354[7] , \n1354[8] }) );
    VMW_PULLDOWN U63 ( .Z(n1536) );
    VMW_FD \cOutput_reg[3]  ( .D(\result60[3] ), .CP(Clk), .Q(cOutput[3]) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW01_add_8_9 add_48_3 ( .A({
        \result285[7] , \result285[6] , \result285[5] , \result285[4] , 
        \result285[3] , \result285[2] , \result285[1] , \result285[0] }), .B({
        \n375[1] , \n375[2] , \n375[3] , \n375[4] , \n375[5] , \n375[6] , 
        \n375[7] , \n375[8] }), .CI(n1551), .SUM({\result374[7] , 
        \result374[6] , \result374[5] , \result374[4] , \result374[3] , 
        \result374[2] , \result374[1] , \result374[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8_DW02_mult_8_8_11 mul_48_4 ( .A(
        vectorAInput[39:32]), .B(vectorBInput[39:32]), .TC(n1553), .PRODUCT({
        UNCONNECTED_121, UNCONNECTED_122, UNCONNECTED_123, UNCONNECTED_124, 
        UNCONNECTED_125, UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
        \n464[1] , \n464[2] , \n464[3] , \n464[4] , \n464[5] , \n464[6] , 
        \n464[7] , \n464[8] }) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \matrixInput[1879] , \matrixInput[954] , \matrixInput[1860] , 
        \matrixInput[1853] , \matrixInput[53] , \vectorInput[83] , 
        \matrixInput[1724] , \matrixInput[1687] , \matrixInput[1584] , 
        \matrixInput[1230] , \matrixInput[1229] , \matrixInput[1133] , 
        \matrixInput[967] , \matrixInput[79] , \matrixInput[60] , 
        \cOutput[67] , \cOutput[54] , \matrixInput[799] , \matrixInput[483] , 
        \matrixInput[780] , \matrixInput[304] , \matrixInput[1203] , 
        \matrixInput[1119] , \matrixInput[1100] , \matrixInput[337] , 
        \matrixInput[610] , \matrixInput[609] , \matrixInput[1717] , 
        \matrixInput[1427] , \matrixInput[513] , \matrixInput[294] , 
        \matrixInput[197] , \matrixInput[1393] , \vectorInput[51] , 
        \matrixInput[2032] , \matrixInput[1922] , \matrixInput[1911] , 
        \matrixInput[1898] , \matrixInput[1881] , \matrixInput[1414] , 
        \matrixInput[623] , \matrixInput[1090] , \matrixInput[539] , 
        \matrixInput[520] , \matrixInput[1089] , \matrixInput[986] , 
        \matrixInput[98] , \matrixInput[81] , \matrixInput[1908] , 
        \matrixInput[825] , \matrixInput[816] , \cOutput[86] , 
        \matrixInput[1655] , \matrixInput[778] , \matrixInput[761] , 
        \matrixInput[2018] , \matrixInput[2001] , \matrixInput[1666] , 
        \matrixInput[1556] , \matrixInput[752] , \matrixInput[462] , 
        \matrixInput[1565] , \matrixInput[451] , \matrixInput[448] , 
        \matrixInput[1042] , \matrixInput[176] , \vectorInput[48] , 
        \matrixInput[1358] , \matrixInput[1341] , \matrixInput[275] , 
        \matrixInput[145] , \vectorInput[93] , \vectorInput[72] , 
        \vectorInput[62] , \matrixInput[1372] , \matrixInput[1071] , 
        \matrixInput[1068] , \matrixInput[246] , \matrixInput[1932] , 
        \matrixInput[1918] , \matrixInput[835] , \matrixInput[806] , 
        \matrixInput[1901] , \matrixInput[1891] , \matrixInput[1888] , 
        \matrixInput[996] , \matrixInput[91] , \cOutput[96] , 
        \matrixInput[88] , \matrixInput[1362] , \matrixInput[1078] , 
        \matrixInput[1061] , \matrixInput[155] , \matrixInput[256] , 
        \vectorInput[58] , \matrixInput[1052] , \matrixInput[166] , 
        \vectorInput[41] , \matrixInput[2022] , \matrixInput[2011] , 
        \matrixInput[2008] , \matrixInput[1676] , \matrixInput[1351] , 
        \matrixInput[1348] , \matrixInput[265] , \matrixInput[1575] , 
        \matrixInput[742] , \matrixInput[458] , \matrixInput[441] , 
        \matrixInput[1645] , \matrixInput[771] , \matrixInput[768] , 
        \matrixInput[1870] , \matrixInput[1843] , \matrixInput[1546] , 
        \matrixInput[472] , \matrixInput[977] , \cOutput[77] , \cOutput[44] , 
        \matrixInput[70] , \matrixInput[69] , \matrixInput[1869] , 
        \matrixInput[1383] , \matrixInput[944] , \matrixInput[43] , 
        \matrixInput[633] , \matrixInput[1734] , \matrixInput[1707] , 
        \matrixInput[1404] , \matrixInput[530] , \matrixInput[529] , 
        \matrixInput[1099] , \matrixInput[1080] , \cOutput[6] , 
        \matrixInput[619] , \matrixInput[600] , \vectorInput[66] , 
        \vectorInput[55] , \matrixInput[1697] , \matrixInput[1594] , 
        \matrixInput[1437] , \matrixInput[284] , \matrixInput[187] , 
        \matrixInput[503] , \matrixInput[1213] , \matrixInput[1110] , 
        \matrixInput[1109] , \matrixInput[327] , \matrixInput[1345] , 
        \matrixInput[1239] , \matrixInput[1220] , \matrixInput[1123] , 
        \matrixInput[790] , \matrixInput[493] , \matrixInput[789] , 
        \matrixInput[314] , \matrixInput[271] , \matrixInput[268] , 
        \matrixInput[1046] , \matrixInput[172] , \matrixInput[1376] , 
        \matrixInput[1075] , \matrixInput[242] , \vectorInput[87] , 
        \matrixInput[2036] , \matrixInput[1552] , \matrixInput[466] , 
        \matrixInput[158] , \matrixInput[141] , \matrixInput[2005] , 
        \matrixInput[1651] , \matrixInput[765] , \matrixInput[1648] , 
        \matrixInput[1926] , \matrixInput[1915] , \matrixInput[1662] , 
        \matrixInput[1578] , \matrixInput[1561] , \matrixInput[455] , 
        \matrixInput[838] , \matrixInput[821] , \matrixInput[756] , 
        \cOutput[82] , \matrixInput[1885] , \matrixInput[812] , 
        \matrixInput[1739] , \matrixInput[1423] , \matrixInput[982] , 
        \matrixInput[85] , \matrixInput[517] , \matrixInput[290] , 
        \matrixInput[289] , \matrixInput[193] , \matrixInput[1720] , 
        \matrixInput[1410] , \matrixInput[1094] , \matrixInput[614] , 
        \matrixInput[524] , \matrixInput[1409] , \matrixInput[627] , 
        \matrixInput[1864] , \matrixInput[1713] , \matrixInput[1683] , 
        \matrixInput[1397] , \matrixInput[1234] , \matrixInput[1137] , 
        \matrixInput[784] , \matrixInput[319] , \matrixInput[300] , 
        \matrixInput[487] , \matrixInput[1599] , \matrixInput[1580] , 
        \matrixInput[1207] , \matrixInput[333] , \matrixInput[1104] , 
        \matrixInput[57] , \cOutput[63] , \cOutput[50] , \cOutput[49] , 
        \matrixInput[1857] , \matrixInput[963] , \matrixInput[950] , 
        \matrixInput[949] , \matrixInput[64] , \vectorInput[97] , 
        \matrixInput[1703] , \matrixInput[1693] , \matrixInput[1590] , 
        \matrixInput[1589] , \matrixInput[1217] , \matrixInput[1114] , 
        \matrixInput[323] , \matrixInput[1419] , \matrixInput[1224] , 
        \matrixInput[310] , \matrixInput[309] , \matrixInput[1127] , 
        \matrixInput[794] , \matrixInput[497] , \matrixInput[1084] , 
        \matrixInput[1400] , \matrixInput[534] , \matrixInput[1730] , 
        \matrixInput[1433] , \matrixInput[1387] , \matrixInput[637] , 
        \matrixInput[507] , \matrixInput[604] , \matrixInput[299] , 
        \matrixInput[280] , \matrixInput[183] , \matrixInput[1729] , 
        \cOutput[2] , \matrixInput[74] , \vectorInput[76] , 
        \matrixInput[2026] , \matrixInput[2015] , \matrixInput[1874] , 
        \matrixInput[1847] , \matrixInput[973] , \matrixInput[959] , 
        \matrixInput[940] , \matrixInput[47] , \cOutput[73] , \cOutput[59] , 
        \cOutput[40] , \matrixInput[1672] , \matrixInput[1571] , 
        \matrixInput[445] , \matrixInput[1568] , \matrixInput[746] , 
        \matrixInput[1542] , \matrixInput[476] , \matrixInput[1658] , 
        \matrixInput[1641] , \matrixInput[775] , \matrixInput[1366] , 
        \matrixInput[252] , \vectorInput[95] , \vectorInput[74] , 
        \vectorInput[45] , \matrixInput[1355] , \matrixInput[1065] , 
        \matrixInput[151] , \matrixInput[148] , \matrixInput[278] , 
        \matrixInput[261] , \matrixInput[2024] , \matrixInput[2017] , 
        \matrixInput[1936] , \matrixInput[1895] , \matrixInput[1056] , 
        \matrixInput[992] , \matrixInput[162] , \matrixInput[95] , 
        \matrixInput[802] , \matrixInput[1905] , \cOutput[92] , 
        \matrixInput[1670] , \matrixInput[1669] , \matrixInput[831] , 
        \matrixInput[828] , \matrixInput[1573] , \matrixInput[744] , 
        \matrixInput[447] , \matrixInput[1643] , \matrixInput[777] , 
        \matrixInput[1559] , \matrixInput[1540] , \matrixInput[474] , 
        \matrixInput[1364] , \matrixInput[1067] , \matrixInput[153] , 
        \matrixInput[250] , \matrixInput[249] , \vectorInput[47] , 
        \matrixInput[1054] , \matrixInput[179] , \matrixInput[160] , 
        \matrixInput[1934] , \matrixInput[1897] , \matrixInput[1357] , 
        \matrixInput[263] , \matrixInput[990] , \matrixInput[989] , 
        \matrixInput[97] , \matrixInput[1907] , \matrixInput[833] , 
        \matrixInput[819] , \matrixInput[800] , \matrixInput[1701] , 
        \matrixInput[1691] , \matrixInput[1592] , \cOutput[90] , \cOutput[89] , 
        \matrixInput[1215] , \matrixInput[1116] , \matrixInput[338] , 
        \matrixInput[321] , \matrixInput[1688] , \matrixInput[1385] , 
        \matrixInput[1226] , \matrixInput[1125] , \matrixInput[796] , 
        \matrixInput[495] , \matrixInput[312] , \matrixInput[635] , 
        \matrixInput[1845] , \matrixInput[1732] , \matrixInput[1718] , 
        \matrixInput[1402] , \matrixInput[536] , \matrixInput[1086] , 
        \matrixInput[1431] , \matrixInput[1428] , \matrixInput[606] , 
        \cOutput[0] , \matrixInput[282] , \matrixInput[198] , 
        \matrixInput[181] , \matrixInput[971] , \matrixInput[505] , 
        \matrixInput[968] , \matrixInput[76] , \matrixInput[1876] , 
        \vectorInput[85] , \matrixInput[1722] , \matrixInput[942] , 
        \matrixInput[616] , \matrixInput[45] , \cOutput[71] , \cOutput[42] , 
        \cOutput[68] , \cOutput[9] , \matrixInput[1438] , \matrixInput[1421] , 
        \matrixInput[515] , \matrixInput[292] , \matrixInput[191] , 
        \matrixInput[188] , \matrixInput[1395] , \matrixInput[1866] , 
        \matrixInput[1711] , \matrixInput[1708] , \matrixInput[1698] , 
        \matrixInput[1582] , \matrixInput[1412] , \matrixInput[625] , 
        \matrixInput[1236] , \matrixInput[1135] , \matrixInput[1096] , 
        \matrixInput[526] , \matrixInput[786] , \matrixInput[485] , 
        \matrixInput[302] , \matrixInput[1205] , \matrixInput[1106] , 
        \matrixInput[331] , \matrixInput[328] , \matrixInput[1681] , 
        \matrixInput[952] , \cOutput[78] , \cOutput[61] , \cOutput[52] , 
        \matrixInput[1855] , \matrixInput[55] , \vectorInput[57] , 
        \matrixInput[1044] , \matrixInput[978] , \matrixInput[961] , 
        \matrixInput[66] , \matrixInput[170] , \matrixInput[169] , 
        \matrixInput[1347] , \matrixInput[273] , \vectorInput[91] , 
        \vectorInput[64] , \matrixInput[1374] , \matrixInput[1077] , 
        \matrixInput[143] , \matrixInput[259] , \matrixInput[240] , 
        \matrixInput[2034] , \matrixInput[1653] , \matrixInput[767] , 
        \matrixInput[2007] , \matrixInput[1679] , \matrixInput[1660] , 
        \matrixInput[1550] , \matrixInput[1549] , \matrixInput[754] , 
        \matrixInput[464] , \matrixInput[1563] , \matrixInput[457] , 
        \matrixInput[1924] , \matrixInput[1917] , \matrixInput[823] , 
        \matrixInput[810] , \cOutput[99] , \cOutput[80] , \matrixInput[809] , 
        \matrixInput[1887] , \matrixInput[1872] , \matrixInput[1858] , 
        \matrixInput[1841] , \matrixInput[999] , \matrixInput[980] , 
        \matrixInput[87] , \matrixInput[72] , \cOutput[75] , \cOutput[46] , 
        \matrixInput[975] , \matrixInput[946] , \matrixInput[58] , 
        \matrixInput[41] , \matrixInput[1406] , \matrixInput[1082] , 
        \matrixInput[532] , \vectorInput[88] , \matrixInput[1705] , 
        \matrixInput[1435] , \matrixInput[1398] , \matrixInput[1381] , 
        \matrixInput[631] , \matrixInput[628] , \matrixInput[518] , 
        \matrixInput[501] , \matrixInput[185] , \vectorInput[79] , 
        \vectorInput[70] , \vectorInput[69] , \matrixInput[1930] , 
        \matrixInput[1929] , \matrixInput[1736] , \matrixInput[602] , 
        \matrixInput[286] , \cOutput[4] , \matrixInput[1695] , 
        \matrixInput[1596] , \matrixInput[1211] , \matrixInput[1208] , 
        \matrixInput[1112] , \matrixInput[325] , \matrixInput[1222] , 
        \matrixInput[316] , \matrixInput[1138] , \matrixInput[792] , 
        \matrixInput[491] , \matrixInput[488] , \matrixInput[1121] , 
        \matrixInput[804] , \matrixInput[1903] , \cOutput[94] , 
        \matrixInput[1893] , \matrixInput[994] , \matrixInput[837] , 
        \matrixInput[93] , \vectorInput[60] , \vectorInput[53] , 
        \vectorInput[43] , \matrixInput[1379] , \matrixInput[254] , 
        \matrixInput[1360] , \matrixInput[1353] , \matrixInput[1063] , 
        \matrixInput[157] , \matrixInput[267] , \matrixInput[2039] , 
        \matrixInput[2013] , \matrixInput[1050] , \matrixInput[1049] , 
        \matrixInput[164] , \matrixInput[1674] , \matrixInput[1577] , 
        \matrixInput[443] , \matrixInput[759] , \matrixInput[740] , 
        \matrixInput[1544] , \matrixInput[470] , \matrixInput[469] , 
        \matrixInput[2030] , \matrixInput[2020] , \matrixInput[1939] , 
        \matrixInput[1920] , \matrixInput[1913] , \matrixInput[1883] , 
        \matrixInput[1647] , \matrixInput[773] , \matrixInput[984] , 
        \matrixInput[827] , \matrixInput[83] , \cOutput[84] , 
        \matrixInput[1554] , \matrixInput[814] , \matrixInput[479] , 
        \matrixInput[460] , \matrixInput[2029] , \matrixInput[2003] , 
        \matrixInput[1657] , \matrixInput[763] , \matrixInput[1664] , 
        \matrixInput[1567] , \matrixInput[453] , \matrixInput[1343] , 
        \matrixInput[750] , \matrixInput[749] , \matrixInput[277] , 
        \matrixInput[1059] , \matrixInput[174] , \matrixInput[1040] , 
        \matrixInput[1370] , \matrixInput[1369] , \matrixInput[1073] , 
        \matrixInput[244] , \matrixInput[147] , \matrixInput[1862] , 
        \matrixInput[51] , \matrixInput[48] , \matrixInput[1851] , 
        \matrixInput[1848] , \matrixInput[965] , \matrixInput[956] , 
        \matrixInput[62] , \vectorInput[98] , \matrixInput[1726] , 
        \matrixInput[1685] , \matrixInput[1232] , \cOutput[65] , \cOutput[56] , 
        \matrixInput[1131] , \matrixInput[782] , \matrixInput[306] , 
        \matrixInput[498] , \matrixInput[481] , \matrixInput[1128] , 
        \matrixInput[1586] , \matrixInput[1218] , \matrixInput[335] , 
        \matrixInput[1201] , \matrixInput[1102] , \matrixInput[1425] , 
        \matrixInput[511] , \matrixInput[508] , \matrixInput[296] , 
        \matrixInput[195] , \matrixInput[1416] , \matrixInput[1092] , 
        \matrixInput[612] , \matrixInput[522] , \matrixInput[638] , 
        \matrixInput[621] , \vectorInput[81] , \matrixInput[1715] , 
        \vectorInput[36] , \matrixInput[1391] , \matrixInput[1388] , 
        \matrixInput[696] , \matrixInput[1976] , \matrixInput[1791] , 
        \matrixInput[1326] , \matrixInput[1315] , \matrixInput[1025] , 
        \matrixInput[212] , \matrixInput[595] , \matrixInput[111] , 
        \matrixInput[108] , \matrixInput[238] , \matrixInput[221] , 
        \matrixInput[1788] , \matrixInput[1632] , \matrixInput[1531] , 
        \matrixInput[1528] , \matrixInput[1492] , \matrixInput[1016] , 
        \matrixInput[122] , \matrixInput[405] , \matrixInput[1618] , 
        \matrixInput[1601] , \matrixInput[1502] , \matrixInput[706] , 
        \matrixInput[436] , \matrixInput[382] , \matrixInput[1285] , 
        \matrixInput[1186] , \matrixInput[735] , \cOutput[106] , 
        \matrixInput[1945] , \matrixInput[871] , \matrixInput[842] , 
        \matrixInput[868] , \vectorInput[102] , \matrixInput[1770] , 
        \matrixInput[1769] , \matrixInput[1743] , \matrixInput[1459] , 
        \matrixInput[1440] , \matrixInput[574] , \matrixInput[677] , 
        \matrixInput[1473] , \matrixInput[547] , \matrixInput[1264] , 
        \matrixInput[1257] , \matrixInput[644] , \matrixInput[363] , 
        \matrixInput[1154] , \matrixInput[350] , \matrixInput[349] , 
        \matrixInput[1997] , \matrixInput[1167] , \matrixInput[889] , 
        \cOutput[19] , \vectorInput[3] , \matrixInput[1834] , 
        \matrixInput[1807] , \matrixInput[933] , \matrixInput[890] , 
        \matrixInput[34] , \matrixInput[7] , \cOutput[33] , 
        \matrixInput[1824] , \matrixInput[1779] , \matrixInput[1760] , 
        \matrixInput[1463] , \matrixInput[1274] , \matrixInput[919] , 
        \matrixInput[900] , \matrixInput[359] , \matrixInput[340] , 
        \matrixInput[1247] , \matrixInput[1177] , \matrixInput[1144] , 
        \matrixInput[373] , \matrixInput[557] , \matrixInput[654] , 
        \matrixInput[1753] , \matrixInput[1450] , \matrixInput[1449] , 
        \matrixInput[564] , \matrixInput[910] , \matrixInput[667] , 
        \matrixInput[17] , \matrixInput[909] , \matrixInput[1817] , 
        \matrixInput[24] , \matrixInput[923] , \matrixInput[899] , 
        \matrixInput[880] , \matrixInput[1987] , \cOutput[23] , \cOutput[10] , 
        \vectorInput[121] , \vectorInput[112] , \vectorInput[26] , 
        \vectorInput[15] , \matrixInput[2045] , \matrixInput[1611] , 
        \matrixInput[1608] , \matrixInput[1512] , \matrixInput[1295] , 
        \matrixInput[1196] , \matrixInput[426] , \matrixInput[725] , 
        \matrixInput[1798] , \matrixInput[1622] , \matrixInput[1538] , 
        \matrixInput[1521] , \matrixInput[415] , \matrixInput[716] , 
        \matrixInput[1305] , \matrixInput[392] , \matrixInput[231] , 
        \matrixInput[228] , \matrixInput[1781] , \matrixInput[1482] , 
        \matrixInput[1006] , \matrixInput[132] , \matrixInput[1336] , 
        \matrixInput[686] , \matrixInput[202] , \matrixInput[1035] , 
        \matrixInput[118] , \matrixInput[101] , \matrixInput[585] , 
        \matrixInput[1966] , \matrixInput[1955] , \cOutput[125] , 
        \matrixInput[878] , \matrixInput[861] , \matrixInput[852] , 
        \cOutput[116] , \matrixInput[1830] , \matrixInput[1829] , 
        \matrixInput[1803] , \matrixInput[937] , \matrixInput[904] , 
        \matrixInput[30] , \matrixInput[29] , \matrixInput[3] , 
        \matrixInput[1993] , \cOutput[37] , \vectorInput[106] , 
        \matrixInput[1774] , \matrixInput[1747] , \matrixInput[1279] , 
        \matrixInput[1253] , \matrixInput[1150] , \matrixInput[894] , 
        \matrixInput[1149] , \matrixInput[1163] , \matrixInput[367] , 
        \matrixInput[354] , \matrixInput[1260] , \matrixInput[1444] , 
        \matrixInput[673] , \matrixInput[659] , \matrixInput[570] , 
        \matrixInput[569] , \matrixInput[640] , \matrixInput[1477] , 
        \matrixInput[543] , \vectorInput[125] , \vectorInput[116] , 
        \vectorInput[32] , \matrixInput[1972] , \matrixInput[846] , 
        \matrixInput[1958] , \matrixInput[1941] , \cOutput[102] , 
        \matrixInput[1636] , \matrixInput[875] , \matrixInput[702] , 
        \matrixInput[386] , \matrixInput[1605] , \matrixInput[1535] , 
        \matrixInput[418] , \matrixInput[401] , \matrixInput[1506] , 
        \matrixInput[1298] , \matrixInput[1281] , \matrixInput[731] , 
        \matrixInput[728] , \matrixInput[1182] , \matrixInput[1322] , 
        \matrixInput[1038] , \matrixInput[591] , \matrixInput[588] , 
        \matrixInput[432] , \matrixInput[115] , \matrixInput[1021] , 
        \matrixInput[216] , \vectorInput[18] , \matrixInput[1795] , 
        \matrixInput[1496] , \matrixInput[1012] , \matrixInput[692] , 
        \matrixInput[126] , \matrixInput[1962] , \matrixInput[1951] , 
        \matrixInput[1948] , \matrixInput[1311] , \matrixInput[1308] , 
        \matrixInput[865] , \matrixInput[225] , \cOutput[121] , 
        \matrixInput[856] , \cOutput[112] , \vectorInput[22] , 
        \vectorInput[11] , \matrixInput[1785] , \matrixInput[1486] , 
        \matrixInput[1002] , \matrixInput[136] , \matrixInput[1332] , 
        \matrixInput[1318] , \matrixInput[235] , \matrixInput[1301] , 
        \matrixInput[1031] , \matrixInput[598] , \matrixInput[581] , 
        \matrixInput[1028] , \matrixInput[105] , \matrixInput[682] , 
        \matrixInput[206] , \matrixInput[2041] , \matrixInput[1626] , 
        \matrixInput[1615] , \matrixInput[738] , \matrixInput[721] , 
        \matrixInput[1516] , \matrixInput[1291] , \matrixInput[1288] , 
        \matrixInput[1192] , \matrixInput[422] , \matrixInput[396] , 
        \matrixInput[1525] , \matrixInput[712] , \matrixInput[411] , 
        \matrixInput[408] , \matrixInput[884] , \cOutput[27] , 
        \vectorInput[7] , \matrixInput[1983] , \cOutput[14] , 
        \matrixInput[1839] , \matrixInput[1820] , \matrixInput[914] , 
        \matrixInput[13] , \matrixInput[1813] , \matrixInput[927] , 
        \matrixInput[1764] , \matrixInput[39] , \matrixInput[20] , 
        \matrixInput[650] , \matrixInput[649] , \matrixInput[1998] , 
        \matrixInput[1981] , \matrixInput[1757] , \matrixInput[1467] , 
        \matrixInput[663] , \matrixInput[553] , \matrixInput[1454] , 
        \matrixInput[579] , \matrixInput[560] , \matrixInput[1270] , 
        \matrixInput[1173] , \matrixInput[1269] , \matrixInput[1243] , 
        \matrixInput[1159] , \matrixInput[344] , \matrixInput[1140] , 
        \matrixInput[377] , \matrixInput[886] , \cOutput[25] , 
        \vectorInput[5] , \matrixInput[1822] , \matrixInput[916] , 
        \matrixInput[11] , \cOutput[16] , \matrixInput[1811] , 
        \matrixInput[22] , \matrixInput[8] , \matrixInput[1808] , 
        \matrixInput[925] , \matrixInput[1979] , \matrixInput[1953] , 
        \matrixInput[1766] , \matrixInput[1465] , \matrixInput[551] , 
        \matrixInput[548] , \matrixInput[652] , \matrixInput[1755] , 
        \matrixInput[1456] , \matrixInput[562] , \matrixInput[1272] , 
        \matrixInput[678] , \matrixInput[661] , \matrixInput[346] , 
        \matrixInput[1258] , \matrixInput[1241] , \matrixInput[1171] , 
        \matrixInput[1168] , \matrixInput[1142] , \matrixInput[375] , 
        \cOutput[123] , \matrixInput[867] , \matrixInput[854] , \cOutput[110] , 
        \cOutput[109] , \matrixInput[1960] , \vectorInput[127] , 
        \vectorInput[114] , \vectorInput[39] , \vectorInput[13] , 
        \matrixInput[1787] , \matrixInput[1303] , \matrixInput[237] , 
        \matrixInput[1484] , \matrixInput[1019] , \matrixInput[1000] , 
        \matrixInput[134] , \vectorInput[20] , \matrixInput[2043] , 
        \matrixInput[1617] , \matrixInput[1514] , \matrixInput[1330] , 
        \matrixInput[1329] , \matrixInput[699] , \matrixInput[680] , 
        \matrixInput[204] , \matrixInput[1033] , \matrixInput[107] , 
        \matrixInput[583] , \matrixInput[1293] , \matrixInput[1190] , 
        \matrixInput[439] , \matrixInput[420] , \matrixInput[1189] , 
        \matrixInput[723] , \matrixInput[1624] , \matrixInput[1527] , 
        \matrixInput[413] , \matrixInput[710] , \matrixInput[709] , 
        \matrixInput[394] , \vectorInput[104] , \matrixInput[1970] , 
        \cOutput[119] , \cOutput[100] , \matrixInput[1969] , 
        \matrixInput[844] , \vectorInput[30] , \matrixInput[1943] , 
        \matrixInput[877] , \matrixInput[1634] , \matrixInput[1537] , 
        \matrixInput[403] , \matrixInput[1607] , \matrixInput[1504] , 
        \matrixInput[719] , \matrixInput[700] , \matrixInput[430] , 
        \matrixInput[429] , \matrixInput[384] , \matrixInput[1283] , 
        \matrixInput[1199] , \matrixInput[1180] , \matrixInput[733] , 
        \matrixInput[690] , \matrixInput[689] , \vectorInput[29] , 
        \matrixInput[1991] , \matrixInput[1988] , \matrixInput[1832] , 
        \matrixInput[1818] , \matrixInput[1797] , \matrixInput[1339] , 
        \matrixInput[1320] , \matrixInput[1313] , \matrixInput[1023] , 
        \matrixInput[214] , \matrixInput[593] , \matrixInput[117] , 
        \matrixInput[227] , \matrixInput[1494] , \matrixInput[1010] , 
        \matrixInput[1009] , \matrixInput[124] , \matrixInput[935] , 
        \matrixInput[32] , \matrixInput[1] , \matrixInput[1801] , 
        \matrixInput[18] , \matrixInput[906] , \matrixInput[896] , 
        \vectorInput[123] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[24] , \vectorInput[17] , \matrixInput[2047] , 
        \matrixInput[1776] , \matrixInput[1745] , \matrixInput[1446] , 
        \matrixInput[1262] , \matrixInput[1251] , \matrixInput[1248] , 
        \matrixInput[365] , \cOutput[35] , \matrixInput[1152] , 
        \matrixInput[1178] , \matrixInput[1161] , \matrixInput[356] , 
        \matrixInput[572] , \matrixInput[671] , \matrixInput[668] , 
        \matrixInput[1475] , \matrixInput[558] , \matrixInput[541] , 
        \matrixInput[1639] , \matrixInput[1613] , \matrixInput[727] , 
        \matrixInput[642] , \matrixInput[1510] , \matrixInput[1297] , 
        \matrixInput[1194] , \matrixInput[424] , \matrixInput[1509] , 
        \matrixInput[390] , \matrixInput[389] , \matrixInput[1620] , 
        \matrixInput[1523] , \matrixInput[714] , \matrixInput[417] , 
        \matrixInput[1499] , \matrixInput[1480] , \matrixInput[1004] , 
        \matrixInput[130] , \matrixInput[129] , \matrixInput[1783] , 
        \matrixInput[1334] , \matrixInput[1307] , \matrixInput[233] , 
        \matrixInput[1037] , \matrixInput[587] , \matrixInput[103] , 
        \matrixInput[684] , \matrixInput[219] , \matrixInput[200] , 
        \vectorInput[1] , \matrixInput[1964] , \matrixInput[1957] , 
        \matrixInput[863] , \cOutput[127] , \matrixInput[1826] , 
        \matrixInput[1762] , \matrixInput[1276] , \matrixInput[1175] , 
        \matrixInput[850] , \matrixInput[849] , \cOutput[114] , 
        \matrixInput[1245] , \matrixInput[1146] , \matrixInput[342] , 
        \matrixInput[371] , \matrixInput[368] , \matrixInput[1751] , 
        \matrixInput[1478] , \matrixInput[656] , \matrixInput[1461] , 
        \matrixInput[665] , \matrixInput[555] , \matrixInput[1748] , 
        \matrixInput[1452] , \matrixInput[566] , \matrixInput[912] , 
        \matrixInput[15] , \matrixInput[1815] , \matrixInput[938] , 
        \matrixInput[921] , \matrixInput[882] , \matrixInput[26] , 
        \cOutput[38] , \cOutput[21] , \cOutput[12] , \matrixInput[1985] , 
        \matrixInput[1772] , \matrixInput[1758] , \matrixInput[1741] , 
        \matrixInput[1442] , \matrixInput[675] , \matrixInput[646] , 
        \matrixInput[576] , \matrixInput[1471] , \matrixInput[545] , 
        \matrixInput[1468] , \matrixInput[1266] , \matrixInput[1255] , 
        \matrixInput[1156] , \matrixInput[1165] , \matrixInput[378] , 
        \matrixInput[361] , \matrixInput[352] , \matrixInput[1995] , 
        \matrixInput[892] , \cOutput[31] , \cOutput[28] , \vectorInput[119] , 
        \vectorInput[100] , \vectorInput[34] , \vectorInput[8] , 
        \matrixInput[1836] , \matrixInput[1805] , \matrixInput[931] , 
        \matrixInput[928] , \matrixInput[902] , \matrixInput[36] , 
        \matrixInput[5] , \matrixInput[1324] , \matrixInput[1027] , 
        \matrixInput[597] , \matrixInput[113] , \matrixInput[210] , 
        \matrixInput[209] , \matrixInput[1974] , \matrixInput[1793] , 
        \matrixInput[1490] , \matrixInput[1489] , \matrixInput[1014] , 
        \matrixInput[694] , \matrixInput[139] , \matrixInput[120] , 
        \matrixInput[1630] , \matrixInput[1317] , \matrixInput[704] , 
        \matrixInput[399] , \matrixInput[380] , \matrixInput[223] , 
        \matrixInput[1629] , \matrixInput[1603] , \matrixInput[1533] , 
        \matrixInput[407] , \matrixInput[1519] , \matrixInput[1287] , 
        \matrixInput[737] , \matrixInput[1184] , \matrixInput[1500] , 
        \matrixInput[859] , \matrixInput[840] , \matrixInput[434] , 
        \matrixInput[1947] , \cOutput[104] , \matrixInput[873] , 
        \vectorInput[122] , \vectorInput[111] , \vectorInput[25] , 
        \vectorInput[16] , \matrixInput[1782] , \matrixInput[1498] , 
        \matrixInput[1306] , \matrixInput[1005] , \matrixInput[232] , 
        \matrixInput[131] , \matrixInput[128] , \matrixInput[1481] , 
        \matrixInput[1335] , \matrixInput[218] , \matrixInput[201] , 
        \matrixInput[2046] , \matrixInput[1612] , \matrixInput[1511] , 
        \matrixInput[1508] , \matrixInput[1195] , \matrixInput[1036] , 
        \matrixInput[685] , \matrixInput[586] , \matrixInput[102] , 
        \matrixInput[425] , \matrixInput[1522] , \matrixInput[1296] , 
        \matrixInput[726] , \matrixInput[416] , \matrixInput[1965] , 
        \matrixInput[1956] , \matrixInput[1638] , \matrixInput[1621] , 
        \matrixInput[715] , \matrixInput[391] , \matrixInput[388] , 
        \cOutput[126] , \matrixInput[862] , \matrixInput[851] , \cOutput[115] , 
        \matrixInput[848] , \vectorInput[108] , \matrixInput[1763] , 
        \matrixInput[1479] , \matrixInput[1460] , \matrixInput[554] , 
        \matrixInput[657] , \matrixInput[1750] , \matrixInput[1749] , 
        \matrixInput[1453] , \matrixInput[567] , \matrixInput[1277] , 
        \matrixInput[664] , \matrixInput[343] , \matrixInput[1244] , 
        \matrixInput[1174] , \matrixInput[1147] , \matrixInput[370] , 
        \matrixInput[369] , \matrixInput[883] , \cOutput[39] , \cOutput[20] , 
        \matrixInput[1984] , \vectorInput[9] , \vectorInput[0] , 
        \matrixInput[1827] , \matrixInput[913] , \matrixInput[14] , 
        \cOutput[13] , \matrixInput[27] , \matrixInput[1814] , 
        \matrixInput[1773] , \matrixInput[1759] , \matrixInput[1740] , 
        \matrixInput[1443] , \matrixInput[1267] , \matrixInput[1254] , 
        \matrixInput[939] , \matrixInput[920] , \matrixInput[379] , 
        \matrixInput[360] , \matrixInput[1157] , \matrixInput[1164] , 
        \matrixInput[353] , \matrixInput[577] , \matrixInput[674] , 
        \matrixInput[1470] , \matrixInput[1469] , \matrixInput[544] , 
        \matrixInput[647] , \matrixInput[37] , \matrixInput[4] , 
        \matrixInput[1994] , \matrixInput[1837] , \matrixInput[1804] , 
        \matrixInput[930] , \matrixInput[929] , \matrixInput[903] , 
        \matrixInput[893] , \vectorInput[35] , \matrixInput[1631] , 
        \matrixInput[1628] , \matrixInput[1532] , \cOutput[30] , \cOutput[29] , 
        \matrixInput[406] , \matrixInput[398] , \matrixInput[381] , 
        \matrixInput[1602] , \matrixInput[1518] , \matrixInput[1501] , 
        \matrixInput[1185] , \matrixInput[705] , \matrixInput[435] , 
        \matrixInput[736] , \matrixInput[1325] , \matrixInput[1286] , 
        \matrixInput[695] , \matrixInput[211] , \matrixInput[208] , 
        \matrixInput[1792] , \matrixInput[1026] , \matrixInput[596] , 
        \matrixInput[112] , \matrixInput[1491] , \matrixInput[1316] , 
        \matrixInput[222] , \matrixInput[1015] , \matrixInput[138] , 
        \matrixInput[121] , \matrixInput[1488] , \vectorInput[118] , 
        \vectorInput[101] , \vectorInput[4] , \matrixInput[1975] , 
        \cOutput[105] , \matrixInput[1946] , \matrixInput[872] , 
        \matrixInput[858] , \matrixInput[841] , \matrixInput[1823] , 
        \matrixInput[1810] , \matrixInput[1809] , \matrixInput[924] , 
        \matrixInput[917] , \matrixInput[10] , \matrixInput[887] , 
        \matrixInput[23] , \matrixInput[9] , \cOutput[24] , \cOutput[17] , 
        \vectorInput[115] , \matrixInput[1999] , \matrixInput[1980] , 
        \matrixInput[1767] , \matrixInput[1273] , \matrixInput[1170] , 
        \matrixInput[1169] , \matrixInput[1259] , \matrixInput[1143] , 
        \matrixInput[347] , \matrixInput[374] , \matrixInput[1240] , 
        \matrixInput[1754] , \matrixInput[1464] , \matrixInput[653] , 
        \matrixInput[679] , \matrixInput[550] , \matrixInput[549] , 
        \matrixInput[660] , \matrixInput[1457] , \matrixInput[563] , 
        \vectorInput[126] , \vectorInput[105] , \vectorInput[38] , 
        \vectorInput[21] , \vectorInput[12] , \matrixInput[2042] , 
        \matrixInput[1978] , \matrixInput[1961] , \matrixInput[1952] , 
        \matrixInput[866] , \cOutput[122] , \matrixInput[1625] , 
        \matrixInput[1616] , \matrixInput[1292] , \matrixInput[855] , 
        \cOutput[111] , \cOutput[108] , \matrixInput[722] , 
        \matrixInput[1515] , \matrixInput[438] , \matrixInput[421] , 
        \matrixInput[1191] , \matrixInput[1188] , \matrixInput[711] , 
        \matrixInput[708] , \matrixInput[395] , \matrixInput[1526] , 
        \matrixInput[1485] , \matrixInput[412] , \matrixInput[1302] , 
        \matrixInput[1018] , \matrixInput[135] , \matrixInput[1001] , 
        \matrixInput[236] , \matrixInput[1786] , \matrixInput[1032] , 
        \matrixInput[698] , \matrixInput[681] , \matrixInput[582] , 
        \matrixInput[106] , \matrixInput[1971] , \matrixInput[1968] , 
        \matrixInput[1331] , \matrixInput[1328] , \matrixInput[845] , 
        \matrixInput[205] , \matrixInput[1942] , \cOutput[118] , 
        \cOutput[101] , \matrixInput[876] , \vectorInput[31] , 
        \vectorInput[28] , \matrixInput[1022] , \matrixInput[116] , 
        \matrixInput[592] , \matrixInput[1796] , \matrixInput[1495] , 
        \matrixInput[1338] , \matrixInput[691] , \matrixInput[688] , 
        \matrixInput[215] , \matrixInput[1321] , \matrixInput[1312] , 
        \matrixInput[1011] , \matrixInput[1008] , \matrixInput[125] , 
        \matrixInput[226] , \matrixInput[1635] , \matrixInput[718] , 
        \matrixInput[701] , \matrixInput[1606] , \matrixInput[1536] , 
        \matrixInput[402] , \matrixInput[385] , \matrixInput[1282] , 
        \matrixInput[1505] , \matrixInput[732] , \matrixInput[1198] , 
        \matrixInput[1181] , \matrixInput[431] , \matrixInput[428] , 
        \matrixInput[1990] , \matrixInput[1989] , \matrixInput[897] , 
        \cOutput[34] , \matrixInput[1992] , \matrixInput[1833] , 
        \matrixInput[1819] , \matrixInput[1800] , \matrixInput[934] , 
        \matrixInput[907] , \matrixInput[33] , \matrixInput[0] , 
        \matrixInput[1777] , \matrixInput[1744] , \matrixInput[19] , 
        \matrixInput[1447] , \matrixInput[670] , \matrixInput[669] , 
        \matrixInput[643] , \matrixInput[573] , \matrixInput[1474] , 
        \matrixInput[559] , \matrixInput[540] , \matrixInput[1263] , 
        \matrixInput[1250] , \matrixInput[1153] , \matrixInput[1249] , 
        \matrixInput[1179] , \matrixInput[364] , \matrixInput[1160] , 
        \matrixInput[357] , \matrixInput[1973] , \matrixInput[1831] , 
        \matrixInput[1802] , \matrixInput[936] , \matrixInput[895] , 
        \matrixInput[31] , \matrixInput[28] , \cOutput[36] , \matrixInput[2] , 
        \matrixInput[1828] , \matrixInput[1775] , \matrixInput[1746] , 
        \matrixInput[1445] , \matrixInput[905] , \matrixInput[571] , 
        \matrixInput[568] , \matrixInput[672] , \matrixInput[1476] , 
        \matrixInput[542] , \matrixInput[1278] , \matrixInput[1261] , 
        \matrixInput[1252] , \matrixInput[658] , \matrixInput[641] , 
        \matrixInput[366] , \matrixInput[1151] , \matrixInput[1148] , 
        \matrixInput[1162] , \matrixInput[355] , \cOutput[103] , 
        \matrixInput[1959] , \matrixInput[874] , \matrixInput[847] , 
        \matrixInput[1940] , \vectorInput[124] , \vectorInput[117] , 
        \vectorInput[107] , \vectorInput[33] , \matrixInput[1323] , 
        \matrixInput[693] , \matrixInput[217] , \vectorInput[19] , 
        \matrixInput[1794] , \matrixInput[1039] , \matrixInput[1020] , 
        \matrixInput[590] , \matrixInput[589] , \matrixInput[114] , 
        \matrixInput[1637] , \matrixInput[1534] , \matrixInput[1497] , 
        \matrixInput[1310] , \matrixInput[1309] , \matrixInput[224] , 
        \matrixInput[1013] , \matrixInput[127] , \matrixInput[419] , 
        \matrixInput[400] , \matrixInput[387] , \matrixInput[1604] , 
        \matrixInput[1507] , \matrixInput[1183] , \matrixInput[703] , 
        \matrixInput[433] , \matrixInput[730] , \matrixInput[729] , 
        \matrixInput[1299] , \matrixInput[1280] , \vectorInput[23] , 
        \vectorInput[10] , \matrixInput[2040] , \matrixInput[1963] , 
        \matrixInput[1950] , \cOutput[120] , \matrixInput[1949] , 
        \matrixInput[864] , \matrixInput[857] , \cOutput[113] , 
        \matrixInput[1614] , \matrixInput[1517] , \matrixInput[1193] , 
        \matrixInput[423] , \matrixInput[1524] , \matrixInput[1290] , 
        \matrixInput[739] , \matrixInput[720] , \matrixInput[1289] , 
        \matrixInput[410] , \matrixInput[409] , \matrixInput[1627] , 
        \matrixInput[713] , \matrixInput[397] , \matrixInput[1784] , 
        \matrixInput[1487] , \matrixInput[1319] , \matrixInput[1300] , 
        \matrixInput[1003] , \matrixInput[234] , \matrixInput[137] , 
        \matrixInput[1333] , \matrixInput[207] , \matrixInput[1838] , 
        \matrixInput[1030] , \matrixInput[1029] , \matrixInput[683] , 
        \matrixInput[599] , \matrixInput[580] , \matrixInput[104] , 
        \matrixInput[915] , \matrixInput[12] , \matrixInput[1821] , 
        \vectorInput[6] , \matrixInput[38] , \matrixInput[21] , 
        \matrixInput[1982] , \matrixInput[1812] , \matrixInput[926] , 
        \matrixInput[885] , \cOutput[26] , \cOutput[15] , \vectorInput[103] , 
        \vectorInput[37] , \matrixInput[1765] , \matrixInput[1466] , 
        \matrixInput[1271] , \matrixInput[1268] , \matrixInput[345] , 
        \matrixInput[1242] , \matrixInput[1172] , \matrixInput[1158] , 
        \matrixInput[1141] , \matrixInput[376] , \matrixInput[552] , 
        \matrixInput[651] , \matrixInput[648] , \matrixInput[1756] , 
        \matrixInput[1455] , \matrixInput[578] , \matrixInput[561] , 
        \matrixInput[1633] , \matrixInput[707] , \matrixInput[662] , 
        \matrixInput[1619] , \matrixInput[1530] , \matrixInput[404] , 
        \matrixInput[383] , \matrixInput[1529] , \matrixInput[1284] , 
        \matrixInput[1600] , \matrixInput[1503] , \matrixInput[734] , 
        \matrixInput[1187] , \matrixInput[437] , \matrixInput[1024] , 
        \matrixInput[110] , \matrixInput[109] , \matrixInput[594] , 
        \matrixInput[1790] , \matrixInput[1789] , \matrixInput[1493] , 
        \matrixInput[1327] , \matrixInput[697] , \matrixInput[213] , 
        \matrixInput[1314] , \matrixInput[1017] , \matrixInput[123] , 
        \matrixInput[239] , \matrixInput[220] , \matrixInput[1977] , 
        \matrixInput[843] , \matrixInput[1944] , \cOutput[107] , 
        \matrixInput[1835] , \matrixInput[1806] , \matrixInput[1771] , 
        \matrixInput[1742] , \matrixInput[1265] , \matrixInput[1256] , 
        \matrixInput[1155] , \matrixInput[870] , \matrixInput[869] , 
        \matrixInput[1166] , \matrixInput[362] , \matrixInput[351] , 
        \matrixInput[348] , \matrixInput[1458] , \matrixInput[676] , 
        \matrixInput[1441] , \matrixInput[645] , \matrixInput[575] , 
        \matrixInput[1768] , \matrixInput[1472] , \matrixInput[546] , 
        \matrixInput[932] , \matrixInput[918] , \matrixInput[901] , 
        \matrixInput[35] , \matrixInput[6] , \cOutput[18] , 
        \matrixInput[1996] , \cOutput[32] , \matrixInput[1778] , 
        \matrixInput[891] , \matrixInput[888] , \matrixInput[1761] , 
        \matrixInput[1752] , \matrixInput[1462] , \matrixInput[655] , 
        \matrixInput[666] , \matrixInput[556] , \matrixInput[1451] , 
        \matrixInput[565] , \matrixInput[1448] , \matrixInput[1275] , 
        \matrixInput[1176] , \matrixInput[1246] , \matrixInput[1145] , 
        \matrixInput[358] , \matrixInput[341] , \matrixInput[372] , 
        \matrixInput[898] , \cOutput[22] , \matrixInput[881] , 
        \vectorInput[120] , \vectorInput[113] , \vectorInput[27] , 
        \vectorInput[14] , \vectorInput[2] , \matrixInput[1986] , 
        \cOutput[11] , \matrixInput[1825] , \matrixInput[1816] , 
        \matrixInput[922] , \matrixInput[911] , \matrixInput[908] , 
        \matrixInput[16] , \matrixInput[1799] , \matrixInput[1780] , 
        \matrixInput[1483] , \matrixInput[25] , \matrixInput[1304] , 
        \matrixInput[1007] , \matrixInput[133] , \matrixInput[230] , 
        \matrixInput[229] , \matrixInput[1034] , \matrixInput[687] , 
        \matrixInput[584] , \matrixInput[119] , \matrixInput[100] , 
        \matrixInput[2044] , \matrixInput[1623] , \matrixInput[1610] , 
        \matrixInput[1337] , \matrixInput[1294] , \matrixInput[203] , 
        \matrixInput[724] , \matrixInput[1609] , \matrixInput[1513] , 
        \matrixInput[427] , \matrixInput[1197] , \matrixInput[717] , 
        \matrixInput[393] , \matrixInput[1967] , \matrixInput[1954] , 
        \matrixInput[1539] , \matrixInput[1520] , \matrixInput[879] , 
        \matrixInput[860] , \matrixInput[414] , \cOutput[124] , 
        \matrixInput[853] , \cOutput[117] , \vectorInput[90] , 
        \vectorInput[89] , \matrixInput[1873] , \matrixInput[1859] , 
        \matrixInput[974] , \matrixInput[1840] , \matrixInput[73] , 
        \matrixInput[1694] , \matrixInput[1597] , \matrixInput[1113] , 
        \matrixInput[947] , \matrixInput[59] , \matrixInput[40] , 
        \cOutput[74] , \cOutput[47] , \matrixInput[1223] , \matrixInput[1210] , 
        \matrixInput[1209] , \matrixInput[324] , \matrixInput[1139] , 
        \matrixInput[1120] , \matrixInput[490] , \matrixInput[489] , 
        \matrixInput[793] , \matrixInput[317] , \matrixInput[630] , 
        \matrixInput[629] , \matrixInput[1704] , \matrixInput[1407] , 
        \matrixInput[1399] , \matrixInput[1380] , \matrixInput[1083] , 
        \matrixInput[533] , \matrixInput[287] , \vectorInput[71] , 
        \matrixInput[2038] , \matrixInput[2021] , \matrixInput[2012] , 
        \matrixInput[1931] , \matrixInput[1892] , \matrixInput[1737] , 
        \matrixInput[1434] , \matrixInput[603] , \cOutput[5] , 
        \matrixInput[995] , \matrixInput[519] , \matrixInput[500] , 
        \matrixInput[184] , \matrixInput[92] , \matrixInput[1928] , 
        \matrixInput[1902] , \matrixInput[836] , \matrixInput[805] , 
        \matrixInput[1675] , \cOutput[95] , \matrixInput[758] , 
        \matrixInput[741] , \matrixInput[1646] , \matrixInput[1576] , 
        \matrixInput[772] , \matrixInput[442] , \matrixInput[1545] , 
        \matrixInput[471] , \matrixInput[468] , \matrixInput[1062] , 
        \matrixInput[156] , \vectorInput[68] , \vectorInput[52] , 
        \vectorInput[42] , \matrixInput[1378] , \matrixInput[1361] , 
        \matrixInput[1352] , \matrixInput[1051] , \matrixInput[1048] , 
        \matrixInput[255] , \matrixInput[165] , \matrixInput[266] , 
        \matrixInput[1938] , \matrixInput[1912] , \matrixInput[826] , 
        \matrixInput[815] , \cOutput[85] , \matrixInput[1921] , 
        \matrixInput[1882] , \matrixInput[1342] , \matrixInput[1058] , 
        \matrixInput[1041] , \matrixInput[985] , \matrixInput[82] , 
        \matrixInput[175] , \matrixInput[276] , \vectorInput[78] , 
        \matrixInput[1072] , \matrixInput[146] , \vectorInput[61] , 
        \matrixInput[2031] , \matrixInput[2028] , \matrixInput[1656] , 
        \matrixInput[1371] , \matrixInput[1368] , \matrixInput[245] , 
        \matrixInput[1555] , \matrixInput[762] , \matrixInput[478] , 
        \matrixInput[461] , \matrixInput[2002] , \matrixInput[1665] , 
        \matrixInput[751] , \matrixInput[748] , \matrixInput[1566] , 
        \matrixInput[452] , \matrixInput[957] , \cOutput[64] , \cOutput[57] , 
        \matrixInput[1863] , \matrixInput[50] , \matrixInput[49] , 
        \vectorInput[99] , \vectorInput[80] , \matrixInput[1850] , 
        \matrixInput[1849] , \matrixInput[1727] , \matrixInput[964] , 
        \matrixInput[613] , \matrixInput[297] , \matrixInput[63] , 
        \matrixInput[1424] , \matrixInput[510] , \matrixInput[509] , 
        \matrixInput[194] , \vectorInput[94] , \vectorInput[75] , 
        \matrixInput[1714] , \matrixInput[1684] , \matrixInput[1587] , 
        \matrixInput[1417] , \matrixInput[1390] , \matrixInput[639] , 
        \matrixInput[620] , \matrixInput[1389] , \matrixInput[1093] , 
        \matrixInput[1233] , \matrixInput[1130] , \matrixInput[1129] , 
        \matrixInput[523] , \matrixInput[499] , \matrixInput[480] , 
        \matrixInput[307] , \matrixInput[1103] , \matrixInput[783] , 
        \matrixInput[1365] , \matrixInput[1219] , \matrixInput[1200] , 
        \matrixInput[334] , \matrixInput[251] , \matrixInput[248] , 
        \vectorInput[46] , \matrixInput[1066] , \matrixInput[152] , 
        \matrixInput[2025] , \matrixInput[2016] , \matrixInput[1572] , 
        \matrixInput[1356] , \matrixInput[1055] , \matrixInput[262] , 
        \matrixInput[446] , \matrixInput[178] , \matrixInput[161] , 
        \matrixInput[1671] , \matrixInput[745] , \matrixInput[1668] , 
        \matrixInput[1935] , \matrixInput[1642] , \matrixInput[1558] , 
        \matrixInput[1541] , \matrixInput[475] , \matrixInput[818] , 
        \matrixInput[801] , \matrixInput[776] , \matrixInput[1906] , 
        \cOutput[91] , \cOutput[88] , \matrixInput[1896] , \matrixInput[991] , 
        \matrixInput[832] , \matrixInput[988] , \matrixInput[96] , 
        \matrixInput[1403] , \matrixInput[1384] , \matrixInput[1087] , 
        \matrixInput[537] , \matrixInput[1733] , \matrixInput[1719] , 
        \matrixInput[1700] , \matrixInput[1430] , \matrixInput[634] , 
        \matrixInput[504] , \matrixInput[199] , \matrixInput[180] , 
        \matrixInput[1429] , \matrixInput[607] , \cOutput[1] , 
        \matrixInput[1844] , \matrixInput[1690] , \matrixInput[1689] , 
        \matrixInput[1214] , \matrixInput[283] , \matrixInput[339] , 
        \matrixInput[320] , \matrixInput[1593] , \matrixInput[1227] , 
        \matrixInput[1117] , \matrixInput[797] , \matrixInput[313] , 
        \matrixInput[1124] , \matrixInput[494] , \matrixInput[77] , 
        \cOutput[70] , \cOutput[69] , \cOutput[43] , \matrixInput[970] , 
        \matrixInput[969] , \matrixInput[943] , \matrixInput[44] , 
        \matrixInput[1877] , \vectorInput[84] , \matrixInput[1723] , 
        \matrixInput[1699] , \matrixInput[1680] , \matrixInput[1237] , 
        \matrixInput[787] , \matrixInput[1204] , \matrixInput[1134] , 
        \matrixInput[303] , \matrixInput[484] , \matrixInput[330] , 
        \matrixInput[329] , \matrixInput[1583] , \matrixInput[1439] , 
        \matrixInput[1107] , \matrixInput[190] , \matrixInput[189] , 
        \matrixInput[1420] , \matrixInput[514] , \matrixInput[1710] , 
        \matrixInput[1413] , \matrixInput[617] , \cOutput[8] , 
        \matrixInput[527] , \matrixInput[293] , \matrixInput[1394] , 
        \matrixInput[1097] , \matrixInput[624] , \matrixInput[1709] , 
        \matrixInput[54] , \matrixInput[1867] , \matrixInput[979] , 
        \matrixInput[960] , \matrixInput[953] , \matrixInput[67] , 
        \vectorInput[65] , \vectorInput[56] , \matrixInput[2035] , 
        \matrixInput[1854] , \cOutput[79] , \cOutput[60] , \cOutput[53] , 
        \matrixInput[2006] , \matrixInput[1652] , \matrixInput[1551] , 
        \matrixInput[465] , \matrixInput[1548] , \matrixInput[766] , 
        \matrixInput[1562] , \matrixInput[456] , \matrixInput[1678] , 
        \matrixInput[1661] , \matrixInput[755] , \matrixInput[1375] , 
        \matrixInput[1346] , \matrixInput[272] , \matrixInput[1045] , 
        \matrixInput[171] , \matrixInput[168] , \matrixInput[258] , 
        \matrixInput[241] , \matrixInput[1076] , \matrixInput[142] , 
        \vectorInput[54] , \matrixInput[2037] , \matrixInput[1925] , 
        \matrixInput[1916] , \matrixInput[1886] , \matrixInput[998] , 
        \matrixInput[981] , \matrixInput[822] , \matrixInput[86] , 
        \cOutput[98] , \cOutput[81] , \matrixInput[1650] , \matrixInput[1649] , 
        \matrixInput[811] , \matrixInput[808] , \matrixInput[1553] , 
        \matrixInput[764] , \matrixInput[467] , \matrixInput[2004] , 
        \matrixInput[1663] , \matrixInput[757] , \matrixInput[1579] , 
        \matrixInput[1560] , \matrixInput[454] , \matrixInput[1344] , 
        \matrixInput[1047] , \matrixInput[173] , \matrixInput[270] , 
        \matrixInput[269] , \matrixInput[140] , \vectorInput[86] , 
        \vectorInput[67] , \matrixInput[1074] , \matrixInput[159] , 
        \matrixInput[1927] , \matrixInput[1914] , \matrixInput[1884] , 
        \matrixInput[1377] , \matrixInput[243] , \matrixInput[983] , 
        \matrixInput[84] , \matrixInput[839] , \matrixInput[820] , 
        \matrixInput[813] , \cOutput[83] , \matrixInput[1738] , 
        \matrixInput[1721] , \matrixInput[1682] , \matrixInput[1598] , 
        \matrixInput[1235] , \matrixInput[1136] , \matrixInput[486] , 
        \matrixInput[318] , \matrixInput[301] , \matrixInput[1105] , 
        \matrixInput[785] , \matrixInput[1581] , \matrixInput[1206] , 
        \matrixInput[615] , \matrixInput[332] , \matrixInput[291] , 
        \matrixInput[288] , \matrixInput[1712] , \matrixInput[1422] , 
        \matrixInput[516] , \matrixInput[192] , \matrixInput[1411] , 
        \matrixInput[1408] , \matrixInput[1396] , \matrixInput[626] , 
        \matrixInput[1095] , \matrixInput[951] , \matrixInput[525] , 
        \matrixInput[948] , \matrixInput[1865] , \matrixInput[56] , 
        \vectorInput[96] , \matrixInput[1856] , \matrixInput[962] , 
        \matrixInput[636] , \matrixInput[65] , \cOutput[62] , \cOutput[51] , 
        \cOutput[48] , \matrixInput[1846] , \matrixInput[1731] , 
        \matrixInput[1728] , \matrixInput[1702] , \matrixInput[1418] , 
        \matrixInput[1401] , \matrixInput[1386] , \matrixInput[1085] , 
        \matrixInput[535] , \matrixInput[298] , \matrixInput[281] , 
        \cOutput[3] , \matrixInput[1692] , \matrixInput[1591] , 
        \matrixInput[1432] , \matrixInput[605] , \matrixInput[1115] , 
        \matrixInput[506] , \matrixInput[182] , \matrixInput[1588] , 
        \matrixInput[1225] , \matrixInput[1216] , \matrixInput[322] , 
        \matrixInput[1126] , \matrixInput[496] , \matrixInput[972] , 
        \matrixInput[795] , \matrixInput[311] , \matrixInput[308] , 
        \cOutput[72] , \cOutput[58] , \cOutput[41] , \matrixInput[1875] , 
        \matrixInput[75] , \matrixInput[1064] , \matrixInput[958] , 
        \matrixInput[941] , \matrixInput[46] , \matrixInput[149] , 
        \vectorInput[77] , \matrixInput[150] , \vectorInput[44] , 
        \matrixInput[1367] , \matrixInput[1354] , \matrixInput[1057] , 
        \matrixInput[253] , \matrixInput[163] , \matrixInput[279] , 
        \matrixInput[260] , \matrixInput[2027] , \matrixInput[2014] , 
        \matrixInput[1673] , \matrixInput[747] , \matrixInput[1659] , 
        \matrixInput[1640] , \matrixInput[1570] , \matrixInput[1569] , 
        \matrixInput[774] , \matrixInput[444] , \matrixInput[1543] , 
        \matrixInput[477] , \matrixInput[1937] , \matrixInput[1904] , 
        \matrixInput[830] , \matrixInput[803] , \matrixInput[829] , 
        \matrixInput[1894] , \matrixInput[993] , \matrixInput[94] , 
        \cOutput[93] , \matrixInput[52] , \cOutput[66] , \cOutput[55] , 
        \matrixInput[1878] , \matrixInput[1861] , \matrixInput[966] , 
        \matrixInput[955] , \matrixInput[78] , \matrixInput[61] , 
        \vectorInput[82] , \matrixInput[1852] , \matrixInput[1725] , 
        \matrixInput[1426] , \matrixInput[196] , \matrixInput[512] , 
        \matrixInput[1415] , \matrixInput[611] , \matrixInput[608] , 
        \matrixInput[538] , \matrixInput[295] , \matrixInput[521] , 
        \matrixInput[1392] , \matrixInput[1091] , \matrixInput[1088] , 
        \matrixInput[622] , \vectorInput[63] , \vectorInput[50] , 
        \vectorInput[49] , \matrixInput[1923] , \matrixInput[1910] , 
        \matrixInput[1909] , \matrixInput[1716] , \matrixInput[1686] , 
        \matrixInput[1231] , \matrixInput[798] , \matrixInput[781] , 
        \matrixInput[1228] , \matrixInput[1202] , \matrixInput[1132] , 
        \matrixInput[305] , \matrixInput[482] , \matrixInput[336] , 
        \matrixInput[1585] , \matrixInput[1118] , \matrixInput[1101] , 
        \matrixInput[824] , \cOutput[87] , \matrixInput[1899] , 
        \matrixInput[817] , \matrixInput[1880] , \matrixInput[987] , 
        \matrixInput[99] , \matrixInput[80] , \matrixInput[1373] , 
        \matrixInput[1359] , \matrixInput[274] , \matrixInput[1340] , 
        \matrixInput[1043] , \matrixInput[177] , \matrixInput[247] , 
        \matrixInput[1070] , \matrixInput[1069] , \vectorInput[92] , 
        \vectorInput[73] , \matrixInput[2033] , \matrixInput[144] , 
        \matrixInput[2023] , \matrixInput[2019] , \matrixInput[1654] , 
        \matrixInput[1557] , \matrixInput[463] , \matrixInput[779] , 
        \matrixInput[760] , \matrixInput[1564] , \matrixInput[450] , 
        \matrixInput[449] , \matrixInput[2010] , \matrixInput[2000] , 
        \matrixInput[1933] , \matrixInput[1890] , \matrixInput[1667] , 
        \matrixInput[997] , \matrixInput[753] , \matrixInput[90] , 
        \matrixInput[89] , \matrixInput[1889] , \matrixInput[807] , 
        \matrixInput[1919] , \matrixInput[1900] , \cOutput[97] , 
        \matrixInput[1574] , \matrixInput[834] , \matrixInput[459] , 
        \matrixInput[440] , \matrixInput[2009] , \matrixInput[1677] , 
        \matrixInput[743] , \matrixInput[1644] , \matrixInput[1547] , 
        \matrixInput[473] , \matrixInput[1363] , \matrixInput[770] , 
        \matrixInput[769] , \matrixInput[257] , \vectorInput[59] , 
        \vectorInput[40] , \matrixInput[1079] , \matrixInput[154] , 
        \matrixInput[1060] , \matrixInput[1871] , \matrixInput[1868] , 
        \matrixInput[1842] , \matrixInput[1350] , \matrixInput[1349] , 
        \matrixInput[1053] , \matrixInput[264] , \matrixInput[167] , 
        \matrixInput[71] , \matrixInput[68] , \matrixInput[976] , 
        \matrixInput[945] , \matrixInput[42] , \matrixInput[1706] , 
        \matrixInput[1696] , \matrixInput[1212] , \cOutput[76] , \cOutput[45] , 
        \matrixInput[326] , \matrixInput[1595] , \matrixInput[1405] , 
        \matrixInput[1238] , \matrixInput[1111] , \matrixInput[1108] , 
        \matrixInput[791] , \matrixInput[788] , \matrixInput[315] , 
        \matrixInput[1221] , \matrixInput[1122] , \matrixInput[492] , 
        \matrixInput[1382] , \matrixInput[1098] , \matrixInput[1081] , 
        \matrixInput[531] , \matrixInput[528] , \matrixInput[1735] , 
        \matrixInput[1436] , \matrixInput[632] , \matrixInput[502] , 
        \matrixInput[186] , \matrixInput[618] , \matrixInput[601] , 
        \matrixInput[285] , \cOutput[7] ;
    IntMatMul_Control_pVectorSize16_pWordSize8_pScan1 U_IntMatMul_Control ( 
        .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(
        DataIn), .DataOut(DataOut), .vectorInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .matrixInput({
        \matrixInput[2047] , \matrixInput[2046] , \matrixInput[2045] , 
        \matrixInput[2044] , \matrixInput[2043] , \matrixInput[2042] , 
        \matrixInput[2041] , \matrixInput[2040] , \matrixInput[2039] , 
        \matrixInput[2038] , \matrixInput[2037] , \matrixInput[2036] , 
        \matrixInput[2035] , \matrixInput[2034] , \matrixInput[2033] , 
        \matrixInput[2032] , \matrixInput[2031] , \matrixInput[2030] , 
        \matrixInput[2029] , \matrixInput[2028] , \matrixInput[2027] , 
        \matrixInput[2026] , \matrixInput[2025] , \matrixInput[2024] , 
        \matrixInput[2023] , \matrixInput[2022] , \matrixInput[2021] , 
        \matrixInput[2020] , \matrixInput[2019] , \matrixInput[2018] , 
        \matrixInput[2017] , \matrixInput[2016] , \matrixInput[2015] , 
        \matrixInput[2014] , \matrixInput[2013] , \matrixInput[2012] , 
        \matrixInput[2011] , \matrixInput[2010] , \matrixInput[2009] , 
        \matrixInput[2008] , \matrixInput[2007] , \matrixInput[2006] , 
        \matrixInput[2005] , \matrixInput[2004] , \matrixInput[2003] , 
        \matrixInput[2002] , \matrixInput[2001] , \matrixInput[2000] , 
        \matrixInput[1999] , \matrixInput[1998] , \matrixInput[1997] , 
        \matrixInput[1996] , \matrixInput[1995] , \matrixInput[1994] , 
        \matrixInput[1993] , \matrixInput[1992] , \matrixInput[1991] , 
        \matrixInput[1990] , \matrixInput[1989] , \matrixInput[1988] , 
        \matrixInput[1987] , \matrixInput[1986] , \matrixInput[1985] , 
        \matrixInput[1984] , \matrixInput[1983] , \matrixInput[1982] , 
        \matrixInput[1981] , \matrixInput[1980] , \matrixInput[1979] , 
        \matrixInput[1978] , \matrixInput[1977] , \matrixInput[1976] , 
        \matrixInput[1975] , \matrixInput[1974] , \matrixInput[1973] , 
        \matrixInput[1972] , \matrixInput[1971] , \matrixInput[1970] , 
        \matrixInput[1969] , \matrixInput[1968] , \matrixInput[1967] , 
        \matrixInput[1966] , \matrixInput[1965] , \matrixInput[1964] , 
        \matrixInput[1963] , \matrixInput[1962] , \matrixInput[1961] , 
        \matrixInput[1960] , \matrixInput[1959] , \matrixInput[1958] , 
        \matrixInput[1957] , \matrixInput[1956] , \matrixInput[1955] , 
        \matrixInput[1954] , \matrixInput[1953] , \matrixInput[1952] , 
        \matrixInput[1951] , \matrixInput[1950] , \matrixInput[1949] , 
        \matrixInput[1948] , \matrixInput[1947] , \matrixInput[1946] , 
        \matrixInput[1945] , \matrixInput[1944] , \matrixInput[1943] , 
        \matrixInput[1942] , \matrixInput[1941] , \matrixInput[1940] , 
        \matrixInput[1939] , \matrixInput[1938] , \matrixInput[1937] , 
        \matrixInput[1936] , \matrixInput[1935] , \matrixInput[1934] , 
        \matrixInput[1933] , \matrixInput[1932] , \matrixInput[1931] , 
        \matrixInput[1930] , \matrixInput[1929] , \matrixInput[1928] , 
        \matrixInput[1927] , \matrixInput[1926] , \matrixInput[1925] , 
        \matrixInput[1924] , \matrixInput[1923] , \matrixInput[1922] , 
        \matrixInput[1921] , \matrixInput[1920] , \matrixInput[1919] , 
        \matrixInput[1918] , \matrixInput[1917] , \matrixInput[1916] , 
        \matrixInput[1915] , \matrixInput[1914] , \matrixInput[1913] , 
        \matrixInput[1912] , \matrixInput[1911] , \matrixInput[1910] , 
        \matrixInput[1909] , \matrixInput[1908] , \matrixInput[1907] , 
        \matrixInput[1906] , \matrixInput[1905] , \matrixInput[1904] , 
        \matrixInput[1903] , \matrixInput[1902] , \matrixInput[1901] , 
        \matrixInput[1900] , \matrixInput[1899] , \matrixInput[1898] , 
        \matrixInput[1897] , \matrixInput[1896] , \matrixInput[1895] , 
        \matrixInput[1894] , \matrixInput[1893] , \matrixInput[1892] , 
        \matrixInput[1891] , \matrixInput[1890] , \matrixInput[1889] , 
        \matrixInput[1888] , \matrixInput[1887] , \matrixInput[1886] , 
        \matrixInput[1885] , \matrixInput[1884] , \matrixInput[1883] , 
        \matrixInput[1882] , \matrixInput[1881] , \matrixInput[1880] , 
        \matrixInput[1879] , \matrixInput[1878] , \matrixInput[1877] , 
        \matrixInput[1876] , \matrixInput[1875] , \matrixInput[1874] , 
        \matrixInput[1873] , \matrixInput[1872] , \matrixInput[1871] , 
        \matrixInput[1870] , \matrixInput[1869] , \matrixInput[1868] , 
        \matrixInput[1867] , \matrixInput[1866] , \matrixInput[1865] , 
        \matrixInput[1864] , \matrixInput[1863] , \matrixInput[1862] , 
        \matrixInput[1861] , \matrixInput[1860] , \matrixInput[1859] , 
        \matrixInput[1858] , \matrixInput[1857] , \matrixInput[1856] , 
        \matrixInput[1855] , \matrixInput[1854] , \matrixInput[1853] , 
        \matrixInput[1852] , \matrixInput[1851] , \matrixInput[1850] , 
        \matrixInput[1849] , \matrixInput[1848] , \matrixInput[1847] , 
        \matrixInput[1846] , \matrixInput[1845] , \matrixInput[1844] , 
        \matrixInput[1843] , \matrixInput[1842] , \matrixInput[1841] , 
        \matrixInput[1840] , \matrixInput[1839] , \matrixInput[1838] , 
        \matrixInput[1837] , \matrixInput[1836] , \matrixInput[1835] , 
        \matrixInput[1834] , \matrixInput[1833] , \matrixInput[1832] , 
        \matrixInput[1831] , \matrixInput[1830] , \matrixInput[1829] , 
        \matrixInput[1828] , \matrixInput[1827] , \matrixInput[1826] , 
        \matrixInput[1825] , \matrixInput[1824] , \matrixInput[1823] , 
        \matrixInput[1822] , \matrixInput[1821] , \matrixInput[1820] , 
        \matrixInput[1819] , \matrixInput[1818] , \matrixInput[1817] , 
        \matrixInput[1816] , \matrixInput[1815] , \matrixInput[1814] , 
        \matrixInput[1813] , \matrixInput[1812] , \matrixInput[1811] , 
        \matrixInput[1810] , \matrixInput[1809] , \matrixInput[1808] , 
        \matrixInput[1807] , \matrixInput[1806] , \matrixInput[1805] , 
        \matrixInput[1804] , \matrixInput[1803] , \matrixInput[1802] , 
        \matrixInput[1801] , \matrixInput[1800] , \matrixInput[1799] , 
        \matrixInput[1798] , \matrixInput[1797] , \matrixInput[1796] , 
        \matrixInput[1795] , \matrixInput[1794] , \matrixInput[1793] , 
        \matrixInput[1792] , \matrixInput[1791] , \matrixInput[1790] , 
        \matrixInput[1789] , \matrixInput[1788] , \matrixInput[1787] , 
        \matrixInput[1786] , \matrixInput[1785] , \matrixInput[1784] , 
        \matrixInput[1783] , \matrixInput[1782] , \matrixInput[1781] , 
        \matrixInput[1780] , \matrixInput[1779] , \matrixInput[1778] , 
        \matrixInput[1777] , \matrixInput[1776] , \matrixInput[1775] , 
        \matrixInput[1774] , \matrixInput[1773] , \matrixInput[1772] , 
        \matrixInput[1771] , \matrixInput[1770] , \matrixInput[1769] , 
        \matrixInput[1768] , \matrixInput[1767] , \matrixInput[1766] , 
        \matrixInput[1765] , \matrixInput[1764] , \matrixInput[1763] , 
        \matrixInput[1762] , \matrixInput[1761] , \matrixInput[1760] , 
        \matrixInput[1759] , \matrixInput[1758] , \matrixInput[1757] , 
        \matrixInput[1756] , \matrixInput[1755] , \matrixInput[1754] , 
        \matrixInput[1753] , \matrixInput[1752] , \matrixInput[1751] , 
        \matrixInput[1750] , \matrixInput[1749] , \matrixInput[1748] , 
        \matrixInput[1747] , \matrixInput[1746] , \matrixInput[1745] , 
        \matrixInput[1744] , \matrixInput[1743] , \matrixInput[1742] , 
        \matrixInput[1741] , \matrixInput[1740] , \matrixInput[1739] , 
        \matrixInput[1738] , \matrixInput[1737] , \matrixInput[1736] , 
        \matrixInput[1735] , \matrixInput[1734] , \matrixInput[1733] , 
        \matrixInput[1732] , \matrixInput[1731] , \matrixInput[1730] , 
        \matrixInput[1729] , \matrixInput[1728] , \matrixInput[1727] , 
        \matrixInput[1726] , \matrixInput[1725] , \matrixInput[1724] , 
        \matrixInput[1723] , \matrixInput[1722] , \matrixInput[1721] , 
        \matrixInput[1720] , \matrixInput[1719] , \matrixInput[1718] , 
        \matrixInput[1717] , \matrixInput[1716] , \matrixInput[1715] , 
        \matrixInput[1714] , \matrixInput[1713] , \matrixInput[1712] , 
        \matrixInput[1711] , \matrixInput[1710] , \matrixInput[1709] , 
        \matrixInput[1708] , \matrixInput[1707] , \matrixInput[1706] , 
        \matrixInput[1705] , \matrixInput[1704] , \matrixInput[1703] , 
        \matrixInput[1702] , \matrixInput[1701] , \matrixInput[1700] , 
        \matrixInput[1699] , \matrixInput[1698] , \matrixInput[1697] , 
        \matrixInput[1696] , \matrixInput[1695] , \matrixInput[1694] , 
        \matrixInput[1693] , \matrixInput[1692] , \matrixInput[1691] , 
        \matrixInput[1690] , \matrixInput[1689] , \matrixInput[1688] , 
        \matrixInput[1687] , \matrixInput[1686] , \matrixInput[1685] , 
        \matrixInput[1684] , \matrixInput[1683] , \matrixInput[1682] , 
        \matrixInput[1681] , \matrixInput[1680] , \matrixInput[1679] , 
        \matrixInput[1678] , \matrixInput[1677] , \matrixInput[1676] , 
        \matrixInput[1675] , \matrixInput[1674] , \matrixInput[1673] , 
        \matrixInput[1672] , \matrixInput[1671] , \matrixInput[1670] , 
        \matrixInput[1669] , \matrixInput[1668] , \matrixInput[1667] , 
        \matrixInput[1666] , \matrixInput[1665] , \matrixInput[1664] , 
        \matrixInput[1663] , \matrixInput[1662] , \matrixInput[1661] , 
        \matrixInput[1660] , \matrixInput[1659] , \matrixInput[1658] , 
        \matrixInput[1657] , \matrixInput[1656] , \matrixInput[1655] , 
        \matrixInput[1654] , \matrixInput[1653] , \matrixInput[1652] , 
        \matrixInput[1651] , \matrixInput[1650] , \matrixInput[1649] , 
        \matrixInput[1648] , \matrixInput[1647] , \matrixInput[1646] , 
        \matrixInput[1645] , \matrixInput[1644] , \matrixInput[1643] , 
        \matrixInput[1642] , \matrixInput[1641] , \matrixInput[1640] , 
        \matrixInput[1639] , \matrixInput[1638] , \matrixInput[1637] , 
        \matrixInput[1636] , \matrixInput[1635] , \matrixInput[1634] , 
        \matrixInput[1633] , \matrixInput[1632] , \matrixInput[1631] , 
        \matrixInput[1630] , \matrixInput[1629] , \matrixInput[1628] , 
        \matrixInput[1627] , \matrixInput[1626] , \matrixInput[1625] , 
        \matrixInput[1624] , \matrixInput[1623] , \matrixInput[1622] , 
        \matrixInput[1621] , \matrixInput[1620] , \matrixInput[1619] , 
        \matrixInput[1618] , \matrixInput[1617] , \matrixInput[1616] , 
        \matrixInput[1615] , \matrixInput[1614] , \matrixInput[1613] , 
        \matrixInput[1612] , \matrixInput[1611] , \matrixInput[1610] , 
        \matrixInput[1609] , \matrixInput[1608] , \matrixInput[1607] , 
        \matrixInput[1606] , \matrixInput[1605] , \matrixInput[1604] , 
        \matrixInput[1603] , \matrixInput[1602] , \matrixInput[1601] , 
        \matrixInput[1600] , \matrixInput[1599] , \matrixInput[1598] , 
        \matrixInput[1597] , \matrixInput[1596] , \matrixInput[1595] , 
        \matrixInput[1594] , \matrixInput[1593] , \matrixInput[1592] , 
        \matrixInput[1591] , \matrixInput[1590] , \matrixInput[1589] , 
        \matrixInput[1588] , \matrixInput[1587] , \matrixInput[1586] , 
        \matrixInput[1585] , \matrixInput[1584] , \matrixInput[1583] , 
        \matrixInput[1582] , \matrixInput[1581] , \matrixInput[1580] , 
        \matrixInput[1579] , \matrixInput[1578] , \matrixInput[1577] , 
        \matrixInput[1576] , \matrixInput[1575] , \matrixInput[1574] , 
        \matrixInput[1573] , \matrixInput[1572] , \matrixInput[1571] , 
        \matrixInput[1570] , \matrixInput[1569] , \matrixInput[1568] , 
        \matrixInput[1567] , \matrixInput[1566] , \matrixInput[1565] , 
        \matrixInput[1564] , \matrixInput[1563] , \matrixInput[1562] , 
        \matrixInput[1561] , \matrixInput[1560] , \matrixInput[1559] , 
        \matrixInput[1558] , \matrixInput[1557] , \matrixInput[1556] , 
        \matrixInput[1555] , \matrixInput[1554] , \matrixInput[1553] , 
        \matrixInput[1552] , \matrixInput[1551] , \matrixInput[1550] , 
        \matrixInput[1549] , \matrixInput[1548] , \matrixInput[1547] , 
        \matrixInput[1546] , \matrixInput[1545] , \matrixInput[1544] , 
        \matrixInput[1543] , \matrixInput[1542] , \matrixInput[1541] , 
        \matrixInput[1540] , \matrixInput[1539] , \matrixInput[1538] , 
        \matrixInput[1537] , \matrixInput[1536] , \matrixInput[1535] , 
        \matrixInput[1534] , \matrixInput[1533] , \matrixInput[1532] , 
        \matrixInput[1531] , \matrixInput[1530] , \matrixInput[1529] , 
        \matrixInput[1528] , \matrixInput[1527] , \matrixInput[1526] , 
        \matrixInput[1525] , \matrixInput[1524] , \matrixInput[1523] , 
        \matrixInput[1522] , \matrixInput[1521] , \matrixInput[1520] , 
        \matrixInput[1519] , \matrixInput[1518] , \matrixInput[1517] , 
        \matrixInput[1516] , \matrixInput[1515] , \matrixInput[1514] , 
        \matrixInput[1513] , \matrixInput[1512] , \matrixInput[1511] , 
        \matrixInput[1510] , \matrixInput[1509] , \matrixInput[1508] , 
        \matrixInput[1507] , \matrixInput[1506] , \matrixInput[1505] , 
        \matrixInput[1504] , \matrixInput[1503] , \matrixInput[1502] , 
        \matrixInput[1501] , \matrixInput[1500] , \matrixInput[1499] , 
        \matrixInput[1498] , \matrixInput[1497] , \matrixInput[1496] , 
        \matrixInput[1495] , \matrixInput[1494] , \matrixInput[1493] , 
        \matrixInput[1492] , \matrixInput[1491] , \matrixInput[1490] , 
        \matrixInput[1489] , \matrixInput[1488] , \matrixInput[1487] , 
        \matrixInput[1486] , \matrixInput[1485] , \matrixInput[1484] , 
        \matrixInput[1483] , \matrixInput[1482] , \matrixInput[1481] , 
        \matrixInput[1480] , \matrixInput[1479] , \matrixInput[1478] , 
        \matrixInput[1477] , \matrixInput[1476] , \matrixInput[1475] , 
        \matrixInput[1474] , \matrixInput[1473] , \matrixInput[1472] , 
        \matrixInput[1471] , \matrixInput[1470] , \matrixInput[1469] , 
        \matrixInput[1468] , \matrixInput[1467] , \matrixInput[1466] , 
        \matrixInput[1465] , \matrixInput[1464] , \matrixInput[1463] , 
        \matrixInput[1462] , \matrixInput[1461] , \matrixInput[1460] , 
        \matrixInput[1459] , \matrixInput[1458] , \matrixInput[1457] , 
        \matrixInput[1456] , \matrixInput[1455] , \matrixInput[1454] , 
        \matrixInput[1453] , \matrixInput[1452] , \matrixInput[1451] , 
        \matrixInput[1450] , \matrixInput[1449] , \matrixInput[1448] , 
        \matrixInput[1447] , \matrixInput[1446] , \matrixInput[1445] , 
        \matrixInput[1444] , \matrixInput[1443] , \matrixInput[1442] , 
        \matrixInput[1441] , \matrixInput[1440] , \matrixInput[1439] , 
        \matrixInput[1438] , \matrixInput[1437] , \matrixInput[1436] , 
        \matrixInput[1435] , \matrixInput[1434] , \matrixInput[1433] , 
        \matrixInput[1432] , \matrixInput[1431] , \matrixInput[1430] , 
        \matrixInput[1429] , \matrixInput[1428] , \matrixInput[1427] , 
        \matrixInput[1426] , \matrixInput[1425] , \matrixInput[1424] , 
        \matrixInput[1423] , \matrixInput[1422] , \matrixInput[1421] , 
        \matrixInput[1420] , \matrixInput[1419] , \matrixInput[1418] , 
        \matrixInput[1417] , \matrixInput[1416] , \matrixInput[1415] , 
        \matrixInput[1414] , \matrixInput[1413] , \matrixInput[1412] , 
        \matrixInput[1411] , \matrixInput[1410] , \matrixInput[1409] , 
        \matrixInput[1408] , \matrixInput[1407] , \matrixInput[1406] , 
        \matrixInput[1405] , \matrixInput[1404] , \matrixInput[1403] , 
        \matrixInput[1402] , \matrixInput[1401] , \matrixInput[1400] , 
        \matrixInput[1399] , \matrixInput[1398] , \matrixInput[1397] , 
        \matrixInput[1396] , \matrixInput[1395] , \matrixInput[1394] , 
        \matrixInput[1393] , \matrixInput[1392] , \matrixInput[1391] , 
        \matrixInput[1390] , \matrixInput[1389] , \matrixInput[1388] , 
        \matrixInput[1387] , \matrixInput[1386] , \matrixInput[1385] , 
        \matrixInput[1384] , \matrixInput[1383] , \matrixInput[1382] , 
        \matrixInput[1381] , \matrixInput[1380] , \matrixInput[1379] , 
        \matrixInput[1378] , \matrixInput[1377] , \matrixInput[1376] , 
        \matrixInput[1375] , \matrixInput[1374] , \matrixInput[1373] , 
        \matrixInput[1372] , \matrixInput[1371] , \matrixInput[1370] , 
        \matrixInput[1369] , \matrixInput[1368] , \matrixInput[1367] , 
        \matrixInput[1366] , \matrixInput[1365] , \matrixInput[1364] , 
        \matrixInput[1363] , \matrixInput[1362] , \matrixInput[1361] , 
        \matrixInput[1360] , \matrixInput[1359] , \matrixInput[1358] , 
        \matrixInput[1357] , \matrixInput[1356] , \matrixInput[1355] , 
        \matrixInput[1354] , \matrixInput[1353] , \matrixInput[1352] , 
        \matrixInput[1351] , \matrixInput[1350] , \matrixInput[1349] , 
        \matrixInput[1348] , \matrixInput[1347] , \matrixInput[1346] , 
        \matrixInput[1345] , \matrixInput[1344] , \matrixInput[1343] , 
        \matrixInput[1342] , \matrixInput[1341] , \matrixInput[1340] , 
        \matrixInput[1339] , \matrixInput[1338] , \matrixInput[1337] , 
        \matrixInput[1336] , \matrixInput[1335] , \matrixInput[1334] , 
        \matrixInput[1333] , \matrixInput[1332] , \matrixInput[1331] , 
        \matrixInput[1330] , \matrixInput[1329] , \matrixInput[1328] , 
        \matrixInput[1327] , \matrixInput[1326] , \matrixInput[1325] , 
        \matrixInput[1324] , \matrixInput[1323] , \matrixInput[1322] , 
        \matrixInput[1321] , \matrixInput[1320] , \matrixInput[1319] , 
        \matrixInput[1318] , \matrixInput[1317] , \matrixInput[1316] , 
        \matrixInput[1315] , \matrixInput[1314] , \matrixInput[1313] , 
        \matrixInput[1312] , \matrixInput[1311] , \matrixInput[1310] , 
        \matrixInput[1309] , \matrixInput[1308] , \matrixInput[1307] , 
        \matrixInput[1306] , \matrixInput[1305] , \matrixInput[1304] , 
        \matrixInput[1303] , \matrixInput[1302] , \matrixInput[1301] , 
        \matrixInput[1300] , \matrixInput[1299] , \matrixInput[1298] , 
        \matrixInput[1297] , \matrixInput[1296] , \matrixInput[1295] , 
        \matrixInput[1294] , \matrixInput[1293] , \matrixInput[1292] , 
        \matrixInput[1291] , \matrixInput[1290] , \matrixInput[1289] , 
        \matrixInput[1288] , \matrixInput[1287] , \matrixInput[1286] , 
        \matrixInput[1285] , \matrixInput[1284] , \matrixInput[1283] , 
        \matrixInput[1282] , \matrixInput[1281] , \matrixInput[1280] , 
        \matrixInput[1279] , \matrixInput[1278] , \matrixInput[1277] , 
        \matrixInput[1276] , \matrixInput[1275] , \matrixInput[1274] , 
        \matrixInput[1273] , \matrixInput[1272] , \matrixInput[1271] , 
        \matrixInput[1270] , \matrixInput[1269] , \matrixInput[1268] , 
        \matrixInput[1267] , \matrixInput[1266] , \matrixInput[1265] , 
        \matrixInput[1264] , \matrixInput[1263] , \matrixInput[1262] , 
        \matrixInput[1261] , \matrixInput[1260] , \matrixInput[1259] , 
        \matrixInput[1258] , \matrixInput[1257] , \matrixInput[1256] , 
        \matrixInput[1255] , \matrixInput[1254] , \matrixInput[1253] , 
        \matrixInput[1252] , \matrixInput[1251] , \matrixInput[1250] , 
        \matrixInput[1249] , \matrixInput[1248] , \matrixInput[1247] , 
        \matrixInput[1246] , \matrixInput[1245] , \matrixInput[1244] , 
        \matrixInput[1243] , \matrixInput[1242] , \matrixInput[1241] , 
        \matrixInput[1240] , \matrixInput[1239] , \matrixInput[1238] , 
        \matrixInput[1237] , \matrixInput[1236] , \matrixInput[1235] , 
        \matrixInput[1234] , \matrixInput[1233] , \matrixInput[1232] , 
        \matrixInput[1231] , \matrixInput[1230] , \matrixInput[1229] , 
        \matrixInput[1228] , \matrixInput[1227] , \matrixInput[1226] , 
        \matrixInput[1225] , \matrixInput[1224] , \matrixInput[1223] , 
        \matrixInput[1222] , \matrixInput[1221] , \matrixInput[1220] , 
        \matrixInput[1219] , \matrixInput[1218] , \matrixInput[1217] , 
        \matrixInput[1216] , \matrixInput[1215] , \matrixInput[1214] , 
        \matrixInput[1213] , \matrixInput[1212] , \matrixInput[1211] , 
        \matrixInput[1210] , \matrixInput[1209] , \matrixInput[1208] , 
        \matrixInput[1207] , \matrixInput[1206] , \matrixInput[1205] , 
        \matrixInput[1204] , \matrixInput[1203] , \matrixInput[1202] , 
        \matrixInput[1201] , \matrixInput[1200] , \matrixInput[1199] , 
        \matrixInput[1198] , \matrixInput[1197] , \matrixInput[1196] , 
        \matrixInput[1195] , \matrixInput[1194] , \matrixInput[1193] , 
        \matrixInput[1192] , \matrixInput[1191] , \matrixInput[1190] , 
        \matrixInput[1189] , \matrixInput[1188] , \matrixInput[1187] , 
        \matrixInput[1186] , \matrixInput[1185] , \matrixInput[1184] , 
        \matrixInput[1183] , \matrixInput[1182] , \matrixInput[1181] , 
        \matrixInput[1180] , \matrixInput[1179] , \matrixInput[1178] , 
        \matrixInput[1177] , \matrixInput[1176] , \matrixInput[1175] , 
        \matrixInput[1174] , \matrixInput[1173] , \matrixInput[1172] , 
        \matrixInput[1171] , \matrixInput[1170] , \matrixInput[1169] , 
        \matrixInput[1168] , \matrixInput[1167] , \matrixInput[1166] , 
        \matrixInput[1165] , \matrixInput[1164] , \matrixInput[1163] , 
        \matrixInput[1162] , \matrixInput[1161] , \matrixInput[1160] , 
        \matrixInput[1159] , \matrixInput[1158] , \matrixInput[1157] , 
        \matrixInput[1156] , \matrixInput[1155] , \matrixInput[1154] , 
        \matrixInput[1153] , \matrixInput[1152] , \matrixInput[1151] , 
        \matrixInput[1150] , \matrixInput[1149] , \matrixInput[1148] , 
        \matrixInput[1147] , \matrixInput[1146] , \matrixInput[1145] , 
        \matrixInput[1144] , \matrixInput[1143] , \matrixInput[1142] , 
        \matrixInput[1141] , \matrixInput[1140] , \matrixInput[1139] , 
        \matrixInput[1138] , \matrixInput[1137] , \matrixInput[1136] , 
        \matrixInput[1135] , \matrixInput[1134] , \matrixInput[1133] , 
        \matrixInput[1132] , \matrixInput[1131] , \matrixInput[1130] , 
        \matrixInput[1129] , \matrixInput[1128] , \matrixInput[1127] , 
        \matrixInput[1126] , \matrixInput[1125] , \matrixInput[1124] , 
        \matrixInput[1123] , \matrixInput[1122] , \matrixInput[1121] , 
        \matrixInput[1120] , \matrixInput[1119] , \matrixInput[1118] , 
        \matrixInput[1117] , \matrixInput[1116] , \matrixInput[1115] , 
        \matrixInput[1114] , \matrixInput[1113] , \matrixInput[1112] , 
        \matrixInput[1111] , \matrixInput[1110] , \matrixInput[1109] , 
        \matrixInput[1108] , \matrixInput[1107] , \matrixInput[1106] , 
        \matrixInput[1105] , \matrixInput[1104] , \matrixInput[1103] , 
        \matrixInput[1102] , \matrixInput[1101] , \matrixInput[1100] , 
        \matrixInput[1099] , \matrixInput[1098] , \matrixInput[1097] , 
        \matrixInput[1096] , \matrixInput[1095] , \matrixInput[1094] , 
        \matrixInput[1093] , \matrixInput[1092] , \matrixInput[1091] , 
        \matrixInput[1090] , \matrixInput[1089] , \matrixInput[1088] , 
        \matrixInput[1087] , \matrixInput[1086] , \matrixInput[1085] , 
        \matrixInput[1084] , \matrixInput[1083] , \matrixInput[1082] , 
        \matrixInput[1081] , \matrixInput[1080] , \matrixInput[1079] , 
        \matrixInput[1078] , \matrixInput[1077] , \matrixInput[1076] , 
        \matrixInput[1075] , \matrixInput[1074] , \matrixInput[1073] , 
        \matrixInput[1072] , \matrixInput[1071] , \matrixInput[1070] , 
        \matrixInput[1069] , \matrixInput[1068] , \matrixInput[1067] , 
        \matrixInput[1066] , \matrixInput[1065] , \matrixInput[1064] , 
        \matrixInput[1063] , \matrixInput[1062] , \matrixInput[1061] , 
        \matrixInput[1060] , \matrixInput[1059] , \matrixInput[1058] , 
        \matrixInput[1057] , \matrixInput[1056] , \matrixInput[1055] , 
        \matrixInput[1054] , \matrixInput[1053] , \matrixInput[1052] , 
        \matrixInput[1051] , \matrixInput[1050] , \matrixInput[1049] , 
        \matrixInput[1048] , \matrixInput[1047] , \matrixInput[1046] , 
        \matrixInput[1045] , \matrixInput[1044] , \matrixInput[1043] , 
        \matrixInput[1042] , \matrixInput[1041] , \matrixInput[1040] , 
        \matrixInput[1039] , \matrixInput[1038] , \matrixInput[1037] , 
        \matrixInput[1036] , \matrixInput[1035] , \matrixInput[1034] , 
        \matrixInput[1033] , \matrixInput[1032] , \matrixInput[1031] , 
        \matrixInput[1030] , \matrixInput[1029] , \matrixInput[1028] , 
        \matrixInput[1027] , \matrixInput[1026] , \matrixInput[1025] , 
        \matrixInput[1024] , \matrixInput[1023] , \matrixInput[1022] , 
        \matrixInput[1021] , \matrixInput[1020] , \matrixInput[1019] , 
        \matrixInput[1018] , \matrixInput[1017] , \matrixInput[1016] , 
        \matrixInput[1015] , \matrixInput[1014] , \matrixInput[1013] , 
        \matrixInput[1012] , \matrixInput[1011] , \matrixInput[1010] , 
        \matrixInput[1009] , \matrixInput[1008] , \matrixInput[1007] , 
        \matrixInput[1006] , \matrixInput[1005] , \matrixInput[1004] , 
        \matrixInput[1003] , \matrixInput[1002] , \matrixInput[1001] , 
        \matrixInput[1000] , \matrixInput[999] , \matrixInput[998] , 
        \matrixInput[997] , \matrixInput[996] , \matrixInput[995] , 
        \matrixInput[994] , \matrixInput[993] , \matrixInput[992] , 
        \matrixInput[991] , \matrixInput[990] , \matrixInput[989] , 
        \matrixInput[988] , \matrixInput[987] , \matrixInput[986] , 
        \matrixInput[985] , \matrixInput[984] , \matrixInput[983] , 
        \matrixInput[982] , \matrixInput[981] , \matrixInput[980] , 
        \matrixInput[979] , \matrixInput[978] , \matrixInput[977] , 
        \matrixInput[976] , \matrixInput[975] , \matrixInput[974] , 
        \matrixInput[973] , \matrixInput[972] , \matrixInput[971] , 
        \matrixInput[970] , \matrixInput[969] , \matrixInput[968] , 
        \matrixInput[967] , \matrixInput[966] , \matrixInput[965] , 
        \matrixInput[964] , \matrixInput[963] , \matrixInput[962] , 
        \matrixInput[961] , \matrixInput[960] , \matrixInput[959] , 
        \matrixInput[958] , \matrixInput[957] , \matrixInput[956] , 
        \matrixInput[955] , \matrixInput[954] , \matrixInput[953] , 
        \matrixInput[952] , \matrixInput[951] , \matrixInput[950] , 
        \matrixInput[949] , \matrixInput[948] , \matrixInput[947] , 
        \matrixInput[946] , \matrixInput[945] , \matrixInput[944] , 
        \matrixInput[943] , \matrixInput[942] , \matrixInput[941] , 
        \matrixInput[940] , \matrixInput[939] , \matrixInput[938] , 
        \matrixInput[937] , \matrixInput[936] , \matrixInput[935] , 
        \matrixInput[934] , \matrixInput[933] , \matrixInput[932] , 
        \matrixInput[931] , \matrixInput[930] , \matrixInput[929] , 
        \matrixInput[928] , \matrixInput[927] , \matrixInput[926] , 
        \matrixInput[925] , \matrixInput[924] , \matrixInput[923] , 
        \matrixInput[922] , \matrixInput[921] , \matrixInput[920] , 
        \matrixInput[919] , \matrixInput[918] , \matrixInput[917] , 
        \matrixInput[916] , \matrixInput[915] , \matrixInput[914] , 
        \matrixInput[913] , \matrixInput[912] , \matrixInput[911] , 
        \matrixInput[910] , \matrixInput[909] , \matrixInput[908] , 
        \matrixInput[907] , \matrixInput[906] , \matrixInput[905] , 
        \matrixInput[904] , \matrixInput[903] , \matrixInput[902] , 
        \matrixInput[901] , \matrixInput[900] , \matrixInput[899] , 
        \matrixInput[898] , \matrixInput[897] , \matrixInput[896] , 
        \matrixInput[895] , \matrixInput[894] , \matrixInput[893] , 
        \matrixInput[892] , \matrixInput[891] , \matrixInput[890] , 
        \matrixInput[889] , \matrixInput[888] , \matrixInput[887] , 
        \matrixInput[886] , \matrixInput[885] , \matrixInput[884] , 
        \matrixInput[883] , \matrixInput[882] , \matrixInput[881] , 
        \matrixInput[880] , \matrixInput[879] , \matrixInput[878] , 
        \matrixInput[877] , \matrixInput[876] , \matrixInput[875] , 
        \matrixInput[874] , \matrixInput[873] , \matrixInput[872] , 
        \matrixInput[871] , \matrixInput[870] , \matrixInput[869] , 
        \matrixInput[868] , \matrixInput[867] , \matrixInput[866] , 
        \matrixInput[865] , \matrixInput[864] , \matrixInput[863] , 
        \matrixInput[862] , \matrixInput[861] , \matrixInput[860] , 
        \matrixInput[859] , \matrixInput[858] , \matrixInput[857] , 
        \matrixInput[856] , \matrixInput[855] , \matrixInput[854] , 
        \matrixInput[853] , \matrixInput[852] , \matrixInput[851] , 
        \matrixInput[850] , \matrixInput[849] , \matrixInput[848] , 
        \matrixInput[847] , \matrixInput[846] , \matrixInput[845] , 
        \matrixInput[844] , \matrixInput[843] , \matrixInput[842] , 
        \matrixInput[841] , \matrixInput[840] , \matrixInput[839] , 
        \matrixInput[838] , \matrixInput[837] , \matrixInput[836] , 
        \matrixInput[835] , \matrixInput[834] , \matrixInput[833] , 
        \matrixInput[832] , \matrixInput[831] , \matrixInput[830] , 
        \matrixInput[829] , \matrixInput[828] , \matrixInput[827] , 
        \matrixInput[826] , \matrixInput[825] , \matrixInput[824] , 
        \matrixInput[823] , \matrixInput[822] , \matrixInput[821] , 
        \matrixInput[820] , \matrixInput[819] , \matrixInput[818] , 
        \matrixInput[817] , \matrixInput[816] , \matrixInput[815] , 
        \matrixInput[814] , \matrixInput[813] , \matrixInput[812] , 
        \matrixInput[811] , \matrixInput[810] , \matrixInput[809] , 
        \matrixInput[808] , \matrixInput[807] , \matrixInput[806] , 
        \matrixInput[805] , \matrixInput[804] , \matrixInput[803] , 
        \matrixInput[802] , \matrixInput[801] , \matrixInput[800] , 
        \matrixInput[799] , \matrixInput[798] , \matrixInput[797] , 
        \matrixInput[796] , \matrixInput[795] , \matrixInput[794] , 
        \matrixInput[793] , \matrixInput[792] , \matrixInput[791] , 
        \matrixInput[790] , \matrixInput[789] , \matrixInput[788] , 
        \matrixInput[787] , \matrixInput[786] , \matrixInput[785] , 
        \matrixInput[784] , \matrixInput[783] , \matrixInput[782] , 
        \matrixInput[781] , \matrixInput[780] , \matrixInput[779] , 
        \matrixInput[778] , \matrixInput[777] , \matrixInput[776] , 
        \matrixInput[775] , \matrixInput[774] , \matrixInput[773] , 
        \matrixInput[772] , \matrixInput[771] , \matrixInput[770] , 
        \matrixInput[769] , \matrixInput[768] , \matrixInput[767] , 
        \matrixInput[766] , \matrixInput[765] , \matrixInput[764] , 
        \matrixInput[763] , \matrixInput[762] , \matrixInput[761] , 
        \matrixInput[760] , \matrixInput[759] , \matrixInput[758] , 
        \matrixInput[757] , \matrixInput[756] , \matrixInput[755] , 
        \matrixInput[754] , \matrixInput[753] , \matrixInput[752] , 
        \matrixInput[751] , \matrixInput[750] , \matrixInput[749] , 
        \matrixInput[748] , \matrixInput[747] , \matrixInput[746] , 
        \matrixInput[745] , \matrixInput[744] , \matrixInput[743] , 
        \matrixInput[742] , \matrixInput[741] , \matrixInput[740] , 
        \matrixInput[739] , \matrixInput[738] , \matrixInput[737] , 
        \matrixInput[736] , \matrixInput[735] , \matrixInput[734] , 
        \matrixInput[733] , \matrixInput[732] , \matrixInput[731] , 
        \matrixInput[730] , \matrixInput[729] , \matrixInput[728] , 
        \matrixInput[727] , \matrixInput[726] , \matrixInput[725] , 
        \matrixInput[724] , \matrixInput[723] , \matrixInput[722] , 
        \matrixInput[721] , \matrixInput[720] , \matrixInput[719] , 
        \matrixInput[718] , \matrixInput[717] , \matrixInput[716] , 
        \matrixInput[715] , \matrixInput[714] , \matrixInput[713] , 
        \matrixInput[712] , \matrixInput[711] , \matrixInput[710] , 
        \matrixInput[709] , \matrixInput[708] , \matrixInput[707] , 
        \matrixInput[706] , \matrixInput[705] , \matrixInput[704] , 
        \matrixInput[703] , \matrixInput[702] , \matrixInput[701] , 
        \matrixInput[700] , \matrixInput[699] , \matrixInput[698] , 
        \matrixInput[697] , \matrixInput[696] , \matrixInput[695] , 
        \matrixInput[694] , \matrixInput[693] , \matrixInput[692] , 
        \matrixInput[691] , \matrixInput[690] , \matrixInput[689] , 
        \matrixInput[688] , \matrixInput[687] , \matrixInput[686] , 
        \matrixInput[685] , \matrixInput[684] , \matrixInput[683] , 
        \matrixInput[682] , \matrixInput[681] , \matrixInput[680] , 
        \matrixInput[679] , \matrixInput[678] , \matrixInput[677] , 
        \matrixInput[676] , \matrixInput[675] , \matrixInput[674] , 
        \matrixInput[673] , \matrixInput[672] , \matrixInput[671] , 
        \matrixInput[670] , \matrixInput[669] , \matrixInput[668] , 
        \matrixInput[667] , \matrixInput[666] , \matrixInput[665] , 
        \matrixInput[664] , \matrixInput[663] , \matrixInput[662] , 
        \matrixInput[661] , \matrixInput[660] , \matrixInput[659] , 
        \matrixInput[658] , \matrixInput[657] , \matrixInput[656] , 
        \matrixInput[655] , \matrixInput[654] , \matrixInput[653] , 
        \matrixInput[652] , \matrixInput[651] , \matrixInput[650] , 
        \matrixInput[649] , \matrixInput[648] , \matrixInput[647] , 
        \matrixInput[646] , \matrixInput[645] , \matrixInput[644] , 
        \matrixInput[643] , \matrixInput[642] , \matrixInput[641] , 
        \matrixInput[640] , \matrixInput[639] , \matrixInput[638] , 
        \matrixInput[637] , \matrixInput[636] , \matrixInput[635] , 
        \matrixInput[634] , \matrixInput[633] , \matrixInput[632] , 
        \matrixInput[631] , \matrixInput[630] , \matrixInput[629] , 
        \matrixInput[628] , \matrixInput[627] , \matrixInput[626] , 
        \matrixInput[625] , \matrixInput[624] , \matrixInput[623] , 
        \matrixInput[622] , \matrixInput[621] , \matrixInput[620] , 
        \matrixInput[619] , \matrixInput[618] , \matrixInput[617] , 
        \matrixInput[616] , \matrixInput[615] , \matrixInput[614] , 
        \matrixInput[613] , \matrixInput[612] , \matrixInput[611] , 
        \matrixInput[610] , \matrixInput[609] , \matrixInput[608] , 
        \matrixInput[607] , \matrixInput[606] , \matrixInput[605] , 
        \matrixInput[604] , \matrixInput[603] , \matrixInput[602] , 
        \matrixInput[601] , \matrixInput[600] , \matrixInput[599] , 
        \matrixInput[598] , \matrixInput[597] , \matrixInput[596] , 
        \matrixInput[595] , \matrixInput[594] , \matrixInput[593] , 
        \matrixInput[592] , \matrixInput[591] , \matrixInput[590] , 
        \matrixInput[589] , \matrixInput[588] , \matrixInput[587] , 
        \matrixInput[586] , \matrixInput[585] , \matrixInput[584] , 
        \matrixInput[583] , \matrixInput[582] , \matrixInput[581] , 
        \matrixInput[580] , \matrixInput[579] , \matrixInput[578] , 
        \matrixInput[577] , \matrixInput[576] , \matrixInput[575] , 
        \matrixInput[574] , \matrixInput[573] , \matrixInput[572] , 
        \matrixInput[571] , \matrixInput[570] , \matrixInput[569] , 
        \matrixInput[568] , \matrixInput[567] , \matrixInput[566] , 
        \matrixInput[565] , \matrixInput[564] , \matrixInput[563] , 
        \matrixInput[562] , \matrixInput[561] , \matrixInput[560] , 
        \matrixInput[559] , \matrixInput[558] , \matrixInput[557] , 
        \matrixInput[556] , \matrixInput[555] , \matrixInput[554] , 
        \matrixInput[553] , \matrixInput[552] , \matrixInput[551] , 
        \matrixInput[550] , \matrixInput[549] , \matrixInput[548] , 
        \matrixInput[547] , \matrixInput[546] , \matrixInput[545] , 
        \matrixInput[544] , \matrixInput[543] , \matrixInput[542] , 
        \matrixInput[541] , \matrixInput[540] , \matrixInput[539] , 
        \matrixInput[538] , \matrixInput[537] , \matrixInput[536] , 
        \matrixInput[535] , \matrixInput[534] , \matrixInput[533] , 
        \matrixInput[532] , \matrixInput[531] , \matrixInput[530] , 
        \matrixInput[529] , \matrixInput[528] , \matrixInput[527] , 
        \matrixInput[526] , \matrixInput[525] , \matrixInput[524] , 
        \matrixInput[523] , \matrixInput[522] , \matrixInput[521] , 
        \matrixInput[520] , \matrixInput[519] , \matrixInput[518] , 
        \matrixInput[517] , \matrixInput[516] , \matrixInput[515] , 
        \matrixInput[514] , \matrixInput[513] , \matrixInput[512] , 
        \matrixInput[511] , \matrixInput[510] , \matrixInput[509] , 
        \matrixInput[508] , \matrixInput[507] , \matrixInput[506] , 
        \matrixInput[505] , \matrixInput[504] , \matrixInput[503] , 
        \matrixInput[502] , \matrixInput[501] , \matrixInput[500] , 
        \matrixInput[499] , \matrixInput[498] , \matrixInput[497] , 
        \matrixInput[496] , \matrixInput[495] , \matrixInput[494] , 
        \matrixInput[493] , \matrixInput[492] , \matrixInput[491] , 
        \matrixInput[490] , \matrixInput[489] , \matrixInput[488] , 
        \matrixInput[487] , \matrixInput[486] , \matrixInput[485] , 
        \matrixInput[484] , \matrixInput[483] , \matrixInput[482] , 
        \matrixInput[481] , \matrixInput[480] , \matrixInput[479] , 
        \matrixInput[478] , \matrixInput[477] , \matrixInput[476] , 
        \matrixInput[475] , \matrixInput[474] , \matrixInput[473] , 
        \matrixInput[472] , \matrixInput[471] , \matrixInput[470] , 
        \matrixInput[469] , \matrixInput[468] , \matrixInput[467] , 
        \matrixInput[466] , \matrixInput[465] , \matrixInput[464] , 
        \matrixInput[463] , \matrixInput[462] , \matrixInput[461] , 
        \matrixInput[460] , \matrixInput[459] , \matrixInput[458] , 
        \matrixInput[457] , \matrixInput[456] , \matrixInput[455] , 
        \matrixInput[454] , \matrixInput[453] , \matrixInput[452] , 
        \matrixInput[451] , \matrixInput[450] , \matrixInput[449] , 
        \matrixInput[448] , \matrixInput[447] , \matrixInput[446] , 
        \matrixInput[445] , \matrixInput[444] , \matrixInput[443] , 
        \matrixInput[442] , \matrixInput[441] , \matrixInput[440] , 
        \matrixInput[439] , \matrixInput[438] , \matrixInput[437] , 
        \matrixInput[436] , \matrixInput[435] , \matrixInput[434] , 
        \matrixInput[433] , \matrixInput[432] , \matrixInput[431] , 
        \matrixInput[430] , \matrixInput[429] , \matrixInput[428] , 
        \matrixInput[427] , \matrixInput[426] , \matrixInput[425] , 
        \matrixInput[424] , \matrixInput[423] , \matrixInput[422] , 
        \matrixInput[421] , \matrixInput[420] , \matrixInput[419] , 
        \matrixInput[418] , \matrixInput[417] , \matrixInput[416] , 
        \matrixInput[415] , \matrixInput[414] , \matrixInput[413] , 
        \matrixInput[412] , \matrixInput[411] , \matrixInput[410] , 
        \matrixInput[409] , \matrixInput[408] , \matrixInput[407] , 
        \matrixInput[406] , \matrixInput[405] , \matrixInput[404] , 
        \matrixInput[403] , \matrixInput[402] , \matrixInput[401] , 
        \matrixInput[400] , \matrixInput[399] , \matrixInput[398] , 
        \matrixInput[397] , \matrixInput[396] , \matrixInput[395] , 
        \matrixInput[394] , \matrixInput[393] , \matrixInput[392] , 
        \matrixInput[391] , \matrixInput[390] , \matrixInput[389] , 
        \matrixInput[388] , \matrixInput[387] , \matrixInput[386] , 
        \matrixInput[385] , \matrixInput[384] , \matrixInput[383] , 
        \matrixInput[382] , \matrixInput[381] , \matrixInput[380] , 
        \matrixInput[379] , \matrixInput[378] , \matrixInput[377] , 
        \matrixInput[376] , \matrixInput[375] , \matrixInput[374] , 
        \matrixInput[373] , \matrixInput[372] , \matrixInput[371] , 
        \matrixInput[370] , \matrixInput[369] , \matrixInput[368] , 
        \matrixInput[367] , \matrixInput[366] , \matrixInput[365] , 
        \matrixInput[364] , \matrixInput[363] , \matrixInput[362] , 
        \matrixInput[361] , \matrixInput[360] , \matrixInput[359] , 
        \matrixInput[358] , \matrixInput[357] , \matrixInput[356] , 
        \matrixInput[355] , \matrixInput[354] , \matrixInput[353] , 
        \matrixInput[352] , \matrixInput[351] , \matrixInput[350] , 
        \matrixInput[349] , \matrixInput[348] , \matrixInput[347] , 
        \matrixInput[346] , \matrixInput[345] , \matrixInput[344] , 
        \matrixInput[343] , \matrixInput[342] , \matrixInput[341] , 
        \matrixInput[340] , \matrixInput[339] , \matrixInput[338] , 
        \matrixInput[337] , \matrixInput[336] , \matrixInput[335] , 
        \matrixInput[334] , \matrixInput[333] , \matrixInput[332] , 
        \matrixInput[331] , \matrixInput[330] , \matrixInput[329] , 
        \matrixInput[328] , \matrixInput[327] , \matrixInput[326] , 
        \matrixInput[325] , \matrixInput[324] , \matrixInput[323] , 
        \matrixInput[322] , \matrixInput[321] , \matrixInput[320] , 
        \matrixInput[319] , \matrixInput[318] , \matrixInput[317] , 
        \matrixInput[316] , \matrixInput[315] , \matrixInput[314] , 
        \matrixInput[313] , \matrixInput[312] , \matrixInput[311] , 
        \matrixInput[310] , \matrixInput[309] , \matrixInput[308] , 
        \matrixInput[307] , \matrixInput[306] , \matrixInput[305] , 
        \matrixInput[304] , \matrixInput[303] , \matrixInput[302] , 
        \matrixInput[301] , \matrixInput[300] , \matrixInput[299] , 
        \matrixInput[298] , \matrixInput[297] , \matrixInput[296] , 
        \matrixInput[295] , \matrixInput[294] , \matrixInput[293] , 
        \matrixInput[292] , \matrixInput[291] , \matrixInput[290] , 
        \matrixInput[289] , \matrixInput[288] , \matrixInput[287] , 
        \matrixInput[286] , \matrixInput[285] , \matrixInput[284] , 
        \matrixInput[283] , \matrixInput[282] , \matrixInput[281] , 
        \matrixInput[280] , \matrixInput[279] , \matrixInput[278] , 
        \matrixInput[277] , \matrixInput[276] , \matrixInput[275] , 
        \matrixInput[274] , \matrixInput[273] , \matrixInput[272] , 
        \matrixInput[271] , \matrixInput[270] , \matrixInput[269] , 
        \matrixInput[268] , \matrixInput[267] , \matrixInput[266] , 
        \matrixInput[265] , \matrixInput[264] , \matrixInput[263] , 
        \matrixInput[262] , \matrixInput[261] , \matrixInput[260] , 
        \matrixInput[259] , \matrixInput[258] , \matrixInput[257] , 
        \matrixInput[256] , \matrixInput[255] , \matrixInput[254] , 
        \matrixInput[253] , \matrixInput[252] , \matrixInput[251] , 
        \matrixInput[250] , \matrixInput[249] , \matrixInput[248] , 
        \matrixInput[247] , \matrixInput[246] , \matrixInput[245] , 
        \matrixInput[244] , \matrixInput[243] , \matrixInput[242] , 
        \matrixInput[241] , \matrixInput[240] , \matrixInput[239] , 
        \matrixInput[238] , \matrixInput[237] , \matrixInput[236] , 
        \matrixInput[235] , \matrixInput[234] , \matrixInput[233] , 
        \matrixInput[232] , \matrixInput[231] , \matrixInput[230] , 
        \matrixInput[229] , \matrixInput[228] , \matrixInput[227] , 
        \matrixInput[226] , \matrixInput[225] , \matrixInput[224] , 
        \matrixInput[223] , \matrixInput[222] , \matrixInput[221] , 
        \matrixInput[220] , \matrixInput[219] , \matrixInput[218] , 
        \matrixInput[217] , \matrixInput[216] , \matrixInput[215] , 
        \matrixInput[214] , \matrixInput[213] , \matrixInput[212] , 
        \matrixInput[211] , \matrixInput[210] , \matrixInput[209] , 
        \matrixInput[208] , \matrixInput[207] , \matrixInput[206] , 
        \matrixInput[205] , \matrixInput[204] , \matrixInput[203] , 
        \matrixInput[202] , \matrixInput[201] , \matrixInput[200] , 
        \matrixInput[199] , \matrixInput[198] , \matrixInput[197] , 
        \matrixInput[196] , \matrixInput[195] , \matrixInput[194] , 
        \matrixInput[193] , \matrixInput[192] , \matrixInput[191] , 
        \matrixInput[190] , \matrixInput[189] , \matrixInput[188] , 
        \matrixInput[187] , \matrixInput[186] , \matrixInput[185] , 
        \matrixInput[184] , \matrixInput[183] , \matrixInput[182] , 
        \matrixInput[181] , \matrixInput[180] , \matrixInput[179] , 
        \matrixInput[178] , \matrixInput[177] , \matrixInput[176] , 
        \matrixInput[175] , \matrixInput[174] , \matrixInput[173] , 
        \matrixInput[172] , \matrixInput[171] , \matrixInput[170] , 
        \matrixInput[169] , \matrixInput[168] , \matrixInput[167] , 
        \matrixInput[166] , \matrixInput[165] , \matrixInput[164] , 
        \matrixInput[163] , \matrixInput[162] , \matrixInput[161] , 
        \matrixInput[160] , \matrixInput[159] , \matrixInput[158] , 
        \matrixInput[157] , \matrixInput[156] , \matrixInput[155] , 
        \matrixInput[154] , \matrixInput[153] , \matrixInput[152] , 
        \matrixInput[151] , \matrixInput[150] , \matrixInput[149] , 
        \matrixInput[148] , \matrixInput[147] , \matrixInput[146] , 
        \matrixInput[145] , \matrixInput[144] , \matrixInput[143] , 
        \matrixInput[142] , \matrixInput[141] , \matrixInput[140] , 
        \matrixInput[139] , \matrixInput[138] , \matrixInput[137] , 
        \matrixInput[136] , \matrixInput[135] , \matrixInput[134] , 
        \matrixInput[133] , \matrixInput[132] , \matrixInput[131] , 
        \matrixInput[130] , \matrixInput[129] , \matrixInput[128] , 
        \matrixInput[127] , \matrixInput[126] , \matrixInput[125] , 
        \matrixInput[124] , \matrixInput[123] , \matrixInput[122] , 
        \matrixInput[121] , \matrixInput[120] , \matrixInput[119] , 
        \matrixInput[118] , \matrixInput[117] , \matrixInput[116] , 
        \matrixInput[115] , \matrixInput[114] , \matrixInput[113] , 
        \matrixInput[112] , \matrixInput[111] , \matrixInput[110] , 
        \matrixInput[109] , \matrixInput[108] , \matrixInput[107] , 
        \matrixInput[106] , \matrixInput[105] , \matrixInput[104] , 
        \matrixInput[103] , \matrixInput[102] , \matrixInput[101] , 
        \matrixInput[100] , \matrixInput[99] , \matrixInput[98] , 
        \matrixInput[97] , \matrixInput[96] , \matrixInput[95] , 
        \matrixInput[94] , \matrixInput[93] , \matrixInput[92] , 
        \matrixInput[91] , \matrixInput[90] , \matrixInput[89] , 
        \matrixInput[88] , \matrixInput[87] , \matrixInput[86] , 
        \matrixInput[85] , \matrixInput[84] , \matrixInput[83] , 
        \matrixInput[82] , \matrixInput[81] , \matrixInput[80] , 
        \matrixInput[79] , \matrixInput[78] , \matrixInput[77] , 
        \matrixInput[76] , \matrixInput[75] , \matrixInput[74] , 
        \matrixInput[73] , \matrixInput[72] , \matrixInput[71] , 
        \matrixInput[70] , \matrixInput[69] , \matrixInput[68] , 
        \matrixInput[67] , \matrixInput[66] , \matrixInput[65] , 
        \matrixInput[64] , \matrixInput[63] , \matrixInput[62] , 
        \matrixInput[61] , \matrixInput[60] , \matrixInput[59] , 
        \matrixInput[58] , \matrixInput[57] , \matrixInput[56] , 
        \matrixInput[55] , \matrixInput[54] , \matrixInput[53] , 
        \matrixInput[52] , \matrixInput[51] , \matrixInput[50] , 
        \matrixInput[49] , \matrixInput[48] , \matrixInput[47] , 
        \matrixInput[46] , \matrixInput[45] , \matrixInput[44] , 
        \matrixInput[43] , \matrixInput[42] , \matrixInput[41] , 
        \matrixInput[40] , \matrixInput[39] , \matrixInput[38] , 
        \matrixInput[37] , \matrixInput[36] , \matrixInput[35] , 
        \matrixInput[34] , \matrixInput[33] , \matrixInput[32] , 
        \matrixInput[31] , \matrixInput[30] , \matrixInput[29] , 
        \matrixInput[28] , \matrixInput[27] , \matrixInput[26] , 
        \matrixInput[25] , \matrixInput[24] , \matrixInput[23] , 
        \matrixInput[22] , \matrixInput[21] , \matrixInput[20] , 
        \matrixInput[19] , \matrixInput[18] , \matrixInput[17] , 
        \matrixInput[16] , \matrixInput[15] , \matrixInput[14] , 
        \matrixInput[13] , \matrixInput[12] , \matrixInput[11] , 
        \matrixInput[10] , \matrixInput[9] , \matrixInput[8] , 
        \matrixInput[7] , \matrixInput[6] , \matrixInput[5] , \matrixInput[4] , 
        \matrixInput[3] , \matrixInput[2] , \matrixInput[1] , \matrixInput[0] 
        }), .cOutput({\cOutput[127] , \cOutput[126] , \cOutput[125] , 
        \cOutput[124] , \cOutput[123] , \cOutput[122] , \cOutput[121] , 
        \cOutput[120] , \cOutput[119] , \cOutput[118] , \cOutput[117] , 
        \cOutput[116] , \cOutput[115] , \cOutput[114] , \cOutput[113] , 
        \cOutput[112] , \cOutput[111] , \cOutput[110] , \cOutput[109] , 
        \cOutput[108] , \cOutput[107] , \cOutput[106] , \cOutput[105] , 
        \cOutput[104] , \cOutput[103] , \cOutput[102] , \cOutput[101] , 
        \cOutput[100] , \cOutput[99] , \cOutput[98] , \cOutput[97] , 
        \cOutput[96] , \cOutput[95] , \cOutput[94] , \cOutput[93] , 
        \cOutput[92] , \cOutput[91] , \cOutput[90] , \cOutput[89] , 
        \cOutput[88] , \cOutput[87] , \cOutput[86] , \cOutput[85] , 
        \cOutput[84] , \cOutput[83] , \cOutput[82] , \cOutput[81] , 
        \cOutput[80] , \cOutput[79] , \cOutput[78] , \cOutput[77] , 
        \cOutput[76] , \cOutput[75] , \cOutput[74] , \cOutput[73] , 
        \cOutput[72] , \cOutput[71] , \cOutput[70] , \cOutput[69] , 
        \cOutput[68] , \cOutput[67] , \cOutput[66] , \cOutput[65] , 
        \cOutput[64] , \cOutput[63] , \cOutput[62] , \cOutput[61] , 
        \cOutput[60] , \cOutput[59] , \cOutput[58] , \cOutput[57] , 
        \cOutput[56] , \cOutput[55] , \cOutput[54] , \cOutput[53] , 
        \cOutput[52] , \cOutput[51] , \cOutput[50] , \cOutput[49] , 
        \cOutput[48] , \cOutput[47] , \cOutput[46] , \cOutput[45] , 
        \cOutput[44] , \cOutput[43] , \cOutput[42] , \cOutput[41] , 
        \cOutput[40] , \cOutput[39] , \cOutput[38] , \cOutput[37] , 
        \cOutput[36] , \cOutput[35] , \cOutput[34] , \cOutput[33] , 
        \cOutput[32] , \cOutput[31] , \cOutput[30] , \cOutput[29] , 
        \cOutput[28] , \cOutput[27] , \cOutput[26] , \cOutput[25] , 
        \cOutput[24] , \cOutput[23] , \cOutput[22] , \cOutput[21] , 
        \cOutput[20] , \cOutput[19] , \cOutput[18] , \cOutput[17] , 
        \cOutput[16] , \cOutput[15] , \cOutput[14] , \cOutput[13] , 
        \cOutput[12] , \cOutput[11] , \cOutput[10] , \cOutput[9] , 
        \cOutput[8] , \cOutput[7] , \cOutput[6] , \cOutput[5] , \cOutput[4] , 
        \cOutput[3] , \cOutput[2] , \cOutput[1] , \cOutput[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[255] , \matrixInput[254] , \matrixInput[253] , 
        \matrixInput[252] , \matrixInput[251] , \matrixInput[250] , 
        \matrixInput[249] , \matrixInput[248] , \matrixInput[247] , 
        \matrixInput[246] , \matrixInput[245] , \matrixInput[244] , 
        \matrixInput[243] , \matrixInput[242] , \matrixInput[241] , 
        \matrixInput[240] , \matrixInput[239] , \matrixInput[238] , 
        \matrixInput[237] , \matrixInput[236] , \matrixInput[235] , 
        \matrixInput[234] , \matrixInput[233] , \matrixInput[232] , 
        \matrixInput[231] , \matrixInput[230] , \matrixInput[229] , 
        \matrixInput[228] , \matrixInput[227] , \matrixInput[226] , 
        \matrixInput[225] , \matrixInput[224] , \matrixInput[223] , 
        \matrixInput[222] , \matrixInput[221] , \matrixInput[220] , 
        \matrixInput[219] , \matrixInput[218] , \matrixInput[217] , 
        \matrixInput[216] , \matrixInput[215] , \matrixInput[214] , 
        \matrixInput[213] , \matrixInput[212] , \matrixInput[211] , 
        \matrixInput[210] , \matrixInput[209] , \matrixInput[208] , 
        \matrixInput[207] , \matrixInput[206] , \matrixInput[205] , 
        \matrixInput[204] , \matrixInput[203] , \matrixInput[202] , 
        \matrixInput[201] , \matrixInput[200] , \matrixInput[199] , 
        \matrixInput[198] , \matrixInput[197] , \matrixInput[196] , 
        \matrixInput[195] , \matrixInput[194] , \matrixInput[193] , 
        \matrixInput[192] , \matrixInput[191] , \matrixInput[190] , 
        \matrixInput[189] , \matrixInput[188] , \matrixInput[187] , 
        \matrixInput[186] , \matrixInput[185] , \matrixInput[184] , 
        \matrixInput[183] , \matrixInput[182] , \matrixInput[181] , 
        \matrixInput[180] , \matrixInput[179] , \matrixInput[178] , 
        \matrixInput[177] , \matrixInput[176] , \matrixInput[175] , 
        \matrixInput[174] , \matrixInput[173] , \matrixInput[172] , 
        \matrixInput[171] , \matrixInput[170] , \matrixInput[169] , 
        \matrixInput[168] , \matrixInput[167] , \matrixInput[166] , 
        \matrixInput[165] , \matrixInput[164] , \matrixInput[163] , 
        \matrixInput[162] , \matrixInput[161] , \matrixInput[160] , 
        \matrixInput[159] , \matrixInput[158] , \matrixInput[157] , 
        \matrixInput[156] , \matrixInput[155] , \matrixInput[154] , 
        \matrixInput[153] , \matrixInput[152] , \matrixInput[151] , 
        \matrixInput[150] , \matrixInput[149] , \matrixInput[148] , 
        \matrixInput[147] , \matrixInput[146] , \matrixInput[145] , 
        \matrixInput[144] , \matrixInput[143] , \matrixInput[142] , 
        \matrixInput[141] , \matrixInput[140] , \matrixInput[139] , 
        \matrixInput[138] , \matrixInput[137] , \matrixInput[136] , 
        \matrixInput[135] , \matrixInput[134] , \matrixInput[133] , 
        \matrixInput[132] , \matrixInput[131] , \matrixInput[130] , 
        \matrixInput[129] , \matrixInput[128] }), .cOutput({\cOutput[15] , 
        \cOutput[14] , \cOutput[13] , \cOutput[12] , \cOutput[11] , 
        \cOutput[10] , \cOutput[9] , \cOutput[8] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[383] , \matrixInput[382] , \matrixInput[381] , 
        \matrixInput[380] , \matrixInput[379] , \matrixInput[378] , 
        \matrixInput[377] , \matrixInput[376] , \matrixInput[375] , 
        \matrixInput[374] , \matrixInput[373] , \matrixInput[372] , 
        \matrixInput[371] , \matrixInput[370] , \matrixInput[369] , 
        \matrixInput[368] , \matrixInput[367] , \matrixInput[366] , 
        \matrixInput[365] , \matrixInput[364] , \matrixInput[363] , 
        \matrixInput[362] , \matrixInput[361] , \matrixInput[360] , 
        \matrixInput[359] , \matrixInput[358] , \matrixInput[357] , 
        \matrixInput[356] , \matrixInput[355] , \matrixInput[354] , 
        \matrixInput[353] , \matrixInput[352] , \matrixInput[351] , 
        \matrixInput[350] , \matrixInput[349] , \matrixInput[348] , 
        \matrixInput[347] , \matrixInput[346] , \matrixInput[345] , 
        \matrixInput[344] , \matrixInput[343] , \matrixInput[342] , 
        \matrixInput[341] , \matrixInput[340] , \matrixInput[339] , 
        \matrixInput[338] , \matrixInput[337] , \matrixInput[336] , 
        \matrixInput[335] , \matrixInput[334] , \matrixInput[333] , 
        \matrixInput[332] , \matrixInput[331] , \matrixInput[330] , 
        \matrixInput[329] , \matrixInput[328] , \matrixInput[327] , 
        \matrixInput[326] , \matrixInput[325] , \matrixInput[324] , 
        \matrixInput[323] , \matrixInput[322] , \matrixInput[321] , 
        \matrixInput[320] , \matrixInput[319] , \matrixInput[318] , 
        \matrixInput[317] , \matrixInput[316] , \matrixInput[315] , 
        \matrixInput[314] , \matrixInput[313] , \matrixInput[312] , 
        \matrixInput[311] , \matrixInput[310] , \matrixInput[309] , 
        \matrixInput[308] , \matrixInput[307] , \matrixInput[306] , 
        \matrixInput[305] , \matrixInput[304] , \matrixInput[303] , 
        \matrixInput[302] , \matrixInput[301] , \matrixInput[300] , 
        \matrixInput[299] , \matrixInput[298] , \matrixInput[297] , 
        \matrixInput[296] , \matrixInput[295] , \matrixInput[294] , 
        \matrixInput[293] , \matrixInput[292] , \matrixInput[291] , 
        \matrixInput[290] , \matrixInput[289] , \matrixInput[288] , 
        \matrixInput[287] , \matrixInput[286] , \matrixInput[285] , 
        \matrixInput[284] , \matrixInput[283] , \matrixInput[282] , 
        \matrixInput[281] , \matrixInput[280] , \matrixInput[279] , 
        \matrixInput[278] , \matrixInput[277] , \matrixInput[276] , 
        \matrixInput[275] , \matrixInput[274] , \matrixInput[273] , 
        \matrixInput[272] , \matrixInput[271] , \matrixInput[270] , 
        \matrixInput[269] , \matrixInput[268] , \matrixInput[267] , 
        \matrixInput[266] , \matrixInput[265] , \matrixInput[264] , 
        \matrixInput[263] , \matrixInput[262] , \matrixInput[261] , 
        \matrixInput[260] , \matrixInput[259] , \matrixInput[258] , 
        \matrixInput[257] , \matrixInput[256] }), .cOutput({\cOutput[23] , 
        \cOutput[22] , \cOutput[21] , \cOutput[20] , \cOutput[19] , 
        \cOutput[18] , \cOutput[17] , \cOutput[16] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1919] , \matrixInput[1918] , \matrixInput[1917] , 
        \matrixInput[1916] , \matrixInput[1915] , \matrixInput[1914] , 
        \matrixInput[1913] , \matrixInput[1912] , \matrixInput[1911] , 
        \matrixInput[1910] , \matrixInput[1909] , \matrixInput[1908] , 
        \matrixInput[1907] , \matrixInput[1906] , \matrixInput[1905] , 
        \matrixInput[1904] , \matrixInput[1903] , \matrixInput[1902] , 
        \matrixInput[1901] , \matrixInput[1900] , \matrixInput[1899] , 
        \matrixInput[1898] , \matrixInput[1897] , \matrixInput[1896] , 
        \matrixInput[1895] , \matrixInput[1894] , \matrixInput[1893] , 
        \matrixInput[1892] , \matrixInput[1891] , \matrixInput[1890] , 
        \matrixInput[1889] , \matrixInput[1888] , \matrixInput[1887] , 
        \matrixInput[1886] , \matrixInput[1885] , \matrixInput[1884] , 
        \matrixInput[1883] , \matrixInput[1882] , \matrixInput[1881] , 
        \matrixInput[1880] , \matrixInput[1879] , \matrixInput[1878] , 
        \matrixInput[1877] , \matrixInput[1876] , \matrixInput[1875] , 
        \matrixInput[1874] , \matrixInput[1873] , \matrixInput[1872] , 
        \matrixInput[1871] , \matrixInput[1870] , \matrixInput[1869] , 
        \matrixInput[1868] , \matrixInput[1867] , \matrixInput[1866] , 
        \matrixInput[1865] , \matrixInput[1864] , \matrixInput[1863] , 
        \matrixInput[1862] , \matrixInput[1861] , \matrixInput[1860] , 
        \matrixInput[1859] , \matrixInput[1858] , \matrixInput[1857] , 
        \matrixInput[1856] , \matrixInput[1855] , \matrixInput[1854] , 
        \matrixInput[1853] , \matrixInput[1852] , \matrixInput[1851] , 
        \matrixInput[1850] , \matrixInput[1849] , \matrixInput[1848] , 
        \matrixInput[1847] , \matrixInput[1846] , \matrixInput[1845] , 
        \matrixInput[1844] , \matrixInput[1843] , \matrixInput[1842] , 
        \matrixInput[1841] , \matrixInput[1840] , \matrixInput[1839] , 
        \matrixInput[1838] , \matrixInput[1837] , \matrixInput[1836] , 
        \matrixInput[1835] , \matrixInput[1834] , \matrixInput[1833] , 
        \matrixInput[1832] , \matrixInput[1831] , \matrixInput[1830] , 
        \matrixInput[1829] , \matrixInput[1828] , \matrixInput[1827] , 
        \matrixInput[1826] , \matrixInput[1825] , \matrixInput[1824] , 
        \matrixInput[1823] , \matrixInput[1822] , \matrixInput[1821] , 
        \matrixInput[1820] , \matrixInput[1819] , \matrixInput[1818] , 
        \matrixInput[1817] , \matrixInput[1816] , \matrixInput[1815] , 
        \matrixInput[1814] , \matrixInput[1813] , \matrixInput[1812] , 
        \matrixInput[1811] , \matrixInput[1810] , \matrixInput[1809] , 
        \matrixInput[1808] , \matrixInput[1807] , \matrixInput[1806] , 
        \matrixInput[1805] , \matrixInput[1804] , \matrixInput[1803] , 
        \matrixInput[1802] , \matrixInput[1801] , \matrixInput[1800] , 
        \matrixInput[1799] , \matrixInput[1798] , \matrixInput[1797] , 
        \matrixInput[1796] , \matrixInput[1795] , \matrixInput[1794] , 
        \matrixInput[1793] , \matrixInput[1792] }), .cOutput({\cOutput[119] , 
        \cOutput[118] , \cOutput[117] , \cOutput[116] , \cOutput[115] , 
        \cOutput[114] , \cOutput[113] , \cOutput[112] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[511] , \matrixInput[510] , \matrixInput[509] , 
        \matrixInput[508] , \matrixInput[507] , \matrixInput[506] , 
        \matrixInput[505] , \matrixInput[504] , \matrixInput[503] , 
        \matrixInput[502] , \matrixInput[501] , \matrixInput[500] , 
        \matrixInput[499] , \matrixInput[498] , \matrixInput[497] , 
        \matrixInput[496] , \matrixInput[495] , \matrixInput[494] , 
        \matrixInput[493] , \matrixInput[492] , \matrixInput[491] , 
        \matrixInput[490] , \matrixInput[489] , \matrixInput[488] , 
        \matrixInput[487] , \matrixInput[486] , \matrixInput[485] , 
        \matrixInput[484] , \matrixInput[483] , \matrixInput[482] , 
        \matrixInput[481] , \matrixInput[480] , \matrixInput[479] , 
        \matrixInput[478] , \matrixInput[477] , \matrixInput[476] , 
        \matrixInput[475] , \matrixInput[474] , \matrixInput[473] , 
        \matrixInput[472] , \matrixInput[471] , \matrixInput[470] , 
        \matrixInput[469] , \matrixInput[468] , \matrixInput[467] , 
        \matrixInput[466] , \matrixInput[465] , \matrixInput[464] , 
        \matrixInput[463] , \matrixInput[462] , \matrixInput[461] , 
        \matrixInput[460] , \matrixInput[459] , \matrixInput[458] , 
        \matrixInput[457] , \matrixInput[456] , \matrixInput[455] , 
        \matrixInput[454] , \matrixInput[453] , \matrixInput[452] , 
        \matrixInput[451] , \matrixInput[450] , \matrixInput[449] , 
        \matrixInput[448] , \matrixInput[447] , \matrixInput[446] , 
        \matrixInput[445] , \matrixInput[444] , \matrixInput[443] , 
        \matrixInput[442] , \matrixInput[441] , \matrixInput[440] , 
        \matrixInput[439] , \matrixInput[438] , \matrixInput[437] , 
        \matrixInput[436] , \matrixInput[435] , \matrixInput[434] , 
        \matrixInput[433] , \matrixInput[432] , \matrixInput[431] , 
        \matrixInput[430] , \matrixInput[429] , \matrixInput[428] , 
        \matrixInput[427] , \matrixInput[426] , \matrixInput[425] , 
        \matrixInput[424] , \matrixInput[423] , \matrixInput[422] , 
        \matrixInput[421] , \matrixInput[420] , \matrixInput[419] , 
        \matrixInput[418] , \matrixInput[417] , \matrixInput[416] , 
        \matrixInput[415] , \matrixInput[414] , \matrixInput[413] , 
        \matrixInput[412] , \matrixInput[411] , \matrixInput[410] , 
        \matrixInput[409] , \matrixInput[408] , \matrixInput[407] , 
        \matrixInput[406] , \matrixInput[405] , \matrixInput[404] , 
        \matrixInput[403] , \matrixInput[402] , \matrixInput[401] , 
        \matrixInput[400] , \matrixInput[399] , \matrixInput[398] , 
        \matrixInput[397] , \matrixInput[396] , \matrixInput[395] , 
        \matrixInput[394] , \matrixInput[393] , \matrixInput[392] , 
        \matrixInput[391] , \matrixInput[390] , \matrixInput[389] , 
        \matrixInput[388] , \matrixInput[387] , \matrixInput[386] , 
        \matrixInput[385] , \matrixInput[384] }), .cOutput({\cOutput[31] , 
        \cOutput[30] , \cOutput[29] , \cOutput[28] , \cOutput[27] , 
        \cOutput[26] , \cOutput[25] , \cOutput[24] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[639] , \matrixInput[638] , \matrixInput[637] , 
        \matrixInput[636] , \matrixInput[635] , \matrixInput[634] , 
        \matrixInput[633] , \matrixInput[632] , \matrixInput[631] , 
        \matrixInput[630] , \matrixInput[629] , \matrixInput[628] , 
        \matrixInput[627] , \matrixInput[626] , \matrixInput[625] , 
        \matrixInput[624] , \matrixInput[623] , \matrixInput[622] , 
        \matrixInput[621] , \matrixInput[620] , \matrixInput[619] , 
        \matrixInput[618] , \matrixInput[617] , \matrixInput[616] , 
        \matrixInput[615] , \matrixInput[614] , \matrixInput[613] , 
        \matrixInput[612] , \matrixInput[611] , \matrixInput[610] , 
        \matrixInput[609] , \matrixInput[608] , \matrixInput[607] , 
        \matrixInput[606] , \matrixInput[605] , \matrixInput[604] , 
        \matrixInput[603] , \matrixInput[602] , \matrixInput[601] , 
        \matrixInput[600] , \matrixInput[599] , \matrixInput[598] , 
        \matrixInput[597] , \matrixInput[596] , \matrixInput[595] , 
        \matrixInput[594] , \matrixInput[593] , \matrixInput[592] , 
        \matrixInput[591] , \matrixInput[590] , \matrixInput[589] , 
        \matrixInput[588] , \matrixInput[587] , \matrixInput[586] , 
        \matrixInput[585] , \matrixInput[584] , \matrixInput[583] , 
        \matrixInput[582] , \matrixInput[581] , \matrixInput[580] , 
        \matrixInput[579] , \matrixInput[578] , \matrixInput[577] , 
        \matrixInput[576] , \matrixInput[575] , \matrixInput[574] , 
        \matrixInput[573] , \matrixInput[572] , \matrixInput[571] , 
        \matrixInput[570] , \matrixInput[569] , \matrixInput[568] , 
        \matrixInput[567] , \matrixInput[566] , \matrixInput[565] , 
        \matrixInput[564] , \matrixInput[563] , \matrixInput[562] , 
        \matrixInput[561] , \matrixInput[560] , \matrixInput[559] , 
        \matrixInput[558] , \matrixInput[557] , \matrixInput[556] , 
        \matrixInput[555] , \matrixInput[554] , \matrixInput[553] , 
        \matrixInput[552] , \matrixInput[551] , \matrixInput[550] , 
        \matrixInput[549] , \matrixInput[548] , \matrixInput[547] , 
        \matrixInput[546] , \matrixInput[545] , \matrixInput[544] , 
        \matrixInput[543] , \matrixInput[542] , \matrixInput[541] , 
        \matrixInput[540] , \matrixInput[539] , \matrixInput[538] , 
        \matrixInput[537] , \matrixInput[536] , \matrixInput[535] , 
        \matrixInput[534] , \matrixInput[533] , \matrixInput[532] , 
        \matrixInput[531] , \matrixInput[530] , \matrixInput[529] , 
        \matrixInput[528] , \matrixInput[527] , \matrixInput[526] , 
        \matrixInput[525] , \matrixInput[524] , \matrixInput[523] , 
        \matrixInput[522] , \matrixInput[521] , \matrixInput[520] , 
        \matrixInput[519] , \matrixInput[518] , \matrixInput[517] , 
        \matrixInput[516] , \matrixInput[515] , \matrixInput[514] , 
        \matrixInput[513] , \matrixInput[512] }), .cOutput({\cOutput[39] , 
        \cOutput[38] , \cOutput[37] , \cOutput[36] , \cOutput[35] , 
        \cOutput[34] , \cOutput[33] , \cOutput[32] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[767] , \matrixInput[766] , \matrixInput[765] , 
        \matrixInput[764] , \matrixInput[763] , \matrixInput[762] , 
        \matrixInput[761] , \matrixInput[760] , \matrixInput[759] , 
        \matrixInput[758] , \matrixInput[757] , \matrixInput[756] , 
        \matrixInput[755] , \matrixInput[754] , \matrixInput[753] , 
        \matrixInput[752] , \matrixInput[751] , \matrixInput[750] , 
        \matrixInput[749] , \matrixInput[748] , \matrixInput[747] , 
        \matrixInput[746] , \matrixInput[745] , \matrixInput[744] , 
        \matrixInput[743] , \matrixInput[742] , \matrixInput[741] , 
        \matrixInput[740] , \matrixInput[739] , \matrixInput[738] , 
        \matrixInput[737] , \matrixInput[736] , \matrixInput[735] , 
        \matrixInput[734] , \matrixInput[733] , \matrixInput[732] , 
        \matrixInput[731] , \matrixInput[730] , \matrixInput[729] , 
        \matrixInput[728] , \matrixInput[727] , \matrixInput[726] , 
        \matrixInput[725] , \matrixInput[724] , \matrixInput[723] , 
        \matrixInput[722] , \matrixInput[721] , \matrixInput[720] , 
        \matrixInput[719] , \matrixInput[718] , \matrixInput[717] , 
        \matrixInput[716] , \matrixInput[715] , \matrixInput[714] , 
        \matrixInput[713] , \matrixInput[712] , \matrixInput[711] , 
        \matrixInput[710] , \matrixInput[709] , \matrixInput[708] , 
        \matrixInput[707] , \matrixInput[706] , \matrixInput[705] , 
        \matrixInput[704] , \matrixInput[703] , \matrixInput[702] , 
        \matrixInput[701] , \matrixInput[700] , \matrixInput[699] , 
        \matrixInput[698] , \matrixInput[697] , \matrixInput[696] , 
        \matrixInput[695] , \matrixInput[694] , \matrixInput[693] , 
        \matrixInput[692] , \matrixInput[691] , \matrixInput[690] , 
        \matrixInput[689] , \matrixInput[688] , \matrixInput[687] , 
        \matrixInput[686] , \matrixInput[685] , \matrixInput[684] , 
        \matrixInput[683] , \matrixInput[682] , \matrixInput[681] , 
        \matrixInput[680] , \matrixInput[679] , \matrixInput[678] , 
        \matrixInput[677] , \matrixInput[676] , \matrixInput[675] , 
        \matrixInput[674] , \matrixInput[673] , \matrixInput[672] , 
        \matrixInput[671] , \matrixInput[670] , \matrixInput[669] , 
        \matrixInput[668] , \matrixInput[667] , \matrixInput[666] , 
        \matrixInput[665] , \matrixInput[664] , \matrixInput[663] , 
        \matrixInput[662] , \matrixInput[661] , \matrixInput[660] , 
        \matrixInput[659] , \matrixInput[658] , \matrixInput[657] , 
        \matrixInput[656] , \matrixInput[655] , \matrixInput[654] , 
        \matrixInput[653] , \matrixInput[652] , \matrixInput[651] , 
        \matrixInput[650] , \matrixInput[649] , \matrixInput[648] , 
        \matrixInput[647] , \matrixInput[646] , \matrixInput[645] , 
        \matrixInput[644] , \matrixInput[643] , \matrixInput[642] , 
        \matrixInput[641] , \matrixInput[640] }), .cOutput({\cOutput[47] , 
        \cOutput[46] , \cOutput[45] , \cOutput[44] , \cOutput[43] , 
        \cOutput[42] , \cOutput[41] , \cOutput[40] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1663] , \matrixInput[1662] , \matrixInput[1661] , 
        \matrixInput[1660] , \matrixInput[1659] , \matrixInput[1658] , 
        \matrixInput[1657] , \matrixInput[1656] , \matrixInput[1655] , 
        \matrixInput[1654] , \matrixInput[1653] , \matrixInput[1652] , 
        \matrixInput[1651] , \matrixInput[1650] , \matrixInput[1649] , 
        \matrixInput[1648] , \matrixInput[1647] , \matrixInput[1646] , 
        \matrixInput[1645] , \matrixInput[1644] , \matrixInput[1643] , 
        \matrixInput[1642] , \matrixInput[1641] , \matrixInput[1640] , 
        \matrixInput[1639] , \matrixInput[1638] , \matrixInput[1637] , 
        \matrixInput[1636] , \matrixInput[1635] , \matrixInput[1634] , 
        \matrixInput[1633] , \matrixInput[1632] , \matrixInput[1631] , 
        \matrixInput[1630] , \matrixInput[1629] , \matrixInput[1628] , 
        \matrixInput[1627] , \matrixInput[1626] , \matrixInput[1625] , 
        \matrixInput[1624] , \matrixInput[1623] , \matrixInput[1622] , 
        \matrixInput[1621] , \matrixInput[1620] , \matrixInput[1619] , 
        \matrixInput[1618] , \matrixInput[1617] , \matrixInput[1616] , 
        \matrixInput[1615] , \matrixInput[1614] , \matrixInput[1613] , 
        \matrixInput[1612] , \matrixInput[1611] , \matrixInput[1610] , 
        \matrixInput[1609] , \matrixInput[1608] , \matrixInput[1607] , 
        \matrixInput[1606] , \matrixInput[1605] , \matrixInput[1604] , 
        \matrixInput[1603] , \matrixInput[1602] , \matrixInput[1601] , 
        \matrixInput[1600] , \matrixInput[1599] , \matrixInput[1598] , 
        \matrixInput[1597] , \matrixInput[1596] , \matrixInput[1595] , 
        \matrixInput[1594] , \matrixInput[1593] , \matrixInput[1592] , 
        \matrixInput[1591] , \matrixInput[1590] , \matrixInput[1589] , 
        \matrixInput[1588] , \matrixInput[1587] , \matrixInput[1586] , 
        \matrixInput[1585] , \matrixInput[1584] , \matrixInput[1583] , 
        \matrixInput[1582] , \matrixInput[1581] , \matrixInput[1580] , 
        \matrixInput[1579] , \matrixInput[1578] , \matrixInput[1577] , 
        \matrixInput[1576] , \matrixInput[1575] , \matrixInput[1574] , 
        \matrixInput[1573] , \matrixInput[1572] , \matrixInput[1571] , 
        \matrixInput[1570] , \matrixInput[1569] , \matrixInput[1568] , 
        \matrixInput[1567] , \matrixInput[1566] , \matrixInput[1565] , 
        \matrixInput[1564] , \matrixInput[1563] , \matrixInput[1562] , 
        \matrixInput[1561] , \matrixInput[1560] , \matrixInput[1559] , 
        \matrixInput[1558] , \matrixInput[1557] , \matrixInput[1556] , 
        \matrixInput[1555] , \matrixInput[1554] , \matrixInput[1553] , 
        \matrixInput[1552] , \matrixInput[1551] , \matrixInput[1550] , 
        \matrixInput[1549] , \matrixInput[1548] , \matrixInput[1547] , 
        \matrixInput[1546] , \matrixInput[1545] , \matrixInput[1544] , 
        \matrixInput[1543] , \matrixInput[1542] , \matrixInput[1541] , 
        \matrixInput[1540] , \matrixInput[1539] , \matrixInput[1538] , 
        \matrixInput[1537] , \matrixInput[1536] }), .cOutput({\cOutput[103] , 
        \cOutput[102] , \cOutput[101] , \cOutput[100] , \cOutput[99] , 
        \cOutput[98] , \cOutput[97] , \cOutput[96] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1791] , \matrixInput[1790] , \matrixInput[1789] , 
        \matrixInput[1788] , \matrixInput[1787] , \matrixInput[1786] , 
        \matrixInput[1785] , \matrixInput[1784] , \matrixInput[1783] , 
        \matrixInput[1782] , \matrixInput[1781] , \matrixInput[1780] , 
        \matrixInput[1779] , \matrixInput[1778] , \matrixInput[1777] , 
        \matrixInput[1776] , \matrixInput[1775] , \matrixInput[1774] , 
        \matrixInput[1773] , \matrixInput[1772] , \matrixInput[1771] , 
        \matrixInput[1770] , \matrixInput[1769] , \matrixInput[1768] , 
        \matrixInput[1767] , \matrixInput[1766] , \matrixInput[1765] , 
        \matrixInput[1764] , \matrixInput[1763] , \matrixInput[1762] , 
        \matrixInput[1761] , \matrixInput[1760] , \matrixInput[1759] , 
        \matrixInput[1758] , \matrixInput[1757] , \matrixInput[1756] , 
        \matrixInput[1755] , \matrixInput[1754] , \matrixInput[1753] , 
        \matrixInput[1752] , \matrixInput[1751] , \matrixInput[1750] , 
        \matrixInput[1749] , \matrixInput[1748] , \matrixInput[1747] , 
        \matrixInput[1746] , \matrixInput[1745] , \matrixInput[1744] , 
        \matrixInput[1743] , \matrixInput[1742] , \matrixInput[1741] , 
        \matrixInput[1740] , \matrixInput[1739] , \matrixInput[1738] , 
        \matrixInput[1737] , \matrixInput[1736] , \matrixInput[1735] , 
        \matrixInput[1734] , \matrixInput[1733] , \matrixInput[1732] , 
        \matrixInput[1731] , \matrixInput[1730] , \matrixInput[1729] , 
        \matrixInput[1728] , \matrixInput[1727] , \matrixInput[1726] , 
        \matrixInput[1725] , \matrixInput[1724] , \matrixInput[1723] , 
        \matrixInput[1722] , \matrixInput[1721] , \matrixInput[1720] , 
        \matrixInput[1719] , \matrixInput[1718] , \matrixInput[1717] , 
        \matrixInput[1716] , \matrixInput[1715] , \matrixInput[1714] , 
        \matrixInput[1713] , \matrixInput[1712] , \matrixInput[1711] , 
        \matrixInput[1710] , \matrixInput[1709] , \matrixInput[1708] , 
        \matrixInput[1707] , \matrixInput[1706] , \matrixInput[1705] , 
        \matrixInput[1704] , \matrixInput[1703] , \matrixInput[1702] , 
        \matrixInput[1701] , \matrixInput[1700] , \matrixInput[1699] , 
        \matrixInput[1698] , \matrixInput[1697] , \matrixInput[1696] , 
        \matrixInput[1695] , \matrixInput[1694] , \matrixInput[1693] , 
        \matrixInput[1692] , \matrixInput[1691] , \matrixInput[1690] , 
        \matrixInput[1689] , \matrixInput[1688] , \matrixInput[1687] , 
        \matrixInput[1686] , \matrixInput[1685] , \matrixInput[1684] , 
        \matrixInput[1683] , \matrixInput[1682] , \matrixInput[1681] , 
        \matrixInput[1680] , \matrixInput[1679] , \matrixInput[1678] , 
        \matrixInput[1677] , \matrixInput[1676] , \matrixInput[1675] , 
        \matrixInput[1674] , \matrixInput[1673] , \matrixInput[1672] , 
        \matrixInput[1671] , \matrixInput[1670] , \matrixInput[1669] , 
        \matrixInput[1668] , \matrixInput[1667] , \matrixInput[1666] , 
        \matrixInput[1665] , \matrixInput[1664] }), .cOutput({\cOutput[111] , 
        \cOutput[110] , \cOutput[109] , \cOutput[108] , \cOutput[107] , 
        \cOutput[106] , \cOutput[105] , \cOutput[104] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[2047] , \matrixInput[2046] , \matrixInput[2045] , 
        \matrixInput[2044] , \matrixInput[2043] , \matrixInput[2042] , 
        \matrixInput[2041] , \matrixInput[2040] , \matrixInput[2039] , 
        \matrixInput[2038] , \matrixInput[2037] , \matrixInput[2036] , 
        \matrixInput[2035] , \matrixInput[2034] , \matrixInput[2033] , 
        \matrixInput[2032] , \matrixInput[2031] , \matrixInput[2030] , 
        \matrixInput[2029] , \matrixInput[2028] , \matrixInput[2027] , 
        \matrixInput[2026] , \matrixInput[2025] , \matrixInput[2024] , 
        \matrixInput[2023] , \matrixInput[2022] , \matrixInput[2021] , 
        \matrixInput[2020] , \matrixInput[2019] , \matrixInput[2018] , 
        \matrixInput[2017] , \matrixInput[2016] , \matrixInput[2015] , 
        \matrixInput[2014] , \matrixInput[2013] , \matrixInput[2012] , 
        \matrixInput[2011] , \matrixInput[2010] , \matrixInput[2009] , 
        \matrixInput[2008] , \matrixInput[2007] , \matrixInput[2006] , 
        \matrixInput[2005] , \matrixInput[2004] , \matrixInput[2003] , 
        \matrixInput[2002] , \matrixInput[2001] , \matrixInput[2000] , 
        \matrixInput[1999] , \matrixInput[1998] , \matrixInput[1997] , 
        \matrixInput[1996] , \matrixInput[1995] , \matrixInput[1994] , 
        \matrixInput[1993] , \matrixInput[1992] , \matrixInput[1991] , 
        \matrixInput[1990] , \matrixInput[1989] , \matrixInput[1988] , 
        \matrixInput[1987] , \matrixInput[1986] , \matrixInput[1985] , 
        \matrixInput[1984] , \matrixInput[1983] , \matrixInput[1982] , 
        \matrixInput[1981] , \matrixInput[1980] , \matrixInput[1979] , 
        \matrixInput[1978] , \matrixInput[1977] , \matrixInput[1976] , 
        \matrixInput[1975] , \matrixInput[1974] , \matrixInput[1973] , 
        \matrixInput[1972] , \matrixInput[1971] , \matrixInput[1970] , 
        \matrixInput[1969] , \matrixInput[1968] , \matrixInput[1967] , 
        \matrixInput[1966] , \matrixInput[1965] , \matrixInput[1964] , 
        \matrixInput[1963] , \matrixInput[1962] , \matrixInput[1961] , 
        \matrixInput[1960] , \matrixInput[1959] , \matrixInput[1958] , 
        \matrixInput[1957] , \matrixInput[1956] , \matrixInput[1955] , 
        \matrixInput[1954] , \matrixInput[1953] , \matrixInput[1952] , 
        \matrixInput[1951] , \matrixInput[1950] , \matrixInput[1949] , 
        \matrixInput[1948] , \matrixInput[1947] , \matrixInput[1946] , 
        \matrixInput[1945] , \matrixInput[1944] , \matrixInput[1943] , 
        \matrixInput[1942] , \matrixInput[1941] , \matrixInput[1940] , 
        \matrixInput[1939] , \matrixInput[1938] , \matrixInput[1937] , 
        \matrixInput[1936] , \matrixInput[1935] , \matrixInput[1934] , 
        \matrixInput[1933] , \matrixInput[1932] , \matrixInput[1931] , 
        \matrixInput[1930] , \matrixInput[1929] , \matrixInput[1928] , 
        \matrixInput[1927] , \matrixInput[1926] , \matrixInput[1925] , 
        \matrixInput[1924] , \matrixInput[1923] , \matrixInput[1922] , 
        \matrixInput[1921] , \matrixInput[1920] }), .cOutput({\cOutput[127] , 
        \cOutput[126] , \cOutput[125] , \cOutput[124] , \cOutput[123] , 
        \cOutput[122] , \cOutput[121] , \cOutput[120] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[895] , \matrixInput[894] , \matrixInput[893] , 
        \matrixInput[892] , \matrixInput[891] , \matrixInput[890] , 
        \matrixInput[889] , \matrixInput[888] , \matrixInput[887] , 
        \matrixInput[886] , \matrixInput[885] , \matrixInput[884] , 
        \matrixInput[883] , \matrixInput[882] , \matrixInput[881] , 
        \matrixInput[880] , \matrixInput[879] , \matrixInput[878] , 
        \matrixInput[877] , \matrixInput[876] , \matrixInput[875] , 
        \matrixInput[874] , \matrixInput[873] , \matrixInput[872] , 
        \matrixInput[871] , \matrixInput[870] , \matrixInput[869] , 
        \matrixInput[868] , \matrixInput[867] , \matrixInput[866] , 
        \matrixInput[865] , \matrixInput[864] , \matrixInput[863] , 
        \matrixInput[862] , \matrixInput[861] , \matrixInput[860] , 
        \matrixInput[859] , \matrixInput[858] , \matrixInput[857] , 
        \matrixInput[856] , \matrixInput[855] , \matrixInput[854] , 
        \matrixInput[853] , \matrixInput[852] , \matrixInput[851] , 
        \matrixInput[850] , \matrixInput[849] , \matrixInput[848] , 
        \matrixInput[847] , \matrixInput[846] , \matrixInput[845] , 
        \matrixInput[844] , \matrixInput[843] , \matrixInput[842] , 
        \matrixInput[841] , \matrixInput[840] , \matrixInput[839] , 
        \matrixInput[838] , \matrixInput[837] , \matrixInput[836] , 
        \matrixInput[835] , \matrixInput[834] , \matrixInput[833] , 
        \matrixInput[832] , \matrixInput[831] , \matrixInput[830] , 
        \matrixInput[829] , \matrixInput[828] , \matrixInput[827] , 
        \matrixInput[826] , \matrixInput[825] , \matrixInput[824] , 
        \matrixInput[823] , \matrixInput[822] , \matrixInput[821] , 
        \matrixInput[820] , \matrixInput[819] , \matrixInput[818] , 
        \matrixInput[817] , \matrixInput[816] , \matrixInput[815] , 
        \matrixInput[814] , \matrixInput[813] , \matrixInput[812] , 
        \matrixInput[811] , \matrixInput[810] , \matrixInput[809] , 
        \matrixInput[808] , \matrixInput[807] , \matrixInput[806] , 
        \matrixInput[805] , \matrixInput[804] , \matrixInput[803] , 
        \matrixInput[802] , \matrixInput[801] , \matrixInput[800] , 
        \matrixInput[799] , \matrixInput[798] , \matrixInput[797] , 
        \matrixInput[796] , \matrixInput[795] , \matrixInput[794] , 
        \matrixInput[793] , \matrixInput[792] , \matrixInput[791] , 
        \matrixInput[790] , \matrixInput[789] , \matrixInput[788] , 
        \matrixInput[787] , \matrixInput[786] , \matrixInput[785] , 
        \matrixInput[784] , \matrixInput[783] , \matrixInput[782] , 
        \matrixInput[781] , \matrixInput[780] , \matrixInput[779] , 
        \matrixInput[778] , \matrixInput[777] , \matrixInput[776] , 
        \matrixInput[775] , \matrixInput[774] , \matrixInput[773] , 
        \matrixInput[772] , \matrixInput[771] , \matrixInput[770] , 
        \matrixInput[769] , \matrixInput[768] }), .cOutput({\cOutput[55] , 
        \cOutput[54] , \cOutput[53] , \cOutput[52] , \cOutput[51] , 
        \cOutput[50] , \cOutput[49] , \cOutput[48] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1151] , \matrixInput[1150] , \matrixInput[1149] , 
        \matrixInput[1148] , \matrixInput[1147] , \matrixInput[1146] , 
        \matrixInput[1145] , \matrixInput[1144] , \matrixInput[1143] , 
        \matrixInput[1142] , \matrixInput[1141] , \matrixInput[1140] , 
        \matrixInput[1139] , \matrixInput[1138] , \matrixInput[1137] , 
        \matrixInput[1136] , \matrixInput[1135] , \matrixInput[1134] , 
        \matrixInput[1133] , \matrixInput[1132] , \matrixInput[1131] , 
        \matrixInput[1130] , \matrixInput[1129] , \matrixInput[1128] , 
        \matrixInput[1127] , \matrixInput[1126] , \matrixInput[1125] , 
        \matrixInput[1124] , \matrixInput[1123] , \matrixInput[1122] , 
        \matrixInput[1121] , \matrixInput[1120] , \matrixInput[1119] , 
        \matrixInput[1118] , \matrixInput[1117] , \matrixInput[1116] , 
        \matrixInput[1115] , \matrixInput[1114] , \matrixInput[1113] , 
        \matrixInput[1112] , \matrixInput[1111] , \matrixInput[1110] , 
        \matrixInput[1109] , \matrixInput[1108] , \matrixInput[1107] , 
        \matrixInput[1106] , \matrixInput[1105] , \matrixInput[1104] , 
        \matrixInput[1103] , \matrixInput[1102] , \matrixInput[1101] , 
        \matrixInput[1100] , \matrixInput[1099] , \matrixInput[1098] , 
        \matrixInput[1097] , \matrixInput[1096] , \matrixInput[1095] , 
        \matrixInput[1094] , \matrixInput[1093] , \matrixInput[1092] , 
        \matrixInput[1091] , \matrixInput[1090] , \matrixInput[1089] , 
        \matrixInput[1088] , \matrixInput[1087] , \matrixInput[1086] , 
        \matrixInput[1085] , \matrixInput[1084] , \matrixInput[1083] , 
        \matrixInput[1082] , \matrixInput[1081] , \matrixInput[1080] , 
        \matrixInput[1079] , \matrixInput[1078] , \matrixInput[1077] , 
        \matrixInput[1076] , \matrixInput[1075] , \matrixInput[1074] , 
        \matrixInput[1073] , \matrixInput[1072] , \matrixInput[1071] , 
        \matrixInput[1070] , \matrixInput[1069] , \matrixInput[1068] , 
        \matrixInput[1067] , \matrixInput[1066] , \matrixInput[1065] , 
        \matrixInput[1064] , \matrixInput[1063] , \matrixInput[1062] , 
        \matrixInput[1061] , \matrixInput[1060] , \matrixInput[1059] , 
        \matrixInput[1058] , \matrixInput[1057] , \matrixInput[1056] , 
        \matrixInput[1055] , \matrixInput[1054] , \matrixInput[1053] , 
        \matrixInput[1052] , \matrixInput[1051] , \matrixInput[1050] , 
        \matrixInput[1049] , \matrixInput[1048] , \matrixInput[1047] , 
        \matrixInput[1046] , \matrixInput[1045] , \matrixInput[1044] , 
        \matrixInput[1043] , \matrixInput[1042] , \matrixInput[1041] , 
        \matrixInput[1040] , \matrixInput[1039] , \matrixInput[1038] , 
        \matrixInput[1037] , \matrixInput[1036] , \matrixInput[1035] , 
        \matrixInput[1034] , \matrixInput[1033] , \matrixInput[1032] , 
        \matrixInput[1031] , \matrixInput[1030] , \matrixInput[1029] , 
        \matrixInput[1028] , \matrixInput[1027] , \matrixInput[1026] , 
        \matrixInput[1025] , \matrixInput[1024] }), .cOutput({\cOutput[71] , 
        \cOutput[70] , \cOutput[69] , \cOutput[68] , \cOutput[67] , 
        \cOutput[66] , \cOutput[65] , \cOutput[64] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1407] , \matrixInput[1406] , \matrixInput[1405] , 
        \matrixInput[1404] , \matrixInput[1403] , \matrixInput[1402] , 
        \matrixInput[1401] , \matrixInput[1400] , \matrixInput[1399] , 
        \matrixInput[1398] , \matrixInput[1397] , \matrixInput[1396] , 
        \matrixInput[1395] , \matrixInput[1394] , \matrixInput[1393] , 
        \matrixInput[1392] , \matrixInput[1391] , \matrixInput[1390] , 
        \matrixInput[1389] , \matrixInput[1388] , \matrixInput[1387] , 
        \matrixInput[1386] , \matrixInput[1385] , \matrixInput[1384] , 
        \matrixInput[1383] , \matrixInput[1382] , \matrixInput[1381] , 
        \matrixInput[1380] , \matrixInput[1379] , \matrixInput[1378] , 
        \matrixInput[1377] , \matrixInput[1376] , \matrixInput[1375] , 
        \matrixInput[1374] , \matrixInput[1373] , \matrixInput[1372] , 
        \matrixInput[1371] , \matrixInput[1370] , \matrixInput[1369] , 
        \matrixInput[1368] , \matrixInput[1367] , \matrixInput[1366] , 
        \matrixInput[1365] , \matrixInput[1364] , \matrixInput[1363] , 
        \matrixInput[1362] , \matrixInput[1361] , \matrixInput[1360] , 
        \matrixInput[1359] , \matrixInput[1358] , \matrixInput[1357] , 
        \matrixInput[1356] , \matrixInput[1355] , \matrixInput[1354] , 
        \matrixInput[1353] , \matrixInput[1352] , \matrixInput[1351] , 
        \matrixInput[1350] , \matrixInput[1349] , \matrixInput[1348] , 
        \matrixInput[1347] , \matrixInput[1346] , \matrixInput[1345] , 
        \matrixInput[1344] , \matrixInput[1343] , \matrixInput[1342] , 
        \matrixInput[1341] , \matrixInput[1340] , \matrixInput[1339] , 
        \matrixInput[1338] , \matrixInput[1337] , \matrixInput[1336] , 
        \matrixInput[1335] , \matrixInput[1334] , \matrixInput[1333] , 
        \matrixInput[1332] , \matrixInput[1331] , \matrixInput[1330] , 
        \matrixInput[1329] , \matrixInput[1328] , \matrixInput[1327] , 
        \matrixInput[1326] , \matrixInput[1325] , \matrixInput[1324] , 
        \matrixInput[1323] , \matrixInput[1322] , \matrixInput[1321] , 
        \matrixInput[1320] , \matrixInput[1319] , \matrixInput[1318] , 
        \matrixInput[1317] , \matrixInput[1316] , \matrixInput[1315] , 
        \matrixInput[1314] , \matrixInput[1313] , \matrixInput[1312] , 
        \matrixInput[1311] , \matrixInput[1310] , \matrixInput[1309] , 
        \matrixInput[1308] , \matrixInput[1307] , \matrixInput[1306] , 
        \matrixInput[1305] , \matrixInput[1304] , \matrixInput[1303] , 
        \matrixInput[1302] , \matrixInput[1301] , \matrixInput[1300] , 
        \matrixInput[1299] , \matrixInput[1298] , \matrixInput[1297] , 
        \matrixInput[1296] , \matrixInput[1295] , \matrixInput[1294] , 
        \matrixInput[1293] , \matrixInput[1292] , \matrixInput[1291] , 
        \matrixInput[1290] , \matrixInput[1289] , \matrixInput[1288] , 
        \matrixInput[1287] , \matrixInput[1286] , \matrixInput[1285] , 
        \matrixInput[1284] , \matrixInput[1283] , \matrixInput[1282] , 
        \matrixInput[1281] , \matrixInput[1280] }), .cOutput({\cOutput[87] , 
        \cOutput[86] , \cOutput[85] , \cOutput[84] , \cOutput[83] , 
        \cOutput[82] , \cOutput[81] , \cOutput[80] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[127] , \matrixInput[126] , \matrixInput[125] , 
        \matrixInput[124] , \matrixInput[123] , \matrixInput[122] , 
        \matrixInput[121] , \matrixInput[120] , \matrixInput[119] , 
        \matrixInput[118] , \matrixInput[117] , \matrixInput[116] , 
        \matrixInput[115] , \matrixInput[114] , \matrixInput[113] , 
        \matrixInput[112] , \matrixInput[111] , \matrixInput[110] , 
        \matrixInput[109] , \matrixInput[108] , \matrixInput[107] , 
        \matrixInput[106] , \matrixInput[105] , \matrixInput[104] , 
        \matrixInput[103] , \matrixInput[102] , \matrixInput[101] , 
        \matrixInput[100] , \matrixInput[99] , \matrixInput[98] , 
        \matrixInput[97] , \matrixInput[96] , \matrixInput[95] , 
        \matrixInput[94] , \matrixInput[93] , \matrixInput[92] , 
        \matrixInput[91] , \matrixInput[90] , \matrixInput[89] , 
        \matrixInput[88] , \matrixInput[87] , \matrixInput[86] , 
        \matrixInput[85] , \matrixInput[84] , \matrixInput[83] , 
        \matrixInput[82] , \matrixInput[81] , \matrixInput[80] , 
        \matrixInput[79] , \matrixInput[78] , \matrixInput[77] , 
        \matrixInput[76] , \matrixInput[75] , \matrixInput[74] , 
        \matrixInput[73] , \matrixInput[72] , \matrixInput[71] , 
        \matrixInput[70] , \matrixInput[69] , \matrixInput[68] , 
        \matrixInput[67] , \matrixInput[66] , \matrixInput[65] , 
        \matrixInput[64] , \matrixInput[63] , \matrixInput[62] , 
        \matrixInput[61] , \matrixInput[60] , \matrixInput[59] , 
        \matrixInput[58] , \matrixInput[57] , \matrixInput[56] , 
        \matrixInput[55] , \matrixInput[54] , \matrixInput[53] , 
        \matrixInput[52] , \matrixInput[51] , \matrixInput[50] , 
        \matrixInput[49] , \matrixInput[48] , \matrixInput[47] , 
        \matrixInput[46] , \matrixInput[45] , \matrixInput[44] , 
        \matrixInput[43] , \matrixInput[42] , \matrixInput[41] , 
        \matrixInput[40] , \matrixInput[39] , \matrixInput[38] , 
        \matrixInput[37] , \matrixInput[36] , \matrixInput[35] , 
        \matrixInput[34] , \matrixInput[33] , \matrixInput[32] , 
        \matrixInput[31] , \matrixInput[30] , \matrixInput[29] , 
        \matrixInput[28] , \matrixInput[27] , \matrixInput[26] , 
        \matrixInput[25] , \matrixInput[24] , \matrixInput[23] , 
        \matrixInput[22] , \matrixInput[21] , \matrixInput[20] , 
        \matrixInput[19] , \matrixInput[18] , \matrixInput[17] , 
        \matrixInput[16] , \matrixInput[15] , \matrixInput[14] , 
        \matrixInput[13] , \matrixInput[12] , \matrixInput[11] , 
        \matrixInput[10] , \matrixInput[9] , \matrixInput[8] , 
        \matrixInput[7] , \matrixInput[6] , \matrixInput[5] , \matrixInput[4] , 
        \matrixInput[3] , \matrixInput[2] , \matrixInput[1] , \matrixInput[0] 
        }), .cOutput({\cOutput[7] , \cOutput[6] , \cOutput[5] , \cOutput[4] , 
        \cOutput[3] , \cOutput[2] , \cOutput[1] , \cOutput[0] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1023] , \matrixInput[1022] , \matrixInput[1021] , 
        \matrixInput[1020] , \matrixInput[1019] , \matrixInput[1018] , 
        \matrixInput[1017] , \matrixInput[1016] , \matrixInput[1015] , 
        \matrixInput[1014] , \matrixInput[1013] , \matrixInput[1012] , 
        \matrixInput[1011] , \matrixInput[1010] , \matrixInput[1009] , 
        \matrixInput[1008] , \matrixInput[1007] , \matrixInput[1006] , 
        \matrixInput[1005] , \matrixInput[1004] , \matrixInput[1003] , 
        \matrixInput[1002] , \matrixInput[1001] , \matrixInput[1000] , 
        \matrixInput[999] , \matrixInput[998] , \matrixInput[997] , 
        \matrixInput[996] , \matrixInput[995] , \matrixInput[994] , 
        \matrixInput[993] , \matrixInput[992] , \matrixInput[991] , 
        \matrixInput[990] , \matrixInput[989] , \matrixInput[988] , 
        \matrixInput[987] , \matrixInput[986] , \matrixInput[985] , 
        \matrixInput[984] , \matrixInput[983] , \matrixInput[982] , 
        \matrixInput[981] , \matrixInput[980] , \matrixInput[979] , 
        \matrixInput[978] , \matrixInput[977] , \matrixInput[976] , 
        \matrixInput[975] , \matrixInput[974] , \matrixInput[973] , 
        \matrixInput[972] , \matrixInput[971] , \matrixInput[970] , 
        \matrixInput[969] , \matrixInput[968] , \matrixInput[967] , 
        \matrixInput[966] , \matrixInput[965] , \matrixInput[964] , 
        \matrixInput[963] , \matrixInput[962] , \matrixInput[961] , 
        \matrixInput[960] , \matrixInput[959] , \matrixInput[958] , 
        \matrixInput[957] , \matrixInput[956] , \matrixInput[955] , 
        \matrixInput[954] , \matrixInput[953] , \matrixInput[952] , 
        \matrixInput[951] , \matrixInput[950] , \matrixInput[949] , 
        \matrixInput[948] , \matrixInput[947] , \matrixInput[946] , 
        \matrixInput[945] , \matrixInput[944] , \matrixInput[943] , 
        \matrixInput[942] , \matrixInput[941] , \matrixInput[940] , 
        \matrixInput[939] , \matrixInput[938] , \matrixInput[937] , 
        \matrixInput[936] , \matrixInput[935] , \matrixInput[934] , 
        \matrixInput[933] , \matrixInput[932] , \matrixInput[931] , 
        \matrixInput[930] , \matrixInput[929] , \matrixInput[928] , 
        \matrixInput[927] , \matrixInput[926] , \matrixInput[925] , 
        \matrixInput[924] , \matrixInput[923] , \matrixInput[922] , 
        \matrixInput[921] , \matrixInput[920] , \matrixInput[919] , 
        \matrixInput[918] , \matrixInput[917] , \matrixInput[916] , 
        \matrixInput[915] , \matrixInput[914] , \matrixInput[913] , 
        \matrixInput[912] , \matrixInput[911] , \matrixInput[910] , 
        \matrixInput[909] , \matrixInput[908] , \matrixInput[907] , 
        \matrixInput[906] , \matrixInput[905] , \matrixInput[904] , 
        \matrixInput[903] , \matrixInput[902] , \matrixInput[901] , 
        \matrixInput[900] , \matrixInput[899] , \matrixInput[898] , 
        \matrixInput[897] , \matrixInput[896] }), .cOutput({\cOutput[63] , 
        \cOutput[62] , \cOutput[61] , \cOutput[60] , \cOutput[59] , 
        \cOutput[58] , \cOutput[57] , \cOutput[56] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1535] , \matrixInput[1534] , \matrixInput[1533] , 
        \matrixInput[1532] , \matrixInput[1531] , \matrixInput[1530] , 
        \matrixInput[1529] , \matrixInput[1528] , \matrixInput[1527] , 
        \matrixInput[1526] , \matrixInput[1525] , \matrixInput[1524] , 
        \matrixInput[1523] , \matrixInput[1522] , \matrixInput[1521] , 
        \matrixInput[1520] , \matrixInput[1519] , \matrixInput[1518] , 
        \matrixInput[1517] , \matrixInput[1516] , \matrixInput[1515] , 
        \matrixInput[1514] , \matrixInput[1513] , \matrixInput[1512] , 
        \matrixInput[1511] , \matrixInput[1510] , \matrixInput[1509] , 
        \matrixInput[1508] , \matrixInput[1507] , \matrixInput[1506] , 
        \matrixInput[1505] , \matrixInput[1504] , \matrixInput[1503] , 
        \matrixInput[1502] , \matrixInput[1501] , \matrixInput[1500] , 
        \matrixInput[1499] , \matrixInput[1498] , \matrixInput[1497] , 
        \matrixInput[1496] , \matrixInput[1495] , \matrixInput[1494] , 
        \matrixInput[1493] , \matrixInput[1492] , \matrixInput[1491] , 
        \matrixInput[1490] , \matrixInput[1489] , \matrixInput[1488] , 
        \matrixInput[1487] , \matrixInput[1486] , \matrixInput[1485] , 
        \matrixInput[1484] , \matrixInput[1483] , \matrixInput[1482] , 
        \matrixInput[1481] , \matrixInput[1480] , \matrixInput[1479] , 
        \matrixInput[1478] , \matrixInput[1477] , \matrixInput[1476] , 
        \matrixInput[1475] , \matrixInput[1474] , \matrixInput[1473] , 
        \matrixInput[1472] , \matrixInput[1471] , \matrixInput[1470] , 
        \matrixInput[1469] , \matrixInput[1468] , \matrixInput[1467] , 
        \matrixInput[1466] , \matrixInput[1465] , \matrixInput[1464] , 
        \matrixInput[1463] , \matrixInput[1462] , \matrixInput[1461] , 
        \matrixInput[1460] , \matrixInput[1459] , \matrixInput[1458] , 
        \matrixInput[1457] , \matrixInput[1456] , \matrixInput[1455] , 
        \matrixInput[1454] , \matrixInput[1453] , \matrixInput[1452] , 
        \matrixInput[1451] , \matrixInput[1450] , \matrixInput[1449] , 
        \matrixInput[1448] , \matrixInput[1447] , \matrixInput[1446] , 
        \matrixInput[1445] , \matrixInput[1444] , \matrixInput[1443] , 
        \matrixInput[1442] , \matrixInput[1441] , \matrixInput[1440] , 
        \matrixInput[1439] , \matrixInput[1438] , \matrixInput[1437] , 
        \matrixInput[1436] , \matrixInput[1435] , \matrixInput[1434] , 
        \matrixInput[1433] , \matrixInput[1432] , \matrixInput[1431] , 
        \matrixInput[1430] , \matrixInput[1429] , \matrixInput[1428] , 
        \matrixInput[1427] , \matrixInput[1426] , \matrixInput[1425] , 
        \matrixInput[1424] , \matrixInput[1423] , \matrixInput[1422] , 
        \matrixInput[1421] , \matrixInput[1420] , \matrixInput[1419] , 
        \matrixInput[1418] , \matrixInput[1417] , \matrixInput[1416] , 
        \matrixInput[1415] , \matrixInput[1414] , \matrixInput[1413] , 
        \matrixInput[1412] , \matrixInput[1411] , \matrixInput[1410] , 
        \matrixInput[1409] , \matrixInput[1408] }), .cOutput({\cOutput[95] , 
        \cOutput[94] , \cOutput[93] , \cOutput[92] , \cOutput[91] , 
        \cOutput[90] , \cOutput[89] , \cOutput[88] }) );
    VectorDotProduct_pVectorSize16_pWordSize8 VectorDotProduct_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .vectorAInput({\vectorInput[127] , 
        \vectorInput[126] , \vectorInput[125] , \vectorInput[124] , 
        \vectorInput[123] , \vectorInput[122] , \vectorInput[121] , 
        \vectorInput[120] , \vectorInput[119] , \vectorInput[118] , 
        \vectorInput[117] , \vectorInput[116] , \vectorInput[115] , 
        \vectorInput[114] , \vectorInput[113] , \vectorInput[112] , 
        \vectorInput[111] , \vectorInput[110] , \vectorInput[109] , 
        \vectorInput[108] , \vectorInput[107] , \vectorInput[106] , 
        \vectorInput[105] , \vectorInput[104] , \vectorInput[103] , 
        \vectorInput[102] , \vectorInput[101] , \vectorInput[100] , 
        \vectorInput[99] , \vectorInput[98] , \vectorInput[97] , 
        \vectorInput[96] , \vectorInput[95] , \vectorInput[94] , 
        \vectorInput[93] , \vectorInput[92] , \vectorInput[91] , 
        \vectorInput[90] , \vectorInput[89] , \vectorInput[88] , 
        \vectorInput[87] , \vectorInput[86] , \vectorInput[85] , 
        \vectorInput[84] , \vectorInput[83] , \vectorInput[82] , 
        \vectorInput[81] , \vectorInput[80] , \vectorInput[79] , 
        \vectorInput[78] , \vectorInput[77] , \vectorInput[76] , 
        \vectorInput[75] , \vectorInput[74] , \vectorInput[73] , 
        \vectorInput[72] , \vectorInput[71] , \vectorInput[70] , 
        \vectorInput[69] , \vectorInput[68] , \vectorInput[67] , 
        \vectorInput[66] , \vectorInput[65] , \vectorInput[64] , 
        \vectorInput[63] , \vectorInput[62] , \vectorInput[61] , 
        \vectorInput[60] , \vectorInput[59] , \vectorInput[58] , 
        \vectorInput[57] , \vectorInput[56] , \vectorInput[55] , 
        \vectorInput[54] , \vectorInput[53] , \vectorInput[52] , 
        \vectorInput[51] , \vectorInput[50] , \vectorInput[49] , 
        \vectorInput[48] , \vectorInput[47] , \vectorInput[46] , 
        \vectorInput[45] , \vectorInput[44] , \vectorInput[43] , 
        \vectorInput[42] , \vectorInput[41] , \vectorInput[40] , 
        \vectorInput[39] , \vectorInput[38] , \vectorInput[37] , 
        \vectorInput[36] , \vectorInput[35] , \vectorInput[34] , 
        \vectorInput[33] , \vectorInput[32] , \vectorInput[31] , 
        \vectorInput[30] , \vectorInput[29] , \vectorInput[28] , 
        \vectorInput[27] , \vectorInput[26] , \vectorInput[25] , 
        \vectorInput[24] , \vectorInput[23] , \vectorInput[22] , 
        \vectorInput[21] , \vectorInput[20] , \vectorInput[19] , 
        \vectorInput[18] , \vectorInput[17] , \vectorInput[16] , 
        \vectorInput[15] , \vectorInput[14] , \vectorInput[13] , 
        \vectorInput[12] , \vectorInput[11] , \vectorInput[10] , 
        \vectorInput[9] , \vectorInput[8] , \vectorInput[7] , \vectorInput[6] , 
        \vectorInput[5] , \vectorInput[4] , \vectorInput[3] , \vectorInput[2] , 
        \vectorInput[1] , \vectorInput[0] }), .vectorBInput({
        \matrixInput[1279] , \matrixInput[1278] , \matrixInput[1277] , 
        \matrixInput[1276] , \matrixInput[1275] , \matrixInput[1274] , 
        \matrixInput[1273] , \matrixInput[1272] , \matrixInput[1271] , 
        \matrixInput[1270] , \matrixInput[1269] , \matrixInput[1268] , 
        \matrixInput[1267] , \matrixInput[1266] , \matrixInput[1265] , 
        \matrixInput[1264] , \matrixInput[1263] , \matrixInput[1262] , 
        \matrixInput[1261] , \matrixInput[1260] , \matrixInput[1259] , 
        \matrixInput[1258] , \matrixInput[1257] , \matrixInput[1256] , 
        \matrixInput[1255] , \matrixInput[1254] , \matrixInput[1253] , 
        \matrixInput[1252] , \matrixInput[1251] , \matrixInput[1250] , 
        \matrixInput[1249] , \matrixInput[1248] , \matrixInput[1247] , 
        \matrixInput[1246] , \matrixInput[1245] , \matrixInput[1244] , 
        \matrixInput[1243] , \matrixInput[1242] , \matrixInput[1241] , 
        \matrixInput[1240] , \matrixInput[1239] , \matrixInput[1238] , 
        \matrixInput[1237] , \matrixInput[1236] , \matrixInput[1235] , 
        \matrixInput[1234] , \matrixInput[1233] , \matrixInput[1232] , 
        \matrixInput[1231] , \matrixInput[1230] , \matrixInput[1229] , 
        \matrixInput[1228] , \matrixInput[1227] , \matrixInput[1226] , 
        \matrixInput[1225] , \matrixInput[1224] , \matrixInput[1223] , 
        \matrixInput[1222] , \matrixInput[1221] , \matrixInput[1220] , 
        \matrixInput[1219] , \matrixInput[1218] , \matrixInput[1217] , 
        \matrixInput[1216] , \matrixInput[1215] , \matrixInput[1214] , 
        \matrixInput[1213] , \matrixInput[1212] , \matrixInput[1211] , 
        \matrixInput[1210] , \matrixInput[1209] , \matrixInput[1208] , 
        \matrixInput[1207] , \matrixInput[1206] , \matrixInput[1205] , 
        \matrixInput[1204] , \matrixInput[1203] , \matrixInput[1202] , 
        \matrixInput[1201] , \matrixInput[1200] , \matrixInput[1199] , 
        \matrixInput[1198] , \matrixInput[1197] , \matrixInput[1196] , 
        \matrixInput[1195] , \matrixInput[1194] , \matrixInput[1193] , 
        \matrixInput[1192] , \matrixInput[1191] , \matrixInput[1190] , 
        \matrixInput[1189] , \matrixInput[1188] , \matrixInput[1187] , 
        \matrixInput[1186] , \matrixInput[1185] , \matrixInput[1184] , 
        \matrixInput[1183] , \matrixInput[1182] , \matrixInput[1181] , 
        \matrixInput[1180] , \matrixInput[1179] , \matrixInput[1178] , 
        \matrixInput[1177] , \matrixInput[1176] , \matrixInput[1175] , 
        \matrixInput[1174] , \matrixInput[1173] , \matrixInput[1172] , 
        \matrixInput[1171] , \matrixInput[1170] , \matrixInput[1169] , 
        \matrixInput[1168] , \matrixInput[1167] , \matrixInput[1166] , 
        \matrixInput[1165] , \matrixInput[1164] , \matrixInput[1163] , 
        \matrixInput[1162] , \matrixInput[1161] , \matrixInput[1160] , 
        \matrixInput[1159] , \matrixInput[1158] , \matrixInput[1157] , 
        \matrixInput[1156] , \matrixInput[1155] , \matrixInput[1154] , 
        \matrixInput[1153] , \matrixInput[1152] }), .cOutput({\cOutput[79] , 
        \cOutput[78] , \cOutput[77] , \cOutput[76] , \cOutput[75] , 
        \cOutput[74] , \cOutput[73] , \cOutput[72] }) );
endmodule

