
module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n185, n182, \ScanOut[1]1 , 
        n184, \ScanOut[0]1 , n183, \ScanOut[6]1 , \ScanOut[3]1 , n176, 
        \ScanOut[2]1 , n181, n186, n178, n179, n177, n180;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO22 U28 ( .A(ScanIn[1]), .B(n176), .C(\ScanOut[1]1 ), .D(n177), .Z(
        n185) );
    VMW_AO22 U33 ( .A(ScanIn[6]), .B(n176), .C(\ScanOut[6]1 ), .D(n177), .Z(
        n180) );
    VMW_AO22 U34 ( .A(ScanIn[7]), .B(n176), .C(\ScanOut[7] ), .D(n177), .Z(
        n179) );
    VMW_NOR2 U35 ( .A(ScanEnable), .B(Reset), .Z(n177) );
    VMW_AO22 U27 ( .A(ScanIn[0]), .B(n176), .C(\ScanOut[0]1 ), .D(n177), .Z(
        n186) );
    VMW_FD \Out_reg[5]  ( .D(n181), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U29 ( .A(ScanIn[2]), .B(n176), .C(\ScanOut[2]1 ), .D(n177), .Z(
        n184) );
    VMW_FD \Out_reg[7]  ( .D(n179), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n183), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n185), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO22 U32 ( .A(ScanIn[5]), .B(n176), .C(\ScanOut[5]1 ), .D(n177), .Z(
        n181) );
    VMW_AO22 U30 ( .A(ScanIn[3]), .B(n176), .C(\ScanOut[3]1 ), .D(n177), .Z(
        n183) );
    VMW_FD \Out_reg[6]  ( .D(n180), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U31 ( .A(ScanIn[4]), .B(n176), .C(\ScanOut[4]1 ), .D(n177), .Z(
        n182) );
    VMW_NOR2 U36 ( .A(n178), .B(Reset), .Z(n176) );
    VMW_INV U37 ( .A(ScanEnable), .Z(n178) );
    VMW_FD \Out_reg[2]  ( .D(n184), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n182), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n186), .CP(Clk), .Q(\ScanOut[0]1 ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n1, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_AND2 U1 ( .A(A[0]), .B(B[0]), .Z(\carry[1] ) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .CO(\carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .CO(\carry[7] ), .S(
        SUM[6]) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .CO(\carry[3] ), .S(
        SUM[2]) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .CO(\carry[4] ), .S(
        SUM[3]) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .CO(\carry[5] ), .S(
        SUM[4]) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .CO(\carry[6] ), .S(
        SUM[5]) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n3, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n3) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n222, n217, n225, n219, 
        n210, \ScanOut[6]1 , n224, \a184[4] , \n161[4] , \ScanOut[1]1 , n218, 
        \n158[4] , \ScanOut[0]1 , n211, n216, \n158[2] , n223, \n161[2] , 
        \n158[6] , \a184[6] , \n161[6] , \ScanOut[3]1 , \n158[7] , n214, 
        \n161[7] , \a184[7] , n206, n221, \n158[3] , \ScanOut[2]1 , \a184[3] , 
        \n161[3] , \n161[1] , \n158[8] , n226, \a184[8] , \n161[8] , \n158[1] , 
        n213, \a184[5] , n208, \n161[5] , \n158[5] , n209, n212, n215, n207, 
        n220;
    wire UNCONNECTED_1 , UNCONNECTED_2 ;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U33 ( .A(\ScanOut[0]1 ), .B(n206), .C(n207), .Z(n223) );
    VMW_AO21 U34 ( .A(\ScanOut[1]1 ), .B(n206), .C(n208), .Z(n222) );
    VMW_NOR2 U41 ( .A(n214), .B(Reset), .Z(n213) );
    VMW_AO22 U46 ( .A(ScanIn[3]), .B(n213), .C(\a184[6] ), .D(n215), .Z(n210)
         );
    VMW_AO21 U35 ( .A(\ScanOut[2]1 ), .B(n206), .C(n209), .Z(n221) );
    VMW_AO22 U48 ( .A(ScanIn[1]), .B(n213), .C(\a184[4] ), .D(n215), .Z(n208)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 add_98 ( .A({
        \n158[1] , \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , 
        \n158[7] , \n158[8] }), .B(WestIn), .CI(n225), .SUM({\a184[8] , 
        \a184[7] , \a184[6] , \a184[5] , \a184[4] , \a184[3] , UNCONNECTED_1, 
        UNCONNECTED_2}) );
    VMW_PULLDOWN U32 ( .Z(n224) );
    VMW_AO22 U40 ( .A(\ScanOut[7] ), .B(n206), .C(ScanIn[7]), .D(n213), .Z(
        n216) );
    VMW_FD \Out_reg[5]  ( .D(n218), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U47 ( .A(ScanIn[2]), .B(n213), .C(\a184[5] ), .D(n215), .Z(n209)
         );
    VMW_AO22 U49 ( .A(ScanIn[0]), .B(n213), .C(\a184[3] ), .D(n215), .Z(n207)
         );
    VMW_FD \Out_reg[1]  ( .D(n222), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_FD \Out_reg[7]  ( .D(n216), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n220), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_PULLDOWN U30 ( .Z(n225) );
    VMW_AO22 U39 ( .A(\ScanOut[6]1 ), .B(n206), .C(ScanIn[6]), .D(n213), .Z(
        n217) );
    VMW_FD \Out_reg[6]  ( .D(n217), .CP(Clk), .Q(\ScanOut[6]1 ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 add_98_2 ( .A(
        NorthIn), .B(SouthIn), .CI(n224), .SUM({\n161[1] , \n161[2] , 
        \n161[3] , \n161[4] , \n161[5] , \n161[6] , \n161[7] , \n161[8] }) );
    VMW_PULLDOWN U31 ( .Z(n226) );
    VMW_AO21 U36 ( .A(\ScanOut[3]1 ), .B(n206), .C(n210), .Z(n220) );
    VMW_AO21 U37 ( .A(\ScanOut[4]1 ), .B(n206), .C(n211), .Z(n219) );
    VMW_NOR3 U42 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n206) );
    VMW_AO22 U45 ( .A(ScanIn[4]), .B(n213), .C(\a184[7] ), .D(n215), .Z(n211)
         );
    VMW_FD \Out_reg[2]  ( .D(n221), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_INV U50 ( .A(ScanEnable), .Z(n214) );
    VMW_FD \Out_reg[4]  ( .D(n219), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n223), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_AO21 U38 ( .A(\ScanOut[5]1 ), .B(n206), .C(n212), .Z(n218) );
    VMW_NOR3 U43 ( .A(Reset), .B(ScanEnable), .C(n206), .Z(n215) );
    VMW_AO22 U44 ( .A(ScanIn[5]), .B(n213), .C(\a184[8] ), .D(n215), .Z(n212)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 add_98_1 ( .A({
        \n161[1] , \n161[2] , \n161[3] , \n161[4] , \n161[5] , \n161[6] , 
        \n161[7] , \n161[8] }), .B(EastIn), .CI(n226), .SUM({\n158[1] , 
        \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , \n158[7] , 
        \n158[8] }) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 ( A, SUM );
input  [6:0] A;
output [6:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[2]), .C(n6), .Z(SUM[2]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n9), .Z(SUM[1]) );
    VMW_INV U6 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO22 U14 ( .A(A[5]), .B(n13), .C(n12), .D(n10), .Z(SUM[5]) );
    VMW_AO21 U7 ( .A(n8), .B(A[4]), .C(n10), .Z(SUM[4]) );
    VMW_AND2 U8 ( .A(n10), .B(n12), .Z(n11) );
    VMW_XOR2 U13 ( .A(A[6]), .B(n11), .Z(SUM[6]) );
    VMW_OR2 U9 ( .A(A[0]), .B(A[1]), .Z(n5) );
    VMW_NOR2 U12 ( .A(n8), .B(A[4]), .Z(n10) );
    VMW_INV U15 ( .A(A[5]), .Z(n12) );
    VMW_INV U17 ( .A(A[3]), .Z(n7) );
    VMW_NOR2 U10 ( .A(n5), .B(A[2]), .Z(n6) );
    VMW_NAND2 U11 ( .A(n6), .B(n7), .Z(n8) );
    VMW_OAI21 U4 ( .A(n6), .B(n7), .C(n8), .Z(SUM[3]) );
    VMW_INV U18 ( .A(n5), .Z(n9) );
    VMW_INV U16 ( .A(n10), .Z(n13) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] ScanIn;
output [7:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n379, \count[2] , n387, n362, n406, n395, \count[6] , n370, n389, 
        n408, n377, n392, \count[4] , n380, n401, n365, \count[0] , n393, n376, 
        \ScanReg[2] , n409, \count260[3] , n388, n364, n400, n381, 
        \ScanReg[6] , n386, n407, \ScanReg[4] , n363, \count260[5] , n378, 
        \count260[1] , \ScanReg[0] , n371, n394, \count260[0] , \ScanReg[1] , 
        \ScanReg[7] , n405, n384, \ScanReg[5] , \count260[4] , n396, n373, 
        n368, n374, \count260[6] , n383, n391, n410, n402, n366, n390, n398, 
        \count260[2] , \ScanReg[3] , n411, n375, \count[1] , n399, n367, n382, 
        n403, n385, \count[5] , n404, n369, \count[3] , n372, n397;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_PULLDOWN U54 ( .Z(n372) );
    VMW_PULLDOWN U73 ( .Z(n399) );
    VMW_INV U113 ( .A(n370), .Z(ScanEnable) );
    VMW_BUFIZ U134 ( .A(n393), .E(n377), .Z(\arr[3] ) );
    VMW_PULLDOWN U68 ( .Z(n391) );
    VMW_AND2 U96 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AO22 U108 ( .A(\count[0] ), .B(n366), .C(\ScanReg[0] ), .D(n365), .Z(
        n373) );
    VMW_BUFIZ U141 ( .A(n400), .E(n377), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n405), .CP(Clk), .Q(\count[6] ) );
    VMW_PULLDOWN U61 ( .Z(n382) );
    VMW_AO22 U84 ( .A(ScanOut[4]), .B(n363), .C(\count260[4] ), .D(n364), .Z(
        n407) );
    VMW_FD \count_reg[2]  ( .D(n409), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U66 ( .Z(n389) );
    VMW_XNOR2 U101 ( .A(Addr[0]), .B(ScanId), .Z(n371) );
    VMW_AO22 U106 ( .A(\count[2] ), .B(n366), .C(\ScanReg[2] ), .D(n365), .Z(
        n388) );
    VMW_BUFIZ U121 ( .A(n380), .E(n377), .Z(\arr[14] ) );
    VMW_BUFIZ U126 ( .A(n385), .E(n377), .Z(\arr[31] ) );
    VMW_PULLDOWN U74 ( .Z(n400) );
    VMW_AO22 U83 ( .A(ScanOut[3]), .B(n363), .C(\count260[3] ), .D(n364), .Z(
        n408) );
    VMW_FD \count_reg[0]  ( .D(n411), .CP(Clk), .Q(\count[0] ) );
    VMW_NOR2 U91 ( .A(n367), .B(n368), .Z(n364) );
    VMW_AND2 U98 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_BUFIZ U128 ( .A(n387), .E(n377), .Z(\arr[28] ) );
    VMW_FD \count_reg[4]  ( .D(n407), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U114 ( .A(n372), .E(n377), .Z(\arr[19] ) );
    VMW_BUFIZ U133 ( .A(n392), .E(n377), .Z(\arr[20] ) );
    VMW_AND2 U99 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_PULLDOWN U55 ( .Z(n374) );
    VMW_PULLDOWN U67 ( .Z(n390) );
    VMW_AO22 U82 ( .A(ScanOut[2]), .B(n363), .C(\count260[2] ), .D(n364), .Z(
        n409) );
    VMW_AO22 U107 ( .A(\count[1] ), .B(n366), .C(\ScanReg[1] ), .D(n365), .Z(
        n403) );
    VMW_BUFIZ U120 ( .A(n379), .E(n377), .Z(\arr[27] ) );
    VMW_PULLDOWN U69 ( .Z(n392) );
    VMW_PULLDOWN U75 ( .Z(n401) );
    VMW_BUFIZ U115 ( .A(n373), .E(n377), .Z(\arr[0] ) );
    VMW_BUFIZ U132 ( .A(n391), .E(n377), .Z(\arr[29] ) );
    VMW_OAI21 U90 ( .A(n368), .B(Enable), .C(n369), .Z(n367) );
    VMW_OR4 U109 ( .A(\count[3] ), .B(\count[4] ), .C(\count[5] ), .D(
        \count[6] ), .Z(n362) );
    VMW_BUFIZ U129 ( .A(n388), .E(n377), .Z(\arr[2] ) );
    VMW_PULLDOWN U72 ( .Z(n398) );
    VMW_AND2 U97 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U140 ( .A(n399), .E(n377), .Z(\arr[15] ) );
    VMW_INV U112 ( .A(Reset), .Z(n369) );
    VMW_BUFIZ U135 ( .A(n394), .E(n377), .Z(\arr[24] ) );
    VMW_PULLDOWN U60 ( .Z(n381) );
    VMW_AO22 U85 ( .A(ScanOut[5]), .B(n363), .C(\count260[5] ), .D(n364), .Z(
        n406) );
    VMW_OAI21 U100 ( .A(WR), .B(RD), .C(n371), .Z(n370) );
    VMW_BUFIZ U127 ( .A(n386), .E(n377), .Z(\arr[21] ) );
    VMW_PULLDOWN U56 ( .Z(n375) );
    VMW_PULLDOWN U57 ( .Z(n376) );
    VMW_BUFIZ U137 ( .A(n396), .E(n377), .Z(\arr[7] ) );
    VMW_PULLDOWN U58 ( .Z(n379) );
    VMW_PULLDOWN U59 ( .Z(n380) );
    VMW_PULLDOWN U62 ( .Z(n383) );
    VMW_PULLDOWN U70 ( .Z(n394) );
    VMW_AND2 U79 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U95 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U110 ( .A(n366), .B(WR), .Z(n368) );
    VMW_BUFIZ U119 ( .A(n378), .E(n377), .Z(\arr[4] ) );
    VMW_BUFIZ U142 ( .A(n401), .E(n377), .Z(\arr[22] ) );
    VMW_AND2 U87 ( .A(\ScanReg[7] ), .B(n365), .Z(n396) );
    VMW_BUFIZ U125 ( .A(n384), .E(n377), .Z(\arr[6] ) );
    VMW_PULLDOWN U65 ( .Z(n387) );
    VMW_AO22 U102 ( .A(\count[6] ), .B(n366), .C(\ScanReg[6] ), .D(n365), .Z(
        n384) );
    VMW_AO22 U105 ( .A(\count[3] ), .B(n366), .C(\ScanReg[3] ), .D(n365), .Z(
        n393) );
    VMW_AO22 U80 ( .A(ScanOut[0]), .B(n363), .C(\count260[0] ), .D(n364), .Z(
        n411) );
    VMW_BUFIZ U122 ( .A(n381), .E(n377), .Z(\arr[25] ) );
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 sub_189 ( .A({
        \count[6] , \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[6] , \count260[5] , \count260[4] , 
        \count260[3] , \count260[2] , \count260[1] , \count260[0] }) );
    VMW_BUFIZ U139 ( .A(n398), .E(n377), .Z(\arr[26] ) );
    VMW_PULLDOWN U77 ( .Z(n404) );
    VMW_XOR2 U89 ( .A(Addr[0]), .B(Id), .Z(n365) );
    VMW_NOR2 U92 ( .A(n367), .B(n365), .Z(n363) );
    VMW_BUFIZ U145 ( .A(n404), .E(n377), .Z(\arr[8] ) );
    VMW_BUFIZ U117 ( .A(n375), .E(n377), .Z(\arr[10] ) );
    VMW_BUFIZ U130 ( .A(n389), .E(n377), .Z(\arr[13] ) );
    VMW_BUFIZ U138 ( .A(n397), .E(n377), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n406), .CP(Clk), .Q(\count[5] ) );
    VMW_PULLDOWN U64 ( .Z(n386) );
    VMW_AO22 U81 ( .A(ScanOut[1]), .B(n363), .C(\count260[1] ), .D(n364), .Z(
        n410) );
    VMW_AO22 U104 ( .A(\count[4] ), .B(n366), .C(\ScanReg[4] ), .D(n365), .Z(
        n378) );
    VMW_PULLDOWN U76 ( .Z(n402) );
    VMW_BUFIZ U116 ( .A(n374), .E(n377), .Z(\arr[23] ) );
    VMW_BUFIZ U123 ( .A(n382), .E(n377), .Z(\arr[16] ) );
    VMW_AO21 U88 ( .A(RD), .B(ScanEnable), .C(n366), .Z(n377) );
    VMW_AND2 U93 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_BUFIZ U131 ( .A(n390), .E(n377), .Z(\arr[30] ) );
    VMW_FD \count_reg[1]  ( .D(n410), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_BUFIZ U143 ( .A(n402), .E(n377), .Z(\arr[11] ) );
    VMW_BUFIZ U144 ( .A(n403), .E(n377), .Z(\arr[1] ) );
    VMW_FD \count_reg[3]  ( .D(n408), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n395), .E(n377), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_PULLDOWN U63 ( .Z(n385) );
    VMW_PULLDOWN U71 ( .Z(n395) );
    VMW_INV U111 ( .A(n365), .Z(n366) );
    VMW_BUFIZ U124 ( .A(n383), .E(n377), .Z(\arr[12] ) );
    VMW_OR4 U78 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n362), 
        .Z(Enable) );
    VMW_AO22 U86 ( .A(ScanOut[6]), .B(n363), .C(\count260[6] ), .D(n364), .Z(
        n405) );
    VMW_AO22 U103 ( .A(\count[5] ), .B(n366), .C(\ScanReg[5] ), .D(n365), .Z(
        n397) );
    VMW_BUFIZ U118 ( .A(n376), .E(n377), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nOut8_10[4] , \nOut2_15[3] , \nScanOut108[0] , \nOut8_13[7] , 
        \nOut0_1[1] , \nOut0_2[2] , \nScanOut4[1] , \nScanOut7[2] , 
        \nScanOut11[1] , \nScanOut12[2] , \nScanOut110[2] , \nOut11_10[4] , 
        \nScanOut113[1] , \nOut1_9[6] , \nOut12_9[3] , \nScanOut52[0] , 
        \nScanOut75[5] , \nOut6_10[0] , \nOut7_9[2] , \nOut11_13[7] , 
        \nScanOut174[6] , \nScanOut214[3] , \nOut14_9[7] , \nScanOut76[6] , 
        \nOut6_13[3] , \nScanOut177[5] , \nScanOut217[0] , \nScanOut181[5] , 
        \nScanOut153[3] , \nScanOut80[6] , \nScanOut150[0] , \nScanOut233[6] , 
        \nScanOut35[7] , \nScanOut36[4] , \nScanOut51[3] , \nScanOut83[5] , 
        \nScanOut230[5] , \nScanOut182[6] , \nOut7_15[0] , \nScanOut137[7] , 
        \nOut10_15[4] , \nOut3_5[0] , \nOut3_6[3] , \nScanOut134[4] , 
        \nOut9_7[6] , \nScanOut148[2] , \nScanOut254[1] , \nScanOut228[7] , 
        \nOut3_13[0] , \nOut10_6[6] , \nScanOut49[1] , \nOut5_6[7] , 
        \nOut10_5[5] , \nScanOut199[7] , \nOut3_10[3] , \nOut5_5[4] , 
        \nOut6_2[6] , \nScanOut98[4] , \nOut9_4[5] , \nOut13_2[7] , 
        \nOut14_13[4] , \nOut15_2[3] , \nOut6_1[5] , \nOut9_15[4] , 
        \nOut14_10[7] , \nOut15_1[0] , \nScanOut9[4] , \nOut1_11[4] , 
        \nOut1_12[7] , \nScanOut38[2] , \nOut13_1[4] , \nScanOut139[1] , 
        \nOut0_14[4] , \nOut2_3[1] , \nScanOut20[0] , \nScanOut23[3] , 
        \nScanOut122[0] , \nScanOut242[5] , \nOut2_0[2] , \nOut3_8[5] , 
        \nOut5_14[7] , \nScanOut121[3] , \nScanOut241[6] , \nScanOut194[2] , 
        \nScanOut44[4] , \nScanOut47[7] , \nOut5_8[1] , \nOut10_8[0] , 
        \nScanOut95[1] , \nOut9_9[0] , \nScanOut146[4] , \nScanOut226[1] , 
        \nScanOut96[2] , \nScanOut145[7] , \nOut12_14[3] , \nScanOut197[1] , 
        \nScanOut225[2] , \nOut4_11[7] , \nScanOut60[2] , \nScanOut161[1] , 
        \nScanOut201[4] , \nOut13_11[3] , \nScanOut63[1] , \nScanOut162[2] , 
        \nScanOut202[7] , \nOut13_12[0] , \nOut4_12[4] , \nScanOut105[5] , 
        \nOut4_0[6] , \nScanOut106[6] , \nOut11_0[7] , \nOut4_3[5] , 
        \nOut8_1[7] , \nOut8_2[4] , \nScanOut179[3] , \nScanOut219[6] , 
        \nScanOut78[0] , \nOut11_3[4] , \nOut1_4[3] , \nOut0_9[0] , 
        \nOut1_7[0] , \nOut7_4[7] , \nOut12_4[6] , \nOut14_4[2] , 
        \nOut12_7[5] , \nScanOut25[4] , \nOut1_14[0] , \nScanOut59[2] , 
        \nScanOut88[7] , \nOut7_7[4] , \nOut14_7[1] , \nScanOut189[4] , 
        \nScanOut158[1] , \nScanOut238[4] , \nScanOut41[0] , \nScanOut42[3] , 
        \nScanOut90[5] , \nScanOut93[6] , \nScanOut192[5] , \nScanOut140[3] , 
        \nScanOut220[6] , \nOut12_11[7] , \nScanOut223[5] , \nScanOut143[0] , 
        \nOut12_12[4] , \nOut5_11[3] , \nScanOut191[6] , \nScanOut244[2] , 
        \nScanOut124[7] , \nScanOut26[7] , \nOut13_9[5] , \nOut0_11[0] , 
        \nOut0_12[3] , \nOut4_14[3] , \nOut5_12[0] , \nOut6_9[4] , 
        \nOut15_9[1] , \nScanOut247[1] , \nScanOut100[1] , \nScanOut103[2] , 
        \nScanOut127[4] , \nScanOut65[6] , \nScanOut66[5] , \nScanOut167[6] , 
        \nScanOut207[3] , \nScanOut118[3] , \nScanOut164[5] , \nOut13_14[7] , 
        \nScanOut204[0] , \nOut1_1[7] , \nOut1_2[4] , \nScanOut19[0] , 
        \nOut7_2[0] , \nOut12_2[1] , \nOut14_2[5] , \nOut7_1[3] , 
        \nOut14_1[6] , \nOut12_1[2] , \nScanOut14[5] , \nScanOut17[6] , 
        \nOut2_5[6] , \nOut2_6[5] , \nOut4_6[1] , \nOut11_6[0] , \nOut8_4[3] , 
        \nOut8_7[0] , \nOut11_5[3] , \nOut2_8[3] , \nOut2_10[7] , 
        \nOut2_13[4] , \nOut4_5[2] , \nScanOut68[3] , \nScanOut169[0] , 
        \nScanOut209[5] , \nOut8_9[6] , \nOut8_15[0] , \nOut15_10[3] , 
        \nOut15_13[0] , \nScanOut172[1] , \nScanOut212[4] , \nOut4_8[7] , 
        \nOut11_8[6] , \nScanOut70[1] , \nScanOut73[2] , \nOut6_15[4] , 
        \nScanOut171[2] , \nScanOut211[7] , \nScanOut115[6] , \nScanOut116[5] , 
        \nOut11_15[0] , \nScanOut30[3] , \nScanOut131[0] , \nScanOut251[5] , 
        \nScanOut33[0] , \nOut10_10[0] , \nScanOut54[7] , \nOut7_10[4] , 
        \nScanOut132[3] , \nOut10_13[3] , \nScanOut252[6] , \nScanOut187[2] , 
        \nScanOut235[1] , \nScanOut1[5] , \nScanOut86[1] , \nScanOut155[4] , 
        \nScanOut2[6] , \nScanOut85[2] , \nScanOut156[7] , \nScanOut236[2] , 
        \nOut0_4[5] , \nScanOut57[4] , \nOut7_13[7] , \nScanOut184[1] , 
        \nOut0_7[6] , \nScanOut28[1] , \nOut6_4[1] , \nOut13_4[0] , 
        \nOut15_4[4] , \nOut14_15[3] , \nScanOut129[2] , \nOut9_10[0] , 
        \nOut9_13[3] , \nScanOut249[7] , \nOut13_7[3] , \nOut2_3[5] , 
        \nOut3_3[7] , \nOut3_0[4] , \nOut3_15[7] , \nOut5_0[0] , \nOut6_7[2] , 
        \nOut9_1[1] , \nOut15_7[7] , \nOut10_0[1] , \nOut5_3[3] , \nOut9_2[2] , 
        \nOut10_3[2] , \nOut11_3[0] , \nOut1_7[4] , \nOut2_0[6] , \nOut4_3[1] , 
        \nScanOut78[4] , \nOut8_1[3] , \nOut8_2[0] , \nScanOut179[7] , 
        \nScanOut219[2] , \nOut4_0[2] , \nOut11_0[3] , \nOut7_7[0] , 
        \nOut14_7[5] , \nOut7_4[3] , \nOut12_7[1] , \nOut14_4[6] , 
        \nOut0_14[0] , \nOut1_4[7] , \nOut12_4[2] , \nOut13_12[4] , 
        \nOut0_1[5] , \nScanOut9[0] , \nScanOut20[4] , \nOut4_11[3] , 
        \nScanOut60[6] , \nScanOut63[5] , \nScanOut162[6] , \nScanOut202[3] , 
        \nOut4_12[0] , \nScanOut106[2] , \nScanOut161[5] , \nScanOut201[0] , 
        \nOut13_11[7] , \nScanOut105[1] , \nOut5_14[3] , \nScanOut241[2] , 
        \nScanOut121[7] , \nScanOut23[7] , \nOut1_11[0] , \nOut3_8[1] , 
        \nScanOut44[0] , \nScanOut122[4] , \nScanOut242[1] , \nScanOut47[3] , 
        \nOut5_8[5] , \nScanOut95[5] , \nScanOut96[6] , \nScanOut197[5] , 
        \nScanOut225[6] , \nScanOut145[3] , \nOut12_14[7] , \nOut9_9[4] , 
        \nScanOut226[5] , \nScanOut146[0] , \nOut10_8[4] , \nScanOut194[6] , 
        \nOut1_12[3] , \nScanOut38[6] , \nScanOut139[5] , \nOut3_5[4] , 
        \nOut3_10[7] , \nScanOut98[0] , \nOut9_4[1] , \nOut5_5[0] , 
        \nScanOut199[3] , \nOut3_6[7] , \nOut3_13[4] , \nScanOut49[5] , 
        \nOut5_6[3] , \nOut10_5[1] , \nOut10_6[2] , \nOut9_7[2] , 
        \nScanOut228[3] , \nScanOut148[6] , \nOut13_1[0] , \nOut0_2[6] , 
        \nOut6_1[1] , \nOut9_15[0] , \nOut14_10[3] , \nOut15_1[4] , 
        \nScanOut4[5] , \nScanOut51[7] , \nOut6_2[2] , \nOut13_2[3] , 
        \nOut14_13[0] , \nOut15_2[7] , \nScanOut83[1] , \nOut7_15[4] , 
        \nScanOut182[2] , \nScanOut150[4] , \nScanOut230[1] , \nScanOut7[6] , 
        \nScanOut80[2] , \nScanOut233[2] , \nScanOut153[7] , \nScanOut11[5] , 
        \nScanOut12[6] , \nOut1_9[2] , \nScanOut35[3] , \nScanOut52[4] , 
        \nScanOut134[0] , \nScanOut181[1] , \nScanOut254[5] , \nScanOut36[0] , 
        \nOut10_15[0] , \nOut7_9[6] , \nScanOut137[3] , \nOut11_13[3] , 
        \nOut14_9[3] , \nOut12_9[7] , \nScanOut110[6] , \nScanOut113[5] , 
        \nOut11_10[0] , \nScanOut75[1] , \nScanOut76[2] , \nScanOut177[1] , 
        \nScanOut217[4] , \nOut6_10[4] , \nOut6_13[7] , \nScanOut108[4] , 
        \nScanOut174[2] , \nScanOut214[7] , \nOut8_13[3] , \nOut8_10[0] , 
        \nScanOut1[1] , \nScanOut2[2] , \nOut0_4[1] , \nOut0_7[2] , 
        \nOut2_15[7] , \nOut6_7[6] , \nOut15_7[3] , \nScanOut28[5] , 
        \nOut13_7[7] , \nOut6_4[5] , \nScanOut129[6] , \nOut9_10[4] , 
        \nOut9_13[7] , \nScanOut249[3] , \nOut13_4[4] , \nOut15_4[0] , 
        \nOut14_15[7] , \nScanOut30[7] , \nScanOut33[4] , \nOut3_3[3] , 
        \nOut9_2[6] , \nOut10_3[6] , \nOut3_0[0] , \nOut5_3[7] , \nOut3_15[3] , 
        \nOut10_0[5] , \nOut5_0[4] , \nOut9_1[5] , \nScanOut132[7] , 
        \nOut10_13[7] , \nScanOut252[2] , \nOut10_10[4] , \nScanOut57[0] , 
        \nScanOut131[4] , \nScanOut184[5] , \nScanOut251[1] , \nOut7_13[3] , 
        \nScanOut156[3] , \nScanOut85[6] , \nScanOut236[6] , \nScanOut155[0] , 
        \nScanOut54[3] , \nScanOut86[5] , \nOut7_10[0] , \nScanOut187[6] , 
        \nScanOut235[5] , \nOut4_8[3] , \nScanOut70[5] , \nScanOut171[6] , 
        \nScanOut211[3] , \nOut6_15[0] , \nScanOut73[6] , \nOut0_11[4] , 
        \nScanOut14[1] , \nOut2_8[7] , \nOut11_8[2] , \nOut8_9[2] , 
        \nScanOut212[0] , \nScanOut172[5] , \nScanOut17[2] , \nScanOut115[2] , 
        \nOut11_15[4] , \nScanOut116[1] , \nOut2_10[3] , \nOut2_13[0] , 
        \nScanOut169[4] , \nScanOut209[1] , \nScanOut68[7] , \nOut8_15[4] , 
        \nOut15_10[7] , \nOut15_13[4] , \nOut0_12[7] , \nOut1_1[3] , 
        \nOut12_1[6] , \nOut1_2[0] , \nOut7_1[7] , \nOut14_1[2] , 
        \nScanOut19[4] , \nOut7_2[4] , \nOut12_2[5] , \nOut14_2[1] , 
        \nOut2_5[2] , \nOut4_5[6] , \nScanOut118[7] , \nOut2_6[1] , 
        \nOut4_6[5] , \nOut8_4[7] , \nOut11_5[7] , \nOut8_7[4] , \nOut11_6[4] , 
        \nOut4_14[7] , \nScanOut100[5] , \nScanOut1[3] , \nOut0_4[3] , 
        \nOut0_9[6] , \nOut0_9[4] , \nScanOut41[4] , \nScanOut42[7] , 
        \nScanOut65[2] , \nScanOut103[6] , \nScanOut164[1] , \nScanOut204[4] , 
        \nOut13_14[3] , \nScanOut66[1] , \nScanOut167[2] , \nScanOut207[7] , 
        \nScanOut191[2] , \nScanOut90[1] , \nScanOut143[4] , \nOut12_12[0] , 
        \nScanOut93[2] , \nScanOut140[7] , \nScanOut223[1] , \nOut12_11[3] , 
        \nScanOut220[2] , \nScanOut192[1] , \nOut5_12[4] , \nScanOut127[0] , 
        \nScanOut247[5] , \nOut6_9[0] , \nOut15_9[5] , \nOut0_11[6] , 
        \nOut0_12[5] , \nScanOut25[0] , \nScanOut26[3] , \nOut13_9[1] , 
        \nOut1_14[4] , \nScanOut59[6] , \nOut5_11[7] , \nScanOut124[3] , 
        \nScanOut244[6] , \nScanOut158[5] , \nScanOut238[0] , \nScanOut88[3] , 
        \nScanOut189[0] , \nScanOut118[5] , \nOut1_1[1] , \nOut1_2[2] , 
        \nOut7_2[6] , \nOut14_2[3] , \nScanOut19[6] , \nOut12_2[7] , 
        \nOut7_1[5] , \nOut12_1[4] , \nOut14_1[0] , \nOut2_5[0] , \nOut2_6[3] , 
        \nOut11_6[6] , \nOut4_6[7] , \nOut8_4[5] , \nOut8_7[6] , 
        \nScanOut25[2] , \nScanOut41[6] , \nOut4_5[4] , \nOut11_5[5] , 
        \nOut4_14[5] , \nScanOut100[7] , \nScanOut103[4] , \nScanOut65[0] , 
        \nScanOut66[3] , \nScanOut167[0] , \nScanOut207[5] , \nScanOut164[3] , 
        \nOut13_14[1] , \nScanOut204[6] , \nScanOut42[5] , \nScanOut90[3] , 
        \nScanOut93[0] , \nScanOut192[3] , \nScanOut220[0] , \nScanOut140[5] , 
        \nOut12_11[1] , \nScanOut143[6] , \nOut12_12[2] , \nScanOut223[3] , 
        \nOut5_11[5] , \nScanOut191[0] , \nScanOut124[1] , \nScanOut244[4] , 
        \nScanOut26[1] , \nOut1_14[6] , \nScanOut59[4] , \nOut5_12[6] , 
        \nOut6_9[2] , \nOut13_9[3] , \nOut15_9[7] , \nScanOut88[1] , 
        \nScanOut127[2] , \nScanOut247[7] , \nScanOut189[2] , \nScanOut158[7] , 
        \nScanOut238[2] , \nOut13_4[6] , \nOut0_7[0] , \nOut6_4[7] , 
        \nScanOut129[4] , \nOut9_10[6] , \nOut15_4[2] , \nOut14_15[5] , 
        \nOut9_13[5] , \nScanOut249[1] , \nScanOut28[7] , \nScanOut30[5] , 
        \nOut3_3[1] , \nOut3_0[2] , \nOut3_15[1] , \nOut6_7[4] , \nOut13_7[5] , 
        \nOut15_7[1] , \nOut9_1[7] , \nOut5_0[6] , \nOut5_3[5] , \nOut10_0[7] , 
        \nOut10_3[4] , \nOut9_2[4] , \nScanOut131[6] , \nScanOut251[3] , 
        \nScanOut33[6] , \nOut10_10[6] , \nScanOut54[1] , \nOut7_10[2] , 
        \nScanOut132[5] , \nOut10_13[5] , \nScanOut252[0] , \nScanOut86[7] , 
        \nScanOut187[4] , \nScanOut235[7] , \nScanOut2[0] , \nScanOut85[4] , 
        \nScanOut155[2] , \nScanOut236[4] , \nOut2_8[5] , \nScanOut57[2] , 
        \nScanOut156[1] , \nOut7_13[1] , \nOut8_9[0] , \nScanOut184[7] , 
        \nOut11_8[0] , \nScanOut172[7] , \nScanOut212[2] , \nOut4_8[1] , 
        \nScanOut73[4] , \nScanOut70[7] , \nOut6_15[2] , \nScanOut171[4] , 
        \nScanOut211[1] , \nScanEnable[0] , \nScanOut14[3] , \nScanOut17[0] , 
        \nScanOut115[0] , \nScanOut116[3] , \nOut11_15[6] , \nOut2_10[1] , 
        \nOut2_13[2] , \nScanOut68[5] , \nScanOut169[6] , \nScanOut209[3] , 
        \nOut3_5[6] , \nOut3_6[5] , \nOut9_7[0] , \nOut8_15[6] , 
        \nOut15_10[5] , \nOut15_13[6] , \nScanOut148[4] , \nOut10_6[0] , 
        \nScanOut228[1] , \nOut3_13[6] , \nScanOut49[7] , \nOut5_6[1] , 
        \nOut3_10[5] , \nOut10_5[3] , \nScanOut199[1] , \nOut0_1[7] , 
        \nOut0_2[4] , \nOut5_5[2] , \nOut6_2[0] , \nScanOut98[2] , 
        \nOut9_4[3] , \nOut14_13[2] , \nOut15_2[5] , \nOut6_1[3] , 
        \nOut9_15[2] , \nOut13_2[1] , \nOut13_1[2] , \nOut14_10[1] , 
        \nOut15_1[6] , \nScanOut4[7] , \nScanOut7[4] , \nScanOut52[6] , 
        \nScanOut181[3] , \nScanOut80[0] , \nScanOut153[5] , \nScanOut233[0] , 
        \nScanOut11[7] , \nScanOut35[1] , \nScanOut36[2] , \nScanOut51[5] , 
        \nScanOut83[3] , \nScanOut150[6] , \nScanOut182[0] , \nScanOut230[3] , 
        \nOut7_15[6] , \nScanOut137[1] , \nOut10_15[2] , \nScanOut134[2] , 
        \nScanOut254[7] , \nScanOut12[4] , \nOut1_9[0] , \nScanOut110[4] , 
        \nOut11_10[2] , \nScanOut113[7] , \nScanOut75[3] , \nOut6_10[6] , 
        \nOut7_9[4] , \nOut12_9[5] , \nOut14_9[1] , \nOut11_13[1] , 
        \nScanOut174[0] , \nScanOut214[5] , \nScanOut76[0] , \nOut6_13[5] , 
        \nOut8_10[2] , \nScanOut177[3] , \nScanOut217[6] , \nOut2_15[5] , 
        \nScanOut108[6] , \nOut8_13[1] , \nOut0_14[2] , \nOut2_3[7] , 
        \nOut2_0[4] , \nOut4_0[0] , \nOut4_3[3] , \nScanOut78[6] , 
        \nOut8_1[1] , \nOut11_0[1] , \nOut8_2[2] , \nScanOut219[0] , 
        \nScanOut179[5] , \nOut11_3[2] , \nOut12_4[0] , \nScanOut1[7] , 
        \nScanOut2[4] , \nScanOut9[2] , \nOut1_4[5] , \nScanOut20[6] , 
        \nOut1_7[6] , \nOut7_4[1] , \nOut14_4[4] , \nScanOut23[5] , 
        \nOut4_11[1] , \nScanOut60[4] , \nOut7_7[2] , \nOut12_7[3] , 
        \nOut14_7[7] , \nScanOut161[7] , \nScanOut201[2] , \nOut13_11[5] , 
        \nScanOut63[7] , \nScanOut162[4] , \nScanOut202[1] , \nOut13_12[6] , 
        \nOut4_12[2] , \nScanOut105[3] , \nScanOut106[0] , \nScanOut122[6] , 
        \nScanOut242[3] , \nOut1_11[2] , \nOut1_12[1] , \nScanOut38[4] , 
        \nOut3_8[3] , \nOut5_14[1] , \nScanOut121[5] , \nOut10_8[6] , 
        \nScanOut241[0] , \nScanOut44[2] , \nScanOut47[1] , \nScanOut194[4] , 
        \nOut5_8[7] , \nScanOut95[7] , \nOut9_9[6] , \nScanOut146[2] , 
        \nScanOut96[4] , \nScanOut145[1] , \nOut12_14[5] , \nScanOut226[7] , 
        \nScanOut225[4] , \nScanOut197[7] , \nScanOut139[7] , \nScanOut14[7] , 
        \nOut2_8[1] , \nOut2_10[5] , \nOut2_13[6] , \nScanOut68[1] , 
        \nScanOut169[2] , \nScanOut209[7] , \nOut4_8[5] , \nScanOut70[3] , 
        \nOut8_15[2] , \nScanOut171[0] , \nScanOut211[5] , \nOut15_10[1] , 
        \nOut15_13[2] , \nScanOut73[0] , \nOut6_15[6] , \nOut8_9[4] , 
        \nOut11_8[4] , \nScanOut172[3] , \nScanOut212[6] , \nScanOut17[4] , 
        \nScanOut115[4] , \nOut11_15[2] , \nScanOut116[7] , \nScanOut30[1] , 
        \nScanOut33[2] , \nScanOut132[1] , \nOut10_13[1] , \nScanOut252[4] , 
        \nOut10_10[2] , \nScanOut57[6] , \nScanOut131[2] , \nScanOut184[3] , 
        \nScanOut251[7] , \nOut7_13[5] , \nScanOut85[0] , \nScanOut156[5] , 
        \nScanOut236[0] , \nScanOut155[6] , \nOut0_4[7] , \nOut0_7[4] , 
        \nScanOut28[3] , \nScanOut54[5] , \nScanOut86[3] , \nScanOut235[3] , 
        \nOut7_10[6] , \nScanOut187[0] , \nOut6_7[0] , \nOut15_7[5] , 
        \nOut13_7[1] , \nOut6_4[3] , \nScanOut129[0] , \nOut9_10[2] , 
        \nOut9_13[1] , \nScanOut249[5] , \nOut15_4[6] , \nOut14_15[1] , 
        \nScanOut9[6] , \nOut0_9[2] , \nScanOut26[5] , \nOut1_14[2] , 
        \nOut3_3[5] , \nOut9_2[0] , \nOut13_4[2] , \nOut3_0[6] , \nOut5_3[1] , 
        \nOut10_3[0] , \nOut10_0[3] , \nScanOut59[0] , \nOut3_15[5] , 
        \nOut5_0[2] , \nOut9_1[3] , \nScanOut158[3] , \nScanOut238[6] , 
        \nScanOut88[5] , \nScanOut189[6] , \nScanOut41[2] , \nScanOut42[1] , 
        \nScanOut191[4] , \nScanOut90[7] , \nScanOut143[2] , \nOut12_12[6] , 
        \nScanOut223[7] , \nScanOut93[4] , \nScanOut140[1] , \nOut12_11[5] , 
        \nScanOut192[7] , \nScanOut220[4] , \nOut5_12[2] , \nScanOut127[6] , 
        \nOut6_9[6] , \nScanOut247[3] , \nOut15_9[3] , \nOut13_9[7] , 
        \nOut0_11[2] , \nScanOut25[6] , \nOut4_14[1] , \nOut5_11[1] , 
        \nScanOut124[5] , \nScanOut244[0] , \nScanOut65[4] , \nScanOut100[3] , 
        \nScanOut103[0] , \nScanOut164[7] , \nScanOut204[2] , \nOut13_14[5] , 
        \nScanOut66[7] , \nScanOut167[4] , \nScanOut207[1] , \nOut0_12[1] , 
        \nOut1_1[5] , \nOut1_2[6] , \nScanOut19[2] , \nOut7_1[1] , 
        \nOut12_1[0] , \nOut14_1[4] , \nOut12_2[3] , \nOut7_2[2] , 
        \nOut14_2[7] , \nOut2_5[4] , \nOut4_5[0] , \nScanOut118[1] , 
        \nOut11_5[1] , \nOut2_6[7] , \nOut4_6[3] , \nOut8_4[1] , \nOut8_7[2] , 
        \nOut1_11[6] , \nOut11_6[2] , \nOut1_12[5] , \nScanOut38[0] , 
        \nScanOut139[3] , \nOut1_4[1] , \nOut2_3[3] , \nScanOut20[2] , 
        \nOut5_14[5] , \nScanOut121[1] , \nScanOut241[4] , \nScanOut23[1] , 
        \nOut3_8[7] , \nScanOut44[6] , \nScanOut122[2] , \nScanOut242[7] , 
        \nScanOut47[5] , \nScanOut95[3] , \nScanOut96[0] , \nScanOut197[3] , 
        \nScanOut145[5] , \nOut12_14[1] , \nScanOut225[0] , \nScanOut226[3] , 
        \nOut9_9[2] , \nScanOut146[6] , \nOut5_8[3] , \nOut4_11[5] , 
        \nScanOut60[0] , \nScanOut63[3] , \nOut10_8[2] , \nScanOut194[0] , 
        \nScanOut162[0] , \nOut13_12[2] , \nScanOut202[5] , \nOut4_12[6] , 
        \nScanOut106[4] , \nScanOut161[3] , \nScanOut201[6] , \nOut13_11[1] , 
        \nScanOut105[7] , \nOut1_7[2] , \nOut2_0[0] , \nOut4_3[7] , 
        \nScanOut78[2] , \nOut11_3[6] , \nOut8_1[5] , \nOut8_2[6] , 
        \nScanOut179[1] , \nScanOut219[4] , \nOut11_0[5] , \nOut4_0[4] , 
        \nOut7_7[6] , \nOut12_7[7] , \nOut14_7[3] , \nOut7_4[5] , 
        \nOut14_4[0] , \nOut12_4[4] , \nOut0_14[6] , \nScanOut108[2] , 
        \nOut8_13[5] , \nOut8_10[6] , \nScanOut0[3] , \nOut0_1[3] , 
        \nScanOut4[3] , \nScanOut11[3] , \nScanOut12[0] , \nOut2_15[1] , 
        \nOut7_9[0] , \nOut11_13[5] , \nOut12_9[1] , \nOut14_9[5] , 
        \nOut1_9[4] , \nScanOut110[0] , \nScanOut113[3] , \nOut11_10[6] , 
        \nScanOut51[1] , \nScanOut75[7] , \nScanOut76[4] , \nScanOut177[7] , 
        \nScanOut217[2] , \nOut6_10[2] , \nOut6_13[1] , \nScanOut174[4] , 
        \nScanOut214[1] , \nScanOut83[7] , \nOut7_15[2] , \nScanOut182[4] , 
        \nScanOut230[7] , \nScanOut7[0] , \nScanOut80[4] , \nScanOut150[2] , 
        \nScanOut233[4] , \nScanOut35[5] , \nScanOut52[2] , \nScanOut153[1] , 
        \nScanOut134[6] , \nScanOut181[7] , \nScanOut254[3] , \nScanOut36[6] , 
        \nOut10_15[6] , \nOut3_5[2] , \nOut3_10[1] , \nOut5_5[6] , 
        \nScanOut98[6] , \nScanOut137[5] , \nOut9_4[7] , \nOut10_5[7] , 
        \nOut3_6[1] , \nOut3_13[2] , \nScanOut199[5] , \nScanOut49[3] , 
        \nOut5_6[5] , \nOut9_7[4] , \nScanOut148[0] , \nOut10_6[4] , 
        \nScanOut228[5] , \nOut0_2[0] , \nOut6_1[7] , \nOut13_1[6] , 
        \nOut14_10[5] , \nOut15_1[2] , \nOut9_15[6] , \nOut13_2[5] , 
        \nScanOut3[0] , \nOut0_5[3] , \nOut0_6[0] , \nOut3_1[2] , \nOut3_2[1] , 
        \nOut5_2[5] , \nOut6_2[4] , \nOut14_13[6] , \nOut15_2[1] , 
        \nOut10_2[4] , \nOut3_14[1] , \nOut9_3[4] , \nOut9_0[7] , \nOut5_1[6] , 
        \nScanOut128[4] , \nOut9_12[5] , \nOut10_1[7] , \nScanOut248[1] , 
        \nScanOut29[7] , \nOut6_6[4] , \nOut13_6[5] , \nOut15_6[1] , 
        \nOut13_5[6] , \nScanOut84[4] , \nOut6_5[7] , \nOut9_11[6] , 
        \nOut14_14[5] , \nOut15_5[2] , \nScanOut237[4] , \nScanOut157[1] , 
        \nScanOut55[1] , \nScanOut56[2] , \nOut7_12[1] , \nScanOut185[7] , 
        \nScanOut87[7] , \nOut7_11[2] , \nScanOut186[4] , \nScanOut154[2] , 
        \nScanOut234[7] , \nScanOut15[3] , \nScanOut31[5] , \nScanOut32[6] , 
        \nScanOut130[6] , \nScanOut133[5] , \nOut10_12[5] , \nScanOut253[0] , 
        \nScanOut250[3] , \nScanOut114[0] , \nOut10_11[6] , \nOut11_14[6] , 
        \nScanOut16[0] , \nOut2_9[5] , \nScanOut71[7] , \nOut6_14[2] , 
        \nScanOut117[3] , \nOut8_8[0] , \nScanOut170[4] , \nScanOut210[1] , 
        \nOut11_9[0] , \nScanOut173[7] , \nScanOut213[2] , \nOut4_9[1] , 
        \nScanOut72[4] , \nOut8_14[6] , \nOut15_11[5] , \nOut15_12[6] , 
        \nOut0_10[6] , \nOut1_0[1] , \nOut2_4[0] , \nOut2_11[1] , 
        \nOut2_12[2] , \nScanOut69[5] , \nOut8_5[5] , \nScanOut168[6] , 
        \nScanOut208[3] , \nOut2_7[3] , \nOut4_4[4] , \nOut11_4[5] , 
        \nOut11_7[6] , \nOut4_7[7] , \nOut7_0[5] , \nOut8_6[6] , \nOut12_0[4] , 
        \nOut14_0[0] , \nOut0_13[5] , \nScanOut119[5] , \nScanOut18[6] , 
        \nOut1_3[2] , \nOut7_3[6] , \nOut14_3[3] , \nOut12_3[7] , 
        \nScanOut64[0] , \nScanOut67[3] , \nScanOut165[3] , \nScanOut166[0] , 
        \nScanOut205[6] , \nOut13_15[1] , \nScanOut206[5] , \nOut4_15[5] , 
        \nScanOut101[7] , \nOut0_8[6] , \nScanOut102[4] , \nScanOut27[1] , 
        \nOut6_8[2] , \nOut13_8[3] , \nOut15_8[7] , \nScanOut24[2] , 
        \nOut5_10[5] , \nOut5_13[6] , \nScanOut126[2] , \nScanOut246[7] , 
        \nScanOut125[1] , \nScanOut245[4] , \nScanOut43[5] , \nScanOut91[3] , 
        \nScanOut142[6] , \nScanOut222[3] , \nOut12_13[2] , \nOut1_6[6] , 
        \nOut1_15[6] , \nScanOut40[6] , \nScanOut190[0] , \nScanOut92[0] , 
        \nScanOut193[3] , \nScanOut221[0] , \nScanOut141[5] , \nOut12_10[1] , 
        \nScanOut58[4] , \nScanOut89[1] , \nScanOut159[7] , \nScanOut239[2] , 
        \nScanOut188[2] , \nOut7_6[2] , \nOut12_6[3] , \nOut14_6[7] , 
        \nOut2_1[4] , \nOut2_2[7] , \nOut1_5[5] , \nOut12_5[0] , \nOut4_2[3] , 
        \nScanOut79[6] , \nOut7_5[1] , \nOut8_3[2] , \nOut14_5[4] , 
        \nScanOut218[0] , \nScanOut178[5] , \nOut11_2[2] , \nOut4_1[0] , 
        \nScanOut21[6] , \nOut3_9[3] , \nScanOut45[2] , \nOut4_10[1] , 
        \nOut4_13[2] , \nOut8_0[1] , \nOut11_1[1] , \nScanOut107[0] , 
        \nScanOut61[4] , \nScanOut62[7] , \nScanOut104[3] , \nScanOut160[7] , 
        \nScanOut163[4] , \nScanOut203[1] , \nScanOut200[2] , \nOut13_13[6] , 
        \nOut13_10[5] , \nScanOut97[4] , \nScanOut144[1] , \nOut12_15[5] , 
        \nScanOut224[4] , \nScanOut196[7] , \nOut10_9[6] , \nScanOut46[1] , 
        \nOut5_9[7] , \nScanOut195[4] , \nScanOut94[7] , \nOut9_8[6] , 
        \nScanOut147[2] , \nScanOut227[7] , \nScanOut22[5] , \nOut5_15[1] , 
        \nScanOut120[5] , \nScanOut123[6] , \nScanOut240[0] , \nScanOut243[3] , 
        \nScanOut8[2] , \nOut1_10[2] , \nOut1_13[1] , \nScanOut39[4] , 
        \nScanOut138[7] , \nOut6_0[3] , \nOut9_14[2] , \nOut13_0[2] , 
        \nOut14_11[1] , \nOut0_3[4] , \nOut6_3[0] , \nOut14_12[2] , 
        \nOut15_3[5] , \nScanOut5[7] , \nScanOut34[1] , \nOut3_4[6] , 
        \nOut13_3[1] , \nOut3_7[5] , \nOut3_11[5] , \nOut10_4[3] , 
        \nScanOut198[1] , \nOut5_4[2] , \nScanOut99[2] , \nOut9_5[3] , 
        \nOut9_6[0] , \nScanOut149[4] , \nOut10_7[0] , \nScanOut229[1] , 
        \nOut3_12[6] , \nScanOut48[7] , \nOut5_7[1] , \nOut10_14[2] , 
        \nScanOut37[2] , \nScanOut135[2] , \nScanOut136[1] , \nScanOut255[7] , 
        \nScanOut256[4] , \nScanOut151[6] , \nScanOut6[4] , \nScanOut50[5] , 
        \nScanOut82[3] , \nOut7_14[6] , \nScanOut183[0] , \nScanOut231[3] , 
        \nScanOut53[6] , \nScanOut180[3] , \nScanOut152[5] , \nScanOut10[7] , 
        \nScanOut13[4] , \nOut1_8[0] , \nScanOut74[3] , \nScanOut77[0] , 
        \nScanOut81[0] , \nScanOut232[0] , \nOut6_12[5] , \nScanOut175[0] , 
        \nScanOut176[3] , \nScanOut216[6] , \nScanOut215[5] , \nOut6_11[6] , 
        \nScanOut112[7] , \nOut7_8[4] , \nOut11_12[1] , \nOut12_8[5] , 
        \nOut14_8[1] , \nScanOut24[6] , \nOut1_15[2] , \nOut2_14[5] , 
        \nScanOut111[4] , \nOut11_11[2] , \nScanOut109[6] , \nOut8_12[1] , 
        \nOut8_11[2] , \nOut15_14[1] , \nScanOut58[0] , \nScanOut89[5] , 
        \nScanOut188[6] , \nScanOut159[3] , \nScanOut239[6] , \nOut5_10[1] , 
        \nScanOut125[5] , \nOut5_13[2] , \nScanOut126[6] , \nScanOut245[0] , 
        \nOut6_8[6] , \nScanOut246[3] , \nOut0_8[2] , \nScanOut27[5] , 
        \nOut15_8[3] , \nOut13_8[7] , \nScanOut40[2] , \nScanOut92[4] , 
        \nScanOut141[1] , \nOut12_10[5] , \nScanOut193[7] , \nScanOut221[4] , 
        \nScanOut190[4] , \nOut0_10[2] , \nOut0_13[1] , \nScanOut18[2] , 
        \nOut2_4[4] , \nOut2_7[7] , \nScanOut43[1] , \nOut4_7[3] , 
        \nScanOut64[4] , \nScanOut67[7] , \nScanOut91[7] , \nScanOut142[2] , 
        \nOut12_13[6] , \nScanOut222[7] , \nScanOut165[7] , \nScanOut166[4] , 
        \nScanOut206[1] , \nScanOut205[2] , \nOut13_15[5] , \nOut4_15[1] , 
        \nScanOut102[0] , \nScanOut101[3] , \nOut8_6[2] , \nOut4_4[0] , 
        \nOut11_7[2] , \nOut11_4[1] , \nOut8_5[1] , \nOut1_3[6] , 
        \nOut12_3[3] , \nOut7_3[2] , \nOut14_3[7] , \nScanOut119[1] , 
        \nOut1_0[5] , \nOut2_12[6] , \nScanOut69[1] , \nOut7_0[1] , 
        \nOut12_0[0] , \nOut14_0[4] , \nOut8_14[2] , \nOut15_12[2] , 
        \nScanOut168[2] , \nScanOut208[7] , \nOut15_11[1] , \nScanOut0[7] , 
        \nScanOut15[7] , \nScanOut16[4] , \nOut2_11[5] , \nScanOut117[7] , 
        \nOut2_9[1] , \nOut4_9[5] , \nScanOut72[0] , \nScanOut114[4] , 
        \nOut11_14[2] , \nScanOut71[3] , \nOut6_14[6] , \nOut8_8[4] , 
        \nOut11_9[4] , \nScanOut173[3] , \nScanOut213[6] , \nScanOut170[0] , 
        \nScanOut210[5] , \nScanOut154[6] , \nScanOut3[4] , \nScanOut55[5] , 
        \nScanOut87[3] , \nScanOut234[3] , \nScanOut186[0] , \nScanOut56[6] , 
        \nOut7_11[6] , \nOut7_12[5] , \nScanOut185[3] , \nScanOut157[5] , 
        \nOut0_3[0] , \nScanOut5[3] , \nOut0_5[7] , \nScanOut31[1] , 
        \nScanOut84[0] , \nOut10_11[2] , \nScanOut237[0] , \nScanOut32[2] , 
        \nScanOut130[2] , \nScanOut133[1] , \nScanOut250[7] , \nOut10_12[1] , 
        \nScanOut253[4] , \nOut3_1[6] , \nOut10_1[3] , \nOut3_2[5] , 
        \nOut3_14[5] , \nOut5_1[2] , \nOut9_3[0] , \nOut9_0[3] , \nOut5_2[1] , 
        \nOut10_2[0] , \nOut6_5[3] , \nOut9_11[2] , \nOut14_14[1] , 
        \nOut15_5[6] , \nScanOut6[0] , \nOut0_6[4] , \nScanOut29[3] , 
        \nOut6_6[0] , \nOut13_5[2] , \nOut15_6[5] , \nOut13_6[1] , 
        \nScanOut10[3] , \nOut2_14[1] , \nScanOut128[0] , \nOut9_12[1] , 
        \nScanOut248[5] , \nScanOut74[7] , \nScanOut109[2] , \nOut8_11[6] , 
        \nOut15_14[5] , \nOut8_12[5] , \nScanOut77[4] , \nOut6_11[2] , 
        \nOut6_12[1] , \nScanOut175[4] , \nScanOut176[7] , \nScanOut215[1] , 
        \nScanOut216[2] , \nScanOut111[0] , \nOut11_11[6] , \nScanOut13[0] , 
        \nOut7_8[0] , \nOut11_12[5] , \nOut12_8[1] , \nOut14_8[5] , 
        \nOut1_8[4] , \nScanOut34[5] , \nScanOut37[6] , \nScanOut112[3] , 
        \nScanOut135[6] , \nScanOut136[5] , \nScanOut256[0] , \nScanOut255[3] , 
        \nScanOut81[4] , \nOut10_14[6] , \nScanOut152[1] , \nScanOut232[4] , 
        \nScanOut50[1] , \nScanOut53[2] , \nOut7_14[2] , \nScanOut180[7] , 
        \nScanOut82[7] , \nScanOut183[4] , \nScanOut231[7] , \nScanOut151[2] , 
        \nOut13_3[5] , \nOut6_3[4] , \nOut14_12[6] , \nOut15_3[1] , 
        \nScanOut8[6] , \nOut3_4[2] , \nOut3_7[1] , \nOut3_12[2] , 
        \nOut6_0[7] , \nOut13_0[6] , \nOut14_11[5] , \nOut9_14[6] , 
        \nScanOut48[3] , \nOut5_7[5] , \nOut3_11[1] , \nOut5_4[6] , 
        \nScanOut99[6] , \nOut9_6[4] , \nScanOut149[0] , \nOut10_7[4] , 
        \nScanOut229[5] , \nOut9_5[7] , \nOut10_4[7] , \nScanOut198[5] , 
        \nOut1_13[5] , \nScanOut39[0] , \nScanOut138[3] , \nScanOut21[2] , 
        \nScanOut22[1] , \nOut1_10[6] , \nOut3_9[7] , \nScanOut46[5] , 
        \nOut5_9[3] , \nScanOut94[3] , \nScanOut227[3] , \nOut9_8[2] , 
        \nScanOut147[6] , \nScanOut45[6] , \nOut10_9[2] , \nScanOut195[0] , 
        \nScanOut97[0] , \nScanOut196[3] , \nScanOut144[5] , \nScanOut224[0] , 
        \nOut12_15[1] , \nOut5_15[5] , \nScanOut123[2] , \nScanOut243[7] , 
        \nScanOut120[1] , \nScanOut240[4] , \nOut4_10[5] , \nScanOut104[7] , 
        \nScanOut8[4] , \nOut1_5[1] , \nScanOut61[0] , \nOut4_13[6] , 
        \nScanOut107[4] , \nScanOut62[3] , \nScanOut160[3] , \nOut13_10[1] , 
        \nScanOut163[0] , \nScanOut200[6] , \nScanOut203[5] , \nOut13_13[2] , 
        \nOut7_5[5] , \nOut14_5[0] , \nOut12_5[4] , \nOut2_1[0] , \nOut1_6[2] , 
        \nOut7_6[6] , \nOut12_6[7] , \nOut14_6[3] , \nOut8_0[5] , 
        \nOut11_1[5] , \nOut2_2[3] , \nOut4_1[4] , \nOut4_2[7] , 
        \nScanOut79[2] , \nOut11_2[6] , \nOut8_3[6] , \nScanOut178[1] , 
        \nScanOut218[4] , \nOut1_10[4] , \nScanOut21[0] , \nOut1_13[7] , 
        \nScanOut39[2] , \nScanOut138[1] , \nOut3_9[5] , \nScanOut45[4] , 
        \nScanOut97[2] , \nScanOut144[7] , \nOut12_15[3] , \nScanOut196[1] , 
        \nScanOut224[2] , \nScanOut195[2] , \nScanOut46[7] , \nOut10_9[0] , 
        \nOut5_9[1] , \nScanOut94[1] , \nOut9_8[0] , \nScanOut147[4] , 
        \nScanOut227[1] , \nOut1_6[0] , \nScanOut22[3] , \nOut5_15[7] , 
        \nScanOut120[3] , \nScanOut240[6] , \nScanOut123[0] , \nScanOut243[5] , 
        \nOut4_10[7] , \nOut4_13[4] , \nScanOut107[6] , \nScanOut61[2] , 
        \nScanOut62[1] , \nScanOut104[5] , \nScanOut160[1] , \nScanOut163[2] , 
        \nScanOut203[7] , \nScanOut200[4] , \nOut13_13[0] , \nOut13_10[3] , 
        \nOut12_6[5] , \nOut7_6[4] , \nOut14_6[1] , \nOut2_1[2] , \nOut2_2[1] , 
        \nOut1_5[3] , \nOut4_2[5] , \nOut7_5[7] , \nOut12_5[6] , \nOut14_5[2] , 
        \nOut8_3[4] , \nScanOut178[3] , \nScanOut218[6] , \nScanOut79[0] , 
        \nOut4_1[6] , \nOut11_2[4] , \nOut11_1[7] , \nOut2_14[3] , 
        \nOut8_0[7] , \nScanOut77[6] , \nOut6_12[3] , \nScanOut109[0] , 
        \nOut8_12[7] , \nOut8_11[4] , \nOut15_14[7] , \nScanOut5[1] , 
        \nScanOut10[1] , \nScanOut13[2] , \nScanOut74[5] , \nScanOut175[6] , 
        \nScanOut176[5] , \nScanOut216[0] , \nScanOut215[3] , \nOut6_11[0] , 
        \nScanOut112[1] , \nOut1_8[6] , \nOut12_8[3] , \nOut7_8[2] , 
        \nOut11_12[7] , \nOut14_8[7] , \nScanOut34[7] , \nScanOut111[2] , 
        \nOut11_11[4] , \nOut10_14[4] , \nScanOut37[4] , \nScanOut135[4] , 
        \nScanOut136[7] , \nScanOut255[1] , \nScanOut256[2] , \nScanOut6[2] , 
        \nScanOut50[3] , \nScanOut82[5] , \nScanOut151[0] , \nScanOut231[5] , 
        \nOut7_14[0] , \nScanOut183[6] , \nScanOut53[0] , \nScanOut180[5] , 
        \nScanOut81[6] , \nScanOut152[3] , \nOut6_0[5] , \nOut9_14[4] , 
        \nScanOut232[6] , \nOut14_11[7] , \nOut0_3[2] , \nOut6_3[6] , 
        \nOut13_0[4] , \nOut13_3[7] , \nOut14_12[4] , \nOut15_3[3] , 
        \nOut3_4[0] , \nOut10_4[5] , \nScanOut198[7] , \nOut3_7[3] , 
        \nOut3_11[3] , \nOut5_4[4] , \nScanOut99[4] , \nOut9_5[5] , 
        \nOut9_6[6] , \nScanOut149[2] , \nScanOut229[7] , \nOut3_12[0] , 
        \nOut10_7[6] , \nScanOut48[1] , \nOut5_7[7] , \nOut8_14[0] , 
        \nOut15_11[3] , \nOut15_12[0] , \nScanOut15[5] , \nOut2_11[7] , 
        \nOut2_12[4] , \nScanOut69[3] , \nScanOut114[6] , \nScanOut168[0] , 
        \nScanOut208[5] , \nOut11_14[0] , \nScanOut16[6] , \nScanOut117[5] , 
        \nScanOut0[5] , \nScanOut3[6] , \nOut2_9[3] , \nScanOut71[1] , 
        \nOut6_14[4] , \nOut8_8[6] , \nScanOut170[2] , \nScanOut173[1] , 
        \nScanOut210[7] , \nScanOut213[4] , \nOut4_9[7] , \nOut11_9[6] , 
        \nScanOut72[2] , \nScanOut84[2] , \nScanOut237[2] , \nScanOut55[7] , 
        \nScanOut56[4] , \nOut7_12[7] , \nScanOut157[7] , \nScanOut185[1] , 
        \nScanOut87[1] , \nOut7_11[4] , \nScanOut186[2] , \nScanOut234[1] , 
        \nOut0_5[5] , \nOut0_6[6] , \nScanOut29[1] , \nScanOut31[3] , 
        \nScanOut32[0] , \nScanOut154[4] , \nScanOut130[0] , \nScanOut133[3] , 
        \nOut10_12[3] , \nScanOut253[6] , \nScanOut250[5] , \nOut3_1[4] , 
        \nOut3_2[7] , \nOut5_2[3] , \nOut10_11[0] , \nOut3_14[7] , 
        \nOut5_1[0] , \nOut9_3[2] , \nOut10_2[2] , \nOut9_0[1] , \nOut10_1[1] , 
        \nScanOut128[2] , \nOut9_12[3] , \nScanOut248[7] , \nOut13_6[3] , 
        \nOut6_6[2] , \nOut15_6[7] , \nOut0_8[0] , \nScanOut27[7] , 
        \nOut1_15[0] , \nOut6_5[1] , \nOut13_5[0] , \nOut14_14[3] , 
        \nOut15_5[4] , \nOut9_11[0] , \nScanOut58[2] , \nScanOut89[7] , 
        \nScanOut159[1] , \nScanOut239[4] , \nScanOut188[4] , \nOut13_8[5] , 
        \nScanOut24[4] , \nOut5_10[3] , \nOut5_13[0] , \nOut6_8[4] , 
        \nOut15_8[1] , \nScanOut246[1] , \nScanOut126[4] , \nScanOut245[2] , 
        \nScanOut125[7] , \nScanOut91[5] , \nScanOut222[5] , \nScanOut142[0] , 
        \nOut12_13[4] , \nOut0_3[6] , \nOut0_10[0] , \nOut1_0[7] , 
        \nOut2_4[6] , \nScanOut40[0] , \nScanOut43[3] , \nScanOut190[6] , 
        \nScanOut64[6] , \nScanOut92[6] , \nScanOut193[5] , \nScanOut141[3] , 
        \nOut12_10[7] , \nScanOut221[6] , \nScanOut67[5] , \nScanOut165[5] , 
        \nScanOut166[6] , \nScanOut205[0] , \nOut13_15[7] , \nScanOut206[3] , 
        \nOut4_15[3] , \nScanOut101[1] , \nScanOut102[2] , \nOut8_5[3] , 
        \nOut11_4[3] , \nOut2_7[5] , \nOut4_4[2] , \nOut4_7[1] , \nOut11_7[0] , 
        \nOut7_0[3] , \nOut8_6[0] , \nOut14_0[6] , \nOut12_0[2] , 
        \nOut0_13[3] , \nScanOut119[3] , \nScanOut18[0] , \nOut7_3[0] , 
        \nOut12_3[1] , \nOut14_3[5] , \nOut1_3[4] , \nOut6_3[2] , 
        \nOut13_3[3] , \nOut14_12[0] , \nOut15_3[7] , \nOut13_0[0] , 
        \nScanOut5[5] , \nScanOut6[6] , \nScanOut34[3] , \nOut3_4[4] , 
        \nOut3_7[7] , \nOut3_12[4] , \nScanOut48[5] , \nOut6_0[1] , 
        \nOut9_14[0] , \nOut14_11[3] , \nOut5_7[3] , \nOut10_7[2] , 
        \nOut3_11[7] , \nScanOut99[0] , \nOut9_6[2] , \nScanOut229[3] , 
        \nScanOut149[6] , \nOut9_5[1] , \nOut5_4[0] , \nScanOut198[3] , 
        \nScanOut37[0] , \nOut10_4[1] , \nScanOut135[0] , \nScanOut136[3] , 
        \nScanOut256[6] , \nScanOut255[5] , \nScanOut81[2] , \nOut10_14[0] , 
        \nScanOut232[2] , \nScanOut50[7] , \nScanOut53[4] , \nScanOut152[7] , 
        \nOut7_14[4] , \nScanOut180[1] , \nScanOut82[1] , \nScanOut183[2] , 
        \nScanOut231[1] , \nScanOut8[0] , \nScanOut10[5] , \nScanOut74[1] , 
        \nScanOut151[4] , \nScanOut77[2] , \nOut6_11[4] , \nOut6_12[7] , 
        \nScanOut175[2] , \nScanOut176[1] , \nScanOut215[7] , \nScanOut216[4] , 
        \nScanOut111[6] , \nOut11_11[0] , \nScanOut13[6] , \nOut1_8[2] , 
        \nOut7_8[6] , \nOut14_8[3] , \nOut11_12[3] , \nOut12_8[7] , 
        \nOut1_5[7] , \nOut2_14[7] , \nScanOut112[5] , \nOut7_5[3] , 
        \nScanOut109[4] , \nOut8_11[0] , \nOut15_14[3] , \nOut8_12[3] , 
        \nOut12_5[2] , \nOut14_5[6] , \nOut2_1[6] , \nOut1_6[4] , \nOut7_6[0] , 
        \nOut14_6[5] , \nOut8_0[3] , \nOut12_6[1] , \nOut2_2[5] , \nOut4_1[2] , 
        \nOut11_1[3] , \nOut11_2[0] , \nScanOut21[4] , \nScanOut22[7] , 
        \nOut3_9[1] , \nScanOut46[3] , \nOut4_2[1] , \nOut4_10[3] , 
        \nScanOut79[4] , \nScanOut104[1] , \nOut8_3[0] , \nScanOut178[7] , 
        \nScanOut218[2] , \nScanOut61[6] , \nOut4_13[0] , \nScanOut107[2] , 
        \nScanOut62[5] , \nScanOut160[5] , \nOut13_10[7] , \nScanOut163[6] , 
        \nScanOut200[0] , \nScanOut203[3] , \nOut13_13[4] , \nScanOut94[5] , 
        \nOut9_8[4] , \nScanOut227[5] , \nScanOut147[0] , \nOut5_9[5] , 
        \nOut10_9[4] , \nScanOut195[6] , \nScanOut45[0] , \nScanOut97[6] , 
        \nScanOut196[5] , \nScanOut224[6] , \nScanOut144[3] , \nOut12_15[7] , 
        \nOut5_15[3] , \nScanOut123[4] , \nScanOut243[1] , \nScanOut240[2] , 
        \nScanOut120[7] , \nOut1_13[3] , \nScanOut39[6] , \nScanOut138[5] , 
        \nOut1_10[0] , \nOut0_10[4] , \nOut0_13[7] , \nScanOut18[4] , 
        \nOut1_3[0] , \nOut2_4[2] , \nOut2_7[1] , \nOut4_7[5] , \nOut8_6[4] , 
        \nOut11_7[4] , \nOut4_4[6] , \nOut8_5[7] , \nOut11_4[7] , \nOut7_3[4] , 
        \nOut12_3[5] , \nOut14_3[1] , \nScanOut119[7] , \nOut1_0[3] , 
        \nOut12_0[6] , \nScanOut24[0] , \nScanOut64[2] , \nScanOut67[1] , 
        \nOut7_0[7] , \nOut14_0[2] , \nScanOut165[1] , \nScanOut166[2] , 
        \nScanOut206[7] , \nScanOut205[4] , \nOut13_15[3] , \nOut4_15[7] , 
        \nScanOut102[6] , \nScanOut101[5] , \nScanOut125[3] , \nOut5_10[7] , 
        \nScanOut245[6] , \nOut5_13[4] , \nScanOut126[0] , \nScanOut246[5] , 
        \nOut15_8[5] , \nOut0_8[4] , \nOut6_8[0] , \nScanOut27[3] , 
        \nOut13_8[1] , \nScanOut40[4] , \nScanOut92[2] , \nScanOut141[7] , 
        \nOut12_10[3] , \nScanOut221[2] , \nScanOut193[1] , \nScanOut43[7] , 
        \nScanOut190[2] , \nScanOut0[1] , \nOut0_5[1] , \nOut1_15[4] , 
        \nScanOut91[1] , \nScanOut142[4] , \nOut12_13[0] , \nScanOut222[1] , 
        \nOut3_1[0] , \nScanOut58[6] , \nScanOut89[3] , \nScanOut188[0] , 
        \nScanOut159[5] , \nScanOut239[0] , \nOut3_2[3] , \nOut3_14[3] , 
        \nOut10_1[5] , \nOut5_1[4] , \nOut9_3[6] , \nOut9_0[5] , \nOut10_2[6] , 
        \nOut5_2[7] , \nOut6_5[5] , \nOut9_11[4] , \nOut13_5[4] , 
        \nOut14_14[7] , \nOut15_5[0] , \nOut0_6[2] , \nOut6_6[6] , 
        \nOut15_6[3] , \nScanOut29[5] , \nOut13_6[7] , \nScanOut128[6] , 
        \nOut9_12[7] , \nScanOut248[3] , \nScanOut3[2] , \nScanOut55[3] , 
        \nScanOut87[5] , \nScanOut154[0] , \nScanOut186[6] , \nScanOut234[5] , 
        \nScanOut56[0] , \nOut7_11[0] , \nOut7_12[3] , \nScanOut185[5] , 
        \nScanOut15[1] , \nScanOut16[2] , \nScanOut31[7] , \nScanOut84[6] , 
        \nScanOut157[3] , \nScanOut237[6] , \nOut10_11[4] , \nScanOut32[4] , 
        \nScanOut130[4] , \nScanOut133[7] , \nScanOut250[1] , \nOut10_12[7] , 
        \nScanOut253[2] , \nScanOut117[1] , \nOut2_9[7] , \nOut4_9[3] , 
        \nScanOut114[2] , \nOut11_14[4] , \nScanOut72[6] , \nOut11_9[2] , 
        \nOut2_12[0] , \nScanOut71[5] , \nOut6_14[0] , \nOut8_8[2] , 
        \nScanOut213[0] , \nScanOut170[6] , \nScanOut173[5] , \nScanOut210[3] , 
        \nOut8_14[4] , \nOut15_12[4] , \nScanOut168[4] , \nScanOut208[1] , 
        \nOut15_11[7] , \nScanOut69[7] , \nScanOut5[4] , \nOut2_11[3] , 
        \nScanOut34[2] , \nScanOut135[1] , \nOut10_14[1] , \nScanOut255[4] , 
        \nScanOut37[1] , \nScanOut50[6] , \nScanOut136[2] , \nScanOut183[3] , 
        \nScanOut256[7] , \nOut7_14[5] , \nScanOut151[5] , \nScanOut6[7] , 
        \nScanOut82[0] , \nScanOut231[0] , \nScanOut152[6] , \nScanOut53[5] , 
        \nScanOut81[3] , \nScanOut180[0] , \nScanOut232[3] , \nOut6_0[0] , 
        \nOut14_11[2] , \nOut0_3[7] , \nOut6_3[3] , \nOut9_14[1] , 
        \nOut13_0[1] , \nOut13_3[2] , \nOut14_12[1] , \nOut15_3[6] , 
        \nScanOut8[1] , \nScanOut10[4] , \nScanOut13[7] , \nOut2_14[6] , 
        \nOut3_4[5] , \nScanOut99[1] , \nOut9_5[0] , \nOut10_4[0] , 
        \nScanOut198[2] , \nOut3_7[6] , \nOut3_11[6] , \nOut5_4[1] , 
        \nOut3_12[5] , \nOut10_7[3] , \nScanOut48[4] , \nOut5_7[2] , 
        \nOut9_6[3] , \nScanOut149[7] , \nScanOut229[2] , \nScanOut74[0] , 
        \nScanOut77[3] , \nScanOut109[5] , \nOut8_12[2] , \nOut8_11[1] , 
        \nOut15_14[2] , \nScanOut176[0] , \nScanOut216[5] , \nOut6_11[5] , 
        \nOut6_12[6] , \nScanOut175[3] , \nScanOut215[6] , \nOut1_8[3] , 
        \nOut12_8[6] , \nOut7_8[7] , \nOut11_12[2] , \nScanOut111[7] , 
        \nScanOut112[4] , \nOut14_8[2] , \nOut1_5[6] , \nOut1_6[5] , 
        \nOut4_10[2] , \nOut4_13[1] , \nOut11_11[1] , \nScanOut107[3] , 
        \nScanOut61[7] , \nScanOut62[4] , \nScanOut104[0] , \nScanOut163[7] , 
        \nScanOut203[2] , \nOut13_13[5] , \nScanOut160[4] , \nScanOut200[1] , 
        \nOut12_6[0] , \nOut13_10[6] , \nOut7_6[1] , \nOut14_6[4] , 
        \nOut7_5[2] , \nOut12_5[3] , \nOut14_5[7] , \nOut2_1[7] , \nOut2_2[4] , 
        \nOut4_2[0] , \nScanOut79[5] , \nOut4_1[3] , \nOut8_3[1] , 
        \nOut11_2[1] , \nScanOut178[6] , \nScanOut218[3] , \nOut8_0[2] , 
        \nOut11_1[2] , \nOut1_10[1] , \nOut1_13[2] , \nScanOut138[4] , 
        \nOut0_8[5] , \nOut0_10[5] , \nOut2_4[3] , \nScanOut21[5] , 
        \nScanOut39[7] , \nOut3_9[0] , \nScanOut45[1] , \nScanOut196[4] , 
        \nScanOut94[4] , \nScanOut97[7] , \nScanOut144[2] , \nOut12_15[6] , 
        \nOut9_8[5] , \nScanOut147[1] , \nScanOut224[7] , \nScanOut227[4] , 
        \nScanOut195[7] , \nScanOut46[2] , \nOut5_9[4] , \nOut10_9[5] , 
        \nOut5_15[2] , \nScanOut120[6] , \nScanOut240[3] , \nScanOut22[6] , 
        \nScanOut64[3] , \nScanOut123[5] , \nScanOut165[0] , \nOut13_15[2] , 
        \nScanOut243[0] , \nScanOut205[5] , \nScanOut67[0] , \nOut4_15[6] , 
        \nScanOut101[4] , \nScanOut166[3] , \nScanOut206[6] , \nScanOut102[7] , 
        \nOut11_4[6] , \nOut2_7[0] , \nOut4_4[7] , \nOut8_5[6] , \nOut8_6[5] , 
        \nOut4_7[4] , \nOut11_7[5] , \nOut0_13[6] , \nOut1_0[2] , \nOut7_0[6] , 
        \nOut14_0[3] , \nScanOut18[5] , \nOut7_3[5] , \nOut12_0[7] , 
        \nOut12_3[4] , \nOut14_3[0] , \nOut1_3[1] , \nScanOut119[6] , 
        \nScanOut27[2] , \nOut1_15[5] , \nScanOut58[7] , \nScanOut159[4] , 
        \nScanOut239[1] , \nOut5_13[5] , \nScanOut89[2] , \nScanOut188[1] , 
        \nScanOut246[4] , \nScanOut126[1] , \nOut13_8[0] , \nScanOut24[1] , 
        \nOut6_8[1] , \nOut15_8[4] , \nOut5_10[6] , \nScanOut245[7] , 
        \nScanOut125[2] , \nScanOut0[0] , \nScanOut3[3] , \nScanOut40[5] , 
        \nScanOut43[6] , \nScanOut91[0] , \nScanOut190[3] , \nScanOut222[0] , 
        \nScanOut92[3] , \nScanOut142[5] , \nOut12_13[1] , \nScanOut141[6] , 
        \nScanOut221[3] , \nOut12_10[2] , \nScanOut56[1] , \nScanOut193[0] , 
        \nScanOut84[7] , \nOut7_12[2] , \nScanOut185[4] , \nScanOut157[2] , 
        \nScanOut237[7] , \nScanOut87[4] , \nScanOut234[4] , \nScanOut154[1] , 
        \nOut0_5[0] , \nOut0_6[3] , \nScanOut29[4] , \nScanOut31[6] , 
        \nScanOut32[5] , \nScanOut55[2] , \nOut7_11[1] , \nScanOut133[6] , 
        \nScanOut186[7] , \nScanOut253[3] , \nOut10_12[6] , \nOut3_1[1] , 
        \nOut3_2[2] , \nOut5_2[6] , \nScanOut130[5] , \nOut10_11[5] , 
        \nScanOut250[0] , \nOut9_3[7] , \nOut3_14[2] , \nOut5_1[5] , 
        \nOut10_2[7] , \nOut10_1[4] , \nOut9_0[4] , \nOut13_6[6] , 
        \nOut6_6[7] , \nScanOut128[7] , \nOut9_12[6] , \nOut15_6[2] , 
        \nScanOut248[2] , \nOut9_11[5] , \nOut2_11[2] , \nOut6_5[4] , 
        \nOut13_5[5] , \nOut14_14[6] , \nOut15_5[1] , \nOut8_14[5] , 
        \nOut15_11[6] , \nOut15_12[5] , \nScanOut8[5] , \nScanOut15[0] , 
        \nOut2_12[1] , \nScanOut69[6] , \nScanOut168[5] , \nScanOut208[0] , 
        \nOut11_14[5] , \nScanOut16[3] , \nScanOut114[3] , \nScanOut117[0] , 
        \nScanOut21[1] , \nScanOut22[2] , \nOut2_9[6] , \nScanOut71[4] , 
        \nScanOut170[7] , \nScanOut210[2] , \nOut6_14[1] , \nOut3_9[4] , 
        \nScanOut46[6] , \nOut4_9[2] , \nOut11_9[3] , \nScanOut72[7] , 
        \nOut5_9[0] , \nOut8_8[3] , \nScanOut173[4] , \nScanOut213[1] , 
        \nOut10_9[1] , \nScanOut195[3] , \nScanOut45[5] , \nScanOut94[0] , 
        \nScanOut97[3] , \nOut9_8[1] , \nScanOut227[0] , \nScanOut147[5] , 
        \nScanOut224[3] , \nScanOut144[6] , \nOut12_15[2] , \nScanOut123[1] , 
        \nScanOut196[0] , \nScanOut243[4] , \nOut5_15[6] , \nScanOut240[7] , 
        \nScanOut120[2] , \nScanOut39[3] , \nOut1_10[5] , \nOut1_13[6] , 
        \nScanOut138[0] , \nOut2_1[3] , \nOut1_5[2] , \nOut7_5[6] , 
        \nOut12_5[7] , \nOut14_5[3] , \nOut1_6[1] , \nOut7_6[5] , 
        \nOut14_6[0] , \nOut12_6[4] , \nOut2_2[0] , \nOut4_1[7] , 
        \nOut11_1[6] , \nOut8_3[5] , \nOut8_0[6] , \nOut11_2[5] , 
        \nScanOut178[2] , \nScanOut218[7] , \nOut4_2[4] , \nOut4_10[6] , 
        \nScanOut79[1] , \nScanOut104[4] , \nScanOut61[3] , \nOut4_13[5] , 
        \nScanOut107[7] , \nScanOut160[0] , \nScanOut200[5] , \nOut13_10[2] , 
        \nScanOut62[0] , \nScanOut74[4] , \nOut6_11[1] , \nScanOut163[3] , 
        \nOut13_13[1] , \nScanOut175[7] , \nScanOut203[6] , \nScanOut215[2] , 
        \nScanOut77[7] , \nOut6_12[2] , \nScanOut176[4] , \nOut0_3[3] , 
        \nScanOut10[0] , \nOut11_11[5] , \nScanOut216[1] , \nScanOut13[3] , 
        \nOut1_8[7] , \nOut7_8[3] , \nScanOut111[3] , \nScanOut112[0] , 
        \nOut11_12[6] , \nOut14_8[6] , \nOut12_8[2] , \nOut2_14[2] , 
        \nScanOut109[1] , \nOut8_11[5] , \nOut15_14[6] , \nOut8_12[6] , 
        \nOut6_3[7] , \nOut13_3[6] , \nOut14_12[5] , \nOut15_3[2] , 
        \nOut9_14[5] , \nOut13_0[5] , \nScanOut5[0] , \nScanOut6[3] , 
        \nScanOut34[6] , \nOut3_4[1] , \nOut3_7[2] , \nOut3_12[1] , 
        \nScanOut48[0] , \nOut5_7[6] , \nOut6_0[4] , \nOut9_6[7] , 
        \nOut14_11[6] , \nScanOut229[6] , \nScanOut149[3] , \nOut10_7[7] , 
        \nOut3_11[2] , \nOut5_4[5] , \nScanOut198[6] , \nScanOut37[5] , 
        \nScanOut99[5] , \nOut10_4[4] , \nOut9_5[4] , \nScanOut136[6] , 
        \nScanOut256[3] , \nScanOut53[1] , \nScanOut135[5] , \nOut10_14[5] , 
        \nScanOut255[0] , \nScanOut81[7] , \nScanOut180[4] , \nScanOut232[7] , 
        \nScanOut152[2] , \nScanOut82[4] , \nScanOut151[1] , \nScanOut231[4] , 
        \nScanOut15[4] , \nScanOut16[7] , \nScanOut50[2] , \nOut7_14[1] , 
        \nScanOut183[7] , \nScanOut114[7] , \nScanOut117[4] , \nOut2_9[2] , 
        \nOut4_9[6] , \nOut8_8[7] , \nOut11_14[1] , \nScanOut213[5] , 
        \nScanOut173[0] , \nScanOut72[3] , \nOut11_9[7] , \nOut2_11[6] , 
        \nOut2_12[5] , \nScanOut71[0] , \nOut6_14[5] , \nOut8_14[1] , 
        \nScanOut170[3] , \nScanOut210[6] , \nOut15_11[2] , \nOut15_12[1] , 
        \nScanOut69[2] , \nScanOut168[1] , \nScanOut208[4] , \nScanOut0[4] , 
        \nOut0_5[4] , \nOut3_1[5] , \nOut9_0[0] , \nOut3_2[6] , \nOut3_14[6] , 
        \nOut10_1[0] , \nOut5_1[1] , \nOut10_2[3] , \nOut5_2[2] , \nOut6_5[0] , 
        \nOut9_3[3] , \nOut13_5[1] , \nOut14_14[2] , \nOut15_5[5] , 
        \nOut0_6[7] , \nOut6_6[3] , \nScanOut128[3] , \nOut9_11[1] , 
        \nOut9_12[2] , \nScanOut248[6] , \nOut15_6[6] , \nScanOut29[0] , 
        \nOut13_6[2] , \nScanOut55[6] , \nOut7_11[5] , \nScanOut186[3] , 
        \nScanOut154[5] , \nScanOut3[7] , \nScanOut87[0] , \nScanOut157[6] , 
        \nScanOut234[0] , \nScanOut24[5] , \nScanOut31[2] , \nScanOut56[5] , 
        \nScanOut84[3] , \nScanOut237[3] , \nScanOut185[0] , \nOut7_12[6] , 
        \nScanOut130[1] , \nOut10_11[1] , \nScanOut250[4] , \nScanOut32[1] , 
        \nOut10_12[2] , \nOut5_10[2] , \nScanOut125[6] , \nScanOut133[2] , 
        \nScanOut253[7] , \nScanOut245[3] , \nOut15_8[0] , \nOut0_8[1] , 
        \nOut6_8[5] , \nScanOut27[6] , \nOut13_8[4] , \nScanOut40[1] , 
        \nOut5_13[1] , \nScanOut126[5] , \nScanOut246[0] , \nScanOut193[4] , 
        \nScanOut43[2] , \nScanOut91[4] , \nScanOut92[7] , \nScanOut141[2] , 
        \nOut12_10[6] , \nScanOut221[7] , \nScanOut142[1] , \nOut12_13[5] , 
        \nScanOut190[7] , \nScanOut222[4] , \nOut0_8[3] , \nOut0_10[1] , 
        \nOut0_13[2] , \nOut2_4[7] , \nOut2_7[4] , \nOut1_15[1] , \nOut4_7[0] , 
        \nScanOut58[3] , \nScanOut89[6] , \nScanOut188[5] , \nScanOut159[0] , 
        \nScanOut239[5] , \nOut11_7[1] , \nOut4_4[3] , \nOut8_5[2] , 
        \nOut8_6[1] , \nOut11_4[2] , \nOut1_0[6] , \nScanOut18[1] , 
        \nOut1_3[5] , \nScanOut119[2] , \nOut7_3[1] , \nOut12_3[0] , 
        \nOut14_3[4] , \nOut12_0[3] , \nOut7_0[2] , \nOut14_0[7] , 
        \nScanOut64[7] , \nScanOut67[4] , \nScanOut166[7] , \nScanOut206[2] , 
        \nOut5_13[3] , \nOut4_15[2] , \nScanOut102[3] , \nScanOut165[4] , 
        \nScanOut205[1] , \nOut13_15[6] , \nScanOut101[0] , \nScanOut126[7] , 
        \nScanOut246[2] , \nScanOut27[4] , \nOut6_8[7] , \nOut13_8[6] , 
        \nOut15_8[2] , \nScanOut24[7] , \nScanOut43[0] , \nOut5_10[0] , 
        \nScanOut125[4] , \nScanOut245[1] , \nOut0_10[3] , \nOut2_4[5] , 
        \nOut1_15[3] , \nScanOut40[3] , \nScanOut91[6] , \nScanOut190[5] , 
        \nScanOut92[5] , \nScanOut142[3] , \nOut12_13[7] , \nScanOut222[6] , 
        \nScanOut221[5] , \nScanOut141[0] , \nOut12_10[4] , \nScanOut193[6] , 
        \nScanOut58[1] , \nScanOut159[2] , \nScanOut239[7] , \nScanOut89[4] , 
        \nScanOut188[7] , \nOut2_7[6] , \nOut4_4[1] , \nOut11_4[0] , 
        \nOut8_5[0] , \nOut8_6[3] , \nOut11_7[3] , \nOut4_7[2] , \nOut0_13[0] , 
        \nOut1_0[4] , \nOut7_0[0] , \nOut12_0[1] , \nOut14_0[5] , 
        \nScanOut18[3] , \nOut1_3[7] , \nOut7_3[3] , \nOut14_3[6] , 
        \nOut12_3[2] , \nScanOut119[0] , \nScanOut15[6] , \nScanOut64[5] , 
        \nScanOut165[6] , \nOut13_15[4] , \nScanOut205[3] , \nScanOut67[6] , 
        \nOut4_15[0] , \nScanOut101[2] , \nScanOut166[5] , \nScanOut206[0] , 
        \nScanOut102[1] , \nOut11_14[3] , \nScanOut16[5] , \nScanOut114[5] , 
        \nScanOut117[6] , \nOut2_9[0] , \nScanOut71[2] , \nScanOut170[1] , 
        \nScanOut210[4] , \nOut6_14[7] , \nOut11_9[5] , \nOut2_11[4] , 
        \nOut4_9[4] , \nScanOut72[1] , \nOut8_8[5] , \nOut8_14[3] , 
        \nScanOut173[2] , \nScanOut213[7] , \nOut15_11[0] , \nOut15_12[3] , 
        \nScanOut0[6] , \nScanOut3[5] , \nOut0_5[6] , \nOut0_6[5] , 
        \nOut2_12[7] , \nScanOut168[3] , \nScanOut208[6] , \nOut3_1[7] , 
        \nOut3_2[4] , \nOut5_2[0] , \nScanOut69[0] , \nOut9_3[1] , 
        \nOut10_2[1] , \nOut3_14[4] , \nOut5_1[3] , \nOut9_0[2] , 
        \nOut10_1[2] , \nScanOut29[2] , \nOut6_6[1] , \nOut13_6[0] , 
        \nOut15_6[4] , \nScanOut128[1] , \nOut9_12[0] , \nScanOut248[4] , 
        \nOut9_11[3] , \nOut13_5[3] , \nScanOut56[7] , \nOut6_5[2] , 
        \nOut14_14[0] , \nOut15_5[7] , \nScanOut84[1] , \nOut7_12[4] , 
        \nScanOut185[2] , \nScanOut237[1] , \nScanOut87[2] , \nScanOut157[4] , 
        \nScanOut234[2] , \nScanOut10[2] , \nScanOut13[1] , \nOut1_8[5] , 
        \nScanOut31[0] , \nScanOut32[3] , \nScanOut55[4] , \nOut7_11[7] , 
        \nScanOut154[7] , \nScanOut133[0] , \nScanOut186[1] , \nScanOut253[5] , 
        \nOut10_12[0] , \nScanOut74[6] , \nScanOut77[5] , \nScanOut130[3] , 
        \nOut10_11[3] , \nScanOut250[6] , \nScanOut176[6] , \nScanOut216[3] , 
        \nOut6_11[3] , \nOut6_12[0] , \nScanOut175[5] , \nScanOut215[0] , 
        \nOut7_8[1] , \nOut12_8[0] , \nOut14_8[4] , \nScanOut111[1] , 
        \nScanOut112[2] , \nOut11_12[4] , \nOut2_14[0] , \nOut11_11[7] , 
        \nOut6_0[6] , \nScanOut109[3] , \nOut8_12[4] , \nOut8_11[7] , 
        \nOut15_14[4] , \nOut13_0[7] , \nOut14_11[4] , \nOut0_3[1] , 
        \nOut6_3[5] , \nOut9_14[7] , \nOut14_12[7] , \nOut15_3[0] , 
        \nScanOut5[2] , \nScanOut34[4] , \nOut3_4[3] , \nScanOut99[7] , 
        \nOut9_5[6] , \nOut13_3[4] , \nOut3_7[0] , \nOut3_11[0] , 
        \nOut10_4[6] , \nScanOut198[4] , \nOut5_4[7] , \nOut10_7[5] , 
        \nOut3_12[3] , \nScanOut48[2] , \nOut5_7[4] , \nOut9_6[5] , 
        \nScanOut135[7] , \nScanOut149[1] , \nScanOut229[4] , \nOut10_14[7] , 
        \nScanOut255[2] , \nScanOut37[7] , \nScanOut50[0] , \nScanOut136[4] , 
        \nScanOut183[5] , \nScanOut256[1] , \nOut7_14[3] , \nScanOut6[1] , 
        \nScanOut82[6] , \nScanOut151[3] , \nScanOut231[6] , \nScanOut45[7] , 
        \nScanOut53[3] , \nScanOut81[5] , \nScanOut152[0] , \nScanOut232[5] , 
        \nScanOut180[6] , \nScanOut196[2] , \nScanOut94[2] , \nScanOut97[1] , 
        \nScanOut144[4] , \nOut12_15[0] , \nScanOut224[1] , \nOut9_8[3] , 
        \nScanOut147[7] , \nScanOut227[2] , \nScanOut8[7] , \nScanOut21[3] , 
        \nOut3_9[6] , \nOut10_9[3] , \nScanOut46[4] , \nScanOut195[1] , 
        \nOut5_9[2] , \nOut5_15[4] , \nScanOut120[0] , \nScanOut240[5] , 
        \nScanOut22[0] , \nScanOut123[3] , \nScanOut243[6] , \nOut1_10[7] , 
        \nOut1_13[4] , \nScanOut138[2] , \nScanOut0[2] , \nOut1_5[0] , 
        \nOut1_6[3] , \nScanOut39[1] , \nOut7_6[7] , \nOut12_6[6] , 
        \nOut14_6[2] , \nOut12_5[5] , \nOut7_5[4] , \nOut14_5[1] , 
        \nOut2_1[1] , \nOut2_2[2] , \nOut4_2[6] , \nScanOut79[3] , 
        \nOut11_2[7] , \nOut4_1[5] , \nOut8_3[7] , \nScanOut218[5] , 
        \nOut8_0[4] , \nScanOut178[0] , \nScanOut55[0] , \nOut4_10[4] , 
        \nOut4_13[7] , \nOut11_1[4] , \nScanOut107[5] , \nScanOut61[1] , 
        \nScanOut62[2] , \nScanOut104[6] , \nScanOut163[1] , \nScanOut203[4] , 
        \nOut13_13[3] , \nOut7_11[3] , \nScanOut160[2] , \nScanOut200[7] , 
        \nScanOut186[5] , \nOut13_10[0] , \nScanOut3[1] , \nScanOut87[6] , 
        \nScanOut154[3] , \nScanOut234[6] , \nOut0_5[2] , \nScanOut31[4] , 
        \nScanOut56[3] , \nScanOut84[5] , \nScanOut157[0] , \nScanOut185[6] , 
        \nScanOut237[5] , \nOut7_12[0] , \nScanOut130[7] , \nOut10_11[7] , 
        \nScanOut250[2] , \nScanOut32[7] , \nOut10_12[4] , \nOut3_1[3] , 
        \nScanOut133[4] , \nOut9_0[6] , \nScanOut253[1] , \nOut10_1[6] , 
        \nOut3_2[0] , \nOut3_14[0] , \nOut5_1[7] , \nOut5_2[4] , \nOut10_2[5] , 
        \nOut6_5[6] , \nOut9_3[5] , \nOut14_14[4] , \nOut15_5[3] , 
        \nOut0_6[1] , \nScanOut29[6] , \nOut6_6[5] , \nScanOut128[5] , 
        \nOut9_11[7] , \nOut13_5[7] , \nOut9_12[4] , \nScanOut248[0] , 
        \nOut15_6[0] , \nOut13_6[4] , \nOut2_11[0] , \nOut2_12[3] , 
        \nScanOut69[4] , \nOut8_14[7] , \nOut15_11[4] , \nOut15_12[7] , 
        \nScanOut168[7] , \nScanOut208[2] , \nOut0_10[7] , \nOut0_13[4] , 
        \nScanOut15[2] , \nScanOut16[1] , \nScanOut114[1] , \nScanOut117[2] , 
        \nOut2_4[1] , \nOut2_7[2] , \nOut2_9[4] , \nOut4_9[0] , 
        \nScanOut72[5] , \nOut8_8[1] , \nScanOut173[6] , \nOut11_14[7] , 
        \nScanOut213[3] , \nOut4_7[6] , \nScanOut64[1] , \nScanOut67[2] , 
        \nScanOut71[6] , \nOut11_9[1] , \nOut6_14[3] , \nScanOut166[1] , 
        \nScanOut170[5] , \nScanOut210[0] , \nScanOut206[4] , \nOut4_15[4] , 
        \nScanOut102[5] , \nScanOut165[2] , \nScanOut205[7] , \nOut13_15[0] , 
        \nScanOut101[6] , \nOut4_4[5] , \nOut8_5[4] , \nOut8_6[7] , 
        \nOut11_7[7] , \nOut11_4[4] , \nOut1_0[0] , \nScanOut18[7] , 
        \nScanOut119[4] , \nOut1_3[3] , \nOut12_3[6] , \nOut7_3[7] , 
        \nOut14_3[2] , \nOut7_0[4] , \nOut12_0[5] , \nOut14_0[1] , 
        \nScanOut24[3] , \nOut1_15[7] , \nScanOut58[5] , \nScanOut89[0] , 
        \nScanOut188[3] , \nOut5_10[4] , \nScanOut125[0] , \nScanOut159[6] , 
        \nScanOut239[3] , \nScanOut245[5] , \nOut6_8[3] , \nOut0_8[7] , 
        \nScanOut27[0] , \nOut15_8[6] , \nOut13_8[2] , \nScanOut40[7] , 
        \nOut5_13[7] , \nScanOut126[3] , \nScanOut193[2] , \nScanOut246[6] , 
        \nScanOut91[2] , \nScanOut92[1] , \nScanOut141[4] , \nOut12_10[0] , 
        \nScanOut142[7] , \nOut12_13[3] , \nScanOut221[1] , \nScanOut222[2] , 
        \nScanOut190[1] , \nScanOut8[3] , \nScanOut43[4] , \nOut4_10[0] , 
        \nScanOut104[2] , \nScanOut61[5] , \nOut4_13[3] , \nScanOut107[1] , 
        \nScanOut160[6] , \nScanOut200[3] , \nOut13_10[4] , \nScanOut62[6] , 
        \nScanOut163[5] , \nOut13_13[7] , \nScanOut203[0] , \nOut2_1[5] , 
        \nOut1_5[4] , \nOut7_5[0] , \nOut14_5[5] , \nOut1_6[7] , \nOut7_6[3] , 
        \nOut12_5[1] , \nOut12_6[2] , \nOut14_6[6] , \nOut11_1[0] , 
        \nOut2_2[6] , \nOut4_1[1] , \nOut8_3[3] , \nOut8_0[0] , 
        \nScanOut178[4] , \nScanOut218[1] , \nOut4_2[2] , \nScanOut79[7] , 
        \nOut11_2[3] , \nScanOut39[5] , \nOut0_3[5] , \nScanOut5[6] , 
        \nScanOut6[5] , \nScanOut21[7] , \nScanOut22[4] , \nOut1_10[3] , 
        \nOut1_13[0] , \nScanOut138[6] , \nOut3_9[2] , \nScanOut46[0] , 
        \nOut5_9[6] , \nScanOut45[3] , \nScanOut94[6] , \nOut10_9[7] , 
        \nScanOut195[5] , \nScanOut227[6] , \nScanOut97[5] , \nOut9_8[7] , 
        \nScanOut147[3] , \nScanOut144[0] , \nOut12_15[4] , \nScanOut224[5] , 
        \nScanOut123[7] , \nScanOut196[6] , \nScanOut243[2] , \nScanOut34[0] , 
        \nScanOut37[3] , \nOut5_15[0] , \nScanOut120[4] , \nScanOut240[1] , 
        \nScanOut136[0] , \nScanOut256[5] , \nScanOut53[7] , \nScanOut135[3] , 
        \nOut10_14[3] , \nScanOut255[6] , \nScanOut81[1] , \nScanOut180[2] , 
        \nScanOut232[1] , \nScanOut82[2] , \nScanOut152[4] , \nScanOut231[2] , 
        \nScanOut50[4] , \nScanOut151[7] , \nOut7_14[7] , \nScanOut183[1] , 
        \nOut13_3[0] , \nOut6_3[1] , \nOut9_14[3] , \nOut14_12[3] , 
        \nOut15_3[4] , \nOut0_4[6] , \nScanOut10[6] , \nOut2_14[4] , 
        \nOut3_4[7] , \nOut3_7[4] , \nOut3_12[7] , \nOut6_0[2] , \nOut13_0[3] , 
        \nOut14_11[0] , \nOut9_6[1] , \nScanOut149[5] , \nScanOut229[0] , 
        \nScanOut48[6] , \nOut5_7[0] , \nOut3_11[4] , \nOut5_4[3] , 
        \nOut10_7[1] , \nOut10_4[2] , \nScanOut99[3] , \nScanOut198[0] , 
        \nOut9_5[2] , \nScanOut74[2] , \nOut6_11[7] , \nScanOut109[7] , 
        \nOut8_11[3] , \nOut15_14[0] , \nOut8_12[0] , \nScanOut175[1] , 
        \nScanOut215[4] , \nScanOut77[1] , \nOut6_12[4] , \nOut11_11[3] , 
        \nScanOut176[2] , \nScanOut216[7] , \nScanOut13[5] , \nOut7_8[5] , 
        \nScanOut111[5] , \nScanOut112[6] , \nOut11_12[0] , \nOut12_8[4] , 
        \nOut14_8[0] , \nScanOut14[6] , \nScanOut17[5] , \nOut1_8[1] , 
        \nOut2_8[0] , \nOut11_8[5] , \nOut4_8[4] , \nScanOut73[1] , 
        \nScanOut70[2] , \nOut6_15[7] , \nOut8_9[5] , \nScanOut171[1] , 
        \nScanOut172[2] , \nScanOut212[7] , \nScanOut211[4] , \nScanOut116[6] , 
        \nOut11_15[3] , \nOut2_10[4] , \nOut2_13[7] , \nScanOut115[5] , 
        \nScanOut169[3] , \nScanOut209[6] , \nScanOut68[0] , \nOut9_10[3] , 
        \nOut8_15[3] , \nOut15_13[3] , \nOut15_10[0] , \nOut13_4[3] , 
        \nOut0_7[5] , \nOut6_4[2] , \nOut15_4[7] , \nOut14_15[0] , 
        \nScanOut28[2] , \nScanOut30[0] , \nOut3_3[4] , \nOut3_0[7] , 
        \nOut3_15[4] , \nOut6_7[1] , \nOut13_7[0] , \nOut15_7[4] , 
        \nScanOut129[1] , \nOut9_13[0] , \nScanOut249[4] , \nOut5_0[3] , 
        \nOut5_3[0] , \nOut9_1[2] , \nOut10_0[2] , \nOut9_2[1] , \nOut10_3[1] , 
        \nScanOut33[3] , \nScanOut131[3] , \nOut10_10[3] , \nScanOut251[6] , 
        \nScanOut132[0] , \nScanOut252[5] , \nScanOut86[2] , \nOut10_13[0] , 
        \nScanOut1[6] , \nScanOut155[7] , \nScanOut235[2] , \nScanOut2[5] , 
        \nScanOut54[4] , \nScanOut57[7] , \nOut7_10[7] , \nOut7_13[4] , 
        \nScanOut187[1] , \nScanOut85[1] , \nScanOut184[2] , \nScanOut236[1] , 
        \nScanOut156[4] , \nScanOut9[7] , \nOut0_9[3] , \nScanOut25[7] , 
        \nScanOut41[3] , \nScanOut93[5] , \nScanOut220[5] , \nScanOut140[0] , 
        \nOut12_11[4] , \nScanOut42[0] , \nScanOut192[6] , \nScanOut90[6] , 
        \nScanOut191[5] , \nScanOut143[3] , \nScanOut223[6] , \nOut12_12[7] , 
        \nOut5_11[0] , \nOut5_12[3] , \nScanOut124[4] , \nScanOut244[1] , 
        \nScanOut127[7] , \nScanOut247[2] , \nOut0_11[3] , \nOut0_12[0] , 
        \nOut1_2[7] , \nScanOut26[4] , \nOut1_14[3] , \nScanOut59[1] , 
        \nScanOut88[4] , \nOut6_9[7] , \nOut13_9[6] , \nOut15_9[2] , 
        \nScanOut189[7] , \nScanOut158[2] , \nScanOut238[7] , \nOut7_2[3] , 
        \nOut14_2[6] , \nScanOut19[3] , \nOut12_2[2] , \nScanOut118[0] , 
        \nOut1_1[4] , \nOut7_1[0] , \nOut12_1[1] , \nOut14_1[5] , 
        \nScanOut20[3] , \nOut2_5[5] , \nOut2_6[6] , \nOut8_7[3] , 
        \nOut11_6[3] , \nOut4_6[2] , \nScanOut23[0] , \nOut4_5[1] , 
        \nOut11_5[0] , \nOut4_14[0] , \nScanOut100[2] , \nScanOut103[1] , 
        \nOut8_4[0] , \nScanOut65[5] , \nScanOut66[6] , \nScanOut164[6] , 
        \nScanOut167[5] , \nScanOut207[0] , \nScanOut204[3] , \nOut13_14[4] , 
        \nOut5_14[4] , \nScanOut121[0] , \nScanOut122[3] , \nScanOut242[6] , 
        \nScanOut241[5] , \nOut1_11[7] , \nOut1_12[4] , \nOut3_8[6] , 
        \nScanOut95[2] , \nOut9_9[3] , \nScanOut146[7] , \nOut10_8[3] , 
        \nScanOut226[2] , \nScanOut44[7] , \nScanOut47[4] , \nOut5_8[2] , 
        \nScanOut194[1] , \nScanOut197[2] , \nScanOut96[1] , \nScanOut145[4] , 
        \nOut12_14[0] , \nScanOut225[1] , \nScanOut139[2] , \nScanOut38[1] , 
        \nOut2_3[2] , \nOut2_0[1] , \nOut4_0[5] , \nOut8_1[4] , \nOut4_3[6] , 
        \nScanOut78[3] , \nOut11_0[4] , \nOut11_3[7] , \nOut8_2[7] , 
        \nScanOut219[5] , \nScanOut179[0] , \nOut12_4[5] , \nScanOut11[2] , 
        \nOut0_14[7] , \nOut1_4[0] , \nOut7_4[4] , \nOut14_4[1] , \nOut1_7[3] , 
        \nOut4_11[4] , \nScanOut60[1] , \nOut7_7[7] , \nOut12_7[6] , 
        \nOut14_7[2] , \nScanOut63[2] , \nScanOut161[2] , \nScanOut201[7] , 
        \nOut13_11[0] , \nScanOut162[1] , \nScanOut202[4] , \nOut13_12[3] , 
        \nOut4_12[7] , \nScanOut105[6] , \nScanOut106[5] , \nScanOut110[1] , 
        \nScanOut12[1] , \nOut1_9[5] , \nOut11_10[7] , \nScanOut75[6] , 
        \nOut7_9[1] , \nOut11_13[4] , \nOut12_9[0] , \nOut14_9[4] , 
        \nScanOut113[2] , \nScanOut76[5] , \nOut6_10[3] , \nOut6_13[0] , 
        \nScanOut174[5] , \nScanOut214[0] , \nScanOut177[6] , \nScanOut217[3] , 
        \nOut8_10[7] , \nScanOut108[3] , \nOut8_13[4] , \nScanOut1[2] , 
        \nOut0_1[2] , \nOut0_2[1] , \nOut3_5[3] , \nOut3_6[0] , \nOut2_15[0] , 
        \nOut10_6[5] , \nOut3_13[3] , \nScanOut49[2] , \nOut5_6[4] , 
        \nScanOut98[7] , \nOut9_4[6] , \nOut9_7[5] , \nScanOut148[1] , 
        \nScanOut228[4] , \nOut3_10[0] , \nOut10_5[6] , \nScanOut199[4] , 
        \nOut5_5[7] , \nOut6_2[5] , \nOut14_13[7] , \nOut15_2[0] , 
        \nOut6_1[6] , \nOut13_2[4] , \nOut13_1[7] , \nOut14_10[4] , 
        \nOut15_1[3] , \nScanOut2[1] , \nScanOut4[2] , \nScanOut7[1] , 
        \nScanOut153[0] , \nOut9_15[7] , \nScanOut51[0] , \nScanOut52[3] , 
        \nScanOut80[5] , \nScanOut233[5] , \nScanOut181[6] , \nOut7_15[3] , 
        \nScanOut182[5] , \nScanOut150[3] , \nOut0_9[7] , \nOut0_11[7] , 
        \nOut1_1[0] , \nScanOut35[4] , \nScanOut36[7] , \nScanOut83[6] , 
        \nScanOut230[6] , \nScanOut134[7] , \nScanOut137[4] , \nOut10_15[7] , 
        \nScanOut254[2] , \nOut4_14[4] , \nScanOut65[1] , \nScanOut100[6] , 
        \nScanOut103[5] , \nScanOut66[2] , \nScanOut164[2] , \nScanOut204[7] , 
        \nScanOut167[1] , \nOut13_14[0] , \nScanOut207[4] , \nOut7_1[4] , 
        \nOut12_1[5] , \nOut14_1[1] , \nOut0_12[4] , \nOut1_2[3] , 
        \nScanOut19[7] , \nScanOut118[4] , \nOut12_2[6] , \nOut2_5[1] , 
        \nOut4_5[5] , \nOut7_2[7] , \nOut8_4[4] , \nOut14_2[2] , \nOut11_5[4] , 
        \nOut2_6[2] , \nOut4_6[6] , \nScanOut26[0] , \nOut1_14[7] , 
        \nScanOut59[5] , \nOut8_7[7] , \nOut11_6[7] , \nScanOut88[0] , 
        \nScanOut158[6] , \nScanOut238[3] , \nScanOut189[3] , \nScanOut41[7] , 
        \nScanOut42[4] , \nScanOut90[2] , \nScanOut143[7] , \nOut12_12[3] , 
        \nScanOut223[2] , \nScanOut191[1] , \nScanOut192[2] , \nOut6_9[3] , 
        \nScanOut93[1] , \nScanOut140[4] , \nOut12_11[0] , \nScanOut220[1] , 
        \nOut15_9[6] , \nOut13_9[2] , \nScanOut25[3] , \nOut5_11[4] , 
        \nOut5_12[7] , \nScanOut127[3] , \nScanOut124[0] , \nScanOut247[6] , 
        \nScanOut244[5] , \nScanOut30[4] , \nScanOut33[7] , \nOut10_13[4] , 
        \nScanOut131[7] , \nScanOut132[4] , \nScanOut252[1] , \nOut10_10[7] , 
        \nScanOut251[2] , \nScanOut156[0] , \nScanOut54[0] , \nScanOut57[3] , 
        \nScanOut85[5] , \nOut7_13[0] , \nScanOut184[6] , \nScanOut236[5] , 
        \nScanOut187[5] , \nOut7_10[3] , \nScanOut155[3] , \nOut0_4[2] , 
        \nOut0_7[1] , \nScanOut28[6] , \nScanOut86[6] , \nScanOut235[6] , 
        \nOut6_7[5] , \nScanOut129[5] , \nOut9_13[4] , \nScanOut249[0] , 
        \nOut15_7[0] , \nOut13_7[4] , \nOut6_4[6] , \nOut15_4[3] , 
        \nOut14_15[4] , \nScanOut14[2] , \nOut2_8[4] , \nOut2_10[0] , 
        \nOut3_3[0] , \nOut9_10[7] , \nOut13_4[7] , \nOut3_0[3] , \nOut5_3[4] , 
        \nOut10_3[5] , \nOut9_1[6] , \nOut9_2[5] , \nOut10_0[6] , 
        \nOut3_15[0] , \nOut5_0[7] , \nOut2_13[3] , \nScanOut68[4] , 
        \nOut4_8[0] , \nScanOut70[6] , \nOut6_15[3] , \nOut8_15[7] , 
        \nScanOut169[7] , \nScanOut209[2] , \nOut15_10[4] , \nOut15_13[7] , 
        \nScanOut73[5] , \nOut8_9[1] , \nScanOut171[5] , \nScanOut211[0] , 
        \nScanOut172[6] , \nScanOut212[3] , \nScanOut115[1] , \nOut11_8[1] , 
        \nScanOut17[1] , \nOut11_15[7] , \nOut0_1[6] , \nScanOut4[6] , 
        \nScanOut83[2] , \nScanOut116[2] , \nScanOut230[2] , \nScanOut150[7] , 
        \nScanOut7[5] , \nScanOut51[4] , \nOut7_15[7] , \nScanOut52[7] , 
        \nScanOut182[1] , \nScanOut80[1] , \nScanOut181[2] , \nScanOut153[4] , 
        \nScanOut233[1] , \nScanOut35[0] , \nScanOut36[3] , \nScanOut134[3] , 
        \nOut10_15[3] , \nScanOut254[6] , \nScanOut137[0] , \nOut3_5[7] , 
        \nOut3_10[4] , \nOut5_5[3] , \nOut10_5[2] , \nOut3_6[4] , 
        \nOut3_13[7] , \nScanOut98[3] , \nScanOut199[0] , \nOut9_4[2] , 
        \nOut9_7[1] , \nScanOut148[5] , \nScanOut228[0] , \nScanOut49[6] , 
        \nOut5_6[0] , \nOut10_6[1] , \nOut9_15[3] , \nOut0_2[5] , \nOut6_1[2] , 
        \nOut13_1[3] , \nOut14_10[0] , \nOut15_1[7] , \nOut13_2[0] , 
        \nOut6_2[1] , \nScanOut108[7] , \nOut14_13[3] , \nOut15_2[4] , 
        \nOut8_13[0] , \nOut2_15[4] , \nOut8_10[3] , \nScanOut11[6] , 
        \nScanOut12[5] , \nOut7_9[5] , \nScanOut113[6] , \nOut11_13[0] , 
        \nOut12_9[4] , \nOut14_9[0] , \nOut1_9[1] , \nOut11_10[3] , 
        \nOut0_14[3] , \nOut2_3[6] , \nOut4_11[0] , \nScanOut60[5] , 
        \nScanOut63[6] , \nScanOut75[2] , \nScanOut76[1] , \nOut6_13[4] , 
        \nScanOut110[5] , \nScanOut174[1] , \nScanOut177[2] , \nScanOut217[7] , 
        \nScanOut214[4] , \nOut6_10[7] , \nScanOut161[6] , \nScanOut162[5] , 
        \nScanOut202[0] , \nOut13_12[7] , \nOut13_11[4] , \nScanOut201[3] , 
        \nOut4_12[3] , \nScanOut106[1] , \nScanOut105[2] , \nOut8_2[3] , 
        \nScanOut179[4] , \nScanOut219[1] , \nOut1_7[7] , \nOut2_0[5] , 
        \nOut4_3[2] , \nScanOut78[7] , \nOut11_3[3] , \nOut11_0[0] , 
        \nOut4_0[1] , \nOut7_7[3] , \nOut8_1[0] , \nOut12_7[2] , \nOut14_7[6] , 
        \nOut1_4[4] , \nOut7_4[0] , \nOut14_4[5] , \nOut12_4[1] , 
        \nScanOut9[3] , \nOut1_11[3] , \nOut1_12[0] , \nScanOut38[5] , 
        \nScanOut139[6] , \nOut1_4[6] , \nOut2_3[4] , \nScanOut20[7] , 
        \nScanOut23[4] , \nOut5_14[0] , \nScanOut121[4] , \nScanOut241[1] , 
        \nScanOut122[7] , \nScanOut242[2] , \nOut2_0[7] , \nOut3_8[2] , 
        \nScanOut44[3] , \nScanOut96[5] , \nScanOut145[0] , \nScanOut225[5] , 
        \nOut12_14[4] , \nScanOut47[0] , \nOut5_8[6] , \nScanOut197[6] , 
        \nOut4_11[2] , \nScanOut60[7] , \nScanOut95[6] , \nOut10_8[7] , 
        \nScanOut194[5] , \nScanOut226[6] , \nOut9_9[7] , \nScanOut146[3] , 
        \nScanOut63[4] , \nScanOut161[4] , \nScanOut201[1] , \nOut13_11[6] , 
        \nScanOut162[7] , \nScanOut202[2] , \nOut13_12[5] , \nOut4_12[1] , 
        \nScanOut105[0] , \nOut4_0[3] , \nScanOut106[3] , \nOut8_1[2] , 
        \nOut11_0[2] , \nOut4_3[0] , \nScanOut78[5] , \nOut8_2[1] , 
        \nOut11_3[1] , \nScanOut179[6] , \nScanOut219[3] , \nOut0_1[4] , 
        \nOut0_2[7] , \nScanOut4[4] , \nScanOut7[7] , \nScanOut9[1] , 
        \nOut0_14[1] , \nOut7_4[2] , \nOut12_4[3] , \nOut14_4[7] , 
        \nOut1_7[5] , \nOut12_7[0] , \nOut1_11[1] , \nOut1_12[2] , 
        \nOut7_7[1] , \nScanOut139[4] , \nOut14_7[4] , \nScanOut38[7] , 
        \nScanOut20[5] , \nScanOut23[6] , \nOut5_14[2] , \nScanOut121[6] , 
        \nScanOut122[5] , \nScanOut242[0] , \nScanOut241[3] , \nOut3_8[0] , 
        \nScanOut95[4] , \nOut9_9[5] , \nScanOut146[1] , \nScanOut226[4] , 
        \nScanOut194[7] , \nScanOut44[1] , \nScanOut47[2] , \nOut10_8[5] , 
        \nOut5_8[4] , \nScanOut197[4] , \nScanOut96[7] , \nScanOut145[2] , 
        \nOut12_14[6] , \nScanOut225[7] , \nScanOut51[6] , \nScanOut52[5] , 
        \nScanOut80[3] , \nScanOut153[6] , \nScanOut181[0] , \nScanOut233[3] , 
        \nOut7_15[5] , \nScanOut182[3] , \nScanOut35[2] , \nScanOut36[1] , 
        \nScanOut83[0] , \nScanOut150[5] , \nScanOut230[0] , \nScanOut134[1] , 
        \nScanOut137[2] , \nOut10_15[1] , \nScanOut254[4] , \nOut3_5[5] , 
        \nOut3_6[6] , \nOut3_13[5] , \nOut10_6[3] , \nScanOut49[4] , 
        \nOut5_6[2] , \nScanOut98[1] , \nOut9_4[0] , \nOut9_7[3] , 
        \nScanOut148[7] , \nScanOut228[2] , \nOut10_5[0] , \nScanOut199[2] , 
        \nOut3_10[6] , \nOut5_5[1] , \nOut6_2[3] , \nOut13_2[2] , 
        \nOut14_13[1] , \nOut15_2[6] , \nOut6_1[0] , \nOut14_10[2] , 
        \nOut15_1[5] , \nOut8_10[1] , \nOut9_15[1] , \nOut13_1[1] , 
        \nScanOut108[5] , \nOut8_13[2] , \nScanOut1[0] , \nScanOut11[4] , 
        \nOut2_15[6] , \nScanOut110[7] , \nScanOut12[7] , \nOut11_10[1] , 
        \nOut1_9[3] , \nOut12_9[6] , \nScanOut30[6] , \nScanOut75[0] , 
        \nOut7_9[7] , \nScanOut113[4] , \nOut11_13[2] , \nOut14_9[2] , 
        \nScanOut76[3] , \nOut6_10[5] , \nOut6_13[6] , \nScanOut174[3] , 
        \nScanOut214[6] , \nScanOut177[0] , \nScanOut217[5] , \nScanOut33[5] , 
        \nScanOut131[5] , \nOut10_10[5] , \nScanOut251[0] , \nScanOut132[6] , 
        \nScanOut252[3] , \nScanOut86[4] , \nOut10_13[6] , \nScanOut235[4] , 
        \nScanOut2[3] , \nScanOut54[2] , \nScanOut155[1] , \nScanOut57[1] , 
        \nOut7_10[1] , \nOut7_13[2] , \nScanOut187[7] , \nScanOut85[7] , 
        \nScanOut184[4] , \nScanOut236[7] , \nOut0_4[0] , \nOut9_10[5] , 
        \nScanOut156[2] , \nOut0_7[3] , \nScanOut28[4] , \nOut6_4[4] , 
        \nOut13_4[5] , \nOut15_4[1] , \nOut14_15[6] , \nOut13_7[6] , 
        \nOut2_8[6] , \nOut2_10[2] , \nOut2_13[1] , \nOut3_3[2] , \nOut3_0[1] , 
        \nOut3_15[2] , \nOut5_0[5] , \nOut6_7[7] , \nScanOut129[7] , 
        \nOut9_13[6] , \nOut15_7[2] , \nScanOut249[2] , \nOut10_0[4] , 
        \nOut5_3[6] , \nOut9_1[4] , \nOut9_2[7] , \nScanOut68[6] , 
        \nOut10_3[7] , \nScanOut169[5] , \nScanOut209[0] , \nOut8_15[5] , 
        \nOut15_13[5] , \nOut15_10[6] , \nOut4_8[2] , \nOut11_8[3] , 
        \nScanOut73[7] , \nScanOut14[0] , \nScanOut17[3] , \nScanOut70[4] , 
        \nOut6_15[1] , \nOut8_9[3] , \nScanOut172[4] , \nScanOut171[7] , 
        \nScanOut212[1] , \nScanOut211[2] , \nScanOut116[0] , \nOut11_15[5] , 
        \nScanOut103[7] , \nScanOut115[3] , \nOut0_9[5] , \nOut0_11[5] , 
        \nOut0_12[6] , \nOut1_2[1] , \nScanOut19[5] , \nOut4_14[6] , 
        \nScanOut100[4] , \nScanOut65[3] , \nScanOut66[0] , \nScanOut164[0] , 
        \nScanOut167[3] , \nScanOut207[6] , \nScanOut204[5] , \nOut13_14[2] , 
        \nOut7_2[5] , \nOut12_2[4] , \nOut14_2[0] , \nScanOut118[6] , 
        \nEnable[0] , \nOut1_1[2] , \nOut7_1[6] , \nOut14_1[3] , \nOut2_5[3] , 
        \nOut2_6[0] , \nOut8_7[5] , \nOut12_1[7] , \nOut4_6[4] , \nOut11_6[5] , 
        \nOut11_5[6] , \nOut4_5[7] , \nOut8_4[6] , \nScanOut25[1] , 
        \nOut1_14[5] , \nScanOut59[7] , \nScanOut88[2] , \nScanOut189[1] , 
        \nScanOut158[4] , \nScanOut238[1] , \nScanOut41[5] , \nScanOut93[3] , 
        \nScanOut140[6] , \nOut12_11[2] , \nScanOut220[3] , \nScanOut42[6] , 
        \nScanOut192[0] , \nScanOut90[0] , \nScanOut191[3] , \nScanOut223[0] , 
        \nScanOut143[5] , \nOut12_12[1] , \nScanOut26[2] , \nOut5_11[6] , 
        \nScanOut244[7] , \nOut5_12[5] , \nScanOut124[2] , \nScanOut247[4] , 
        \nScanOut127[1] , \nOut13_9[0] , \nScanOut11[0] , \nScanOut12[3] , 
        \nOut1_9[7] , \nOut6_9[1] , \nOut7_9[3] , \nScanOut113[0] , 
        \nOut15_9[4] , \nOut14_9[6] , \nOut11_13[6] , \nOut12_9[2] , 
        \nOut11_10[5] , \nScanOut75[4] , \nScanOut76[7] , \nOut6_13[2] , 
        \nScanOut110[3] , \nScanOut174[7] , \nScanOut177[4] , \nScanOut217[1] , 
        \nScanOut214[2] , \nOut6_10[1] , \nScanOut108[1] , \nOut8_13[6] , 
        \nOut2_15[2] , \nOut8_10[5] , \nOut0_1[0] , \nOut3_5[1] , 
        \nOut3_10[2] , \nOut5_5[5] , \nScanOut199[6] , \nOut3_6[2] , 
        \nOut3_13[1] , \nScanOut49[0] , \nScanOut98[5] , \nOut10_5[4] , 
        \nOut9_4[4] , \nOut9_7[7] , \nScanOut228[6] , \nScanOut148[3] , 
        \nOut5_6[6] , \nOut10_6[7] , \nOut9_15[5] , \nOut13_1[5] , 
        \nOut0_2[3] , \nOut6_1[4] , \nOut14_10[6] , \nOut15_1[1] , 
        \nScanOut4[0] , \nOut6_2[7] , \nOut13_2[6] , \nOut14_13[5] , 
        \nOut15_2[2] , \nScanOut83[4] , \nScanOut230[4] , \nScanOut7[3] , 
        \nScanOut51[2] , \nOut7_15[1] , \nScanOut150[1] , \nScanOut52[1] , 
        \nScanOut182[7] , \nScanOut80[7] , \nScanOut181[4] , \nScanOut233[7] , 
        \nScanOut9[5] , \nScanOut20[1] , \nScanOut35[6] , \nScanOut153[2] , 
        \nScanOut36[5] , \nScanOut134[5] , \nOut10_15[5] , \nScanOut254[0] , 
        \nScanOut137[6] , \nScanOut23[2] , \nOut5_14[6] , \nScanOut241[7] , 
        \nScanOut121[2] , \nScanOut122[1] , \nScanOut242[4] , \nOut1_11[5] , 
        \nOut3_8[4] , \nScanOut44[5] , \nScanOut96[3] , \nScanOut225[3] , 
        \nScanOut145[6] , \nOut12_14[2] , \nScanOut47[6] , \nScanOut197[0] , 
        \nOut5_8[0] , \nOut10_8[1] , \nScanOut194[3] , \nScanOut95[0] , 
        \nOut9_9[1] , \nScanOut226[0] , \nScanOut146[5] , \nOut1_12[6] , 
        \nScanOut38[3] , \nScanOut139[0] , \nOut0_14[5] , \nOut2_3[0] , 
        \nOut8_2[5] , \nOut11_3[5] , \nScanOut179[2] , \nScanOut219[7] , 
        \nOut1_7[1] , \nOut2_0[3] , \nOut4_3[4] , \nScanOut78[1] , 
        \nOut4_0[7] , \nOut11_0[6] , \nOut7_7[5] , \nOut8_1[6] , \nOut14_7[0] , 
        \nOut12_7[4] , \nOut7_4[6] , \nOut14_4[3] , \nScanOut1[4] , 
        \nScanOut2[7] , \nOut0_4[4] , \nOut0_7[7] , \nOut0_9[1] , \nOut1_4[2] , 
        \nOut12_4[7] , \nScanOut41[1] , \nScanOut42[2] , \nOut4_11[6] , 
        \nScanOut60[3] , \nScanOut63[0] , \nScanOut161[0] , \nScanOut162[3] , 
        \nScanOut202[6] , \nOut13_12[1] , \nOut13_11[2] , \nScanOut201[5] , 
        \nOut4_12[5] , \nScanOut106[7] , \nScanOut105[4] , \nScanOut90[4] , 
        \nScanOut143[1] , \nOut12_12[5] , \nScanOut191[7] , \nScanOut223[4] , 
        \nScanOut192[4] , \nOut6_9[5] , \nScanOut93[7] , \nScanOut140[2] , 
        \nOut12_11[6] , \nScanOut220[7] , \nOut15_9[0] , \nOut0_11[1] , 
        \nOut1_1[6] , \nScanOut25[5] , \nScanOut26[6] , \nOut13_9[4] , 
        \nOut5_11[2] , \nOut5_12[1] , \nScanOut127[5] , \nScanOut247[0] , 
        \nScanOut124[6] , \nScanOut244[3] , \nOut1_14[1] , \nScanOut59[3] , 
        \nScanOut88[6] , \nScanOut158[0] , \nScanOut238[5] , \nScanOut189[5] , 
        \nOut12_1[3] , \nOut7_1[2] , \nOut14_1[7] , \nOut0_12[2] , 
        \nScanOut14[4] , \nOut1_2[5] , \nScanOut118[2] , \nScanOut19[1] , 
        \nOut2_5[7] , \nOut4_5[3] , \nOut7_2[1] , \nOut12_2[0] , \nOut14_2[4] , 
        \nOut8_4[2] , \nOut2_6[4] , \nOut4_6[0] , \nOut11_5[2] , \nOut11_6[1] , 
        \nOut2_8[2] , \nOut4_8[6] , \nOut4_14[2] , \nOut8_7[1] , 
        \nScanOut65[7] , \nScanOut100[0] , \nScanOut103[3] , \nScanOut66[4] , 
        \nScanOut164[4] , \nScanOut204[1] , \nScanOut167[7] , \nOut13_14[6] , 
        \nScanOut207[2] , \nScanOut70[0] , \nOut6_15[5] , \nOut8_9[7] , 
        \nScanOut171[3] , \nScanOut211[6] , \nScanOut212[5] , \nScanOut172[0] , 
        \nScanOut73[3] , \nOut11_8[7] , \nScanOut115[7] , \nScanOut17[7] , 
        \nOut11_15[1] , \nOut2_10[6] , \nScanOut116[4] , \nOut2_13[5] , 
        \nScanOut68[2] , \nOut6_7[3] , \nScanOut129[3] , \nOut8_15[1] , 
        \nScanOut169[1] , \nScanOut209[4] , \nOut15_10[2] , \nOut15_13[1] , 
        \nOut9_13[2] , \nScanOut249[6] , \nOut15_7[6] , \nScanOut28[0] , 
        \nOut13_7[2] , \nOut6_4[0] , \nOut13_4[1] , \nOut15_4[5] , 
        \nOut14_15[2] , \nScanOut30[2] , \nScanOut33[1] , \nOut3_3[6] , 
        \nOut9_10[1] , \nOut10_3[3] , \nOut3_0[5] , \nOut5_3[2] , \nOut9_1[0] , 
        \nOut9_2[3] , \nOut3_15[6] , \nOut10_0[0] , \nOut5_0[1] , 
        \nOut10_13[2] , \nScanOut131[1] , \nScanOut132[2] , \nScanOut252[7] , 
        \nOut10_10[1] , \nScanOut251[4] , \nScanOut54[6] , \nScanOut57[5] , 
        \nScanOut85[3] , \nScanOut156[6] , \nScanOut236[3] , \nOut7_13[6] , 
        \nScanOut184[0] , \nScanOut187[3] , \nOut7_10[5] , \nScanOut86[0] , 
        \nScanOut155[5] , \nScanOut235[0] ;
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_19 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut20[7] , \nScanOut20[6] , 
        \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , 
        \nScanOut20[1] , \nScanOut20[0] }), .ScanOut({\nScanOut19[7] , 
        \nScanOut19[6] , \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , 
        \nScanOut19[2] , \nScanOut19[1] , \nScanOut19[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , 
        \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), .SouthIn({\nOut1_4[7] , 
        \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , 
        \nOut1_4[1] , \nOut1_4[0] }), .EastIn({\nOut2_3[7] , \nOut2_3[6] , 
        \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , 
        \nOut2_3[0] }), .WestIn({\nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , 
        \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), 
        .Out({\nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , 
        \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_25 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut26[7] , \nScanOut26[6] , 
        \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , 
        \nScanOut26[1] , \nScanOut26[0] }), .ScanOut({\nScanOut25[7] , 
        \nScanOut25[6] , \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , 
        \nScanOut25[2] , \nScanOut25[1] , \nScanOut25[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , 
        \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), .SouthIn({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .EastIn({\nOut2_9[7] , 
        \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , 
        \nOut2_9[1] , \nOut2_9[0] }), .WestIn({\nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }), .Out({\nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , 
        \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_89 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut90[7] , \nScanOut90[6] , 
        \nScanOut90[5] , \nScanOut90[4] , \nScanOut90[3] , \nScanOut90[2] , 
        \nScanOut90[1] , \nScanOut90[0] }), .ScanOut({\nScanOut89[7] , 
        \nScanOut89[6] , \nScanOut89[5] , \nScanOut89[4] , \nScanOut89[3] , 
        \nScanOut89[2] , \nScanOut89[1] , \nScanOut89[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , 
        \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }), .SouthIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .EastIn({\nOut6_9[7] , 
        \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , 
        \nOut6_9[1] , \nOut6_9[0] }), .WestIn({\nOut4_9[7] , \nOut4_9[6] , 
        \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , \nOut4_9[1] , 
        \nOut4_9[0] }), .Out({\nOut5_9[7] , \nOut5_9[6] , \nOut5_9[5] , 
        \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , \nOut5_9[1] , \nOut5_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_50 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut51[7] , \nScanOut51[6] , 
        \nScanOut51[5] , \nScanOut51[4] , \nScanOut51[3] , \nScanOut51[2] , 
        \nScanOut51[1] , \nScanOut51[0] }), .ScanOut({\nScanOut50[7] , 
        \nScanOut50[6] , \nScanOut50[5] , \nScanOut50[4] , \nScanOut50[3] , 
        \nScanOut50[2] , \nScanOut50[1] , \nScanOut50[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , 
        \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }), .SouthIn({\nOut3_3[7] , 
        \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , 
        \nOut3_3[1] , \nOut3_3[0] }), .EastIn({\nOut4_2[7] , \nOut4_2[6] , 
        \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , 
        \nOut4_2[0] }), .WestIn({\nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , 
        \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), 
        .Out({\nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , 
        \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_154 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut155[7] , \nScanOut155[6] , 
        \nScanOut155[5] , \nScanOut155[4] , \nScanOut155[3] , \nScanOut155[2] , 
        \nScanOut155[1] , \nScanOut155[0] }), .ScanOut({\nScanOut154[7] , 
        \nScanOut154[6] , \nScanOut154[5] , \nScanOut154[4] , \nScanOut154[3] , 
        \nScanOut154[2] , \nScanOut154[1] , \nScanOut154[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_9[7] , \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , 
        \nOut9_9[2] , \nOut9_9[1] , \nOut9_9[0] }), .SouthIn({\nOut9_11[7] , 
        \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , \nOut9_11[3] , 
        \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .EastIn({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), .WestIn({
        \nOut8_10[7] , \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , 
        \nOut8_10[3] , \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .Out({
        \nOut9_10[7] , \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , 
        \nOut9_10[3] , \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_173 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut174[7] , \nScanOut174[6] , 
        \nScanOut174[5] , \nScanOut174[4] , \nScanOut174[3] , \nScanOut174[2] , 
        \nScanOut174[1] , \nScanOut174[0] }), .ScanOut({\nScanOut173[7] , 
        \nScanOut173[6] , \nScanOut173[5] , \nScanOut173[4] , \nScanOut173[3] , 
        \nScanOut173[2] , \nScanOut173[1] , \nScanOut173[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , 
        \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), 
        .SouthIn({\nOut10_14[7] , \nOut10_14[6] , \nOut10_14[5] , 
        \nOut10_14[4] , \nOut10_14[3] , \nOut10_14[2] , \nOut10_14[1] , 
        \nOut10_14[0] }), .EastIn({\nOut11_13[7] , \nOut11_13[6] , 
        \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , \nOut11_13[2] , 
        \nOut11_13[1] , \nOut11_13[0] }), .WestIn({\nOut9_13[7] , 
        \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , \nOut9_13[3] , 
        \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .Out({\nOut10_13[7] , 
        \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , \nOut10_13[3] , 
        \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_196 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut197[7] , \nScanOut197[6] , 
        \nScanOut197[5] , \nScanOut197[4] , \nScanOut197[3] , \nScanOut197[2] , 
        \nScanOut197[1] , \nScanOut197[0] }), .ScanOut({\nScanOut196[7] , 
        \nScanOut196[6] , \nScanOut196[5] , \nScanOut196[4] , \nScanOut196[3] , 
        \nScanOut196[2] , \nScanOut196[1] , \nScanOut196[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), 
        .SouthIn({\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .EastIn(
        {\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .WestIn(
        {\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .Out({
        \nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }) );
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 U_Jacobi_Control ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanOut({\nScanOut256[7] , 
        \nScanOut256[6] , \nScanOut256[5] , \nScanOut256[4] , \nScanOut256[3] , 
        \nScanOut256[2] , \nScanOut256[1] , \nScanOut256[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b1), .ScanId(1'b0), .Enable(\nEnable[0] ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_243 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut244[7] , \nScanOut244[6] , 
        \nScanOut244[5] , \nScanOut244[4] , \nScanOut244[3] , \nScanOut244[2] , 
        \nScanOut244[1] , \nScanOut244[0] }), .ScanOut({\nScanOut243[7] , 
        \nScanOut243[6] , \nScanOut243[5] , \nScanOut243[4] , \nScanOut243[3] , 
        \nScanOut243[2] , \nScanOut243[1] , \nScanOut243[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_3[7] , \nOut15_3[6] , 
        \nOut15_3[5] , \nOut15_3[4] , \nOut15_3[3] , \nOut15_3[2] , 
        \nOut15_3[1] , \nOut15_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_168 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut169[7] , \nScanOut169[6] , 
        \nScanOut169[5] , \nScanOut169[4] , \nScanOut169[3] , \nScanOut169[2] , 
        \nScanOut169[1] , \nScanOut169[0] }), .ScanOut({\nScanOut168[7] , 
        \nScanOut168[6] , \nScanOut168[5] , \nScanOut168[4] , \nScanOut168[3] , 
        \nScanOut168[2] , \nScanOut168[1] , \nScanOut168[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), 
        .SouthIn({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), .EastIn(
        {\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .WestIn(
        {\nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , 
        \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] }), .Out({\nOut10_8[7] , 
        \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , \nOut10_8[3] , 
        \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_77 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut78[7] , \nScanOut78[6] , 
        \nScanOut78[5] , \nScanOut78[4] , \nScanOut78[3] , \nScanOut78[2] , 
        \nScanOut78[1] , \nScanOut78[0] }), .ScanOut({\nScanOut77[7] , 
        \nScanOut77[6] , \nScanOut77[5] , \nScanOut77[4] , \nScanOut77[3] , 
        \nScanOut77[2] , \nScanOut77[1] , \nScanOut77[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), 
        .SouthIn({\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .EastIn(
        {\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .WestIn(
        {\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .Out({
        \nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_80 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut81[7] , \nScanOut81[6] , 
        \nScanOut81[5] , \nScanOut81[4] , \nScanOut81[3] , \nScanOut81[2] , 
        \nScanOut81[1] , \nScanOut81[0] }), .ScanOut({\nScanOut80[7] , 
        \nScanOut80[6] , \nScanOut80[5] , \nScanOut80[4] , \nScanOut80[3] , 
        \nScanOut80[2] , \nScanOut80[1] , \nScanOut80[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut5_0[7] , \nOut5_0[6] , 
        \nOut5_0[5] , \nOut5_0[4] , \nOut5_0[3] , \nOut5_0[2] , \nOut5_0[1] , 
        \nOut5_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_92 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut93[7] , \nScanOut93[6] , 
        \nScanOut93[5] , \nScanOut93[4] , \nScanOut93[3] , \nScanOut93[2] , 
        \nScanOut93[1] , \nScanOut93[0] }), .ScanOut({\nScanOut92[7] , 
        \nScanOut92[6] , \nScanOut92[5] , \nScanOut92[4] , \nScanOut92[3] , 
        \nScanOut92[2] , \nScanOut92[1] , \nScanOut92[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), 
        .SouthIn({\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .EastIn(
        {\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .WestIn(
        {\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .Out({
        \nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_236 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut237[7] , \nScanOut237[6] , 
        \nScanOut237[5] , \nScanOut237[4] , \nScanOut237[3] , \nScanOut237[2] , 
        \nScanOut237[1] , \nScanOut237[0] }), .ScanOut({\nScanOut236[7] , 
        \nScanOut236[6] , \nScanOut236[5] , \nScanOut236[4] , \nScanOut236[3] , 
        \nScanOut236[2] , \nScanOut236[1] , \nScanOut236[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_11[7] , \nOut14_11[6] , \nOut14_11[5] , \nOut14_11[4] , 
        \nOut14_11[3] , \nOut14_11[2] , \nOut14_11[1] , \nOut14_11[0] }), 
        .SouthIn({\nOut14_13[7] , \nOut14_13[6] , \nOut14_13[5] , 
        \nOut14_13[4] , \nOut14_13[3] , \nOut14_13[2] , \nOut14_13[1] , 
        \nOut14_13[0] }), .EastIn({\nOut15_12[7] , \nOut15_12[6] , 
        \nOut15_12[5] , \nOut15_12[4] , \nOut15_12[3] , \nOut15_12[2] , 
        \nOut15_12[1] , \nOut15_12[0] }), .WestIn({\nOut13_12[7] , 
        \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , 
        \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }), .Out({\nOut14_12[7] , 
        \nOut14_12[6] , \nOut14_12[5] , \nOut14_12[4] , \nOut14_12[3] , 
        \nOut14_12[2] , \nOut14_12[1] , \nOut14_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_106 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut107[7] , \nScanOut107[6] , 
        \nScanOut107[5] , \nScanOut107[4] , \nScanOut107[3] , \nScanOut107[2] , 
        \nScanOut107[1] , \nScanOut107[0] }), .ScanOut({\nScanOut106[7] , 
        \nScanOut106[6] , \nScanOut106[5] , \nScanOut106[4] , \nScanOut106[3] , 
        \nScanOut106[2] , \nScanOut106[1] , \nScanOut106[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_9[7] , \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , 
        \nOut6_9[2] , \nOut6_9[1] , \nOut6_9[0] }), .SouthIn({\nOut6_11[7] , 
        \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , \nOut6_11[3] , 
        \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .EastIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .WestIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .Out({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_121 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut122[7] , \nScanOut122[6] , 
        \nScanOut122[5] , \nScanOut122[4] , \nScanOut122[3] , \nScanOut122[2] , 
        \nScanOut122[1] , \nScanOut122[0] }), .ScanOut({\nScanOut121[7] , 
        \nScanOut121[6] , \nScanOut121[5] , \nScanOut121[4] , \nScanOut121[3] , 
        \nScanOut121[2] , \nScanOut121[1] , \nScanOut121[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , 
        \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }), .SouthIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .EastIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .WestIn({\nOut6_9[7] , \nOut6_9[6] , 
        \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , \nOut6_9[1] , 
        \nOut6_9[0] }), .Out({\nOut7_9[7] , \nOut7_9[6] , \nOut7_9[5] , 
        \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , \nOut7_9[1] , \nOut7_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_211 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut212[7] , \nScanOut212[6] , 
        \nScanOut212[5] , \nScanOut212[4] , \nScanOut212[3] , \nScanOut212[2] , 
        \nScanOut212[1] , \nScanOut212[0] }), .ScanOut({\nScanOut211[7] , 
        \nScanOut211[6] , \nScanOut211[5] , \nScanOut211[4] , \nScanOut211[3] , 
        \nScanOut211[2] , \nScanOut211[1] , \nScanOut211[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), 
        .SouthIn({\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .EastIn(
        {\nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), .WestIn(
        {\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .Out({
        \nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_224 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut225[7] , \nScanOut225[6] , 
        \nScanOut225[5] , \nScanOut225[4] , \nScanOut225[3] , \nScanOut225[2] , 
        \nScanOut225[1] , \nScanOut225[0] }), .ScanOut({\nScanOut224[7] , 
        \nScanOut224[6] , \nScanOut224[5] , \nScanOut224[4] , \nScanOut224[3] , 
        \nScanOut224[2] , \nScanOut224[1] , \nScanOut224[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut14_0[7] , \nOut14_0[6] , 
        \nOut14_0[5] , \nOut14_0[4] , \nOut14_0[3] , \nOut14_0[2] , 
        \nOut14_0[1] , \nOut14_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_114 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut115[7] , \nScanOut115[6] , 
        \nScanOut115[5] , \nScanOut115[4] , \nScanOut115[3] , \nScanOut115[2] , 
        \nScanOut115[1] , \nScanOut115[0] }), .ScanOut({\nScanOut114[7] , 
        \nScanOut114[6] , \nScanOut114[5] , \nScanOut114[4] , \nScanOut114[3] , 
        \nScanOut114[2] , \nScanOut114[1] , \nScanOut114[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , \nOut7_1[4] , \nOut7_1[3] , 
        \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }), .SouthIn({\nOut7_3[7] , 
        \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , 
        \nOut7_3[1] , \nOut7_3[0] }), .EastIn({\nOut8_2[7] , \nOut8_2[6] , 
        \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , 
        \nOut8_2[0] }), .WestIn({\nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , 
        \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }), 
        .Out({\nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , 
        \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1[7] , \nScanOut1[6] , 
        \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , 
        \nScanOut1[1] , \nScanOut1[0] }), .ScanOut({\nScanOut0[7] , 
        \nScanOut0[6] , \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , 
        \nScanOut0[2] , \nScanOut0[1] , \nScanOut0[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut3[7] , \nScanOut3[6] , 
        \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , 
        \nScanOut3[1] , \nScanOut3[0] }), .ScanOut({\nScanOut2[7] , 
        \nScanOut2[6] , \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , 
        \nScanOut2[2] , \nScanOut2[1] , \nScanOut2[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_2[7] , \nOut0_2[6] , 
        \nOut0_2[5] , \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , 
        \nOut0_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut4[7] , \nScanOut4[6] , 
        \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , 
        \nScanOut4[1] , \nScanOut4[0] }), .ScanOut({\nScanOut3[7] , 
        \nScanOut3[6] , \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , 
        \nScanOut3[2] , \nScanOut3[1] , \nScanOut3[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_3[7] , \nOut0_3[6] , 
        \nOut0_3[5] , \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , 
        \nOut0_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut5[7] , \nScanOut5[6] , 
        \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , 
        \nScanOut5[1] , \nScanOut5[0] }), .ScanOut({\nScanOut4[7] , 
        \nScanOut4[6] , \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , 
        \nScanOut4[2] , \nScanOut4[1] , \nScanOut4[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_4[7] , \nOut0_4[6] , 
        \nOut0_4[5] , \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , 
        \nOut0_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_133 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut134[7] , \nScanOut134[6] , 
        \nScanOut134[5] , \nScanOut134[4] , \nScanOut134[3] , \nScanOut134[2] , 
        \nScanOut134[1] , \nScanOut134[0] }), .ScanOut({\nScanOut133[7] , 
        \nScanOut133[6] , \nScanOut133[5] , \nScanOut133[4] , \nScanOut133[3] , 
        \nScanOut133[2] , \nScanOut133[1] , \nScanOut133[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_4[7] , \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , 
        \nOut8_4[2] , \nOut8_4[1] , \nOut8_4[0] }), .SouthIn({\nOut8_6[7] , 
        \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , 
        \nOut8_6[1] , \nOut8_6[0] }), .EastIn({\nOut9_5[7] , \nOut9_5[6] , 
        \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , \nOut9_5[1] , 
        \nOut9_5[0] }), .WestIn({\nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , 
        \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }), 
        .Out({\nOut8_5[7] , \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , 
        \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , \nOut8_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_203 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut204[7] , \nScanOut204[6] , 
        \nScanOut204[5] , \nScanOut204[4] , \nScanOut204[3] , \nScanOut204[2] , 
        \nScanOut204[1] , \nScanOut204[0] }), .ScanOut({\nScanOut203[7] , 
        \nScanOut203[6] , \nScanOut203[5] , \nScanOut203[4] , \nScanOut203[3] , 
        \nScanOut203[2] , \nScanOut203[1] , \nScanOut203[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_10[7] , \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , 
        \nOut12_10[3] , \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }), 
        .SouthIn({\nOut12_12[7] , \nOut12_12[6] , \nOut12_12[5] , 
        \nOut12_12[4] , \nOut12_12[3] , \nOut12_12[2] , \nOut12_12[1] , 
        \nOut12_12[0] }), .EastIn({\nOut13_11[7] , \nOut13_11[6] , 
        \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , \nOut13_11[2] , 
        \nOut13_11[1] , \nOut13_11[0] }), .WestIn({\nOut11_11[7] , 
        \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , 
        \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }), .Out({\nOut12_11[7] , 
        \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , 
        \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut11[7] , \nScanOut11[6] , 
        \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , 
        \nScanOut11[1] , \nScanOut11[0] }), .ScanOut({\nScanOut10[7] , 
        \nScanOut10[6] , \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , 
        \nScanOut10[2] , \nScanOut10[1] , \nScanOut10[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_10[7] , \nOut0_10[6] , 
        \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , \nOut0_10[2] , 
        \nOut0_10[1] , \nOut0_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_37 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut38[7] , \nScanOut38[6] , 
        \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , 
        \nScanOut38[1] , \nScanOut38[0] }), .ScanOut({\nScanOut37[7] , 
        \nScanOut37[6] , \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , 
        \nScanOut37[2] , \nScanOut37[1] , \nScanOut37[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , 
        \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), .SouthIn({\nOut2_6[7] , 
        \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , 
        \nOut2_6[1] , \nOut2_6[0] }), .EastIn({\nOut3_5[7] , \nOut3_5[6] , 
        \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , 
        \nOut3_5[0] }), .WestIn({\nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , 
        \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), 
        .Out({\nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , 
        \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_42 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut43[7] , \nScanOut43[6] , 
        \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , 
        \nScanOut43[1] , \nScanOut43[0] }), .ScanOut({\nScanOut42[7] , 
        \nScanOut42[6] , \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , 
        \nScanOut42[2] , \nScanOut42[1] , \nScanOut42[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_9[7] , \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , 
        \nOut2_9[2] , \nOut2_9[1] , \nOut2_9[0] }), .SouthIn({\nOut2_11[7] , 
        \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , \nOut2_11[3] , 
        \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .EastIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .WestIn({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .Out({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_59 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut60[7] , \nScanOut60[6] , 
        \nScanOut60[5] , \nScanOut60[4] , \nScanOut60[3] , \nScanOut60[2] , 
        \nScanOut60[1] , \nScanOut60[0] }), .ScanOut({\nScanOut59[7] , 
        \nScanOut59[6] , \nScanOut59[5] , \nScanOut59[4] , \nScanOut59[3] , 
        \nScanOut59[2] , \nScanOut59[1] , \nScanOut59[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_10[7] , \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , 
        \nOut3_10[3] , \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), 
        .SouthIn({\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .EastIn(
        {\nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .WestIn(
        {\nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .Out({
        \nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_65 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut66[7] , \nScanOut66[6] , 
        \nScanOut66[5] , \nScanOut66[4] , \nScanOut66[3] , \nScanOut66[2] , 
        \nScanOut66[1] , \nScanOut66[0] }), .ScanOut({\nScanOut65[7] , 
        \nScanOut65[6] , \nScanOut65[5] , \nScanOut65[4] , \nScanOut65[3] , 
        \nScanOut65[2] , \nScanOut65[1] , \nScanOut65[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_0[7] , \nOut4_0[6] , \nOut4_0[5] , \nOut4_0[4] , \nOut4_0[3] , 
        \nOut4_0[2] , \nOut4_0[1] , \nOut4_0[0] }), .SouthIn({\nOut4_2[7] , 
        \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , 
        \nOut4_2[1] , \nOut4_2[0] }), .EastIn({\nOut5_1[7] , \nOut5_1[6] , 
        \nOut5_1[5] , \nOut5_1[4] , \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , 
        \nOut5_1[0] }), .WestIn({\nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , 
        \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }), 
        .Out({\nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , \nOut4_1[4] , 
        \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_146 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut147[7] , \nScanOut147[6] , 
        \nScanOut147[5] , \nScanOut147[4] , \nScanOut147[3] , \nScanOut147[2] , 
        \nScanOut147[1] , \nScanOut147[0] }), .ScanOut({\nScanOut146[7] , 
        \nScanOut146[6] , \nScanOut146[5] , \nScanOut146[4] , \nScanOut146[3] , 
        \nScanOut146[2] , \nScanOut146[1] , \nScanOut146[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , 
        \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] }), .SouthIn({\nOut9_3[7] , 
        \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , 
        \nOut9_3[1] , \nOut9_3[0] }), .EastIn({\nOut10_2[7] , \nOut10_2[6] , 
        \nOut10_2[5] , \nOut10_2[4] , \nOut10_2[3] , \nOut10_2[2] , 
        \nOut10_2[1] , \nOut10_2[0] }), .WestIn({\nOut8_2[7] , \nOut8_2[6] , 
        \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , 
        \nOut8_2[0] }), .Out({\nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , 
        \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_161 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut162[7] , \nScanOut162[6] , 
        \nScanOut162[5] , \nScanOut162[4] , \nScanOut162[3] , \nScanOut162[2] , 
        \nScanOut162[1] , \nScanOut162[0] }), .ScanOut({\nScanOut161[7] , 
        \nScanOut161[6] , \nScanOut161[5] , \nScanOut161[4] , \nScanOut161[3] , 
        \nScanOut161[2] , \nScanOut161[1] , \nScanOut161[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_0[7] , \nOut10_0[6] , \nOut10_0[5] , \nOut10_0[4] , 
        \nOut10_0[3] , \nOut10_0[2] , \nOut10_0[1] , \nOut10_0[0] }), 
        .SouthIn({\nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), .EastIn(
        {\nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), .WestIn(
        {\nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , 
        \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] }), .Out({\nOut10_1[7] , 
        \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , \nOut10_1[3] , 
        \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_251 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut252[7] , \nScanOut252[6] , 
        \nScanOut252[5] , \nScanOut252[4] , \nScanOut252[3] , \nScanOut252[2] , 
        \nScanOut252[1] , \nScanOut252[0] }), .ScanOut({\nScanOut251[7] , 
        \nScanOut251[6] , \nScanOut251[5] , \nScanOut251[4] , \nScanOut251[3] , 
        \nScanOut251[2] , \nScanOut251[1] , \nScanOut251[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_11[7] , \nOut15_11[6] , 
        \nOut15_11[5] , \nOut15_11[4] , \nOut15_11[3] , \nOut15_11[2] , 
        \nOut15_11[1] , \nOut15_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_17 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut18[7] , \nScanOut18[6] , 
        \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , 
        \nScanOut18[1] , \nScanOut18[0] }), .ScanOut({\nScanOut17[7] , 
        \nScanOut17[6] , \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , 
        \nScanOut17[2] , \nScanOut17[1] , \nScanOut17[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_0[7] , \nOut1_0[6] , \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , 
        \nOut1_0[2] , \nOut1_0[1] , \nOut1_0[0] }), .SouthIn({\nOut1_2[7] , 
        \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , 
        \nOut1_2[1] , \nOut1_2[0] }), .EastIn({\nOut2_1[7] , \nOut2_1[6] , 
        \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , 
        \nOut2_1[0] }), .WestIn({\nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , 
        \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), 
        .Out({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , 
        \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_128 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut129[7] , \nScanOut129[6] , 
        \nScanOut129[5] , \nScanOut129[4] , \nScanOut129[3] , \nScanOut129[2] , 
        \nScanOut129[1] , \nScanOut129[0] }), .ScanOut({\nScanOut128[7] , 
        \nScanOut128[6] , \nScanOut128[5] , \nScanOut128[4] , \nScanOut128[3] , 
        \nScanOut128[2] , \nScanOut128[1] , \nScanOut128[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut8_0[7] , \nOut8_0[6] , 
        \nOut8_0[5] , \nOut8_0[4] , \nOut8_0[3] , \nOut8_0[2] , \nOut8_0[1] , 
        \nOut8_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_184 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut185[7] , \nScanOut185[6] , 
        \nScanOut185[5] , \nScanOut185[4] , \nScanOut185[3] , \nScanOut185[2] , 
        \nScanOut185[1] , \nScanOut185[0] }), .ScanOut({\nScanOut184[7] , 
        \nScanOut184[6] , \nScanOut184[5] , \nScanOut184[4] , \nScanOut184[3] , 
        \nScanOut184[2] , \nScanOut184[1] , \nScanOut184[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), 
        .SouthIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , \nOut11_9[4] , 
        \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , \nOut11_9[0] }), .EastIn(
        {\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .WestIn(
        {\nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), .Out({
        \nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_218 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut219[7] , \nScanOut219[6] , 
        \nScanOut219[5] , \nScanOut219[4] , \nScanOut219[3] , \nScanOut219[2] , 
        \nScanOut219[1] , \nScanOut219[0] }), .ScanOut({\nScanOut218[7] , 
        \nScanOut218[6] , \nScanOut218[5] , \nScanOut218[4] , \nScanOut218[3] , 
        \nScanOut218[2] , \nScanOut218[1] , \nScanOut218[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , \nOut13_9[4] , 
        \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , \nOut13_9[0] }), 
        .SouthIn({\nOut13_11[7] , \nOut13_11[6] , \nOut13_11[5] , 
        \nOut13_11[4] , \nOut13_11[3] , \nOut13_11[2] , \nOut13_11[1] , 
        \nOut13_11[0] }), .EastIn({\nOut14_10[7] , \nOut14_10[6] , 
        \nOut14_10[5] , \nOut14_10[4] , \nOut14_10[3] , \nOut14_10[2] , 
        \nOut14_10[1] , \nOut14_10[0] }), .WestIn({\nOut12_10[7] , 
        \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , 
        \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }), .Out({\nOut13_10[7] , 
        \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , 
        \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_183 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut184[7] , \nScanOut184[6] , 
        \nScanOut184[5] , \nScanOut184[4] , \nScanOut184[3] , \nScanOut184[2] , 
        \nScanOut184[1] , \nScanOut184[0] }), .ScanOut({\nScanOut183[7] , 
        \nScanOut183[6] , \nScanOut183[5] , \nScanOut183[4] , \nScanOut183[3] , 
        \nScanOut183[2] , \nScanOut183[1] , \nScanOut183[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), 
        .SouthIn({\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .EastIn(
        {\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .WestIn(
        {\nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), .Out({
        \nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_30 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut31[7] , \nScanOut31[6] , 
        \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , 
        \nScanOut31[1] , \nScanOut31[0] }), .ScanOut({\nScanOut30[7] , 
        \nScanOut30[6] , \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , 
        \nScanOut30[2] , \nScanOut30[1] , \nScanOut30[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), 
        .SouthIn({\nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , 
        \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), .EastIn(
        {\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .WestIn(
        {\nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , 
        \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), .Out({
        \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_45 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut46[7] , \nScanOut46[6] , 
        \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , 
        \nScanOut46[1] , \nScanOut46[0] }), .ScanOut({\nScanOut45[7] , 
        \nScanOut45[6] , \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , 
        \nScanOut45[2] , \nScanOut45[1] , \nScanOut45[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), 
        .SouthIn({\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .EastIn(
        {\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .WestIn(
        {\nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .Out({
        \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_62 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut63[7] , \nScanOut63[6] , 
        \nScanOut63[5] , \nScanOut63[4] , \nScanOut63[3] , \nScanOut63[2] , 
        \nScanOut63[1] , \nScanOut63[0] }), .ScanOut({\nScanOut62[7] , 
        \nScanOut62[6] , \nScanOut62[5] , \nScanOut62[4] , \nScanOut62[3] , 
        \nScanOut62[2] , \nScanOut62[1] , \nScanOut62[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), 
        .SouthIn({\nOut3_15[7] , \nOut3_15[6] , \nOut3_15[5] , \nOut3_15[4] , 
        \nOut3_15[3] , \nOut3_15[2] , \nOut3_15[1] , \nOut3_15[0] }), .EastIn(
        {\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .WestIn(
        {\nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .Out({
        \nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_79 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut80[7] , \nScanOut80[6] , 
        \nScanOut80[5] , \nScanOut80[4] , \nScanOut80[3] , \nScanOut80[2] , 
        \nScanOut80[1] , \nScanOut80[0] }), .ScanOut({\nScanOut79[7] , 
        \nScanOut79[6] , \nScanOut79[5] , \nScanOut79[4] , \nScanOut79[3] , 
        \nScanOut79[2] , \nScanOut79[1] , \nScanOut79[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut4_15[7] , \nOut4_15[6] , 
        \nOut4_15[5] , \nOut4_15[4] , \nOut4_15[3] , \nOut4_15[2] , 
        \nOut4_15[1] , \nOut4_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_108 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut109[7] , \nScanOut109[6] , 
        \nScanOut109[5] , \nScanOut109[4] , \nScanOut109[3] , \nScanOut109[2] , 
        \nScanOut109[1] , \nScanOut109[0] }), .ScanOut({\nScanOut108[7] , 
        \nScanOut108[6] , \nScanOut108[5] , \nScanOut108[4] , \nScanOut108[3] , 
        \nScanOut108[2] , \nScanOut108[1] , \nScanOut108[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), 
        .SouthIn({\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .EastIn(
        {\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .WestIn(
        {\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .Out({
        \nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_238 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut239[7] , \nScanOut239[6] , 
        \nScanOut239[5] , \nScanOut239[4] , \nScanOut239[3] , \nScanOut239[2] , 
        \nScanOut239[1] , \nScanOut239[0] }), .ScanOut({\nScanOut238[7] , 
        \nScanOut238[6] , \nScanOut238[5] , \nScanOut238[4] , \nScanOut238[3] , 
        \nScanOut238[2] , \nScanOut238[1] , \nScanOut238[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_13[7] , \nOut14_13[6] , \nOut14_13[5] , \nOut14_13[4] , 
        \nOut14_13[3] , \nOut14_13[2] , \nOut14_13[1] , \nOut14_13[0] }), 
        .SouthIn({\nOut14_15[7] , \nOut14_15[6] , \nOut14_15[5] , 
        \nOut14_15[4] , \nOut14_15[3] , \nOut14_15[2] , \nOut14_15[1] , 
        \nOut14_15[0] }), .EastIn({\nOut15_14[7] , \nOut15_14[6] , 
        \nOut15_14[5] , \nOut15_14[4] , \nOut15_14[3] , \nOut15_14[2] , 
        \nOut15_14[1] , \nOut15_14[0] }), .WestIn({\nOut13_14[7] , 
        \nOut13_14[6] , \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , 
        \nOut13_14[2] , \nOut13_14[1] , \nOut13_14[0] }), .Out({\nOut14_14[7] , 
        \nOut14_14[6] , \nOut14_14[5] , \nOut14_14[4] , \nOut14_14[3] , 
        \nOut14_14[2] , \nOut14_14[1] , \nOut14_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_141 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut142[7] , \nScanOut142[6] , 
        \nScanOut142[5] , \nScanOut142[4] , \nScanOut142[3] , \nScanOut142[2] , 
        \nScanOut142[1] , \nScanOut142[0] }), .ScanOut({\nScanOut141[7] , 
        \nScanOut141[6] , \nScanOut141[5] , \nScanOut141[4] , \nScanOut141[3] , 
        \nScanOut141[2] , \nScanOut141[1] , \nScanOut141[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), 
        .SouthIn({\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .EastIn(
        {\nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .WestIn(
        {\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .Out({
        \nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_166 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut167[7] , \nScanOut167[6] , 
        \nScanOut167[5] , \nScanOut167[4] , \nScanOut167[3] , \nScanOut167[2] , 
        \nScanOut167[1] , \nScanOut167[0] }), .ScanOut({\nScanOut166[7] , 
        \nScanOut166[6] , \nScanOut166[5] , \nScanOut166[4] , \nScanOut166[3] , 
        \nScanOut166[2] , \nScanOut166[1] , \nScanOut166[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), 
        .SouthIn({\nOut10_7[7] , \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , 
        \nOut10_7[3] , \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }), .EastIn(
        {\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .WestIn(
        {\nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , 
        \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] }), .Out({\nOut10_6[7] , 
        \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , \nOut10_6[3] , 
        \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_22 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut23[7] , \nScanOut23[6] , 
        \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , 
        \nScanOut23[1] , \nScanOut23[0] }), .ScanOut({\nScanOut22[7] , 
        \nScanOut22[6] , \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , 
        \nScanOut22[2] , \nScanOut22[1] , \nScanOut22[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , 
        \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), .SouthIn({\nOut1_7[7] , 
        \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , 
        \nOut1_7[1] , \nOut1_7[0] }), .EastIn({\nOut2_6[7] , \nOut2_6[6] , 
        \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , 
        \nOut2_6[0] }), .WestIn({\nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , 
        \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), 
        .Out({\nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , 
        \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_39 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut40[7] , \nScanOut40[6] , 
        \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , 
        \nScanOut40[1] , \nScanOut40[0] }), .ScanOut({\nScanOut39[7] , 
        \nScanOut39[6] , \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , 
        \nScanOut39[2] , \nScanOut39[1] , \nScanOut39[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , 
        \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), .SouthIn({\nOut2_8[7] , 
        \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , 
        \nOut2_8[1] , \nOut2_8[0] }), .EastIn({\nOut3_7[7] , \nOut3_7[6] , 
        \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , 
        \nOut3_7[0] }), .WestIn({\nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , 
        \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), 
        .Out({\nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , 
        \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_87 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut88[7] , \nScanOut88[6] , 
        \nScanOut88[5] , \nScanOut88[4] , \nScanOut88[3] , \nScanOut88[2] , 
        \nScanOut88[1] , \nScanOut88[0] }), .ScanOut({\nScanOut87[7] , 
        \nScanOut87[6] , \nScanOut87[5] , \nScanOut87[4] , \nScanOut87[3] , 
        \nScanOut87[2] , \nScanOut87[1] , \nScanOut87[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , 
        \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }), .SouthIn({\nOut5_8[7] , 
        \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , 
        \nOut5_8[1] , \nOut5_8[0] }), .EastIn({\nOut6_7[7] , \nOut6_7[6] , 
        \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , 
        \nOut6_7[0] }), .WestIn({\nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , 
        \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }), 
        .Out({\nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , 
        \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_113 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut114[7] , \nScanOut114[6] , 
        \nScanOut114[5] , \nScanOut114[4] , \nScanOut114[3] , \nScanOut114[2] , 
        \nScanOut114[1] , \nScanOut114[0] }), .ScanOut({\nScanOut113[7] , 
        \nScanOut113[6] , \nScanOut113[5] , \nScanOut113[4] , \nScanOut113[3] , 
        \nScanOut113[2] , \nScanOut113[1] , \nScanOut113[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_0[7] , \nOut7_0[6] , \nOut7_0[5] , \nOut7_0[4] , \nOut7_0[3] , 
        \nOut7_0[2] , \nOut7_0[1] , \nOut7_0[0] }), .SouthIn({\nOut7_2[7] , 
        \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , 
        \nOut7_2[1] , \nOut7_2[0] }), .EastIn({\nOut8_1[7] , \nOut8_1[6] , 
        \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , 
        \nOut8_1[0] }), .WestIn({\nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , 
        \nOut6_1[4] , \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }), 
        .Out({\nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , \nOut7_1[4] , 
        \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_134 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut135[7] , \nScanOut135[6] , 
        \nScanOut135[5] , \nScanOut135[4] , \nScanOut135[3] , \nScanOut135[2] , 
        \nScanOut135[1] , \nScanOut135[0] }), .ScanOut({\nScanOut134[7] , 
        \nScanOut134[6] , \nScanOut134[5] , \nScanOut134[4] , \nScanOut134[3] , 
        \nScanOut134[2] , \nScanOut134[1] , \nScanOut134[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_5[7] , \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , 
        \nOut8_5[2] , \nOut8_5[1] , \nOut8_5[0] }), .SouthIn({\nOut8_7[7] , 
        \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , 
        \nOut8_7[1] , \nOut8_7[0] }), .EastIn({\nOut9_6[7] , \nOut9_6[6] , 
        \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , \nOut9_6[1] , 
        \nOut9_6[0] }), .WestIn({\nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , 
        \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }), 
        .Out({\nOut8_6[7] , \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , 
        \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , \nOut8_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_204 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut205[7] , \nScanOut205[6] , 
        \nScanOut205[5] , \nScanOut205[4] , \nScanOut205[3] , \nScanOut205[2] , 
        \nScanOut205[1] , \nScanOut205[0] }), .ScanOut({\nScanOut204[7] , 
        \nScanOut204[6] , \nScanOut204[5] , \nScanOut204[4] , \nScanOut204[3] , 
        \nScanOut204[2] , \nScanOut204[1] , \nScanOut204[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_11[7] , \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , 
        \nOut12_11[3] , \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }), 
        .SouthIn({\nOut12_13[7] , \nOut12_13[6] , \nOut12_13[5] , 
        \nOut12_13[4] , \nOut12_13[3] , \nOut12_13[2] , \nOut12_13[1] , 
        \nOut12_13[0] }), .EastIn({\nOut13_12[7] , \nOut13_12[6] , 
        \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , \nOut13_12[2] , 
        \nOut13_12[1] , \nOut13_12[0] }), .WestIn({\nOut11_12[7] , 
        \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , 
        \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }), .Out({\nOut12_12[7] , 
        \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , 
        \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_198 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut199[7] , \nScanOut199[6] , 
        \nScanOut199[5] , \nScanOut199[4] , \nScanOut199[3] , \nScanOut199[2] , 
        \nScanOut199[1] , \nScanOut199[0] }), .ScanOut({\nScanOut198[7] , 
        \nScanOut198[6] , \nScanOut198[5] , \nScanOut198[4] , \nScanOut198[3] , 
        \nScanOut198[2] , \nScanOut198[1] , \nScanOut198[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), 
        .SouthIn({\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .EastIn(
        {\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .WestIn(
        {\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .Out({
        \nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_223 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut224[7] , \nScanOut224[6] , 
        \nScanOut224[5] , \nScanOut224[4] , \nScanOut224[3] , \nScanOut224[2] , 
        \nScanOut224[1] , \nScanOut224[0] }), .ScanOut({\nScanOut223[7] , 
        \nScanOut223[6] , \nScanOut223[5] , \nScanOut223[4] , \nScanOut223[3] , 
        \nScanOut223[2] , \nScanOut223[1] , \nScanOut223[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut13_15[7] , \nOut13_15[6] , 
        \nOut13_15[5] , \nOut13_15[4] , \nOut13_15[3] , \nOut13_15[2] , 
        \nOut13_15[1] , \nOut13_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_57 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut58[7] , \nScanOut58[6] , 
        \nScanOut58[5] , \nScanOut58[4] , \nScanOut58[3] , \nScanOut58[2] , 
        \nScanOut58[1] , \nScanOut58[0] }), .ScanOut({\nScanOut57[7] , 
        \nScanOut57[6] , \nScanOut57[5] , \nScanOut57[4] , \nScanOut57[3] , 
        \nScanOut57[2] , \nScanOut57[1] , \nScanOut57[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , 
        \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }), .SouthIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .EastIn({\nOut4_9[7] , 
        \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , 
        \nOut4_9[1] , \nOut4_9[0] }), .WestIn({\nOut2_9[7] , \nOut2_9[6] , 
        \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , 
        \nOut2_9[0] }), .Out({\nOut3_9[7] , \nOut3_9[6] , \nOut3_9[5] , 
        \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , \nOut3_9[1] , \nOut3_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_70 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut71[7] , \nScanOut71[6] , 
        \nScanOut71[5] , \nScanOut71[4] , \nScanOut71[3] , \nScanOut71[2] , 
        \nScanOut71[1] , \nScanOut71[0] }), .ScanOut({\nScanOut70[7] , 
        \nScanOut70[6] , \nScanOut70[5] , \nScanOut70[4] , \nScanOut70[3] , 
        \nScanOut70[2] , \nScanOut70[1] , \nScanOut70[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , 
        \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }), .SouthIn({\nOut4_7[7] , 
        \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , 
        \nOut4_7[1] , \nOut4_7[0] }), .EastIn({\nOut5_6[7] , \nOut5_6[6] , 
        \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , 
        \nOut5_6[0] }), .WestIn({\nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , 
        \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }), 
        .Out({\nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , 
        \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_95 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut96[7] , \nScanOut96[6] , 
        \nScanOut96[5] , \nScanOut96[4] , \nScanOut96[3] , \nScanOut96[2] , 
        \nScanOut96[1] , \nScanOut96[0] }), .ScanOut({\nScanOut95[7] , 
        \nScanOut95[6] , \nScanOut95[5] , \nScanOut95[4] , \nScanOut95[3] , 
        \nScanOut95[2] , \nScanOut95[1] , \nScanOut95[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut5_15[7] , \nOut5_15[6] , 
        \nOut5_15[5] , \nOut5_15[4] , \nOut5_15[3] , \nOut5_15[2] , 
        \nOut5_15[1] , \nOut5_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_101 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut102[7] , \nScanOut102[6] , 
        \nScanOut102[5] , \nScanOut102[4] , \nScanOut102[3] , \nScanOut102[2] , 
        \nScanOut102[1] , \nScanOut102[0] }), .ScanOut({\nScanOut101[7] , 
        \nScanOut101[6] , \nScanOut101[5] , \nScanOut101[4] , \nScanOut101[3] , 
        \nScanOut101[2] , \nScanOut101[1] , \nScanOut101[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , 
        \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }), .SouthIn({\nOut6_6[7] , 
        \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , 
        \nOut6_6[1] , \nOut6_6[0] }), .EastIn({\nOut7_5[7] , \nOut7_5[6] , 
        \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , 
        \nOut7_5[0] }), .WestIn({\nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , 
        \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }), 
        .Out({\nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , 
        \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_126 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut127[7] , \nScanOut127[6] , 
        \nScanOut127[5] , \nScanOut127[4] , \nScanOut127[3] , \nScanOut127[2] , 
        \nScanOut127[1] , \nScanOut127[0] }), .ScanOut({\nScanOut126[7] , 
        \nScanOut126[6] , \nScanOut126[5] , \nScanOut126[4] , \nScanOut126[3] , 
        \nScanOut126[2] , \nScanOut126[1] , \nScanOut126[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), 
        .SouthIn({\nOut7_15[7] , \nOut7_15[6] , \nOut7_15[5] , \nOut7_15[4] , 
        \nOut7_15[3] , \nOut7_15[2] , \nOut7_15[1] , \nOut7_15[0] }), .EastIn(
        {\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .WestIn(
        {\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .Out({
        \nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_216 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut217[7] , \nScanOut217[6] , 
        \nScanOut217[5] , \nScanOut217[4] , \nScanOut217[3] , \nScanOut217[2] , 
        \nScanOut217[1] , \nScanOut217[0] }), .ScanOut({\nScanOut216[7] , 
        \nScanOut216[6] , \nScanOut216[5] , \nScanOut216[4] , \nScanOut216[3] , 
        \nScanOut216[2] , \nScanOut216[1] , \nScanOut216[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), 
        .SouthIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , \nOut13_9[4] , 
        \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , \nOut13_9[0] }), .EastIn(
        {\nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), .WestIn(
        {\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .Out({
        \nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_148 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut149[7] , \nScanOut149[6] , 
        \nScanOut149[5] , \nScanOut149[4] , \nScanOut149[3] , \nScanOut149[2] , 
        \nScanOut149[1] , \nScanOut149[0] }), .ScanOut({\nScanOut148[7] , 
        \nScanOut148[6] , \nScanOut148[5] , \nScanOut148[4] , \nScanOut148[3] , 
        \nScanOut148[2] , \nScanOut148[1] , \nScanOut148[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , 
        \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] }), .SouthIn({\nOut9_5[7] , 
        \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , 
        \nOut9_5[1] , \nOut9_5[0] }), .EastIn({\nOut10_4[7] , \nOut10_4[6] , 
        \nOut10_4[5] , \nOut10_4[4] , \nOut10_4[3] , \nOut10_4[2] , 
        \nOut10_4[1] , \nOut10_4[0] }), .WestIn({\nOut8_4[7] , \nOut8_4[6] , 
        \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , 
        \nOut8_4[0] }), .Out({\nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , 
        \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_231 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut232[7] , \nScanOut232[6] , 
        \nScanOut232[5] , \nScanOut232[4] , \nScanOut232[3] , \nScanOut232[2] , 
        \nScanOut232[1] , \nScanOut232[0] }), .ScanOut({\nScanOut231[7] , 
        \nScanOut231[6] , \nScanOut231[5] , \nScanOut231[4] , \nScanOut231[3] , 
        \nScanOut231[2] , \nScanOut231[1] , \nScanOut231[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), 
        .SouthIn({\nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), .EastIn(
        {\nOut15_7[7] , \nOut15_7[6] , \nOut15_7[5] , \nOut15_7[4] , 
        \nOut15_7[3] , \nOut15_7[2] , \nOut15_7[1] , \nOut15_7[0] }), .WestIn(
        {\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .Out({
        \nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_153 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut154[7] , \nScanOut154[6] , 
        \nScanOut154[5] , \nScanOut154[4] , \nScanOut154[3] , \nScanOut154[2] , 
        \nScanOut154[1] , \nScanOut154[0] }), .ScanOut({\nScanOut153[7] , 
        \nScanOut153[6] , \nScanOut153[5] , \nScanOut153[4] , \nScanOut153[3] , 
        \nScanOut153[2] , \nScanOut153[1] , \nScanOut153[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , 
        \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] }), .SouthIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .EastIn({\nOut10_9[7] , 
        \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , \nOut10_9[3] , 
        \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), .WestIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .Out({\nOut9_9[7] , \nOut9_9[6] , 
        \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , \nOut9_9[1] , 
        \nOut9_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_174 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut175[7] , \nScanOut175[6] , 
        \nScanOut175[5] , \nScanOut175[4] , \nScanOut175[3] , \nScanOut175[2] , 
        \nScanOut175[1] , \nScanOut175[0] }), .ScanOut({\nScanOut174[7] , 
        \nScanOut174[6] , \nScanOut174[5] , \nScanOut174[4] , \nScanOut174[3] , 
        \nScanOut174[2] , \nScanOut174[1] , \nScanOut174[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , 
        \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), 
        .SouthIn({\nOut10_15[7] , \nOut10_15[6] , \nOut10_15[5] , 
        \nOut10_15[4] , \nOut10_15[3] , \nOut10_15[2] , \nOut10_15[1] , 
        \nOut10_15[0] }), .EastIn({\nOut11_14[7] , \nOut11_14[6] , 
        \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , \nOut11_14[2] , 
        \nOut11_14[1] , \nOut11_14[0] }), .WestIn({\nOut9_14[7] , 
        \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , \nOut9_14[3] , 
        \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .Out({\nOut10_14[7] , 
        \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , \nOut10_14[3] , 
        \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_244 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut245[7] , \nScanOut245[6] , 
        \nScanOut245[5] , \nScanOut245[4] , \nScanOut245[3] , \nScanOut245[2] , 
        \nScanOut245[1] , \nScanOut245[0] }), .ScanOut({\nScanOut244[7] , 
        \nScanOut244[6] , \nScanOut244[5] , \nScanOut244[4] , \nScanOut244[3] , 
        \nScanOut244[2] , \nScanOut244[1] , \nScanOut244[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_4[7] , \nOut15_4[6] , 
        \nOut15_4[5] , \nOut15_4[4] , \nOut15_4[3] , \nOut15_4[2] , 
        \nOut15_4[1] , \nOut15_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_191 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut192[7] , \nScanOut192[6] , 
        \nScanOut192[5] , \nScanOut192[4] , \nScanOut192[3] , \nScanOut192[2] , 
        \nScanOut192[1] , \nScanOut192[0] }), .ScanOut({\nScanOut191[7] , 
        \nScanOut191[6] , \nScanOut191[5] , \nScanOut191[4] , \nScanOut191[3] , 
        \nScanOut191[2] , \nScanOut191[1] , \nScanOut191[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut11_15[7] , \nOut11_15[6] , 
        \nOut11_15[5] , \nOut11_15[4] , \nOut11_15[3] , \nOut11_15[2] , 
        \nOut11_15[1] , \nOut11_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_63 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut64[7] , \nScanOut64[6] , 
        \nScanOut64[5] , \nScanOut64[4] , \nScanOut64[3] , \nScanOut64[2] , 
        \nScanOut64[1] , \nScanOut64[0] }), .ScanOut({\nScanOut63[7] , 
        \nScanOut63[6] , \nScanOut63[5] , \nScanOut63[4] , \nScanOut63[3] , 
        \nScanOut63[2] , \nScanOut63[1] , \nScanOut63[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_15[7] , \nOut3_15[6] , 
        \nOut3_15[5] , \nOut3_15[4] , \nOut3_15[3] , \nOut3_15[2] , 
        \nOut3_15[1] , \nOut3_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_86 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut87[7] , \nScanOut87[6] , 
        \nScanOut87[5] , \nScanOut87[4] , \nScanOut87[3] , \nScanOut87[2] , 
        \nScanOut87[1] , \nScanOut87[0] }), .ScanOut({\nScanOut86[7] , 
        \nScanOut86[6] , \nScanOut86[5] , \nScanOut86[4] , \nScanOut86[3] , 
        \nScanOut86[2] , \nScanOut86[1] , \nScanOut86[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , 
        \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }), .SouthIn({\nOut5_7[7] , 
        \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , 
        \nOut5_7[1] , \nOut5_7[0] }), .EastIn({\nOut6_6[7] , \nOut6_6[6] , 
        \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , 
        \nOut6_6[0] }), .WestIn({\nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , 
        \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }), 
        .Out({\nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , 
        \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_135 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut136[7] , \nScanOut136[6] , 
        \nScanOut136[5] , \nScanOut136[4] , \nScanOut136[3] , \nScanOut136[2] , 
        \nScanOut136[1] , \nScanOut136[0] }), .ScanOut({\nScanOut135[7] , 
        \nScanOut135[6] , \nScanOut135[5] , \nScanOut135[4] , \nScanOut135[3] , 
        \nScanOut135[2] , \nScanOut135[1] , \nScanOut135[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_6[7] , \nOut8_6[6] , \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , 
        \nOut8_6[2] , \nOut8_6[1] , \nOut8_6[0] }), .SouthIn({\nOut8_8[7] , 
        \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , 
        \nOut8_8[1] , \nOut8_8[0] }), .EastIn({\nOut9_7[7] , \nOut9_7[6] , 
        \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , \nOut9_7[1] , 
        \nOut9_7[0] }), .WestIn({\nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , 
        \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }), 
        .Out({\nOut8_7[7] , \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , 
        \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , \nOut8_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_205 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut206[7] , \nScanOut206[6] , 
        \nScanOut206[5] , \nScanOut206[4] , \nScanOut206[3] , \nScanOut206[2] , 
        \nScanOut206[1] , \nScanOut206[0] }), .ScanOut({\nScanOut205[7] , 
        \nScanOut205[6] , \nScanOut205[5] , \nScanOut205[4] , \nScanOut205[3] , 
        \nScanOut205[2] , \nScanOut205[1] , \nScanOut205[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_12[7] , \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , 
        \nOut12_12[3] , \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }), 
        .SouthIn({\nOut12_14[7] , \nOut12_14[6] , \nOut12_14[5] , 
        \nOut12_14[4] , \nOut12_14[3] , \nOut12_14[2] , \nOut12_14[1] , 
        \nOut12_14[0] }), .EastIn({\nOut13_13[7] , \nOut13_13[6] , 
        \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , \nOut13_13[2] , 
        \nOut13_13[1] , \nOut13_13[0] }), .WestIn({\nOut11_13[7] , 
        \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , 
        \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }), .Out({\nOut12_13[7] , 
        \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , 
        \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_112 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut113[7] , \nScanOut113[6] , 
        \nScanOut113[5] , \nScanOut113[4] , \nScanOut113[3] , \nScanOut113[2] , 
        \nScanOut113[1] , \nScanOut113[0] }), .ScanOut({\nScanOut112[7] , 
        \nScanOut112[6] , \nScanOut112[5] , \nScanOut112[4] , \nScanOut112[3] , 
        \nScanOut112[2] , \nScanOut112[1] , \nScanOut112[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut7_0[7] , \nOut7_0[6] , 
        \nOut7_0[5] , \nOut7_0[4] , \nOut7_0[3] , \nOut7_0[2] , \nOut7_0[1] , 
        \nOut7_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_199 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut200[7] , \nScanOut200[6] , 
        \nScanOut200[5] , \nScanOut200[4] , \nScanOut200[3] , \nScanOut200[2] , 
        \nScanOut200[1] , \nScanOut200[0] }), .ScanOut({\nScanOut199[7] , 
        \nScanOut199[6] , \nScanOut199[5] , \nScanOut199[4] , \nScanOut199[3] , 
        \nScanOut199[2] , \nScanOut199[1] , \nScanOut199[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), 
        .SouthIn({\nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), .EastIn(
        {\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .WestIn(
        {\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .Out({
        \nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_222 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut223[7] , \nScanOut223[6] , 
        \nScanOut223[5] , \nScanOut223[4] , \nScanOut223[3] , \nScanOut223[2] , 
        \nScanOut223[1] , \nScanOut223[0] }), .ScanOut({\nScanOut222[7] , 
        \nScanOut222[6] , \nScanOut222[5] , \nScanOut222[4] , \nScanOut222[3] , 
        \nScanOut222[2] , \nScanOut222[1] , \nScanOut222[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_13[7] , \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , 
        \nOut13_13[3] , \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }), 
        .SouthIn({\nOut13_15[7] , \nOut13_15[6] , \nOut13_15[5] , 
        \nOut13_15[4] , \nOut13_15[3] , \nOut13_15[2] , \nOut13_15[1] , 
        \nOut13_15[0] }), .EastIn({\nOut14_14[7] , \nOut14_14[6] , 
        \nOut14_14[5] , \nOut14_14[4] , \nOut14_14[3] , \nOut14_14[2] , 
        \nOut14_14[1] , \nOut14_14[0] }), .WestIn({\nOut12_14[7] , 
        \nOut12_14[6] , \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , 
        \nOut12_14[2] , \nOut12_14[1] , \nOut12_14[0] }), .Out({\nOut13_14[7] , 
        \nOut13_14[6] , \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , 
        \nOut13_14[2] , \nOut13_14[1] , \nOut13_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut6[7] , \nScanOut6[6] , 
        \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , 
        \nScanOut6[1] , \nScanOut6[0] }), .ScanOut({\nScanOut5[7] , 
        \nScanOut5[6] , \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , 
        \nScanOut5[2] , \nScanOut5[1] , \nScanOut5[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_5[7] , \nOut0_5[6] , 
        \nOut0_5[5] , \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , 
        \nOut0_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut12[7] , \nScanOut12[6] , 
        \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , 
        \nScanOut12[1] , \nScanOut12[0] }), .ScanOut({\nScanOut11[7] , 
        \nScanOut11[6] , \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , 
        \nScanOut11[2] , \nScanOut11[1] , \nScanOut11[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_11[7] , \nOut0_11[6] , 
        \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , \nOut0_11[2] , 
        \nOut0_11[1] , \nOut0_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_16 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut17[7] , \nScanOut17[6] , 
        \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , 
        \nScanOut17[1] , \nScanOut17[0] }), .ScanOut({\nScanOut16[7] , 
        \nScanOut16[6] , \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , 
        \nScanOut16[2] , \nScanOut16[1] , \nScanOut16[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_0[7] , \nOut1_0[6] , 
        \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , 
        \nOut1_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_44 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut45[7] , \nScanOut45[6] , 
        \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , 
        \nScanOut45[1] , \nScanOut45[0] }), .ScanOut({\nScanOut44[7] , 
        \nScanOut44[6] , \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , 
        \nScanOut44[2] , \nScanOut44[1] , \nScanOut44[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), 
        .SouthIn({\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .EastIn(
        {\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .WestIn(
        {\nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .Out({
        \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_78 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut79[7] , \nScanOut79[6] , 
        \nScanOut79[5] , \nScanOut79[4] , \nScanOut79[3] , \nScanOut79[2] , 
        \nScanOut79[1] , \nScanOut79[0] }), .ScanOut({\nScanOut78[7] , 
        \nScanOut78[6] , \nScanOut78[5] , \nScanOut78[4] , \nScanOut78[3] , 
        \nScanOut78[2] , \nScanOut78[1] , \nScanOut78[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), 
        .SouthIn({\nOut4_15[7] , \nOut4_15[6] , \nOut4_15[5] , \nOut4_15[4] , 
        \nOut4_15[3] , \nOut4_15[2] , \nOut4_15[1] , \nOut4_15[0] }), .EastIn(
        {\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .WestIn(
        {\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .Out({
        \nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_140 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut141[7] , \nScanOut141[6] , 
        \nScanOut141[5] , \nScanOut141[4] , \nScanOut141[3] , \nScanOut141[2] , 
        \nScanOut141[1] , \nScanOut141[0] }), .ScanOut({\nScanOut140[7] , 
        \nScanOut140[6] , \nScanOut140[5] , \nScanOut140[4] , \nScanOut140[3] , 
        \nScanOut140[2] , \nScanOut140[1] , \nScanOut140[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), 
        .SouthIn({\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .EastIn(
        {\nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .WestIn(
        {\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .Out({
        \nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_167 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut168[7] , \nScanOut168[6] , 
        \nScanOut168[5] , \nScanOut168[4] , \nScanOut168[3] , \nScanOut168[2] , 
        \nScanOut168[1] , \nScanOut168[0] }), .ScanOut({\nScanOut167[7] , 
        \nScanOut167[6] , \nScanOut167[5] , \nScanOut167[4] , \nScanOut167[3] , 
        \nScanOut167[2] , \nScanOut167[1] , \nScanOut167[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), 
        .SouthIn({\nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), .EastIn(
        {\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .WestIn(
        {\nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , 
        \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] }), .Out({\nOut10_7[7] , 
        \nOut10_7[6] , \nOut10_7[5] , \nOut10_7[4] , \nOut10_7[3] , 
        \nOut10_7[2] , \nOut10_7[1] , \nOut10_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_18 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut19[7] , \nScanOut19[6] , 
        \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , 
        \nScanOut19[1] , \nScanOut19[0] }), .ScanOut({\nScanOut18[7] , 
        \nScanOut18[6] , \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , 
        \nScanOut18[2] , \nScanOut18[1] , \nScanOut18[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , \nOut1_1[3] , 
        \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), .SouthIn({\nOut1_3[7] , 
        \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , 
        \nOut1_3[1] , \nOut1_3[0] }), .EastIn({\nOut2_2[7] , \nOut2_2[6] , 
        \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , 
        \nOut2_2[0] }), .WestIn({\nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , 
        \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), 
        .Out({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , 
        \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_23 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut24[7] , \nScanOut24[6] , 
        \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , 
        \nScanOut24[1] , \nScanOut24[0] }), .ScanOut({\nScanOut23[7] , 
        \nScanOut23[6] , \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , 
        \nScanOut23[2] , \nScanOut23[1] , \nScanOut23[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , 
        \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), .SouthIn({\nOut1_8[7] , 
        \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , 
        \nOut1_8[1] , \nOut1_8[0] }), .EastIn({\nOut2_7[7] , \nOut2_7[6] , 
        \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , 
        \nOut2_7[0] }), .WestIn({\nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , 
        \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), 
        .Out({\nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , 
        \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_31 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut32[7] , \nScanOut32[6] , 
        \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , 
        \nScanOut32[1] , \nScanOut32[0] }), .ScanOut({\nScanOut31[7] , 
        \nScanOut31[6] , \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , 
        \nScanOut31[2] , \nScanOut31[1] , \nScanOut31[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_15[7] , \nOut1_15[6] , 
        \nOut1_15[5] , \nOut1_15[4] , \nOut1_15[3] , \nOut1_15[2] , 
        \nOut1_15[1] , \nOut1_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_182 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut183[7] , \nScanOut183[6] , 
        \nScanOut183[5] , \nScanOut183[4] , \nScanOut183[3] , \nScanOut183[2] , 
        \nScanOut183[1] , \nScanOut183[0] }), .ScanOut({\nScanOut182[7] , 
        \nScanOut182[6] , \nScanOut182[5] , \nScanOut182[4] , \nScanOut182[3] , 
        \nScanOut182[2] , \nScanOut182[1] , \nScanOut182[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), 
        .SouthIn({\nOut11_7[7] , \nOut11_7[6] , \nOut11_7[5] , \nOut11_7[4] , 
        \nOut11_7[3] , \nOut11_7[2] , \nOut11_7[1] , \nOut11_7[0] }), .EastIn(
        {\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .WestIn(
        {\nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), .Out({
        \nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_109 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut110[7] , \nScanOut110[6] , 
        \nScanOut110[5] , \nScanOut110[4] , \nScanOut110[3] , \nScanOut110[2] , 
        \nScanOut110[1] , \nScanOut110[0] }), .ScanOut({\nScanOut109[7] , 
        \nScanOut109[6] , \nScanOut109[5] , \nScanOut109[4] , \nScanOut109[3] , 
        \nScanOut109[2] , \nScanOut109[1] , \nScanOut109[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), 
        .SouthIn({\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .EastIn(
        {\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .WestIn(
        {\nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), .Out({
        \nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_239 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut240[7] , \nScanOut240[6] , 
        \nScanOut240[5] , \nScanOut240[4] , \nScanOut240[3] , \nScanOut240[2] , 
        \nScanOut240[1] , \nScanOut240[0] }), .ScanOut({\nScanOut239[7] , 
        \nScanOut239[6] , \nScanOut239[5] , \nScanOut239[4] , \nScanOut239[3] , 
        \nScanOut239[2] , \nScanOut239[1] , \nScanOut239[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut14_15[7] , \nOut14_15[6] , 
        \nOut14_15[5] , \nOut14_15[4] , \nOut14_15[3] , \nOut14_15[2] , 
        \nOut14_15[1] , \nOut14_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_190 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut191[7] , \nScanOut191[6] , 
        \nScanOut191[5] , \nScanOut191[4] , \nScanOut191[3] , \nScanOut191[2] , 
        \nScanOut191[1] , \nScanOut191[0] }), .ScanOut({\nScanOut190[7] , 
        \nScanOut190[6] , \nScanOut190[5] , \nScanOut190[4] , \nScanOut190[3] , 
        \nScanOut190[2] , \nScanOut190[1] , \nScanOut190[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_13[7] , \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , 
        \nOut11_13[3] , \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }), 
        .SouthIn({\nOut11_15[7] , \nOut11_15[6] , \nOut11_15[5] , 
        \nOut11_15[4] , \nOut11_15[3] , \nOut11_15[2] , \nOut11_15[1] , 
        \nOut11_15[0] }), .EastIn({\nOut12_14[7] , \nOut12_14[6] , 
        \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , \nOut12_14[2] , 
        \nOut12_14[1] , \nOut12_14[0] }), .WestIn({\nOut10_14[7] , 
        \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , \nOut10_14[3] , 
        \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }), .Out({\nOut11_14[7] , 
        \nOut11_14[6] , \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , 
        \nOut11_14[2] , \nOut11_14[1] , \nOut11_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_38 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut39[7] , \nScanOut39[6] , 
        \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , 
        \nScanOut39[1] , \nScanOut39[0] }), .ScanOut({\nScanOut38[7] , 
        \nScanOut38[6] , \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , 
        \nScanOut38[2] , \nScanOut38[1] , \nScanOut38[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , 
        \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), .SouthIn({\nOut2_7[7] , 
        \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , 
        \nOut2_7[1] , \nOut2_7[0] }), .EastIn({\nOut3_6[7] , \nOut3_6[6] , 
        \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , 
        \nOut3_6[0] }), .WestIn({\nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , 
        \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), 
        .Out({\nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , 
        \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_56 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut57[7] , \nScanOut57[6] , 
        \nScanOut57[5] , \nScanOut57[4] , \nScanOut57[3] , \nScanOut57[2] , 
        \nScanOut57[1] , \nScanOut57[0] }), .ScanOut({\nScanOut56[7] , 
        \nScanOut56[6] , \nScanOut56[5] , \nScanOut56[4] , \nScanOut56[3] , 
        \nScanOut56[2] , \nScanOut56[1] , \nScanOut56[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , 
        \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }), .SouthIn({\nOut3_9[7] , 
        \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , 
        \nOut3_9[1] , \nOut3_9[0] }), .EastIn({\nOut4_8[7] , \nOut4_8[6] , 
        \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , 
        \nOut4_8[0] }), .WestIn({\nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , 
        \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), 
        .Out({\nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , 
        \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_71 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut72[7] , \nScanOut72[6] , 
        \nScanOut72[5] , \nScanOut72[4] , \nScanOut72[3] , \nScanOut72[2] , 
        \nScanOut72[1] , \nScanOut72[0] }), .ScanOut({\nScanOut71[7] , 
        \nScanOut71[6] , \nScanOut71[5] , \nScanOut71[4] , \nScanOut71[3] , 
        \nScanOut71[2] , \nScanOut71[1] , \nScanOut71[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_6[7] , \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , 
        \nOut4_6[2] , \nOut4_6[1] , \nOut4_6[0] }), .SouthIn({\nOut4_8[7] , 
        \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , 
        \nOut4_8[1] , \nOut4_8[0] }), .EastIn({\nOut5_7[7] , \nOut5_7[6] , 
        \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , 
        \nOut5_7[0] }), .WestIn({\nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , 
        \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }), 
        .Out({\nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , 
        \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_149 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut150[7] , \nScanOut150[6] , 
        \nScanOut150[5] , \nScanOut150[4] , \nScanOut150[3] , \nScanOut150[2] , 
        \nScanOut150[1] , \nScanOut150[0] }), .ScanOut({\nScanOut149[7] , 
        \nScanOut149[6] , \nScanOut149[5] , \nScanOut149[4] , \nScanOut149[3] , 
        \nScanOut149[2] , \nScanOut149[1] , \nScanOut149[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , 
        \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] }), .SouthIn({\nOut9_6[7] , 
        \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , 
        \nOut9_6[1] , \nOut9_6[0] }), .EastIn({\nOut10_5[7] , \nOut10_5[6] , 
        \nOut10_5[5] , \nOut10_5[4] , \nOut10_5[3] , \nOut10_5[2] , 
        \nOut10_5[1] , \nOut10_5[0] }), .WestIn({\nOut8_5[7] , \nOut8_5[6] , 
        \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , 
        \nOut8_5[0] }), .Out({\nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , 
        \nOut9_5[4] , \nOut9_5[3] , \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_152 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut153[7] , \nScanOut153[6] , 
        \nScanOut153[5] , \nScanOut153[4] , \nScanOut153[3] , \nScanOut153[2] , 
        \nScanOut153[1] , \nScanOut153[0] }), .ScanOut({\nScanOut152[7] , 
        \nScanOut152[6] , \nScanOut152[5] , \nScanOut152[4] , \nScanOut152[3] , 
        \nScanOut152[2] , \nScanOut152[1] , \nScanOut152[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , 
        \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] }), .SouthIn({\nOut9_9[7] , 
        \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , 
        \nOut9_9[1] , \nOut9_9[0] }), .EastIn({\nOut10_8[7] , \nOut10_8[6] , 
        \nOut10_8[5] , \nOut10_8[4] , \nOut10_8[3] , \nOut10_8[2] , 
        \nOut10_8[1] , \nOut10_8[0] }), .WestIn({\nOut8_8[7] , \nOut8_8[6] , 
        \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , 
        \nOut8_8[0] }), .Out({\nOut9_8[7] , \nOut9_8[6] , \nOut9_8[5] , 
        \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , \nOut9_8[1] , \nOut9_8[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_175 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut176[7] , \nScanOut176[6] , 
        \nScanOut176[5] , \nScanOut176[4] , \nScanOut176[3] , \nScanOut176[2] , 
        \nScanOut176[1] , \nScanOut176[0] }), .ScanOut({\nScanOut175[7] , 
        \nScanOut175[6] , \nScanOut175[5] , \nScanOut175[4] , \nScanOut175[3] , 
        \nScanOut175[2] , \nScanOut175[1] , \nScanOut175[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut10_15[7] , \nOut10_15[6] , 
        \nOut10_15[5] , \nOut10_15[4] , \nOut10_15[3] , \nOut10_15[2] , 
        \nOut10_15[1] , \nOut10_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_245 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut246[7] , \nScanOut246[6] , 
        \nScanOut246[5] , \nScanOut246[4] , \nScanOut246[3] , \nScanOut246[2] , 
        \nScanOut246[1] , \nScanOut246[0] }), .ScanOut({\nScanOut245[7] , 
        \nScanOut245[6] , \nScanOut245[5] , \nScanOut245[4] , \nScanOut245[3] , 
        \nScanOut245[2] , \nScanOut245[1] , \nScanOut245[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_5[7] , \nOut15_5[6] , 
        \nOut15_5[5] , \nOut15_5[4] , \nOut15_5[3] , \nOut15_5[2] , 
        \nOut15_5[1] , \nOut15_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_94 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut95[7] , \nScanOut95[6] , 
        \nScanOut95[5] , \nScanOut95[4] , \nScanOut95[3] , \nScanOut95[2] , 
        \nScanOut95[1] , \nScanOut95[0] }), .ScanOut({\nScanOut94[7] , 
        \nScanOut94[6] , \nScanOut94[5] , \nScanOut94[4] , \nScanOut94[3] , 
        \nScanOut94[2] , \nScanOut94[1] , \nScanOut94[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }), 
        .SouthIn({\nOut5_15[7] , \nOut5_15[6] , \nOut5_15[5] , \nOut5_15[4] , 
        \nOut5_15[3] , \nOut5_15[2] , \nOut5_15[1] , \nOut5_15[0] }), .EastIn(
        {\nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }), .WestIn(
        {\nOut4_14[7] , \nOut4_14[6] , \nOut4_14[5] , \nOut4_14[4] , 
        \nOut4_14[3] , \nOut4_14[2] , \nOut4_14[1] , \nOut4_14[0] }), .Out({
        \nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_127 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut128[7] , \nScanOut128[6] , 
        \nScanOut128[5] , \nScanOut128[4] , \nScanOut128[3] , \nScanOut128[2] , 
        \nScanOut128[1] , \nScanOut128[0] }), .ScanOut({\nScanOut127[7] , 
        \nScanOut127[6] , \nScanOut127[5] , \nScanOut127[4] , \nScanOut127[3] , 
        \nScanOut127[2] , \nScanOut127[1] , \nScanOut127[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut7_15[7] , \nOut7_15[6] , 
        \nOut7_15[5] , \nOut7_15[4] , \nOut7_15[3] , \nOut7_15[2] , 
        \nOut7_15[1] , \nOut7_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_217 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut218[7] , \nScanOut218[6] , 
        \nScanOut218[5] , \nScanOut218[4] , \nScanOut218[3] , \nScanOut218[2] , 
        \nScanOut218[1] , \nScanOut218[0] }), .ScanOut({\nScanOut217[7] , 
        \nScanOut217[6] , \nScanOut217[5] , \nScanOut217[4] , \nScanOut217[3] , 
        \nScanOut217[2] , \nScanOut217[1] , \nScanOut217[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), 
        .SouthIn({\nOut13_10[7] , \nOut13_10[6] , \nOut13_10[5] , 
        \nOut13_10[4] , \nOut13_10[3] , \nOut13_10[2] , \nOut13_10[1] , 
        \nOut13_10[0] }), .EastIn({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , 
        \nOut14_9[4] , \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , 
        \nOut14_9[0] }), .WestIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }), .Out({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_100 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut101[7] , \nScanOut101[6] , 
        \nScanOut101[5] , \nScanOut101[4] , \nScanOut101[3] , \nScanOut101[2] , 
        \nScanOut101[1] , \nScanOut101[0] }), .ScanOut({\nScanOut100[7] , 
        \nScanOut100[6] , \nScanOut100[5] , \nScanOut100[4] , \nScanOut100[3] , 
        \nScanOut100[2] , \nScanOut100[1] , \nScanOut100[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , 
        \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }), .SouthIn({\nOut6_5[7] , 
        \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , 
        \nOut6_5[1] , \nOut6_5[0] }), .EastIn({\nOut7_4[7] , \nOut7_4[6] , 
        \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , 
        \nOut7_4[0] }), .WestIn({\nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , 
        \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }), 
        .Out({\nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , 
        \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_230 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut231[7] , \nScanOut231[6] , 
        \nScanOut231[5] , \nScanOut231[4] , \nScanOut231[3] , \nScanOut231[2] , 
        \nScanOut231[1] , \nScanOut231[0] }), .ScanOut({\nScanOut230[7] , 
        \nScanOut230[6] , \nScanOut230[5] , \nScanOut230[4] , \nScanOut230[3] , 
        \nScanOut230[2] , \nScanOut230[1] , \nScanOut230[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), 
        .SouthIn({\nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), .EastIn(
        {\nOut15_6[7] , \nOut15_6[6] , \nOut15_6[5] , \nOut15_6[4] , 
        \nOut15_6[3] , \nOut15_6[2] , \nOut15_6[1] , \nOut15_6[0] }), .WestIn(
        {\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .Out({
        \nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_24 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut25[7] , \nScanOut25[6] , 
        \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , 
        \nScanOut25[1] , \nScanOut25[0] }), .ScanOut({\nScanOut24[7] , 
        \nScanOut24[6] , \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , 
        \nScanOut24[2] , \nScanOut24[1] , \nScanOut24[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , 
        \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), .SouthIn({\nOut1_9[7] , 
        \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , 
        \nOut1_9[1] , \nOut1_9[0] }), .EastIn({\nOut2_8[7] , \nOut2_8[6] , 
        \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , 
        \nOut2_8[0] }), .WestIn({\nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , 
        \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), 
        .Out({\nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , 
        \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_51 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut52[7] , \nScanOut52[6] , 
        \nScanOut52[5] , \nScanOut52[4] , \nScanOut52[3] , \nScanOut52[2] , 
        \nScanOut52[1] , \nScanOut52[0] }), .ScanOut({\nScanOut51[7] , 
        \nScanOut51[6] , \nScanOut51[5] , \nScanOut51[4] , \nScanOut51[3] , 
        \nScanOut51[2] , \nScanOut51[1] , \nScanOut51[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , 
        \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }), .SouthIn({\nOut3_4[7] , 
        \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , 
        \nOut3_4[1] , \nOut3_4[0] }), .EastIn({\nOut4_3[7] , \nOut4_3[6] , 
        \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , 
        \nOut4_3[0] }), .WestIn({\nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , 
        \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), 
        .Out({\nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , 
        \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_93 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut94[7] , \nScanOut94[6] , 
        \nScanOut94[5] , \nScanOut94[4] , \nScanOut94[3] , \nScanOut94[2] , 
        \nScanOut94[1] , \nScanOut94[0] }), .ScanOut({\nScanOut93[7] , 
        \nScanOut93[6] , \nScanOut93[5] , \nScanOut93[4] , \nScanOut93[3] , 
        \nScanOut93[2] , \nScanOut93[1] , \nScanOut93[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), 
        .SouthIn({\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .EastIn(
        {\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .WestIn(
        {\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .Out({
        \nOut5_13[7] , \nOut5_13[6] , \nOut5_13[5] , \nOut5_13[4] , 
        \nOut5_13[3] , \nOut5_13[2] , \nOut5_13[1] , \nOut5_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_107 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut108[7] , \nScanOut108[6] , 
        \nScanOut108[5] , \nScanOut108[4] , \nScanOut108[3] , \nScanOut108[2] , 
        \nScanOut108[1] , \nScanOut108[0] }), .ScanOut({\nScanOut107[7] , 
        \nScanOut107[6] , \nScanOut107[5] , \nScanOut107[4] , \nScanOut107[3] , 
        \nScanOut107[2] , \nScanOut107[1] , \nScanOut107[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_10[7] , \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , 
        \nOut6_10[3] , \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), 
        .SouthIn({\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .EastIn(
        {\nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .WestIn(
        {\nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .Out({
        \nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_237 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut238[7] , \nScanOut238[6] , 
        \nScanOut238[5] , \nScanOut238[4] , \nScanOut238[3] , \nScanOut238[2] , 
        \nScanOut238[1] , \nScanOut238[0] }), .ScanOut({\nScanOut237[7] , 
        \nScanOut237[6] , \nScanOut237[5] , \nScanOut237[4] , \nScanOut237[3] , 
        \nScanOut237[2] , \nScanOut237[1] , \nScanOut237[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_12[7] , \nOut14_12[6] , \nOut14_12[5] , \nOut14_12[4] , 
        \nOut14_12[3] , \nOut14_12[2] , \nOut14_12[1] , \nOut14_12[0] }), 
        .SouthIn({\nOut14_14[7] , \nOut14_14[6] , \nOut14_14[5] , 
        \nOut14_14[4] , \nOut14_14[3] , \nOut14_14[2] , \nOut14_14[1] , 
        \nOut14_14[0] }), .EastIn({\nOut15_13[7] , \nOut15_13[6] , 
        \nOut15_13[5] , \nOut15_13[4] , \nOut15_13[3] , \nOut15_13[2] , 
        \nOut15_13[1] , \nOut15_13[0] }), .WestIn({\nOut13_13[7] , 
        \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , 
        \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }), .Out({\nOut14_13[7] , 
        \nOut14_13[6] , \nOut14_13[5] , \nOut14_13[4] , \nOut14_13[3] , 
        \nOut14_13[2] , \nOut14_13[1] , \nOut14_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_120 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut121[7] , \nScanOut121[6] , 
        \nScanOut121[5] , \nScanOut121[4] , \nScanOut121[3] , \nScanOut121[2] , 
        \nScanOut121[1] , \nScanOut121[0] }), .ScanOut({\nScanOut120[7] , 
        \nScanOut120[6] , \nScanOut120[5] , \nScanOut120[4] , \nScanOut120[3] , 
        \nScanOut120[2] , \nScanOut120[1] , \nScanOut120[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , 
        \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }), .SouthIn({\nOut7_9[7] , 
        \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , 
        \nOut7_9[1] , \nOut7_9[0] }), .EastIn({\nOut8_8[7] , \nOut8_8[6] , 
        \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , 
        \nOut8_8[0] }), .WestIn({\nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , 
        \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }), 
        .Out({\nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , 
        \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_169 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut170[7] , \nScanOut170[6] , 
        \nScanOut170[5] , \nScanOut170[4] , \nScanOut170[3] , \nScanOut170[2] , 
        \nScanOut170[1] , \nScanOut170[0] }), .ScanOut({\nScanOut169[7] , 
        \nScanOut169[6] , \nScanOut169[5] , \nScanOut169[4] , \nScanOut169[3] , 
        \nScanOut169[2] , \nScanOut169[1] , \nScanOut169[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_8[7] , \nOut10_8[6] , \nOut10_8[5] , \nOut10_8[4] , 
        \nOut10_8[3] , \nOut10_8[2] , \nOut10_8[1] , \nOut10_8[0] }), 
        .SouthIn({\nOut10_10[7] , \nOut10_10[6] , \nOut10_10[5] , 
        \nOut10_10[4] , \nOut10_10[3] , \nOut10_10[2] , \nOut10_10[1] , 
        \nOut10_10[0] }), .EastIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }), .WestIn({\nOut9_9[7] , \nOut9_9[6] , \nOut9_9[5] , 
        \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , \nOut9_9[1] , \nOut9_9[0] }), 
        .Out({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_210 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut211[7] , \nScanOut211[6] , 
        \nScanOut211[5] , \nScanOut211[4] , \nScanOut211[3] , \nScanOut211[2] , 
        \nScanOut211[1] , \nScanOut211[0] }), .ScanOut({\nScanOut210[7] , 
        \nScanOut210[6] , \nScanOut210[5] , \nScanOut210[4] , \nScanOut210[3] , 
        \nScanOut210[2] , \nScanOut210[1] , \nScanOut210[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), 
        .SouthIn({\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .EastIn(
        {\nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), .WestIn(
        {\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .Out({
        \nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_76 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut77[7] , \nScanOut77[6] , 
        \nScanOut77[5] , \nScanOut77[4] , \nScanOut77[3] , \nScanOut77[2] , 
        \nScanOut77[1] , \nScanOut77[0] }), .ScanOut({\nScanOut76[7] , 
        \nScanOut76[6] , \nScanOut76[5] , \nScanOut76[4] , \nScanOut76[3] , 
        \nScanOut76[2] , \nScanOut76[1] , \nScanOut76[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), 
        .SouthIn({\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .EastIn(
        {\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .WestIn(
        {\nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), .Out({
        \nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_88 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut89[7] , \nScanOut89[6] , 
        \nScanOut89[5] , \nScanOut89[4] , \nScanOut89[3] , \nScanOut89[2] , 
        \nScanOut89[1] , \nScanOut89[0] }), .ScanOut({\nScanOut88[7] , 
        \nScanOut88[6] , \nScanOut88[5] , \nScanOut88[4] , \nScanOut88[3] , 
        \nScanOut88[2] , \nScanOut88[1] , \nScanOut88[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , \nOut5_7[4] , \nOut5_7[3] , 
        \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }), .SouthIn({\nOut5_9[7] , 
        \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , 
        \nOut5_9[1] , \nOut5_9[0] }), .EastIn({\nOut6_8[7] , \nOut6_8[6] , 
        \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , 
        \nOut6_8[0] }), .WestIn({\nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , 
        \nOut4_8[4] , \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }), 
        .Out({\nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , \nOut5_8[4] , 
        \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_155 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut156[7] , \nScanOut156[6] , 
        \nScanOut156[5] , \nScanOut156[4] , \nScanOut156[3] , \nScanOut156[2] , 
        \nScanOut156[1] , \nScanOut156[0] }), .ScanOut({\nScanOut155[7] , 
        \nScanOut155[6] , \nScanOut155[5] , \nScanOut155[4] , \nScanOut155[3] , 
        \nScanOut155[2] , \nScanOut155[1] , \nScanOut155[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_10[7] , \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , 
        \nOut9_10[3] , \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), 
        .SouthIn({\nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .EastIn(
        {\nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , 
        \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), 
        .WestIn({\nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .Out({
        \nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_172 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut173[7] , \nScanOut173[6] , 
        \nScanOut173[5] , \nScanOut173[4] , \nScanOut173[3] , \nScanOut173[2] , 
        \nScanOut173[1] , \nScanOut173[0] }), .ScanOut({\nScanOut172[7] , 
        \nScanOut172[6] , \nScanOut172[5] , \nScanOut172[4] , \nScanOut172[3] , 
        \nScanOut172[2] , \nScanOut172[1] , \nScanOut172[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , 
        \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), 
        .SouthIn({\nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , 
        \nOut10_13[4] , \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , 
        \nOut10_13[0] }), .EastIn({\nOut11_12[7] , \nOut11_12[6] , 
        \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , \nOut11_12[2] , 
        \nOut11_12[1] , \nOut11_12[0] }), .WestIn({\nOut9_12[7] , 
        \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , \nOut9_12[3] , 
        \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), .Out({\nOut10_12[7] , 
        \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , \nOut10_12[3] , 
        \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_242 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut243[7] , \nScanOut243[6] , 
        \nScanOut243[5] , \nScanOut243[4] , \nScanOut243[3] , \nScanOut243[2] , 
        \nScanOut243[1] , \nScanOut243[0] }), .ScanOut({\nScanOut242[7] , 
        \nScanOut242[6] , \nScanOut242[5] , \nScanOut242[4] , \nScanOut242[3] , 
        \nScanOut242[2] , \nScanOut242[1] , \nScanOut242[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_2[7] , \nOut15_2[6] , 
        \nOut15_2[5] , \nOut15_2[4] , \nOut15_2[3] , \nOut15_2[2] , 
        \nOut15_2[1] , \nOut15_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_36 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut37[7] , \nScanOut37[6] , 
        \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , 
        \nScanOut37[1] , \nScanOut37[0] }), .ScanOut({\nScanOut36[7] , 
        \nScanOut36[6] , \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , 
        \nScanOut36[2] , \nScanOut36[1] , \nScanOut36[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , 
        \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), .SouthIn({\nOut2_5[7] , 
        \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , 
        \nOut2_5[1] , \nOut2_5[0] }), .EastIn({\nOut3_4[7] , \nOut3_4[6] , 
        \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , 
        \nOut3_4[0] }), .WestIn({\nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , 
        \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), 
        .Out({\nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , 
        \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_197 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut198[7] , \nScanOut198[6] , 
        \nScanOut198[5] , \nScanOut198[4] , \nScanOut198[3] , \nScanOut198[2] , 
        \nScanOut198[1] , \nScanOut198[0] }), .ScanOut({\nScanOut197[7] , 
        \nScanOut197[6] , \nScanOut197[5] , \nScanOut197[4] , \nScanOut197[3] , 
        \nScanOut197[2] , \nScanOut197[1] , \nScanOut197[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), 
        .SouthIn({\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .EastIn(
        {\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .WestIn(
        {\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .Out({
        \nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_185 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut186[7] , \nScanOut186[6] , 
        \nScanOut186[5] , \nScanOut186[4] , \nScanOut186[3] , \nScanOut186[2] , 
        \nScanOut186[1] , \nScanOut186[0] }), .ScanOut({\nScanOut185[7] , 
        \nScanOut185[6] , \nScanOut185[5] , \nScanOut185[4] , \nScanOut185[3] , 
        \nScanOut185[2] , \nScanOut185[1] , \nScanOut185[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), 
        .SouthIn({\nOut11_10[7] , \nOut11_10[6] , \nOut11_10[5] , 
        \nOut11_10[4] , \nOut11_10[3] , \nOut11_10[2] , \nOut11_10[1] , 
        \nOut11_10[0] }), .EastIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }), .WestIn({\nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , 
        \nOut10_9[4] , \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , 
        \nOut10_9[0] }), .Out({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_43 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut44[7] , \nScanOut44[6] , 
        \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , 
        \nScanOut44[1] , \nScanOut44[0] }), .ScanOut({\nScanOut43[7] , 
        \nScanOut43[6] , \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , 
        \nScanOut43[2] , \nScanOut43[1] , \nScanOut43[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_10[7] , \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , 
        \nOut2_10[3] , \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), 
        .SouthIn({\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .EastIn(
        {\nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .WestIn(
        {\nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .Out({
        \nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_58 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut59[7] , \nScanOut59[6] , 
        \nScanOut59[5] , \nScanOut59[4] , \nScanOut59[3] , \nScanOut59[2] , 
        \nScanOut59[1] , \nScanOut59[0] }), .ScanOut({\nScanOut58[7] , 
        \nScanOut58[6] , \nScanOut58[5] , \nScanOut58[4] , \nScanOut58[3] , 
        \nScanOut58[2] , \nScanOut58[1] , \nScanOut58[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_9[7] , \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , 
        \nOut3_9[2] , \nOut3_9[1] , \nOut3_9[0] }), .SouthIn({\nOut3_11[7] , 
        \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , \nOut3_11[3] , 
        \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .EastIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .WestIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .Out({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_129 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut130[7] , \nScanOut130[6] , 
        \nScanOut130[5] , \nScanOut130[4] , \nScanOut130[3] , \nScanOut130[2] , 
        \nScanOut130[1] , \nScanOut130[0] }), .ScanOut({\nScanOut129[7] , 
        \nScanOut129[6] , \nScanOut129[5] , \nScanOut129[4] , \nScanOut129[3] , 
        \nScanOut129[2] , \nScanOut129[1] , \nScanOut129[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_0[7] , \nOut8_0[6] , \nOut8_0[5] , \nOut8_0[4] , \nOut8_0[3] , 
        \nOut8_0[2] , \nOut8_0[1] , \nOut8_0[0] }), .SouthIn({\nOut8_2[7] , 
        \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , \nOut8_2[2] , 
        \nOut8_2[1] , \nOut8_2[0] }), .EastIn({\nOut9_1[7] , \nOut9_1[6] , 
        \nOut9_1[5] , \nOut9_1[4] , \nOut9_1[3] , \nOut9_1[2] , \nOut9_1[1] , 
        \nOut9_1[0] }), .WestIn({\nOut7_1[7] , \nOut7_1[6] , \nOut7_1[5] , 
        \nOut7_1[4] , \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , \nOut7_1[0] }), 
        .Out({\nOut8_1[7] , \nOut8_1[6] , \nOut8_1[5] , \nOut8_1[4] , 
        \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , \nOut8_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_219 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut220[7] , \nScanOut220[6] , 
        \nScanOut220[5] , \nScanOut220[4] , \nScanOut220[3] , \nScanOut220[2] , 
        \nScanOut220[1] , \nScanOut220[0] }), .ScanOut({\nScanOut219[7] , 
        \nScanOut219[6] , \nScanOut219[5] , \nScanOut219[4] , \nScanOut219[3] , 
        \nScanOut219[2] , \nScanOut219[1] , \nScanOut219[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_10[7] , \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , 
        \nOut13_10[3] , \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }), 
        .SouthIn({\nOut13_12[7] , \nOut13_12[6] , \nOut13_12[5] , 
        \nOut13_12[4] , \nOut13_12[3] , \nOut13_12[2] , \nOut13_12[1] , 
        \nOut13_12[0] }), .EastIn({\nOut14_11[7] , \nOut14_11[6] , 
        \nOut14_11[5] , \nOut14_11[4] , \nOut14_11[3] , \nOut14_11[2] , 
        \nOut14_11[1] , \nOut14_11[0] }), .WestIn({\nOut12_11[7] , 
        \nOut12_11[6] , \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , 
        \nOut12_11[2] , \nOut12_11[1] , \nOut12_11[0] }), .Out({\nOut13_11[7] , 
        \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , 
        \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_147 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut148[7] , \nScanOut148[6] , 
        \nScanOut148[5] , \nScanOut148[4] , \nScanOut148[3] , \nScanOut148[2] , 
        \nScanOut148[1] , \nScanOut148[0] }), .ScanOut({\nScanOut147[7] , 
        \nScanOut147[6] , \nScanOut147[5] , \nScanOut147[4] , \nScanOut147[3] , 
        \nScanOut147[2] , \nScanOut147[1] , \nScanOut147[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , 
        \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] }), .SouthIn({\nOut9_4[7] , 
        \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , 
        \nOut9_4[1] , \nOut9_4[0] }), .EastIn({\nOut10_3[7] , \nOut10_3[6] , 
        \nOut10_3[5] , \nOut10_3[4] , \nOut10_3[3] , \nOut10_3[2] , 
        \nOut10_3[1] , \nOut10_3[0] }), .WestIn({\nOut8_3[7] , \nOut8_3[6] , 
        \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , 
        \nOut8_3[0] }), .Out({\nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , 
        \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_160 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut161[7] , \nScanOut161[6] , 
        \nScanOut161[5] , \nScanOut161[4] , \nScanOut161[3] , \nScanOut161[2] , 
        \nScanOut161[1] , \nScanOut161[0] }), .ScanOut({\nScanOut160[7] , 
        \nScanOut160[6] , \nScanOut160[5] , \nScanOut160[4] , \nScanOut160[3] , 
        \nScanOut160[2] , \nScanOut160[1] , \nScanOut160[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut10_0[7] , \nOut10_0[6] , 
        \nOut10_0[5] , \nOut10_0[4] , \nOut10_0[3] , \nOut10_0[2] , 
        \nOut10_0[1] , \nOut10_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_250 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut251[7] , \nScanOut251[6] , 
        \nScanOut251[5] , \nScanOut251[4] , \nScanOut251[3] , \nScanOut251[2] , 
        \nScanOut251[1] , \nScanOut251[0] }), .ScanOut({\nScanOut250[7] , 
        \nScanOut250[6] , \nScanOut250[5] , \nScanOut250[4] , \nScanOut250[3] , 
        \nScanOut250[2] , \nScanOut250[1] , \nScanOut250[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_10[7] , \nOut15_10[6] , 
        \nOut15_10[5] , \nOut15_10[4] , \nOut15_10[3] , \nOut15_10[2] , 
        \nOut15_10[1] , \nOut15_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut8[7] , \nScanOut8[6] , 
        \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , 
        \nScanOut8[1] , \nScanOut8[0] }), .ScanOut({\nScanOut7[7] , 
        \nScanOut7[6] , \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , 
        \nScanOut7[2] , \nScanOut7[1] , \nScanOut7[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_7[7] , \nOut0_7[6] , 
        \nOut0_7[5] , \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , 
        \nOut0_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_26 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut27[7] , \nScanOut27[6] , 
        \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , 
        \nScanOut27[1] , \nScanOut27[0] }), .ScanOut({\nScanOut26[7] , 
        \nScanOut26[6] , \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , 
        \nScanOut26[2] , \nScanOut26[1] , \nScanOut26[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , 
        \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] }), .SouthIn({\nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .EastIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .WestIn({\nOut0_10[7] , 
        \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , 
        \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), .Out({\nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_64 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut65[7] , \nScanOut65[6] , 
        \nScanOut65[5] , \nScanOut65[4] , \nScanOut65[3] , \nScanOut65[2] , 
        \nScanOut65[1] , \nScanOut65[0] }), .ScanOut({\nScanOut64[7] , 
        \nScanOut64[6] , \nScanOut64[5] , \nScanOut64[4] , \nScanOut64[3] , 
        \nScanOut64[2] , \nScanOut64[1] , \nScanOut64[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut4_0[7] , \nOut4_0[6] , 
        \nOut4_0[5] , \nOut4_0[4] , \nOut4_0[3] , \nOut4_0[2] , \nOut4_0[1] , 
        \nOut4_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_81 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut82[7] , \nScanOut82[6] , 
        \nScanOut82[5] , \nScanOut82[4] , \nScanOut82[3] , \nScanOut82[2] , 
        \nScanOut82[1] , \nScanOut82[0] }), .ScanOut({\nScanOut81[7] , 
        \nScanOut81[6] , \nScanOut81[5] , \nScanOut81[4] , \nScanOut81[3] , 
        \nScanOut81[2] , \nScanOut81[1] , \nScanOut81[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_0[7] , \nOut5_0[6] , \nOut5_0[5] , \nOut5_0[4] , \nOut5_0[3] , 
        \nOut5_0[2] , \nOut5_0[1] , \nOut5_0[0] }), .SouthIn({\nOut5_2[7] , 
        \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , 
        \nOut5_2[1] , \nOut5_2[0] }), .EastIn({\nOut6_1[7] , \nOut6_1[6] , 
        \nOut6_1[5] , \nOut6_1[4] , \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , 
        \nOut6_1[0] }), .WestIn({\nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , 
        \nOut4_1[4] , \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }), 
        .Out({\nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , \nOut5_1[4] , 
        \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_115 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut116[7] , \nScanOut116[6] , 
        \nScanOut116[5] , \nScanOut116[4] , \nScanOut116[3] , \nScanOut116[2] , 
        \nScanOut116[1] , \nScanOut116[0] }), .ScanOut({\nScanOut115[7] , 
        \nScanOut115[6] , \nScanOut115[5] , \nScanOut115[4] , \nScanOut115[3] , 
        \nScanOut115[2] , \nScanOut115[1] , \nScanOut115[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , 
        \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }), .SouthIn({\nOut7_4[7] , 
        \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , 
        \nOut7_4[1] , \nOut7_4[0] }), .EastIn({\nOut8_3[7] , \nOut8_3[6] , 
        \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , 
        \nOut8_3[0] }), .WestIn({\nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , 
        \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }), 
        .Out({\nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , 
        \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_225 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut226[7] , \nScanOut226[6] , 
        \nScanOut226[5] , \nScanOut226[4] , \nScanOut226[3] , \nScanOut226[2] , 
        \nScanOut226[1] , \nScanOut226[0] }), .ScanOut({\nScanOut225[7] , 
        \nScanOut225[6] , \nScanOut225[5] , \nScanOut225[4] , \nScanOut225[3] , 
        \nScanOut225[2] , \nScanOut225[1] , \nScanOut225[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_0[7] , \nOut14_0[6] , \nOut14_0[5] , \nOut14_0[4] , 
        \nOut14_0[3] , \nOut14_0[2] , \nOut14_0[1] , \nOut14_0[0] }), 
        .SouthIn({\nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), .EastIn(
        {\nOut15_1[7] , \nOut15_1[6] , \nOut15_1[5] , \nOut15_1[4] , 
        \nOut15_1[3] , \nOut15_1[2] , \nOut15_1[1] , \nOut15_1[0] }), .WestIn(
        {\nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), .Out({
        \nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_132 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut133[7] , \nScanOut133[6] , 
        \nScanOut133[5] , \nScanOut133[4] , \nScanOut133[3] , \nScanOut133[2] , 
        \nScanOut133[1] , \nScanOut133[0] }), .ScanOut({\nScanOut132[7] , 
        \nScanOut132[6] , \nScanOut132[5] , \nScanOut132[4] , \nScanOut132[3] , 
        \nScanOut132[2] , \nScanOut132[1] , \nScanOut132[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_3[7] , \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , 
        \nOut8_3[2] , \nOut8_3[1] , \nOut8_3[0] }), .SouthIn({\nOut8_5[7] , 
        \nOut8_5[6] , \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , 
        \nOut8_5[1] , \nOut8_5[0] }), .EastIn({\nOut9_4[7] , \nOut9_4[6] , 
        \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , \nOut9_4[2] , \nOut9_4[1] , 
        \nOut9_4[0] }), .WestIn({\nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , 
        \nOut7_4[4] , \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }), 
        .Out({\nOut8_4[7] , \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , 
        \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , \nOut8_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_195 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut196[7] , \nScanOut196[6] , 
        \nScanOut196[5] , \nScanOut196[4] , \nScanOut196[3] , \nScanOut196[2] , 
        \nScanOut196[1] , \nScanOut196[0] }), .ScanOut({\nScanOut195[7] , 
        \nScanOut195[6] , \nScanOut195[5] , \nScanOut195[4] , \nScanOut195[3] , 
        \nScanOut195[2] , \nScanOut195[1] , \nScanOut195[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), 
        .SouthIn({\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .EastIn(
        {\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .WestIn(
        {\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .Out({
        \nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_202 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut203[7] , \nScanOut203[6] , 
        \nScanOut203[5] , \nScanOut203[4] , \nScanOut203[3] , \nScanOut203[2] , 
        \nScanOut203[1] , \nScanOut203[0] }), .ScanOut({\nScanOut202[7] , 
        \nScanOut202[6] , \nScanOut202[5] , \nScanOut202[4] , \nScanOut202[3] , 
        \nScanOut202[2] , \nScanOut202[1] , \nScanOut202[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , \nOut12_9[4] , 
        \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , \nOut12_9[0] }), 
        .SouthIn({\nOut12_11[7] , \nOut12_11[6] , \nOut12_11[5] , 
        \nOut12_11[4] , \nOut12_11[3] , \nOut12_11[2] , \nOut12_11[1] , 
        \nOut12_11[0] }), .EastIn({\nOut13_10[7] , \nOut13_10[6] , 
        \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , \nOut13_10[2] , 
        \nOut13_10[1] , \nOut13_10[0] }), .WestIn({\nOut11_10[7] , 
        \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , 
        \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }), .Out({\nOut12_10[7] , 
        \nOut12_10[6] , \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , 
        \nOut12_10[2] , \nOut12_10[1] , \nOut12_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_48 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut49[7] , \nScanOut49[6] , 
        \nScanOut49[5] , \nScanOut49[4] , \nScanOut49[3] , \nScanOut49[2] , 
        \nScanOut49[1] , \nScanOut49[0] }), .ScanOut({\nScanOut48[7] , 
        \nScanOut48[6] , \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , 
        \nScanOut48[2] , \nScanOut48[1] , \nScanOut48[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_0[7] , \nOut3_0[6] , 
        \nOut3_0[5] , \nOut3_0[4] , \nOut3_0[3] , \nOut3_0[2] , \nOut3_0[1] , 
        \nOut3_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_139 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut140[7] , \nScanOut140[6] , 
        \nScanOut140[5] , \nScanOut140[4] , \nScanOut140[3] , \nScanOut140[2] , 
        \nScanOut140[1] , \nScanOut140[0] }), .ScanOut({\nScanOut139[7] , 
        \nScanOut139[6] , \nScanOut139[5] , \nScanOut139[4] , \nScanOut139[3] , 
        \nScanOut139[2] , \nScanOut139[1] , \nScanOut139[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_10[7] , \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , 
        \nOut8_10[3] , \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), 
        .SouthIn({\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .EastIn(
        {\nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .WestIn(
        {\nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .Out({
        \nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_209 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut210[7] , \nScanOut210[6] , 
        \nScanOut210[5] , \nScanOut210[4] , \nScanOut210[3] , \nScanOut210[2] , 
        \nScanOut210[1] , \nScanOut210[0] }), .ScanOut({\nScanOut209[7] , 
        \nScanOut209[6] , \nScanOut209[5] , \nScanOut209[4] , \nScanOut209[3] , 
        \nScanOut209[2] , \nScanOut209[1] , \nScanOut209[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_0[7] , \nOut13_0[6] , \nOut13_0[5] , \nOut13_0[4] , 
        \nOut13_0[3] , \nOut13_0[2] , \nOut13_0[1] , \nOut13_0[0] }), 
        .SouthIn({\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .EastIn(
        {\nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }), .WestIn(
        {\nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), .Out({
        \nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_157 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut158[7] , \nScanOut158[6] , 
        \nScanOut158[5] , \nScanOut158[4] , \nScanOut158[3] , \nScanOut158[2] , 
        \nScanOut158[1] , \nScanOut158[0] }), .ScanOut({\nScanOut157[7] , 
        \nScanOut157[6] , \nScanOut157[5] , \nScanOut157[4] , \nScanOut157[3] , 
        \nScanOut157[2] , \nScanOut157[1] , \nScanOut157[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }), 
        .SouthIn({\nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .EastIn(
        {\nOut10_13[7] , \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , 
        \nOut10_13[3] , \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), 
        .WestIn({\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .Out({
        \nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_170 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut171[7] , \nScanOut171[6] , 
        \nScanOut171[5] , \nScanOut171[4] , \nScanOut171[3] , \nScanOut171[2] , 
        \nScanOut171[1] , \nScanOut171[0] }), .ScanOut({\nScanOut170[7] , 
        \nScanOut170[6] , \nScanOut170[5] , \nScanOut170[4] , \nScanOut170[3] , 
        \nScanOut170[2] , \nScanOut170[1] , \nScanOut170[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_9[7] , \nOut10_9[6] , \nOut10_9[5] , \nOut10_9[4] , 
        \nOut10_9[3] , \nOut10_9[2] , \nOut10_9[1] , \nOut10_9[0] }), 
        .SouthIn({\nOut10_11[7] , \nOut10_11[6] , \nOut10_11[5] , 
        \nOut10_11[4] , \nOut10_11[3] , \nOut10_11[2] , \nOut10_11[1] , 
        \nOut10_11[0] }), .EastIn({\nOut11_10[7] , \nOut11_10[6] , 
        \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , \nOut11_10[2] , 
        \nOut11_10[1] , \nOut11_10[0] }), .WestIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .Out({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_240 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut241[7] , \nScanOut241[6] , 
        \nScanOut241[5] , \nScanOut241[4] , \nScanOut241[3] , \nScanOut241[2] , 
        \nScanOut241[1] , \nScanOut241[0] }), .ScanOut({\nScanOut240[7] , 
        \nScanOut240[6] , \nScanOut240[5] , \nScanOut240[4] , \nScanOut240[3] , 
        \nScanOut240[2] , \nScanOut240[1] , \nScanOut240[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_53 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut54[7] , \nScanOut54[6] , 
        \nScanOut54[5] , \nScanOut54[4] , \nScanOut54[3] , \nScanOut54[2] , 
        \nScanOut54[1] , \nScanOut54[0] }), .ScanOut({\nScanOut53[7] , 
        \nScanOut53[6] , \nScanOut53[5] , \nScanOut53[4] , \nScanOut53[3] , 
        \nScanOut53[2] , \nScanOut53[1] , \nScanOut53[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , \nOut3_4[3] , 
        \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }), .SouthIn({\nOut3_6[7] , 
        \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , \nOut3_6[2] , 
        \nOut3_6[1] , \nOut3_6[0] }), .EastIn({\nOut4_5[7] , \nOut4_5[6] , 
        \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , 
        \nOut4_5[0] }), .WestIn({\nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , 
        \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), 
        .Out({\nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , 
        \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_74 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut75[7] , \nScanOut75[6] , 
        \nScanOut75[5] , \nScanOut75[4] , \nScanOut75[3] , \nScanOut75[2] , 
        \nScanOut75[1] , \nScanOut75[0] }), .ScanOut({\nScanOut74[7] , 
        \nScanOut74[6] , \nScanOut74[5] , \nScanOut74[4] , \nScanOut74[3] , 
        \nScanOut74[2] , \nScanOut74[1] , \nScanOut74[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_9[7] , \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , 
        \nOut4_9[2] , \nOut4_9[1] , \nOut4_9[0] }), .SouthIn({\nOut4_11[7] , 
        \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , \nOut4_11[3] , 
        \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .EastIn({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), .WestIn({\nOut3_10[7] , 
        \nOut3_10[6] , \nOut3_10[5] , \nOut3_10[4] , \nOut3_10[3] , 
        \nOut3_10[2] , \nOut3_10[1] , \nOut3_10[0] }), .Out({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_66 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut67[7] , \nScanOut67[6] , 
        \nScanOut67[5] , \nScanOut67[4] , \nScanOut67[3] , \nScanOut67[2] , 
        \nScanOut67[1] , \nScanOut67[0] }), .ScanOut({\nScanOut66[7] , 
        \nScanOut66[6] , \nScanOut66[5] , \nScanOut66[4] , \nScanOut66[3] , 
        \nScanOut66[2] , \nScanOut66[1] , \nScanOut66[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_1[7] , \nOut4_1[6] , \nOut4_1[5] , \nOut4_1[4] , \nOut4_1[3] , 
        \nOut4_1[2] , \nOut4_1[1] , \nOut4_1[0] }), .SouthIn({\nOut4_3[7] , 
        \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , 
        \nOut4_3[1] , \nOut4_3[0] }), .EastIn({\nOut5_2[7] , \nOut5_2[6] , 
        \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , 
        \nOut5_2[0] }), .WestIn({\nOut3_2[7] , \nOut3_2[6] , \nOut3_2[5] , 
        \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , \nOut3_2[0] }), 
        .Out({\nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , 
        \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_83 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut84[7] , \nScanOut84[6] , 
        \nScanOut84[5] , \nScanOut84[4] , \nScanOut84[3] , \nScanOut84[2] , 
        \nScanOut84[1] , \nScanOut84[0] }), .ScanOut({\nScanOut83[7] , 
        \nScanOut83[6] , \nScanOut83[5] , \nScanOut83[4] , \nScanOut83[3] , 
        \nScanOut83[2] , \nScanOut83[1] , \nScanOut83[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , \nOut5_2[3] , 
        \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }), .SouthIn({\nOut5_4[7] , 
        \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , 
        \nOut5_4[1] , \nOut5_4[0] }), .EastIn({\nOut6_3[7] , \nOut6_3[6] , 
        \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , 
        \nOut6_3[0] }), .WestIn({\nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , 
        \nOut4_3[4] , \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }), 
        .Out({\nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , 
        \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_91 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut92[7] , \nScanOut92[6] , 
        \nScanOut92[5] , \nScanOut92[4] , \nScanOut92[3] , \nScanOut92[2] , 
        \nScanOut92[1] , \nScanOut92[0] }), .ScanOut({\nScanOut91[7] , 
        \nScanOut91[6] , \nScanOut91[5] , \nScanOut91[4] , \nScanOut91[3] , 
        \nScanOut91[2] , \nScanOut91[1] , \nScanOut91[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_10[7] , \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , 
        \nOut5_10[3] , \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }), 
        .SouthIn({\nOut5_12[7] , \nOut5_12[6] , \nOut5_12[5] , \nOut5_12[4] , 
        \nOut5_12[3] , \nOut5_12[2] , \nOut5_12[1] , \nOut5_12[0] }), .EastIn(
        {\nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .WestIn(
        {\nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }), .Out({
        \nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_122 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut123[7] , \nScanOut123[6] , 
        \nScanOut123[5] , \nScanOut123[4] , \nScanOut123[3] , \nScanOut123[2] , 
        \nScanOut123[1] , \nScanOut123[0] }), .ScanOut({\nScanOut122[7] , 
        \nScanOut122[6] , \nScanOut122[5] , \nScanOut122[4] , \nScanOut122[3] , 
        \nScanOut122[2] , \nScanOut122[1] , \nScanOut122[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_9[7] , \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , 
        \nOut7_9[2] , \nOut7_9[1] , \nOut7_9[0] }), .SouthIn({\nOut7_11[7] , 
        \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , \nOut7_11[3] , 
        \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), .EastIn({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .WestIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .Out({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_212 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut213[7] , \nScanOut213[6] , 
        \nScanOut213[5] , \nScanOut213[4] , \nScanOut213[3] , \nScanOut213[2] , 
        \nScanOut213[1] , \nScanOut213[0] }), .ScanOut({\nScanOut212[7] , 
        \nScanOut212[6] , \nScanOut212[5] , \nScanOut212[4] , \nScanOut212[3] , 
        \nScanOut212[2] , \nScanOut212[1] , \nScanOut212[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), 
        .SouthIn({\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .EastIn(
        {\nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), .WestIn(
        {\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .Out({
        \nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_235 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut236[7] , \nScanOut236[6] , 
        \nScanOut236[5] , \nScanOut236[4] , \nScanOut236[3] , \nScanOut236[2] , 
        \nScanOut236[1] , \nScanOut236[0] }), .ScanOut({\nScanOut235[7] , 
        \nScanOut235[6] , \nScanOut235[5] , \nScanOut235[4] , \nScanOut235[3] , 
        \nScanOut235[2] , \nScanOut235[1] , \nScanOut235[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_10[7] , \nOut14_10[6] , \nOut14_10[5] , \nOut14_10[4] , 
        \nOut14_10[3] , \nOut14_10[2] , \nOut14_10[1] , \nOut14_10[0] }), 
        .SouthIn({\nOut14_12[7] , \nOut14_12[6] , \nOut14_12[5] , 
        \nOut14_12[4] , \nOut14_12[3] , \nOut14_12[2] , \nOut14_12[1] , 
        \nOut14_12[0] }), .EastIn({\nOut15_11[7] , \nOut15_11[6] , 
        \nOut15_11[5] , \nOut15_11[4] , \nOut15_11[3] , \nOut15_11[2] , 
        \nOut15_11[1] , \nOut15_11[0] }), .WestIn({\nOut13_11[7] , 
        \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , \nOut13_11[3] , 
        \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }), .Out({\nOut14_11[7] , 
        \nOut14_11[6] , \nOut14_11[5] , \nOut14_11[4] , \nOut14_11[3] , 
        \nOut14_11[2] , \nOut14_11[1] , \nOut14_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_105 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut106[7] , \nScanOut106[6] , 
        \nScanOut106[5] , \nScanOut106[4] , \nScanOut106[3] , \nScanOut106[2] , 
        \nScanOut106[1] , \nScanOut106[0] }), .ScanOut({\nScanOut105[7] , 
        \nScanOut105[6] , \nScanOut105[5] , \nScanOut105[4] , \nScanOut105[3] , 
        \nScanOut105[2] , \nScanOut105[1] , \nScanOut105[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , 
        \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }), .SouthIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .EastIn({\nOut7_9[7] , 
        \nOut7_9[6] , \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , 
        \nOut7_9[1] , \nOut7_9[0] }), .WestIn({\nOut5_9[7] , \nOut5_9[6] , 
        \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , \nOut5_9[1] , 
        \nOut5_9[0] }), .Out({\nOut6_9[7] , \nOut6_9[6] , \nOut6_9[5] , 
        \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , \nOut6_9[1] , \nOut6_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_130 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut131[7] , \nScanOut131[6] , 
        \nScanOut131[5] , \nScanOut131[4] , \nScanOut131[3] , \nScanOut131[2] , 
        \nScanOut131[1] , \nScanOut131[0] }), .ScanOut({\nScanOut130[7] , 
        \nScanOut130[6] , \nScanOut130[5] , \nScanOut130[4] , \nScanOut130[3] , 
        \nScanOut130[2] , \nScanOut130[1] , \nScanOut130[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_1[7] , \nOut8_1[6] , \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , 
        \nOut8_1[2] , \nOut8_1[1] , \nOut8_1[0] }), .SouthIn({\nOut8_3[7] , 
        \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , \nOut8_3[3] , \nOut8_3[2] , 
        \nOut8_3[1] , \nOut8_3[0] }), .EastIn({\nOut9_2[7] , \nOut9_2[6] , 
        \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , \nOut9_2[1] , 
        \nOut9_2[0] }), .WestIn({\nOut7_2[7] , \nOut7_2[6] , \nOut7_2[5] , 
        \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , \nOut7_2[0] }), 
        .Out({\nOut8_2[7] , \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , 
        \nOut8_2[3] , \nOut8_2[2] , \nOut8_2[1] , \nOut8_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_200 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut201[7] , \nScanOut201[6] , 
        \nScanOut201[5] , \nScanOut201[4] , \nScanOut201[3] , \nScanOut201[2] , 
        \nScanOut201[1] , \nScanOut201[0] }), .ScanOut({\nScanOut200[7] , 
        \nScanOut200[6] , \nScanOut200[5] , \nScanOut200[4] , \nScanOut200[3] , 
        \nScanOut200[2] , \nScanOut200[1] , \nScanOut200[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), 
        .SouthIn({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , \nOut12_9[4] , 
        \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , \nOut12_9[0] }), .EastIn(
        {\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .WestIn(
        {\nOut11_8[7] , \nOut11_8[6] , \nOut11_8[5] , \nOut11_8[4] , 
        \nOut11_8[3] , \nOut11_8[2] , \nOut11_8[1] , \nOut11_8[0] }), .Out({
        \nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_227 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut228[7] , \nScanOut228[6] , 
        \nScanOut228[5] , \nScanOut228[4] , \nScanOut228[3] , \nScanOut228[2] , 
        \nScanOut228[1] , \nScanOut228[0] }), .ScanOut({\nScanOut227[7] , 
        \nScanOut227[6] , \nScanOut227[5] , \nScanOut227[4] , \nScanOut227[3] , 
        \nScanOut227[2] , \nScanOut227[1] , \nScanOut227[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }), 
        .SouthIn({\nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), .EastIn(
        {\nOut15_3[7] , \nOut15_3[6] , \nOut15_3[5] , \nOut15_3[4] , 
        \nOut15_3[3] , \nOut15_3[2] , \nOut15_3[1] , \nOut15_3[0] }), .WestIn(
        {\nOut13_3[7] , \nOut13_3[6] , \nOut13_3[5] , \nOut13_3[4] , 
        \nOut13_3[3] , \nOut13_3[2] , \nOut13_3[1] , \nOut13_3[0] }), .Out({
        \nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_117 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut118[7] , \nScanOut118[6] , 
        \nScanOut118[5] , \nScanOut118[4] , \nScanOut118[3] , \nScanOut118[2] , 
        \nScanOut118[1] , \nScanOut118[0] }), .ScanOut({\nScanOut117[7] , 
        \nScanOut117[6] , \nScanOut117[5] , \nScanOut117[4] , \nScanOut117[3] , 
        \nScanOut117[2] , \nScanOut117[1] , \nScanOut117[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , \nOut7_4[3] , 
        \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }), .SouthIn({\nOut7_6[7] , 
        \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , 
        \nOut7_6[1] , \nOut7_6[0] }), .EastIn({\nOut8_5[7] , \nOut8_5[6] , 
        \nOut8_5[5] , \nOut8_5[4] , \nOut8_5[3] , \nOut8_5[2] , \nOut8_5[1] , 
        \nOut8_5[0] }), .WestIn({\nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , 
        \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }), 
        .Out({\nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , 
        \nOut7_5[3] , \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_179 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut180[7] , \nScanOut180[6] , 
        \nScanOut180[5] , \nScanOut180[4] , \nScanOut180[3] , \nScanOut180[2] , 
        \nScanOut180[1] , \nScanOut180[0] }), .ScanOut({\nScanOut179[7] , 
        \nScanOut179[6] , \nScanOut179[5] , \nScanOut179[4] , \nScanOut179[3] , 
        \nScanOut179[2] , \nScanOut179[1] , \nScanOut179[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), 
        .SouthIn({\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .EastIn(
        {\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .WestIn(
        {\nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), .Out({
        \nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_249 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut250[7] , \nScanOut250[6] , 
        \nScanOut250[5] , \nScanOut250[4] , \nScanOut250[3] , \nScanOut250[2] , 
        \nScanOut250[1] , \nScanOut250[0] }), .ScanOut({\nScanOut249[7] , 
        \nScanOut249[6] , \nScanOut249[5] , \nScanOut249[4] , \nScanOut249[3] , 
        \nScanOut249[2] , \nScanOut249[1] , \nScanOut249[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_9[7] , \nOut15_9[6] , 
        \nOut15_9[5] , \nOut15_9[4] , \nOut15_9[3] , \nOut15_9[2] , 
        \nOut15_9[1] , \nOut15_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut14[7] , \nScanOut14[6] , 
        \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , 
        \nScanOut14[1] , \nScanOut14[0] }), .ScanOut({\nScanOut13[7] , 
        \nScanOut13[6] , \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , 
        \nScanOut13[2] , \nScanOut13[1] , \nScanOut13[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_13[7] , \nOut0_13[6] , 
        \nOut0_13[5] , \nOut0_13[4] , \nOut0_13[3] , \nOut0_13[2] , 
        \nOut0_13[1] , \nOut0_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_41 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut42[7] , \nScanOut42[6] , 
        \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , 
        \nScanOut42[1] , \nScanOut42[0] }), .ScanOut({\nScanOut41[7] , 
        \nScanOut41[6] , \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , 
        \nScanOut41[2] , \nScanOut41[1] , \nScanOut41[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , 
        \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), .SouthIn({\nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .EastIn({\nOut3_9[7] , 
        \nOut3_9[6] , \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , 
        \nOut3_9[1] , \nOut3_9[0] }), .WestIn({\nOut1_9[7] , \nOut1_9[6] , 
        \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , 
        \nOut1_9[0] }), .Out({\nOut2_9[7] , \nOut2_9[6] , \nOut2_9[5] , 
        \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , \nOut2_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_98 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut99[7] , \nScanOut99[6] , 
        \nScanOut99[5] , \nScanOut99[4] , \nScanOut99[3] , \nScanOut99[2] , 
        \nScanOut99[1] , \nScanOut99[0] }), .ScanOut({\nScanOut98[7] , 
        \nScanOut98[6] , \nScanOut98[5] , \nScanOut98[4] , \nScanOut98[3] , 
        \nScanOut98[2] , \nScanOut98[1] , \nScanOut98[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , \nOut6_1[4] , \nOut6_1[3] , 
        \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }), .SouthIn({\nOut6_3[7] , 
        \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , \nOut6_3[3] , \nOut6_3[2] , 
        \nOut6_3[1] , \nOut6_3[0] }), .EastIn({\nOut7_2[7] , \nOut7_2[6] , 
        \nOut7_2[5] , \nOut7_2[4] , \nOut7_2[3] , \nOut7_2[2] , \nOut7_2[1] , 
        \nOut7_2[0] }), .WestIn({\nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , 
        \nOut5_2[4] , \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }), 
        .Out({\nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , 
        \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_145 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut146[7] , \nScanOut146[6] , 
        \nScanOut146[5] , \nScanOut146[4] , \nScanOut146[3] , \nScanOut146[2] , 
        \nScanOut146[1] , \nScanOut146[0] }), .ScanOut({\nScanOut145[7] , 
        \nScanOut145[6] , \nScanOut145[5] , \nScanOut145[4] , \nScanOut145[3] , 
        \nScanOut145[2] , \nScanOut145[1] , \nScanOut145[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_0[7] , \nOut9_0[6] , \nOut9_0[5] , \nOut9_0[4] , \nOut9_0[3] , 
        \nOut9_0[2] , \nOut9_0[1] , \nOut9_0[0] }), .SouthIn({\nOut9_2[7] , 
        \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , \nOut9_2[2] , 
        \nOut9_2[1] , \nOut9_2[0] }), .EastIn({\nOut10_1[7] , \nOut10_1[6] , 
        \nOut10_1[5] , \nOut10_1[4] , \nOut10_1[3] , \nOut10_1[2] , 
        \nOut10_1[1] , \nOut10_1[0] }), .WestIn({\nOut8_1[7] , \nOut8_1[6] , 
        \nOut8_1[5] , \nOut8_1[4] , \nOut8_1[3] , \nOut8_1[2] , \nOut8_1[1] , 
        \nOut8_1[0] }), .Out({\nOut9_1[7] , \nOut9_1[6] , \nOut9_1[5] , 
        \nOut9_1[4] , \nOut9_1[3] , \nOut9_1[2] , \nOut9_1[1] , \nOut9_1[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_162 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut163[7] , \nScanOut163[6] , 
        \nScanOut163[5] , \nScanOut163[4] , \nScanOut163[3] , \nScanOut163[2] , 
        \nScanOut163[1] , \nScanOut163[0] }), .ScanOut({\nScanOut162[7] , 
        \nScanOut162[6] , \nScanOut162[5] , \nScanOut162[4] , \nScanOut162[3] , 
        \nScanOut162[2] , \nScanOut162[1] , \nScanOut162[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_1[7] , \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , 
        \nOut10_1[3] , \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }), 
        .SouthIn({\nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), .EastIn(
        {\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .WestIn(
        {\nOut9_2[7] , \nOut9_2[6] , \nOut9_2[5] , \nOut9_2[4] , \nOut9_2[3] , 
        \nOut9_2[2] , \nOut9_2[1] , \nOut9_2[0] }), .Out({\nOut10_2[7] , 
        \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , \nOut10_2[3] , 
        \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_252 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut253[7] , \nScanOut253[6] , 
        \nScanOut253[5] , \nScanOut253[4] , \nScanOut253[3] , \nScanOut253[2] , 
        \nScanOut253[1] , \nScanOut253[0] }), .ScanOut({\nScanOut252[7] , 
        \nScanOut252[6] , \nScanOut252[5] , \nScanOut252[4] , \nScanOut252[3] , 
        \nScanOut252[2] , \nScanOut252[1] , \nScanOut252[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_12[7] , \nOut15_12[6] , 
        \nOut15_12[5] , \nOut15_12[4] , \nOut15_12[3] , \nOut15_12[2] , 
        \nOut15_12[1] , \nOut15_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut15[7] , \nScanOut15[6] , 
        \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , 
        \nScanOut15[1] , \nScanOut15[0] }), .ScanOut({\nScanOut14[7] , 
        \nScanOut14[6] , \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , 
        \nScanOut14[2] , \nScanOut14[1] , \nScanOut14[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_14[7] , \nOut0_14[6] , 
        \nOut0_14[5] , \nOut0_14[4] , \nOut0_14[3] , \nOut0_14[2] , 
        \nOut0_14[1] , \nOut0_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_33 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut34[7] , \nScanOut34[6] , 
        \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , 
        \nScanOut34[1] , \nScanOut34[0] }), .ScanOut({\nScanOut33[7] , 
        \nScanOut33[6] , \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , 
        \nScanOut33[2] , \nScanOut33[1] , \nScanOut33[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_0[7] , \nOut2_0[6] , \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , 
        \nOut2_0[2] , \nOut2_0[1] , \nOut2_0[0] }), .SouthIn({\nOut2_2[7] , 
        \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , 
        \nOut2_2[1] , \nOut2_2[0] }), .EastIn({\nOut3_1[7] , \nOut3_1[6] , 
        \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , 
        \nOut3_1[0] }), .WestIn({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , 
        \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), 
        .Out({\nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , 
        \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_34 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut35[7] , \nScanOut35[6] , 
        \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , 
        \nScanOut35[1] , \nScanOut35[0] }), .ScanOut({\nScanOut34[7] , 
        \nScanOut34[6] , \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , 
        \nScanOut34[2] , \nScanOut34[1] , \nScanOut34[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , 
        \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), .SouthIn({\nOut2_3[7] , 
        \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , 
        \nOut2_3[1] , \nOut2_3[0] }), .EastIn({\nOut3_2[7] , \nOut3_2[6] , 
        \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , 
        \nOut3_2[0] }), .WestIn({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , 
        \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), 
        .Out({\nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , 
        \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_187 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut188[7] , \nScanOut188[6] , 
        \nScanOut188[5] , \nScanOut188[4] , \nScanOut188[3] , \nScanOut188[2] , 
        \nScanOut188[1] , \nScanOut188[0] }), .ScanOut({\nScanOut187[7] , 
        \nScanOut187[6] , \nScanOut187[5] , \nScanOut187[4] , \nScanOut187[3] , 
        \nScanOut187[2] , \nScanOut187[1] , \nScanOut187[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_10[7] , \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , 
        \nOut11_10[3] , \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }), 
        .SouthIn({\nOut11_12[7] , \nOut11_12[6] , \nOut11_12[5] , 
        \nOut11_12[4] , \nOut11_12[3] , \nOut11_12[2] , \nOut11_12[1] , 
        \nOut11_12[0] }), .EastIn({\nOut12_11[7] , \nOut12_11[6] , 
        \nOut12_11[5] , \nOut12_11[4] , \nOut12_11[3] , \nOut12_11[2] , 
        \nOut12_11[1] , \nOut12_11[0] }), .WestIn({\nOut10_11[7] , 
        \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , \nOut10_11[3] , 
        \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }), .Out({\nOut11_11[7] , 
        \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , 
        \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_180 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut181[7] , \nScanOut181[6] , 
        \nScanOut181[5] , \nScanOut181[4] , \nScanOut181[3] , \nScanOut181[2] , 
        \nScanOut181[1] , \nScanOut181[0] }), .ScanOut({\nScanOut180[7] , 
        \nScanOut180[6] , \nScanOut180[5] , \nScanOut180[4] , \nScanOut180[3] , 
        \nScanOut180[2] , \nScanOut180[1] , \nScanOut180[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), 
        .SouthIn({\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .EastIn(
        {\nOut12_4[7] , \nOut12_4[6] , \nOut12_4[5] , \nOut12_4[4] , 
        \nOut12_4[3] , \nOut12_4[2] , \nOut12_4[1] , \nOut12_4[0] }), .WestIn(
        {\nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), .Out({
        \nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_46 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut47[7] , \nScanOut47[6] , 
        \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , 
        \nScanOut47[1] , \nScanOut47[0] }), .ScanOut({\nScanOut46[7] , 
        \nScanOut46[6] , \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , 
        \nScanOut46[2] , \nScanOut46[1] , \nScanOut46[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), 
        .SouthIn({\nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , 
        \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), .EastIn(
        {\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .WestIn(
        {\nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .Out({
        \nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_142 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut143[7] , \nScanOut143[6] , 
        \nScanOut143[5] , \nScanOut143[4] , \nScanOut143[3] , \nScanOut143[2] , 
        \nScanOut143[1] , \nScanOut143[0] }), .ScanOut({\nScanOut142[7] , 
        \nScanOut142[6] , \nScanOut142[5] , \nScanOut142[4] , \nScanOut142[3] , 
        \nScanOut142[2] , \nScanOut142[1] , \nScanOut142[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), 
        .SouthIn({\nOut8_15[7] , \nOut8_15[6] , \nOut8_15[5] , \nOut8_15[4] , 
        \nOut8_15[3] , \nOut8_15[2] , \nOut8_15[1] , \nOut8_15[0] }), .EastIn(
        {\nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }), .WestIn(
        {\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .Out({
        \nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_165 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut166[7] , \nScanOut166[6] , 
        \nScanOut166[5] , \nScanOut166[4] , \nScanOut166[3] , \nScanOut166[2] , 
        \nScanOut166[1] , \nScanOut166[0] }), .ScanOut({\nScanOut165[7] , 
        \nScanOut165[6] , \nScanOut165[5] , \nScanOut165[4] , \nScanOut165[3] , 
        \nScanOut165[2] , \nScanOut165[1] , \nScanOut165[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), 
        .SouthIn({\nOut10_6[7] , \nOut10_6[6] , \nOut10_6[5] , \nOut10_6[4] , 
        \nOut10_6[3] , \nOut10_6[2] , \nOut10_6[1] , \nOut10_6[0] }), .EastIn(
        {\nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }), .WestIn(
        {\nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , 
        \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] }), .Out({\nOut10_5[7] , 
        \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , \nOut10_5[3] , 
        \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_255 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut256[7] , \nScanOut256[6] , 
        \nScanOut256[5] , \nScanOut256[4] , \nScanOut256[3] , \nScanOut256[2] , 
        \nScanOut256[1] , \nScanOut256[0] }), .ScanOut({\nScanOut255[7] , 
        \nScanOut255[6] , \nScanOut255[5] , \nScanOut255[4] , \nScanOut255[3] , 
        \nScanOut255[2] , \nScanOut255[1] , \nScanOut255[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_159 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut160[7] , \nScanOut160[6] , 
        \nScanOut160[5] , \nScanOut160[4] , \nScanOut160[3] , \nScanOut160[2] , 
        \nScanOut160[1] , \nScanOut160[0] }), .ScanOut({\nScanOut159[7] , 
        \nScanOut159[6] , \nScanOut159[5] , \nScanOut159[4] , \nScanOut159[3] , 
        \nScanOut159[2] , \nScanOut159[1] , \nScanOut159[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut9_15[7] , \nOut9_15[6] , 
        \nOut9_15[5] , \nOut9_15[4] , \nOut9_15[3] , \nOut9_15[2] , 
        \nOut9_15[1] , \nOut9_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut2[7] , \nScanOut2[6] , 
        \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , 
        \nScanOut2[1] , \nScanOut2[0] }), .ScanOut({\nScanOut1[7] , 
        \nScanOut1[6] , \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , 
        \nScanOut1[2] , \nScanOut1[1] , \nScanOut1[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_1[7] , \nOut0_1[6] , 
        \nOut0_1[5] , \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , 
        \nOut0_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut10[7] , \nScanOut10[6] , 
        \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , 
        \nScanOut10[1] , \nScanOut10[0] }), .ScanOut({\nScanOut9[7] , 
        \nScanOut9[6] , \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , 
        \nScanOut9[2] , \nScanOut9[1] , \nScanOut9[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_28 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut29[7] , \nScanOut29[6] , 
        \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , 
        \nScanOut29[1] , \nScanOut29[0] }), .ScanOut({\nScanOut28[7] , 
        \nScanOut28[6] , \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , 
        \nScanOut28[2] , \nScanOut28[1] , \nScanOut28[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), 
        .SouthIn({\nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .EastIn(
        {\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .WestIn(
        {\nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , 
        \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), .Out({
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_61 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut62[7] , \nScanOut62[6] , 
        \nScanOut62[5] , \nScanOut62[4] , \nScanOut62[3] , \nScanOut62[2] , 
        \nScanOut62[1] , \nScanOut62[0] }), .ScanOut({\nScanOut61[7] , 
        \nScanOut61[6] , \nScanOut61[5] , \nScanOut61[4] , \nScanOut61[3] , 
        \nScanOut61[2] , \nScanOut61[1] , \nScanOut61[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }), 
        .SouthIn({\nOut3_14[7] , \nOut3_14[6] , \nOut3_14[5] , \nOut3_14[4] , 
        \nOut3_14[3] , \nOut3_14[2] , \nOut3_14[1] , \nOut3_14[0] }), .EastIn(
        {\nOut4_13[7] , \nOut4_13[6] , \nOut4_13[5] , \nOut4_13[4] , 
        \nOut4_13[3] , \nOut4_13[2] , \nOut4_13[1] , \nOut4_13[0] }), .WestIn(
        {\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .Out({
        \nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_54 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut55[7] , \nScanOut55[6] , 
        \nScanOut55[5] , \nScanOut55[4] , \nScanOut55[3] , \nScanOut55[2] , 
        \nScanOut55[1] , \nScanOut55[0] }), .ScanOut({\nScanOut54[7] , 
        \nScanOut54[6] , \nScanOut54[5] , \nScanOut54[4] , \nScanOut54[3] , 
        \nScanOut54[2] , \nScanOut54[1] , \nScanOut54[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , 
        \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }), .SouthIn({\nOut3_7[7] , 
        \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , \nOut3_7[3] , \nOut3_7[2] , 
        \nOut3_7[1] , \nOut3_7[0] }), .EastIn({\nOut4_6[7] , \nOut4_6[6] , 
        \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , \nOut4_6[1] , 
        \nOut4_6[0] }), .WestIn({\nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , 
        \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), 
        .Out({\nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , 
        \nOut3_6[3] , \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_84 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut85[7] , \nScanOut85[6] , 
        \nScanOut85[5] , \nScanOut85[4] , \nScanOut85[3] , \nScanOut85[2] , 
        \nScanOut85[1] , \nScanOut85[0] }), .ScanOut({\nScanOut84[7] , 
        \nScanOut84[6] , \nScanOut84[5] , \nScanOut84[4] , \nScanOut84[3] , 
        \nScanOut84[2] , \nScanOut84[1] , \nScanOut84[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , 
        \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }), .SouthIn({\nOut5_5[7] , 
        \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , 
        \nOut5_5[1] , \nOut5_5[0] }), .EastIn({\nOut6_4[7] , \nOut6_4[6] , 
        \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , 
        \nOut6_4[0] }), .WestIn({\nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , 
        \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }), 
        .Out({\nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , 
        \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_110 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut111[7] , \nScanOut111[6] , 
        \nScanOut111[5] , \nScanOut111[4] , \nScanOut111[3] , \nScanOut111[2] , 
        \nScanOut111[1] , \nScanOut111[0] }), .ScanOut({\nScanOut110[7] , 
        \nScanOut110[6] , \nScanOut110[5] , \nScanOut110[4] , \nScanOut110[3] , 
        \nScanOut110[2] , \nScanOut110[1] , \nScanOut110[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), 
        .SouthIn({\nOut6_15[7] , \nOut6_15[6] , \nOut6_15[5] , \nOut6_15[4] , 
        \nOut6_15[3] , \nOut6_15[2] , \nOut6_15[1] , \nOut6_15[0] }), .EastIn(
        {\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .WestIn(
        {\nOut5_14[7] , \nOut5_14[6] , \nOut5_14[5] , \nOut5_14[4] , 
        \nOut5_14[3] , \nOut5_14[2] , \nOut5_14[1] , \nOut5_14[0] }), .Out({
        \nOut6_14[7] , \nOut6_14[6] , \nOut6_14[5] , \nOut6_14[4] , 
        \nOut6_14[3] , \nOut6_14[2] , \nOut6_14[1] , \nOut6_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_96 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut97[7] , \nScanOut97[6] , 
        \nScanOut97[5] , \nScanOut97[4] , \nScanOut97[3] , \nScanOut97[2] , 
        \nScanOut97[1] , \nScanOut97[0] }), .ScanOut({\nScanOut96[7] , 
        \nScanOut96[6] , \nScanOut96[5] , \nScanOut96[4] , \nScanOut96[3] , 
        \nScanOut96[2] , \nScanOut96[1] , \nScanOut96[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut6_0[7] , \nOut6_0[6] , 
        \nOut6_0[5] , \nOut6_0[4] , \nOut6_0[3] , \nOut6_0[2] , \nOut6_0[1] , 
        \nOut6_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_102 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut103[7] , \nScanOut103[6] , 
        \nScanOut103[5] , \nScanOut103[4] , \nScanOut103[3] , \nScanOut103[2] , 
        \nScanOut103[1] , \nScanOut103[0] }), .ScanOut({\nScanOut102[7] , 
        \nScanOut102[6] , \nScanOut102[5] , \nScanOut102[4] , \nScanOut102[3] , 
        \nScanOut102[2] , \nScanOut102[1] , \nScanOut102[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_5[7] , \nOut6_5[6] , \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , 
        \nOut6_5[2] , \nOut6_5[1] , \nOut6_5[0] }), .SouthIn({\nOut6_7[7] , 
        \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , 
        \nOut6_7[1] , \nOut6_7[0] }), .EastIn({\nOut7_6[7] , \nOut7_6[6] , 
        \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , 
        \nOut7_6[0] }), .WestIn({\nOut5_6[7] , \nOut5_6[6] , \nOut5_6[5] , 
        \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , \nOut5_6[1] , \nOut5_6[0] }), 
        .Out({\nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , 
        \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_137 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut138[7] , \nScanOut138[6] , 
        \nScanOut138[5] , \nScanOut138[4] , \nScanOut138[3] , \nScanOut138[2] , 
        \nScanOut138[1] , \nScanOut138[0] }), .ScanOut({\nScanOut137[7] , 
        \nScanOut137[6] , \nScanOut137[5] , \nScanOut137[4] , \nScanOut137[3] , 
        \nScanOut137[2] , \nScanOut137[1] , \nScanOut137[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_8[7] , \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , \nOut8_8[3] , 
        \nOut8_8[2] , \nOut8_8[1] , \nOut8_8[0] }), .SouthIn({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }), .EastIn({\nOut9_9[7] , 
        \nOut9_9[6] , \nOut9_9[5] , \nOut9_9[4] , \nOut9_9[3] , \nOut9_9[2] , 
        \nOut9_9[1] , \nOut9_9[0] }), .WestIn({\nOut7_9[7] , \nOut7_9[6] , 
        \nOut7_9[5] , \nOut7_9[4] , \nOut7_9[3] , \nOut7_9[2] , \nOut7_9[1] , 
        \nOut7_9[0] }), .Out({\nOut8_9[7] , \nOut8_9[6] , \nOut8_9[5] , 
        \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , \nOut8_9[1] , \nOut8_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_207 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut208[7] , \nScanOut208[6] , 
        \nScanOut208[5] , \nScanOut208[4] , \nScanOut208[3] , \nScanOut208[2] , 
        \nScanOut208[1] , \nScanOut208[0] }), .ScanOut({\nScanOut207[7] , 
        \nScanOut207[6] , \nScanOut207[5] , \nScanOut207[4] , \nScanOut207[3] , 
        \nScanOut207[2] , \nScanOut207[1] , \nScanOut207[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut12_15[7] , \nOut12_15[6] , 
        \nOut12_15[5] , \nOut12_15[4] , \nOut12_15[3] , \nOut12_15[2] , 
        \nOut12_15[1] , \nOut12_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_220 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut221[7] , \nScanOut221[6] , 
        \nScanOut221[5] , \nScanOut221[4] , \nScanOut221[3] , \nScanOut221[2] , 
        \nScanOut221[1] , \nScanOut221[0] }), .ScanOut({\nScanOut220[7] , 
        \nScanOut220[6] , \nScanOut220[5] , \nScanOut220[4] , \nScanOut220[3] , 
        \nScanOut220[2] , \nScanOut220[1] , \nScanOut220[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_11[7] , \nOut13_11[6] , \nOut13_11[5] , \nOut13_11[4] , 
        \nOut13_11[3] , \nOut13_11[2] , \nOut13_11[1] , \nOut13_11[0] }), 
        .SouthIn({\nOut13_13[7] , \nOut13_13[6] , \nOut13_13[5] , 
        \nOut13_13[4] , \nOut13_13[3] , \nOut13_13[2] , \nOut13_13[1] , 
        \nOut13_13[0] }), .EastIn({\nOut14_12[7] , \nOut14_12[6] , 
        \nOut14_12[5] , \nOut14_12[4] , \nOut14_12[3] , \nOut14_12[2] , 
        \nOut14_12[1] , \nOut14_12[0] }), .WestIn({\nOut12_12[7] , 
        \nOut12_12[6] , \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , 
        \nOut12_12[2] , \nOut12_12[1] , \nOut12_12[0] }), .Out({\nOut13_12[7] , 
        \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , \nOut13_12[3] , 
        \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_125 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut126[7] , \nScanOut126[6] , 
        \nScanOut126[5] , \nScanOut126[4] , \nScanOut126[3] , \nScanOut126[2] , 
        \nScanOut126[1] , \nScanOut126[0] }), .ScanOut({\nScanOut125[7] , 
        \nScanOut125[6] , \nScanOut125[5] , \nScanOut125[4] , \nScanOut125[3] , 
        \nScanOut125[2] , \nScanOut125[1] , \nScanOut125[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), 
        .SouthIn({\nOut7_14[7] , \nOut7_14[6] , \nOut7_14[5] , \nOut7_14[4] , 
        \nOut7_14[3] , \nOut7_14[2] , \nOut7_14[1] , \nOut7_14[0] }), .EastIn(
        {\nOut8_13[7] , \nOut8_13[6] , \nOut8_13[5] , \nOut8_13[4] , 
        \nOut8_13[3] , \nOut8_13[2] , \nOut8_13[1] , \nOut8_13[0] }), .WestIn(
        {\nOut6_13[7] , \nOut6_13[6] , \nOut6_13[5] , \nOut6_13[4] , 
        \nOut6_13[3] , \nOut6_13[2] , \nOut6_13[1] , \nOut6_13[0] }), .Out({
        \nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_215 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut216[7] , \nScanOut216[6] , 
        \nScanOut216[5] , \nScanOut216[4] , \nScanOut216[3] , \nScanOut216[2] , 
        \nScanOut216[1] , \nScanOut216[0] }), .ScanOut({\nScanOut215[7] , 
        \nScanOut215[6] , \nScanOut215[5] , \nScanOut215[4] , \nScanOut215[3] , 
        \nScanOut215[2] , \nScanOut215[1] , \nScanOut215[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), 
        .SouthIn({\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .EastIn(
        {\nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), .WestIn(
        {\nOut12_7[7] , \nOut12_7[6] , \nOut12_7[5] , \nOut12_7[4] , 
        \nOut12_7[3] , \nOut12_7[2] , \nOut12_7[1] , \nOut12_7[0] }), .Out({
        \nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_232 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut233[7] , \nScanOut233[6] , 
        \nScanOut233[5] , \nScanOut233[4] , \nScanOut233[3] , \nScanOut233[2] , 
        \nScanOut233[1] , \nScanOut233[0] }), .ScanOut({\nScanOut232[7] , 
        \nScanOut232[6] , \nScanOut232[5] , \nScanOut232[4] , \nScanOut232[3] , 
        \nScanOut232[2] , \nScanOut232[1] , \nScanOut232[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_7[7] , \nOut14_7[6] , \nOut14_7[5] , \nOut14_7[4] , 
        \nOut14_7[3] , \nOut14_7[2] , \nOut14_7[1] , \nOut14_7[0] }), 
        .SouthIn({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , \nOut14_9[4] , 
        \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , \nOut14_9[0] }), .EastIn(
        {\nOut15_8[7] , \nOut15_8[6] , \nOut15_8[5] , \nOut15_8[4] , 
        \nOut15_8[3] , \nOut15_8[2] , \nOut15_8[1] , \nOut15_8[0] }), .WestIn(
        {\nOut13_8[7] , \nOut13_8[6] , \nOut13_8[5] , \nOut13_8[4] , 
        \nOut13_8[3] , \nOut13_8[2] , \nOut13_8[1] , \nOut13_8[0] }), .Out({
        \nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_189 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut190[7] , \nScanOut190[6] , 
        \nScanOut190[5] , \nScanOut190[4] , \nScanOut190[3] , \nScanOut190[2] , 
        \nScanOut190[1] , \nScanOut190[0] }), .ScanOut({\nScanOut189[7] , 
        \nScanOut189[6] , \nScanOut189[5] , \nScanOut189[4] , \nScanOut189[3] , 
        \nScanOut189[2] , \nScanOut189[1] , \nScanOut189[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_12[7] , \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , 
        \nOut11_12[3] , \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }), 
        .SouthIn({\nOut11_14[7] , \nOut11_14[6] , \nOut11_14[5] , 
        \nOut11_14[4] , \nOut11_14[3] , \nOut11_14[2] , \nOut11_14[1] , 
        \nOut11_14[0] }), .EastIn({\nOut12_13[7] , \nOut12_13[6] , 
        \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , \nOut12_13[2] , 
        \nOut12_13[1] , \nOut12_13[0] }), .WestIn({\nOut10_13[7] , 
        \nOut10_13[6] , \nOut10_13[5] , \nOut10_13[4] , \nOut10_13[3] , 
        \nOut10_13[2] , \nOut10_13[1] , \nOut10_13[0] }), .Out({\nOut11_13[7] , 
        \nOut11_13[6] , \nOut11_13[5] , \nOut11_13[4] , \nOut11_13[3] , 
        \nOut11_13[2] , \nOut11_13[1] , \nOut11_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_68 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut69[7] , \nScanOut69[6] , 
        \nScanOut69[5] , \nScanOut69[4] , \nScanOut69[3] , \nScanOut69[2] , 
        \nScanOut69[1] , \nScanOut69[0] }), .ScanOut({\nScanOut68[7] , 
        \nScanOut68[6] , \nScanOut68[5] , \nScanOut68[4] , \nScanOut68[3] , 
        \nScanOut68[2] , \nScanOut68[1] , \nScanOut68[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , \nOut4_3[3] , 
        \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }), .SouthIn({\nOut4_5[7] , 
        \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , 
        \nOut4_5[1] , \nOut4_5[0] }), .EastIn({\nOut5_4[7] , \nOut5_4[6] , 
        \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , \nOut5_4[2] , \nOut5_4[1] , 
        \nOut5_4[0] }), .WestIn({\nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , 
        \nOut3_4[4] , \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }), 
        .Out({\nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , 
        \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_73 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut74[7] , \nScanOut74[6] , 
        \nScanOut74[5] , \nScanOut74[4] , \nScanOut74[3] , \nScanOut74[2] , 
        \nScanOut74[1] , \nScanOut74[0] }), .ScanOut({\nScanOut73[7] , 
        \nScanOut73[6] , \nScanOut73[5] , \nScanOut73[4] , \nScanOut73[3] , 
        \nScanOut73[2] , \nScanOut73[1] , \nScanOut73[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , \nOut4_8[3] , 
        \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }), .SouthIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .EastIn({\nOut5_9[7] , 
        \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , \nOut5_9[2] , 
        \nOut5_9[1] , \nOut5_9[0] }), .WestIn({\nOut3_9[7] , \nOut3_9[6] , 
        \nOut3_9[5] , \nOut3_9[4] , \nOut3_9[3] , \nOut3_9[2] , \nOut3_9[1] , 
        \nOut3_9[0] }), .Out({\nOut4_9[7] , \nOut4_9[6] , \nOut4_9[5] , 
        \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , \nOut4_9[1] , \nOut4_9[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_150 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut151[7] , \nScanOut151[6] , 
        \nScanOut151[5] , \nScanOut151[4] , \nScanOut151[3] , \nScanOut151[2] , 
        \nScanOut151[1] , \nScanOut151[0] }), .ScanOut({\nScanOut150[7] , 
        \nScanOut150[6] , \nScanOut150[5] , \nScanOut150[4] , \nScanOut150[3] , 
        \nScanOut150[2] , \nScanOut150[1] , \nScanOut150[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_5[7] , \nOut9_5[6] , \nOut9_5[5] , \nOut9_5[4] , \nOut9_5[3] , 
        \nOut9_5[2] , \nOut9_5[1] , \nOut9_5[0] }), .SouthIn({\nOut9_7[7] , 
        \nOut9_7[6] , \nOut9_7[5] , \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , 
        \nOut9_7[1] , \nOut9_7[0] }), .EastIn({\nOut10_6[7] , \nOut10_6[6] , 
        \nOut10_6[5] , \nOut10_6[4] , \nOut10_6[3] , \nOut10_6[2] , 
        \nOut10_6[1] , \nOut10_6[0] }), .WestIn({\nOut8_6[7] , \nOut8_6[6] , 
        \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , 
        \nOut8_6[0] }), .Out({\nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , 
        \nOut9_6[4] , \nOut9_6[3] , \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_177 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut178[7] , \nScanOut178[6] , 
        \nScanOut178[5] , \nScanOut178[4] , \nScanOut178[3] , \nScanOut178[2] , 
        \nScanOut178[1] , \nScanOut178[0] }), .ScanOut({\nScanOut177[7] , 
        \nScanOut177[6] , \nScanOut177[5] , \nScanOut177[4] , \nScanOut177[3] , 
        \nScanOut177[2] , \nScanOut177[1] , \nScanOut177[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_0[7] , \nOut11_0[6] , \nOut11_0[5] , \nOut11_0[4] , 
        \nOut11_0[3] , \nOut11_0[2] , \nOut11_0[1] , \nOut11_0[0] }), 
        .SouthIn({\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .EastIn(
        {\nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), .WestIn(
        {\nOut10_1[7] , \nOut10_1[6] , \nOut10_1[5] , \nOut10_1[4] , 
        \nOut10_1[3] , \nOut10_1[2] , \nOut10_1[1] , \nOut10_1[0] }), .Out({
        \nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_247 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut248[7] , \nScanOut248[6] , 
        \nScanOut248[5] , \nScanOut248[4] , \nScanOut248[3] , \nScanOut248[2] , 
        \nScanOut248[1] , \nScanOut248[0] }), .ScanOut({\nScanOut247[7] , 
        \nScanOut247[6] , \nScanOut247[5] , \nScanOut247[4] , \nScanOut247[3] , 
        \nScanOut247[2] , \nScanOut247[1] , \nScanOut247[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_7[7] , \nOut15_7[6] , 
        \nOut15_7[5] , \nOut15_7[4] , \nOut15_7[3] , \nOut15_7[2] , 
        \nOut15_7[1] , \nOut15_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_21 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut22[7] , \nScanOut22[6] , 
        \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , 
        \nScanOut22[1] , \nScanOut22[0] }), .ScanOut({\nScanOut21[7] , 
        \nScanOut21[6] , \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , 
        \nScanOut21[2] , \nScanOut21[1] , \nScanOut21[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , 
        \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), .SouthIn({\nOut1_6[7] , 
        \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , 
        \nOut1_6[1] , \nOut1_6[0] }), .EastIn({\nOut2_5[7] , \nOut2_5[6] , 
        \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , 
        \nOut2_5[0] }), .WestIn({\nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , 
        \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), 
        .Out({\nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , 
        \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_29 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut30[7] , \nScanOut30[6] , 
        \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , 
        \nScanOut30[1] , \nScanOut30[0] }), .ScanOut({\nScanOut29[7] , 
        \nScanOut29[6] , \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , 
        \nScanOut29[2] , \nScanOut29[1] , \nScanOut29[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), 
        .SouthIn({\nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .EastIn(
        {\nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .WestIn(
        {\nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , 
        \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), .Out({
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_119 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut120[7] , \nScanOut120[6] , 
        \nScanOut120[5] , \nScanOut120[4] , \nScanOut120[3] , \nScanOut120[2] , 
        \nScanOut120[1] , \nScanOut120[0] }), .ScanOut({\nScanOut119[7] , 
        \nScanOut119[6] , \nScanOut119[5] , \nScanOut119[4] , \nScanOut119[3] , 
        \nScanOut119[2] , \nScanOut119[1] , \nScanOut119[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , \nOut7_6[3] , 
        \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }), .SouthIn({\nOut7_8[7] , 
        \nOut7_8[6] , \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , 
        \nOut7_8[1] , \nOut7_8[0] }), .EastIn({\nOut8_7[7] , \nOut8_7[6] , 
        \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , 
        \nOut8_7[0] }), .WestIn({\nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , 
        \nOut6_7[4] , \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }), 
        .Out({\nOut7_7[7] , \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , 
        \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , \nOut7_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_192 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut193[7] , \nScanOut193[6] , 
        \nScanOut193[5] , \nScanOut193[4] , \nScanOut193[3] , \nScanOut193[2] , 
        \nScanOut193[1] , \nScanOut193[0] }), .ScanOut({\nScanOut192[7] , 
        \nScanOut192[6] , \nScanOut192[5] , \nScanOut192[4] , \nScanOut192[3] , 
        \nScanOut192[2] , \nScanOut192[1] , \nScanOut192[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut12_0[7] , \nOut12_0[6] , 
        \nOut12_0[5] , \nOut12_0[4] , \nOut12_0[3] , \nOut12_0[2] , 
        \nOut12_0[1] , \nOut12_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_229 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut230[7] , \nScanOut230[6] , 
        \nScanOut230[5] , \nScanOut230[4] , \nScanOut230[3] , \nScanOut230[2] , 
        \nScanOut230[1] , \nScanOut230[0] }), .ScanOut({\nScanOut229[7] , 
        \nScanOut229[6] , \nScanOut229[5] , \nScanOut229[4] , \nScanOut229[3] , 
        \nScanOut229[2] , \nScanOut229[1] , \nScanOut229[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }), 
        .SouthIn({\nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), .EastIn(
        {\nOut15_5[7] , \nOut15_5[6] , \nOut15_5[5] , \nOut15_5[4] , 
        \nOut15_5[3] , \nOut15_5[2] , \nOut15_5[1] , \nOut15_5[0] }), .WestIn(
        {\nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), .Out({
        \nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_85 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut86[7] , \nScanOut86[6] , 
        \nScanOut86[5] , \nScanOut86[4] , \nScanOut86[3] , \nScanOut86[2] , 
        \nScanOut86[1] , \nScanOut86[0] }), .ScanOut({\nScanOut85[7] , 
        \nScanOut85[6] , \nScanOut85[5] , \nScanOut85[4] , \nScanOut85[3] , 
        \nScanOut85[2] , \nScanOut85[1] , \nScanOut85[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_4[7] , \nOut5_4[6] , \nOut5_4[5] , \nOut5_4[4] , \nOut5_4[3] , 
        \nOut5_4[2] , \nOut5_4[1] , \nOut5_4[0] }), .SouthIn({\nOut5_6[7] , 
        \nOut5_6[6] , \nOut5_6[5] , \nOut5_6[4] , \nOut5_6[3] , \nOut5_6[2] , 
        \nOut5_6[1] , \nOut5_6[0] }), .EastIn({\nOut6_5[7] , \nOut6_5[6] , 
        \nOut6_5[5] , \nOut6_5[4] , \nOut6_5[3] , \nOut6_5[2] , \nOut6_5[1] , 
        \nOut6_5[0] }), .WestIn({\nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , 
        \nOut4_5[4] , \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }), 
        .Out({\nOut5_5[7] , \nOut5_5[6] , \nOut5_5[5] , \nOut5_5[4] , 
        \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , \nOut5_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_111 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut112[7] , \nScanOut112[6] , 
        \nScanOut112[5] , \nScanOut112[4] , \nScanOut112[3] , \nScanOut112[2] , 
        \nScanOut112[1] , \nScanOut112[0] }), .ScanOut({\nScanOut111[7] , 
        \nScanOut111[6] , \nScanOut111[5] , \nScanOut111[4] , \nScanOut111[3] , 
        \nScanOut111[2] , \nScanOut111[1] , \nScanOut111[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut6_15[7] , \nOut6_15[6] , 
        \nOut6_15[5] , \nOut6_15[4] , \nOut6_15[3] , \nOut6_15[2] , 
        \nOut6_15[1] , \nOut6_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_136 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut137[7] , \nScanOut137[6] , 
        \nScanOut137[5] , \nScanOut137[4] , \nScanOut137[3] , \nScanOut137[2] , 
        \nScanOut137[1] , \nScanOut137[0] }), .ScanOut({\nScanOut136[7] , 
        \nScanOut136[6] , \nScanOut136[5] , \nScanOut136[4] , \nScanOut136[3] , 
        \nScanOut136[2] , \nScanOut136[1] , \nScanOut136[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_7[7] , \nOut8_7[6] , \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , 
        \nOut8_7[2] , \nOut8_7[1] , \nOut8_7[0] }), .SouthIn({\nOut8_9[7] , 
        \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , \nOut8_9[2] , 
        \nOut8_9[1] , \nOut8_9[0] }), .EastIn({\nOut9_8[7] , \nOut9_8[6] , 
        \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , \nOut9_8[1] , 
        \nOut9_8[0] }), .WestIn({\nOut7_8[7] , \nOut7_8[6] , \nOut7_8[5] , 
        \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , \nOut7_8[0] }), 
        .Out({\nOut8_8[7] , \nOut8_8[6] , \nOut8_8[5] , \nOut8_8[4] , 
        \nOut8_8[3] , \nOut8_8[2] , \nOut8_8[1] , \nOut8_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_206 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut207[7] , \nScanOut207[6] , 
        \nScanOut207[5] , \nScanOut207[4] , \nScanOut207[3] , \nScanOut207[2] , 
        \nScanOut207[1] , \nScanOut207[0] }), .ScanOut({\nScanOut206[7] , 
        \nScanOut206[6] , \nScanOut206[5] , \nScanOut206[4] , \nScanOut206[3] , 
        \nScanOut206[2] , \nScanOut206[1] , \nScanOut206[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_13[7] , \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , 
        \nOut12_13[3] , \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }), 
        .SouthIn({\nOut12_15[7] , \nOut12_15[6] , \nOut12_15[5] , 
        \nOut12_15[4] , \nOut12_15[3] , \nOut12_15[2] , \nOut12_15[1] , 
        \nOut12_15[0] }), .EastIn({\nOut13_14[7] , \nOut13_14[6] , 
        \nOut13_14[5] , \nOut13_14[4] , \nOut13_14[3] , \nOut13_14[2] , 
        \nOut13_14[1] , \nOut13_14[0] }), .WestIn({\nOut11_14[7] , 
        \nOut11_14[6] , \nOut11_14[5] , \nOut11_14[4] , \nOut11_14[3] , 
        \nOut11_14[2] , \nOut11_14[1] , \nOut11_14[0] }), .Out({\nOut12_14[7] , 
        \nOut12_14[6] , \nOut12_14[5] , \nOut12_14[4] , \nOut12_14[3] , 
        \nOut12_14[2] , \nOut12_14[1] , \nOut12_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_221 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut222[7] , \nScanOut222[6] , 
        \nScanOut222[5] , \nScanOut222[4] , \nScanOut222[3] , \nScanOut222[2] , 
        \nScanOut222[1] , \nScanOut222[0] }), .ScanOut({\nScanOut221[7] , 
        \nScanOut221[6] , \nScanOut221[5] , \nScanOut221[4] , \nScanOut221[3] , 
        \nScanOut221[2] , \nScanOut221[1] , \nScanOut221[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_12[7] , \nOut13_12[6] , \nOut13_12[5] , \nOut13_12[4] , 
        \nOut13_12[3] , \nOut13_12[2] , \nOut13_12[1] , \nOut13_12[0] }), 
        .SouthIn({\nOut13_14[7] , \nOut13_14[6] , \nOut13_14[5] , 
        \nOut13_14[4] , \nOut13_14[3] , \nOut13_14[2] , \nOut13_14[1] , 
        \nOut13_14[0] }), .EastIn({\nOut14_13[7] , \nOut14_13[6] , 
        \nOut14_13[5] , \nOut14_13[4] , \nOut14_13[3] , \nOut14_13[2] , 
        \nOut14_13[1] , \nOut14_13[0] }), .WestIn({\nOut12_13[7] , 
        \nOut12_13[6] , \nOut12_13[5] , \nOut12_13[4] , \nOut12_13[3] , 
        \nOut12_13[2] , \nOut12_13[1] , \nOut12_13[0] }), .Out({\nOut13_13[7] , 
        \nOut13_13[6] , \nOut13_13[5] , \nOut13_13[4] , \nOut13_13[3] , 
        \nOut13_13[2] , \nOut13_13[1] , \nOut13_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_158 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut159[7] , \nScanOut159[6] , 
        \nScanOut159[5] , \nScanOut159[4] , \nScanOut159[3] , \nScanOut159[2] , 
        \nScanOut159[1] , \nScanOut159[0] }), .ScanOut({\nScanOut158[7] , 
        \nScanOut158[6] , \nScanOut158[5] , \nScanOut158[4] , \nScanOut158[3] , 
        \nScanOut158[2] , \nScanOut158[1] , \nScanOut158[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), 
        .SouthIn({\nOut9_15[7] , \nOut9_15[6] , \nOut9_15[5] , \nOut9_15[4] , 
        \nOut9_15[3] , \nOut9_15[2] , \nOut9_15[1] , \nOut9_15[0] }), .EastIn(
        {\nOut10_14[7] , \nOut10_14[6] , \nOut10_14[5] , \nOut10_14[4] , 
        \nOut10_14[3] , \nOut10_14[2] , \nOut10_14[1] , \nOut10_14[0] }), 
        .WestIn({\nOut8_14[7] , \nOut8_14[6] , \nOut8_14[5] , \nOut8_14[4] , 
        \nOut8_14[3] , \nOut8_14[2] , \nOut8_14[1] , \nOut8_14[0] }), .Out({
        \nOut9_14[7] , \nOut9_14[6] , \nOut9_14[5] , \nOut9_14[4] , 
        \nOut9_14[3] , \nOut9_14[2] , \nOut9_14[1] , \nOut9_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut7[7] , \nScanOut7[6] , 
        \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , 
        \nScanOut7[1] , \nScanOut7[0] }), .ScanOut({\nScanOut6[7] , 
        \nScanOut6[6] , \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , 
        \nScanOut6[2] , \nScanOut6[1] , \nScanOut6[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_6[7] , \nOut0_6[6] , 
        \nOut0_6[5] , \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , 
        \nOut0_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut9[7] , \nScanOut9[6] , 
        \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , 
        \nScanOut9[1] , \nScanOut9[0] }), .ScanOut({\nScanOut8[7] , 
        \nScanOut8[6] , \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , 
        \nScanOut8[2] , \nScanOut8[1] , \nScanOut8[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_8[7] , \nOut0_8[6] , 
        \nOut0_8[5] , \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , 
        \nOut0_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut16[7] , \nScanOut16[6] , 
        \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , 
        \nScanOut16[1] , \nScanOut16[0] }), .ScanOut({\nScanOut15[7] , 
        \nScanOut15[6] , \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , 
        \nScanOut15[2] , \nScanOut15[1] , \nScanOut15[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_32 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut33[7] , \nScanOut33[6] , 
        \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , 
        \nScanOut33[1] , \nScanOut33[0] }), .ScanOut({\nScanOut32[7] , 
        \nScanOut32[6] , \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , 
        \nScanOut32[2] , \nScanOut32[1] , \nScanOut32[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_0[7] , \nOut2_0[6] , 
        \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , \nOut2_0[2] , \nOut2_0[1] , 
        \nOut2_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_47 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut48[7] , \nScanOut48[6] , 
        \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , \nScanOut48[2] , 
        \nScanOut48[1] , \nScanOut48[0] }), .ScanOut({\nScanOut47[7] , 
        \nScanOut47[6] , \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , 
        \nScanOut47[2] , \nScanOut47[1] , \nScanOut47[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_15[7] , \nOut2_15[6] , 
        \nOut2_15[5] , \nOut2_15[4] , \nOut2_15[3] , \nOut2_15[2] , 
        \nOut2_15[1] , \nOut2_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_60 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut61[7] , \nScanOut61[6] , 
        \nScanOut61[5] , \nScanOut61[4] , \nScanOut61[3] , \nScanOut61[2] , 
        \nScanOut61[1] , \nScanOut61[0] }), .ScanOut({\nScanOut60[7] , 
        \nScanOut60[6] , \nScanOut60[5] , \nScanOut60[4] , \nScanOut60[3] , 
        \nScanOut60[2] , \nScanOut60[1] , \nScanOut60[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), 
        .SouthIn({\nOut3_13[7] , \nOut3_13[6] , \nOut3_13[5] , \nOut3_13[4] , 
        \nOut3_13[3] , \nOut3_13[2] , \nOut3_13[1] , \nOut3_13[0] }), .EastIn(
        {\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .WestIn(
        {\nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .Out({
        \nOut3_12[7] , \nOut3_12[6] , \nOut3_12[5] , \nOut3_12[4] , 
        \nOut3_12[3] , \nOut3_12[2] , \nOut3_12[1] , \nOut3_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_143 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut144[7] , \nScanOut144[6] , 
        \nScanOut144[5] , \nScanOut144[4] , \nScanOut144[3] , \nScanOut144[2] , 
        \nScanOut144[1] , \nScanOut144[0] }), .ScanOut({\nScanOut143[7] , 
        \nScanOut143[6] , \nScanOut143[5] , \nScanOut143[4] , \nScanOut143[3] , 
        \nScanOut143[2] , \nScanOut143[1] , \nScanOut143[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut8_15[7] , \nOut8_15[6] , 
        \nOut8_15[5] , \nOut8_15[4] , \nOut8_15[3] , \nOut8_15[2] , 
        \nOut8_15[1] , \nOut8_15[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_164 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut165[7] , \nScanOut165[6] , 
        \nScanOut165[5] , \nScanOut165[4] , \nScanOut165[3] , \nScanOut165[2] , 
        \nScanOut165[1] , \nScanOut165[0] }), .ScanOut({\nScanOut164[7] , 
        \nScanOut164[6] , \nScanOut164[5] , \nScanOut164[4] , \nScanOut164[3] , 
        \nScanOut164[2] , \nScanOut164[1] , \nScanOut164[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_3[7] , \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , 
        \nOut10_3[3] , \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }), 
        .SouthIn({\nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), .EastIn(
        {\nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), .WestIn(
        {\nOut9_4[7] , \nOut9_4[6] , \nOut9_4[5] , \nOut9_4[4] , \nOut9_4[3] , 
        \nOut9_4[2] , \nOut9_4[1] , \nOut9_4[0] }), .Out({\nOut10_4[7] , 
        \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , \nOut10_4[3] , 
        \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_254 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut255[7] , \nScanOut255[6] , 
        \nScanOut255[5] , \nScanOut255[4] , \nScanOut255[3] , \nScanOut255[2] , 
        \nScanOut255[1] , \nScanOut255[0] }), .ScanOut({\nScanOut254[7] , 
        \nScanOut254[6] , \nScanOut254[5] , \nScanOut254[4] , \nScanOut254[3] , 
        \nScanOut254[2] , \nScanOut254[1] , \nScanOut254[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_14[7] , \nOut15_14[6] , 
        \nOut15_14[5] , \nOut15_14[4] , \nOut15_14[3] , \nOut15_14[2] , 
        \nOut15_14[1] , \nOut15_14[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_20 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut21[7] , \nScanOut21[6] , 
        \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , 
        \nScanOut21[1] , \nScanOut21[0] }), .ScanOut({\nScanOut20[7] , 
        \nScanOut20[6] , \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , 
        \nScanOut20[2] , \nScanOut20[1] , \nScanOut20[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , 
        \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), .SouthIn({\nOut1_5[7] , 
        \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , 
        \nOut1_5[1] , \nOut1_5[0] }), .EastIn({\nOut2_4[7] , \nOut2_4[6] , 
        \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , 
        \nOut2_4[0] }), .WestIn({\nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , 
        \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), 
        .Out({\nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , 
        \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_181 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut182[7] , \nScanOut182[6] , 
        \nScanOut182[5] , \nScanOut182[4] , \nScanOut182[3] , \nScanOut182[2] , 
        \nScanOut182[1] , \nScanOut182[0] }), .ScanOut({\nScanOut181[7] , 
        \nScanOut181[6] , \nScanOut181[5] , \nScanOut181[4] , \nScanOut181[3] , 
        \nScanOut181[2] , \nScanOut181[1] , \nScanOut181[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_4[7] , \nOut11_4[6] , \nOut11_4[5] , \nOut11_4[4] , 
        \nOut11_4[3] , \nOut11_4[2] , \nOut11_4[1] , \nOut11_4[0] }), 
        .SouthIn({\nOut11_6[7] , \nOut11_6[6] , \nOut11_6[5] , \nOut11_6[4] , 
        \nOut11_6[3] , \nOut11_6[2] , \nOut11_6[1] , \nOut11_6[0] }), .EastIn(
        {\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .WestIn(
        {\nOut10_5[7] , \nOut10_5[6] , \nOut10_5[5] , \nOut10_5[4] , 
        \nOut10_5[3] , \nOut10_5[2] , \nOut10_5[1] , \nOut10_5[0] }), .Out({
        \nOut11_5[7] , \nOut11_5[6] , \nOut11_5[5] , \nOut11_5[4] , 
        \nOut11_5[3] , \nOut11_5[2] , \nOut11_5[1] , \nOut11_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_69 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut70[7] , \nScanOut70[6] , 
        \nScanOut70[5] , \nScanOut70[4] , \nScanOut70[3] , \nScanOut70[2] , 
        \nScanOut70[1] , \nScanOut70[0] }), .ScanOut({\nScanOut69[7] , 
        \nScanOut69[6] , \nScanOut69[5] , \nScanOut69[4] , \nScanOut69[3] , 
        \nScanOut69[2] , \nScanOut69[1] , \nScanOut69[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_4[7] , \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , 
        \nOut4_4[2] , \nOut4_4[1] , \nOut4_4[0] }), .SouthIn({\nOut4_6[7] , 
        \nOut4_6[6] , \nOut4_6[5] , \nOut4_6[4] , \nOut4_6[3] , \nOut4_6[2] , 
        \nOut4_6[1] , \nOut4_6[0] }), .EastIn({\nOut5_5[7] , \nOut5_5[6] , 
        \nOut5_5[5] , \nOut5_5[4] , \nOut5_5[3] , \nOut5_5[2] , \nOut5_5[1] , 
        \nOut5_5[0] }), .WestIn({\nOut3_5[7] , \nOut3_5[6] , \nOut3_5[5] , 
        \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , \nOut3_5[1] , \nOut3_5[0] }), 
        .Out({\nOut4_5[7] , \nOut4_5[6] , \nOut4_5[5] , \nOut4_5[4] , 
        \nOut4_5[3] , \nOut4_5[2] , \nOut4_5[1] , \nOut4_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_118 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut119[7] , \nScanOut119[6] , 
        \nScanOut119[5] , \nScanOut119[4] , \nScanOut119[3] , \nScanOut119[2] , 
        \nScanOut119[1] , \nScanOut119[0] }), .ScanOut({\nScanOut118[7] , 
        \nScanOut118[6] , \nScanOut118[5] , \nScanOut118[4] , \nScanOut118[3] , 
        \nScanOut118[2] , \nScanOut118[1] , \nScanOut118[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_5[7] , \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , 
        \nOut7_5[2] , \nOut7_5[1] , \nOut7_5[0] }), .SouthIn({\nOut7_7[7] , 
        \nOut7_7[6] , \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , 
        \nOut7_7[1] , \nOut7_7[0] }), .EastIn({\nOut8_6[7] , \nOut8_6[6] , 
        \nOut8_6[5] , \nOut8_6[4] , \nOut8_6[3] , \nOut8_6[2] , \nOut8_6[1] , 
        \nOut8_6[0] }), .WestIn({\nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , 
        \nOut6_6[4] , \nOut6_6[3] , \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }), 
        .Out({\nOut7_6[7] , \nOut7_6[6] , \nOut7_6[5] , \nOut7_6[4] , 
        \nOut7_6[3] , \nOut7_6[2] , \nOut7_6[1] , \nOut7_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_193 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut194[7] , \nScanOut194[6] , 
        \nScanOut194[5] , \nScanOut194[4] , \nScanOut194[3] , \nScanOut194[2] , 
        \nScanOut194[1] , \nScanOut194[0] }), .ScanOut({\nScanOut193[7] , 
        \nScanOut193[6] , \nScanOut193[5] , \nScanOut193[4] , \nScanOut193[3] , 
        \nScanOut193[2] , \nScanOut193[1] , \nScanOut193[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_0[7] , \nOut12_0[6] , \nOut12_0[5] , \nOut12_0[4] , 
        \nOut12_0[3] , \nOut12_0[2] , \nOut12_0[1] , \nOut12_0[0] }), 
        .SouthIn({\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .EastIn(
        {\nOut13_1[7] , \nOut13_1[6] , \nOut13_1[5] , \nOut13_1[4] , 
        \nOut13_1[3] , \nOut13_1[2] , \nOut13_1[1] , \nOut13_1[0] }), .WestIn(
        {\nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), .Out({
        \nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_228 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut229[7] , \nScanOut229[6] , 
        \nScanOut229[5] , \nScanOut229[4] , \nScanOut229[3] , \nScanOut229[2] , 
        \nScanOut229[1] , \nScanOut229[0] }), .ScanOut({\nScanOut228[7] , 
        \nScanOut228[6] , \nScanOut228[5] , \nScanOut228[4] , \nScanOut228[3] , 
        \nScanOut228[2] , \nScanOut228[1] , \nScanOut228[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), 
        .SouthIn({\nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), .EastIn(
        {\nOut15_4[7] , \nOut15_4[6] , \nOut15_4[5] , \nOut15_4[4] , 
        \nOut15_4[3] , \nOut15_4[2] , \nOut15_4[1] , \nOut15_4[0] }), .WestIn(
        {\nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), .Out({
        \nOut14_4[7] , \nOut14_4[6] , \nOut14_4[5] , \nOut14_4[4] , 
        \nOut14_4[3] , \nOut14_4[2] , \nOut14_4[1] , \nOut14_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_151 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut152[7] , \nScanOut152[6] , 
        \nScanOut152[5] , \nScanOut152[4] , \nScanOut152[3] , \nScanOut152[2] , 
        \nScanOut152[1] , \nScanOut152[0] }), .ScanOut({\nScanOut151[7] , 
        \nScanOut151[6] , \nScanOut151[5] , \nScanOut151[4] , \nScanOut151[3] , 
        \nScanOut151[2] , \nScanOut151[1] , \nScanOut151[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_6[7] , \nOut9_6[6] , \nOut9_6[5] , \nOut9_6[4] , \nOut9_6[3] , 
        \nOut9_6[2] , \nOut9_6[1] , \nOut9_6[0] }), .SouthIn({\nOut9_8[7] , 
        \nOut9_8[6] , \nOut9_8[5] , \nOut9_8[4] , \nOut9_8[3] , \nOut9_8[2] , 
        \nOut9_8[1] , \nOut9_8[0] }), .EastIn({\nOut10_7[7] , \nOut10_7[6] , 
        \nOut10_7[5] , \nOut10_7[4] , \nOut10_7[3] , \nOut10_7[2] , 
        \nOut10_7[1] , \nOut10_7[0] }), .WestIn({\nOut8_7[7] , \nOut8_7[6] , 
        \nOut8_7[5] , \nOut8_7[4] , \nOut8_7[3] , \nOut8_7[2] , \nOut8_7[1] , 
        \nOut8_7[0] }), .Out({\nOut9_7[7] , \nOut9_7[6] , \nOut9_7[5] , 
        \nOut9_7[4] , \nOut9_7[3] , \nOut9_7[2] , \nOut9_7[1] , \nOut9_7[0] })
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_176 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut177[7] , \nScanOut177[6] , 
        \nScanOut177[5] , \nScanOut177[4] , \nScanOut177[3] , \nScanOut177[2] , 
        \nScanOut177[1] , \nScanOut177[0] }), .ScanOut({\nScanOut176[7] , 
        \nScanOut176[6] , \nScanOut176[5] , \nScanOut176[4] , \nScanOut176[3] , 
        \nScanOut176[2] , \nScanOut176[1] , \nScanOut176[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut11_0[7] , \nOut11_0[6] , 
        \nOut11_0[5] , \nOut11_0[4] , \nOut11_0[3] , \nOut11_0[2] , 
        \nOut11_0[1] , \nOut11_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_246 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut247[7] , \nScanOut247[6] , 
        \nScanOut247[5] , \nScanOut247[4] , \nScanOut247[3] , \nScanOut247[2] , 
        \nScanOut247[1] , \nScanOut247[0] }), .ScanOut({\nScanOut246[7] , 
        \nScanOut246[6] , \nScanOut246[5] , \nScanOut246[4] , \nScanOut246[3] , 
        \nScanOut246[2] , \nScanOut246[1] , \nScanOut246[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_6[7] , \nOut15_6[6] , 
        \nOut15_6[5] , \nOut15_6[4] , \nOut15_6[3] , \nOut15_6[2] , 
        \nOut15_6[1] , \nOut15_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut13[7] , \nScanOut13[6] , 
        \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , 
        \nScanOut13[1] , \nScanOut13[0] }), .ScanOut({\nScanOut12[7] , 
        \nScanOut12[6] , \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , 
        \nScanOut12[2] , \nScanOut12[1] , \nScanOut12[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_12[7] , \nOut0_12[6] , 
        \nOut0_12[5] , \nOut0_12[4] , \nOut0_12[3] , \nOut0_12[2] , 
        \nOut0_12[1] , \nOut0_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_27 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut28[7] , \nScanOut28[6] , 
        \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , 
        \nScanOut28[1] , \nScanOut28[0] }), .ScanOut({\nScanOut27[7] , 
        \nScanOut27[6] , \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , 
        \nScanOut27[2] , \nScanOut27[1] , \nScanOut27[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , 
        \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), 
        .SouthIn({\nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .EastIn(
        {\nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .WestIn(
        {\nOut0_11[7] , \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , 
        \nOut0_11[3] , \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .Out({
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_49 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut50[7] , \nScanOut50[6] , 
        \nScanOut50[5] , \nScanOut50[4] , \nScanOut50[3] , \nScanOut50[2] , 
        \nScanOut50[1] , \nScanOut50[0] }), .ScanOut({\nScanOut49[7] , 
        \nScanOut49[6] , \nScanOut49[5] , \nScanOut49[4] , \nScanOut49[3] , 
        \nScanOut49[2] , \nScanOut49[1] , \nScanOut49[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_0[7] , \nOut3_0[6] , \nOut3_0[5] , \nOut3_0[4] , \nOut3_0[3] , 
        \nOut3_0[2] , \nOut3_0[1] , \nOut3_0[0] }), .SouthIn({\nOut3_2[7] , 
        \nOut3_2[6] , \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , 
        \nOut3_2[1] , \nOut3_2[0] }), .EastIn({\nOut4_1[7] , \nOut4_1[6] , 
        \nOut4_1[5] , \nOut4_1[4] , \nOut4_1[3] , \nOut4_1[2] , \nOut4_1[1] , 
        \nOut4_1[0] }), .WestIn({\nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , 
        \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), 
        .Out({\nOut3_1[7] , \nOut3_1[6] , \nOut3_1[5] , \nOut3_1[4] , 
        \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , \nOut3_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_52 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut53[7] , \nScanOut53[6] , 
        \nScanOut53[5] , \nScanOut53[4] , \nScanOut53[3] , \nScanOut53[2] , 
        \nScanOut53[1] , \nScanOut53[0] }), .ScanOut({\nScanOut52[7] , 
        \nScanOut52[6] , \nScanOut52[5] , \nScanOut52[4] , \nScanOut52[3] , 
        \nScanOut52[2] , \nScanOut52[1] , \nScanOut52[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , 
        \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }), .SouthIn({\nOut3_5[7] , 
        \nOut3_5[6] , \nOut3_5[5] , \nOut3_5[4] , \nOut3_5[3] , \nOut3_5[2] , 
        \nOut3_5[1] , \nOut3_5[0] }), .EastIn({\nOut4_4[7] , \nOut4_4[6] , 
        \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , \nOut4_4[1] , 
        \nOut4_4[0] }), .WestIn({\nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , 
        \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), 
        .Out({\nOut3_4[7] , \nOut3_4[6] , \nOut3_4[5] , \nOut3_4[4] , 
        \nOut3_4[3] , \nOut3_4[2] , \nOut3_4[1] , \nOut3_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_55 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut56[7] , \nScanOut56[6] , 
        \nScanOut56[5] , \nScanOut56[4] , \nScanOut56[3] , \nScanOut56[2] , 
        \nScanOut56[1] , \nScanOut56[0] }), .ScanOut({\nScanOut55[7] , 
        \nScanOut55[6] , \nScanOut55[5] , \nScanOut55[4] , \nScanOut55[3] , 
        \nScanOut55[2] , \nScanOut55[1] , \nScanOut55[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut3_6[7] , \nOut3_6[6] , \nOut3_6[5] , \nOut3_6[4] , \nOut3_6[3] , 
        \nOut3_6[2] , \nOut3_6[1] , \nOut3_6[0] }), .SouthIn({\nOut3_8[7] , 
        \nOut3_8[6] , \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , 
        \nOut3_8[1] , \nOut3_8[0] }), .EastIn({\nOut4_7[7] , \nOut4_7[6] , 
        \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , \nOut4_7[2] , \nOut4_7[1] , 
        \nOut4_7[0] }), .WestIn({\nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , 
        \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), 
        .Out({\nOut3_7[7] , \nOut3_7[6] , \nOut3_7[5] , \nOut3_7[4] , 
        \nOut3_7[3] , \nOut3_7[2] , \nOut3_7[1] , \nOut3_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_72 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut73[7] , \nScanOut73[6] , 
        \nScanOut73[5] , \nScanOut73[4] , \nScanOut73[3] , \nScanOut73[2] , 
        \nScanOut73[1] , \nScanOut73[0] }), .ScanOut({\nScanOut72[7] , 
        \nScanOut72[6] , \nScanOut72[5] , \nScanOut72[4] , \nScanOut72[3] , 
        \nScanOut72[2] , \nScanOut72[1] , \nScanOut72[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_7[7] , \nOut4_7[6] , \nOut4_7[5] , \nOut4_7[4] , \nOut4_7[3] , 
        \nOut4_7[2] , \nOut4_7[1] , \nOut4_7[0] }), .SouthIn({\nOut4_9[7] , 
        \nOut4_9[6] , \nOut4_9[5] , \nOut4_9[4] , \nOut4_9[3] , \nOut4_9[2] , 
        \nOut4_9[1] , \nOut4_9[0] }), .EastIn({\nOut5_8[7] , \nOut5_8[6] , 
        \nOut5_8[5] , \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , 
        \nOut5_8[0] }), .WestIn({\nOut3_8[7] , \nOut3_8[6] , \nOut3_8[5] , 
        \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , \nOut3_8[0] }), 
        .Out({\nOut4_8[7] , \nOut4_8[6] , \nOut4_8[5] , \nOut4_8[4] , 
        \nOut4_8[3] , \nOut4_8[2] , \nOut4_8[1] , \nOut4_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_75 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut76[7] , \nScanOut76[6] , 
        \nScanOut76[5] , \nScanOut76[4] , \nScanOut76[3] , \nScanOut76[2] , 
        \nScanOut76[1] , \nScanOut76[0] }), .ScanOut({\nScanOut75[7] , 
        \nScanOut75[6] , \nScanOut75[5] , \nScanOut75[4] , \nScanOut75[3] , 
        \nScanOut75[2] , \nScanOut75[1] , \nScanOut75[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_10[7] , \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , 
        \nOut4_10[3] , \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), 
        .SouthIn({\nOut4_12[7] , \nOut4_12[6] , \nOut4_12[5] , \nOut4_12[4] , 
        \nOut4_12[3] , \nOut4_12[2] , \nOut4_12[1] , \nOut4_12[0] }), .EastIn(
        {\nOut5_11[7] , \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , 
        \nOut5_11[3] , \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .WestIn(
        {\nOut3_11[7] , \nOut3_11[6] , \nOut3_11[5] , \nOut3_11[4] , 
        \nOut3_11[3] , \nOut3_11[2] , \nOut3_11[1] , \nOut3_11[0] }), .Out({
        \nOut4_11[7] , \nOut4_11[6] , \nOut4_11[5] , \nOut4_11[4] , 
        \nOut4_11[3] , \nOut4_11[2] , \nOut4_11[1] , \nOut4_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_90 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut91[7] , \nScanOut91[6] , 
        \nScanOut91[5] , \nScanOut91[4] , \nScanOut91[3] , \nScanOut91[2] , 
        \nScanOut91[1] , \nScanOut91[0] }), .ScanOut({\nScanOut90[7] , 
        \nScanOut90[6] , \nScanOut90[5] , \nScanOut90[4] , \nScanOut90[3] , 
        \nScanOut90[2] , \nScanOut90[1] , \nScanOut90[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_9[7] , \nOut5_9[6] , \nOut5_9[5] , \nOut5_9[4] , \nOut5_9[3] , 
        \nOut5_9[2] , \nOut5_9[1] , \nOut5_9[0] }), .SouthIn({\nOut5_11[7] , 
        \nOut5_11[6] , \nOut5_11[5] , \nOut5_11[4] , \nOut5_11[3] , 
        \nOut5_11[2] , \nOut5_11[1] , \nOut5_11[0] }), .EastIn({\nOut6_10[7] , 
        \nOut6_10[6] , \nOut6_10[5] , \nOut6_10[4] , \nOut6_10[3] , 
        \nOut6_10[2] , \nOut6_10[1] , \nOut6_10[0] }), .WestIn({\nOut4_10[7] , 
        \nOut4_10[6] , \nOut4_10[5] , \nOut4_10[4] , \nOut4_10[3] , 
        \nOut4_10[2] , \nOut4_10[1] , \nOut4_10[0] }), .Out({\nOut5_10[7] , 
        \nOut5_10[6] , \nOut5_10[5] , \nOut5_10[4] , \nOut5_10[3] , 
        \nOut5_10[2] , \nOut5_10[1] , \nOut5_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_97 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut98[7] , \nScanOut98[6] , 
        \nScanOut98[5] , \nScanOut98[4] , \nScanOut98[3] , \nScanOut98[2] , 
        \nScanOut98[1] , \nScanOut98[0] }), .ScanOut({\nScanOut97[7] , 
        \nScanOut97[6] , \nScanOut97[5] , \nScanOut97[4] , \nScanOut97[3] , 
        \nScanOut97[2] , \nScanOut97[1] , \nScanOut97[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_0[7] , \nOut6_0[6] , \nOut6_0[5] , \nOut6_0[4] , \nOut6_0[3] , 
        \nOut6_0[2] , \nOut6_0[1] , \nOut6_0[0] }), .SouthIn({\nOut6_2[7] , 
        \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , 
        \nOut6_2[1] , \nOut6_2[0] }), .EastIn({\nOut7_1[7] , \nOut7_1[6] , 
        \nOut7_1[5] , \nOut7_1[4] , \nOut7_1[3] , \nOut7_1[2] , \nOut7_1[1] , 
        \nOut7_1[0] }), .WestIn({\nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , 
        \nOut5_1[4] , \nOut5_1[3] , \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }), 
        .Out({\nOut6_1[7] , \nOut6_1[6] , \nOut6_1[5] , \nOut6_1[4] , 
        \nOut6_1[3] , \nOut6_1[2] , \nOut6_1[1] , \nOut6_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_103 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut104[7] , \nScanOut104[6] , 
        \nScanOut104[5] , \nScanOut104[4] , \nScanOut104[3] , \nScanOut104[2] , 
        \nScanOut104[1] , \nScanOut104[0] }), .ScanOut({\nScanOut103[7] , 
        \nScanOut103[6] , \nScanOut103[5] , \nScanOut103[4] , \nScanOut103[3] , 
        \nScanOut103[2] , \nScanOut103[1] , \nScanOut103[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_6[7] , \nOut6_6[6] , \nOut6_6[5] , \nOut6_6[4] , \nOut6_6[3] , 
        \nOut6_6[2] , \nOut6_6[1] , \nOut6_6[0] }), .SouthIn({\nOut6_8[7] , 
        \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , \nOut6_8[3] , \nOut6_8[2] , 
        \nOut6_8[1] , \nOut6_8[0] }), .EastIn({\nOut7_7[7] , \nOut7_7[6] , 
        \nOut7_7[5] , \nOut7_7[4] , \nOut7_7[3] , \nOut7_7[2] , \nOut7_7[1] , 
        \nOut7_7[0] }), .WestIn({\nOut5_7[7] , \nOut5_7[6] , \nOut5_7[5] , 
        \nOut5_7[4] , \nOut5_7[3] , \nOut5_7[2] , \nOut5_7[1] , \nOut5_7[0] }), 
        .Out({\nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , 
        \nOut6_7[3] , \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_104 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut105[7] , \nScanOut105[6] , 
        \nScanOut105[5] , \nScanOut105[4] , \nScanOut105[3] , \nScanOut105[2] , 
        \nScanOut105[1] , \nScanOut105[0] }), .ScanOut({\nScanOut104[7] , 
        \nScanOut104[6] , \nScanOut104[5] , \nScanOut104[4] , \nScanOut104[3] , 
        \nScanOut104[2] , \nScanOut104[1] , \nScanOut104[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_7[7] , \nOut6_7[6] , \nOut6_7[5] , \nOut6_7[4] , \nOut6_7[3] , 
        \nOut6_7[2] , \nOut6_7[1] , \nOut6_7[0] }), .SouthIn({\nOut6_9[7] , 
        \nOut6_9[6] , \nOut6_9[5] , \nOut6_9[4] , \nOut6_9[3] , \nOut6_9[2] , 
        \nOut6_9[1] , \nOut6_9[0] }), .EastIn({\nOut7_8[7] , \nOut7_8[6] , 
        \nOut7_8[5] , \nOut7_8[4] , \nOut7_8[3] , \nOut7_8[2] , \nOut7_8[1] , 
        \nOut7_8[0] }), .WestIn({\nOut5_8[7] , \nOut5_8[6] , \nOut5_8[5] , 
        \nOut5_8[4] , \nOut5_8[3] , \nOut5_8[2] , \nOut5_8[1] , \nOut5_8[0] }), 
        .Out({\nOut6_8[7] , \nOut6_8[6] , \nOut6_8[5] , \nOut6_8[4] , 
        \nOut6_8[3] , \nOut6_8[2] , \nOut6_8[1] , \nOut6_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_123 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut124[7] , \nScanOut124[6] , 
        \nScanOut124[5] , \nScanOut124[4] , \nScanOut124[3] , \nScanOut124[2] , 
        \nScanOut124[1] , \nScanOut124[0] }), .ScanOut({\nScanOut123[7] , 
        \nScanOut123[6] , \nScanOut123[5] , \nScanOut123[4] , \nScanOut123[3] , 
        \nScanOut123[2] , \nScanOut123[1] , \nScanOut123[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_10[7] , \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , 
        \nOut7_10[3] , \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), 
        .SouthIn({\nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }), .EastIn(
        {\nOut8_11[7] , \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , 
        \nOut8_11[3] , \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .WestIn(
        {\nOut6_11[7] , \nOut6_11[6] , \nOut6_11[5] , \nOut6_11[4] , 
        \nOut6_11[3] , \nOut6_11[2] , \nOut6_11[1] , \nOut6_11[0] }), .Out({
        \nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_124 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut125[7] , \nScanOut125[6] , 
        \nScanOut125[5] , \nScanOut125[4] , \nScanOut125[3] , \nScanOut125[2] , 
        \nScanOut125[1] , \nScanOut125[0] }), .ScanOut({\nScanOut124[7] , 
        \nScanOut124[6] , \nScanOut124[5] , \nScanOut124[4] , \nScanOut124[3] , 
        \nScanOut124[2] , \nScanOut124[1] , \nScanOut124[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_11[7] , \nOut7_11[6] , \nOut7_11[5] , \nOut7_11[4] , 
        \nOut7_11[3] , \nOut7_11[2] , \nOut7_11[1] , \nOut7_11[0] }), 
        .SouthIn({\nOut7_13[7] , \nOut7_13[6] , \nOut7_13[5] , \nOut7_13[4] , 
        \nOut7_13[3] , \nOut7_13[2] , \nOut7_13[1] , \nOut7_13[0] }), .EastIn(
        {\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .WestIn(
        {\nOut6_12[7] , \nOut6_12[6] , \nOut6_12[5] , \nOut6_12[4] , 
        \nOut6_12[3] , \nOut6_12[2] , \nOut6_12[1] , \nOut6_12[0] }), .Out({
        \nOut7_12[7] , \nOut7_12[6] , \nOut7_12[5] , \nOut7_12[4] , 
        \nOut7_12[3] , \nOut7_12[2] , \nOut7_12[1] , \nOut7_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_214 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut215[7] , \nScanOut215[6] , 
        \nScanOut215[5] , \nScanOut215[4] , \nScanOut215[3] , \nScanOut215[2] , 
        \nScanOut215[1] , \nScanOut215[0] }), .ScanOut({\nScanOut214[7] , 
        \nScanOut214[6] , \nScanOut214[5] , \nScanOut214[4] , \nScanOut214[3] , 
        \nScanOut214[2] , \nScanOut214[1] , \nScanOut214[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }), 
        .SouthIn({\nOut13_7[7] , \nOut13_7[6] , \nOut13_7[5] , \nOut13_7[4] , 
        \nOut13_7[3] , \nOut13_7[2] , \nOut13_7[1] , \nOut13_7[0] }), .EastIn(
        {\nOut14_6[7] , \nOut14_6[6] , \nOut14_6[5] , \nOut14_6[4] , 
        \nOut14_6[3] , \nOut14_6[2] , \nOut14_6[1] , \nOut14_6[0] }), .WestIn(
        {\nOut12_6[7] , \nOut12_6[6] , \nOut12_6[5] , \nOut12_6[4] , 
        \nOut12_6[3] , \nOut12_6[2] , \nOut12_6[1] , \nOut12_6[0] }), .Out({
        \nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_233 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut234[7] , \nScanOut234[6] , 
        \nScanOut234[5] , \nScanOut234[4] , \nScanOut234[3] , \nScanOut234[2] , 
        \nScanOut234[1] , \nScanOut234[0] }), .ScanOut({\nScanOut233[7] , 
        \nScanOut233[6] , \nScanOut233[5] , \nScanOut233[4] , \nScanOut233[3] , 
        \nScanOut233[2] , \nScanOut233[1] , \nScanOut233[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_8[7] , \nOut14_8[6] , \nOut14_8[5] , \nOut14_8[4] , 
        \nOut14_8[3] , \nOut14_8[2] , \nOut14_8[1] , \nOut14_8[0] }), 
        .SouthIn({\nOut14_10[7] , \nOut14_10[6] , \nOut14_10[5] , 
        \nOut14_10[4] , \nOut14_10[3] , \nOut14_10[2] , \nOut14_10[1] , 
        \nOut14_10[0] }), .EastIn({\nOut15_9[7] , \nOut15_9[6] , \nOut15_9[5] , 
        \nOut15_9[4] , \nOut15_9[3] , \nOut15_9[2] , \nOut15_9[1] , 
        \nOut15_9[0] }), .WestIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }), .Out({\nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , 
        \nOut14_9[4] , \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , 
        \nOut14_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_188 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut189[7] , \nScanOut189[6] , 
        \nScanOut189[5] , \nScanOut189[4] , \nScanOut189[3] , \nScanOut189[2] , 
        \nScanOut189[1] , \nScanOut189[0] }), .ScanOut({\nScanOut188[7] , 
        \nScanOut188[6] , \nScanOut188[5] , \nScanOut188[4] , \nScanOut188[3] , 
        \nScanOut188[2] , \nScanOut188[1] , \nScanOut188[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_11[7] , \nOut11_11[6] , \nOut11_11[5] , \nOut11_11[4] , 
        \nOut11_11[3] , \nOut11_11[2] , \nOut11_11[1] , \nOut11_11[0] }), 
        .SouthIn({\nOut11_13[7] , \nOut11_13[6] , \nOut11_13[5] , 
        \nOut11_13[4] , \nOut11_13[3] , \nOut11_13[2] , \nOut11_13[1] , 
        \nOut11_13[0] }), .EastIn({\nOut12_12[7] , \nOut12_12[6] , 
        \nOut12_12[5] , \nOut12_12[4] , \nOut12_12[3] , \nOut12_12[2] , 
        \nOut12_12[1] , \nOut12_12[0] }), .WestIn({\nOut10_12[7] , 
        \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , \nOut10_12[3] , 
        \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), .Out({\nOut11_12[7] , 
        \nOut11_12[6] , \nOut11_12[5] , \nOut11_12[4] , \nOut11_12[3] , 
        \nOut11_12[2] , \nOut11_12[1] , \nOut11_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_213 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut214[7] , \nScanOut214[6] , 
        \nScanOut214[5] , \nScanOut214[4] , \nScanOut214[3] , \nScanOut214[2] , 
        \nScanOut214[1] , \nScanOut214[0] }), .ScanOut({\nScanOut213[7] , 
        \nScanOut213[6] , \nScanOut213[5] , \nScanOut213[4] , \nScanOut213[3] , 
        \nScanOut213[2] , \nScanOut213[1] , \nScanOut213[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut13_4[7] , \nOut13_4[6] , \nOut13_4[5] , \nOut13_4[4] , 
        \nOut13_4[3] , \nOut13_4[2] , \nOut13_4[1] , \nOut13_4[0] }), 
        .SouthIn({\nOut13_6[7] , \nOut13_6[6] , \nOut13_6[5] , \nOut13_6[4] , 
        \nOut13_6[3] , \nOut13_6[2] , \nOut13_6[1] , \nOut13_6[0] }), .EastIn(
        {\nOut14_5[7] , \nOut14_5[6] , \nOut14_5[5] , \nOut14_5[4] , 
        \nOut14_5[3] , \nOut14_5[2] , \nOut14_5[1] , \nOut14_5[0] }), .WestIn(
        {\nOut12_5[7] , \nOut12_5[6] , \nOut12_5[5] , \nOut12_5[4] , 
        \nOut12_5[3] , \nOut12_5[2] , \nOut12_5[1] , \nOut12_5[0] }), .Out({
        \nOut13_5[7] , \nOut13_5[6] , \nOut13_5[5] , \nOut13_5[4] , 
        \nOut13_5[3] , \nOut13_5[2] , \nOut13_5[1] , \nOut13_5[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_234 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut235[7] , \nScanOut235[6] , 
        \nScanOut235[5] , \nScanOut235[4] , \nScanOut235[3] , \nScanOut235[2] , 
        \nScanOut235[1] , \nScanOut235[0] }), .ScanOut({\nScanOut234[7] , 
        \nScanOut234[6] , \nScanOut234[5] , \nScanOut234[4] , \nScanOut234[3] , 
        \nScanOut234[2] , \nScanOut234[1] , \nScanOut234[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_9[7] , \nOut14_9[6] , \nOut14_9[5] , \nOut14_9[4] , 
        \nOut14_9[3] , \nOut14_9[2] , \nOut14_9[1] , \nOut14_9[0] }), 
        .SouthIn({\nOut14_11[7] , \nOut14_11[6] , \nOut14_11[5] , 
        \nOut14_11[4] , \nOut14_11[3] , \nOut14_11[2] , \nOut14_11[1] , 
        \nOut14_11[0] }), .EastIn({\nOut15_10[7] , \nOut15_10[6] , 
        \nOut15_10[5] , \nOut15_10[4] , \nOut15_10[3] , \nOut15_10[2] , 
        \nOut15_10[1] , \nOut15_10[0] }), .WestIn({\nOut13_10[7] , 
        \nOut13_10[6] , \nOut13_10[5] , \nOut13_10[4] , \nOut13_10[3] , 
        \nOut13_10[2] , \nOut13_10[1] , \nOut13_10[0] }), .Out({\nOut14_10[7] , 
        \nOut14_10[6] , \nOut14_10[5] , \nOut14_10[4] , \nOut14_10[3] , 
        \nOut14_10[2] , \nOut14_10[1] , \nOut14_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_156 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut157[7] , \nScanOut157[6] , 
        \nScanOut157[5] , \nScanOut157[4] , \nScanOut157[3] , \nScanOut157[2] , 
        \nScanOut157[1] , \nScanOut157[0] }), .ScanOut({\nScanOut156[7] , 
        \nScanOut156[6] , \nScanOut156[5] , \nScanOut156[4] , \nScanOut156[3] , 
        \nScanOut156[2] , \nScanOut156[1] , \nScanOut156[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut9_11[7] , \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , 
        \nOut9_11[3] , \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), 
        .SouthIn({\nOut9_13[7] , \nOut9_13[6] , \nOut9_13[5] , \nOut9_13[4] , 
        \nOut9_13[3] , \nOut9_13[2] , \nOut9_13[1] , \nOut9_13[0] }), .EastIn(
        {\nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , \nOut10_12[4] , 
        \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , \nOut10_12[0] }), 
        .WestIn({\nOut8_12[7] , \nOut8_12[6] , \nOut8_12[5] , \nOut8_12[4] , 
        \nOut8_12[3] , \nOut8_12[2] , \nOut8_12[1] , \nOut8_12[0] }), .Out({
        \nOut9_12[7] , \nOut9_12[6] , \nOut9_12[5] , \nOut9_12[4] , 
        \nOut9_12[3] , \nOut9_12[2] , \nOut9_12[1] , \nOut9_12[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_171 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut172[7] , \nScanOut172[6] , 
        \nScanOut172[5] , \nScanOut172[4] , \nScanOut172[3] , \nScanOut172[2] , 
        \nScanOut172[1] , \nScanOut172[0] }), .ScanOut({\nScanOut171[7] , 
        \nScanOut171[6] , \nScanOut171[5] , \nScanOut171[4] , \nScanOut171[3] , 
        \nScanOut171[2] , \nScanOut171[1] , \nScanOut171[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_10[7] , \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , 
        \nOut10_10[3] , \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), 
        .SouthIn({\nOut10_12[7] , \nOut10_12[6] , \nOut10_12[5] , 
        \nOut10_12[4] , \nOut10_12[3] , \nOut10_12[2] , \nOut10_12[1] , 
        \nOut10_12[0] }), .EastIn({\nOut11_11[7] , \nOut11_11[6] , 
        \nOut11_11[5] , \nOut11_11[4] , \nOut11_11[3] , \nOut11_11[2] , 
        \nOut11_11[1] , \nOut11_11[0] }), .WestIn({\nOut9_11[7] , 
        \nOut9_11[6] , \nOut9_11[5] , \nOut9_11[4] , \nOut9_11[3] , 
        \nOut9_11[2] , \nOut9_11[1] , \nOut9_11[0] }), .Out({\nOut10_11[7] , 
        \nOut10_11[6] , \nOut10_11[5] , \nOut10_11[4] , \nOut10_11[3] , 
        \nOut10_11[2] , \nOut10_11[1] , \nOut10_11[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_241 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut242[7] , \nScanOut242[6] , 
        \nScanOut242[5] , \nScanOut242[4] , \nScanOut242[3] , \nScanOut242[2] , 
        \nScanOut242[1] , \nScanOut242[0] }), .ScanOut({\nScanOut241[7] , 
        \nScanOut241[6] , \nScanOut241[5] , \nScanOut241[4] , \nScanOut241[3] , 
        \nScanOut241[2] , \nScanOut241[1] , \nScanOut241[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_1[7] , \nOut15_1[6] , 
        \nOut15_1[5] , \nOut15_1[4] , \nOut15_1[3] , \nOut15_1[2] , 
        \nOut15_1[1] , \nOut15_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_194 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut195[7] , \nScanOut195[6] , 
        \nScanOut195[5] , \nScanOut195[4] , \nScanOut195[3] , \nScanOut195[2] , 
        \nScanOut195[1] , \nScanOut195[0] }), .ScanOut({\nScanOut194[7] , 
        \nScanOut194[6] , \nScanOut194[5] , \nScanOut194[4] , \nScanOut194[3] , 
        \nScanOut194[2] , \nScanOut194[1] , \nScanOut194[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_1[7] , \nOut12_1[6] , \nOut12_1[5] , \nOut12_1[4] , 
        \nOut12_1[3] , \nOut12_1[2] , \nOut12_1[1] , \nOut12_1[0] }), 
        .SouthIn({\nOut12_3[7] , \nOut12_3[6] , \nOut12_3[5] , \nOut12_3[4] , 
        \nOut12_3[3] , \nOut12_3[2] , \nOut12_3[1] , \nOut12_3[0] }), .EastIn(
        {\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .WestIn(
        {\nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }), .Out({
        \nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_99 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut100[7] , \nScanOut100[6] , 
        \nScanOut100[5] , \nScanOut100[4] , \nScanOut100[3] , \nScanOut100[2] , 
        \nScanOut100[1] , \nScanOut100[0] }), .ScanOut({\nScanOut99[7] , 
        \nScanOut99[6] , \nScanOut99[5] , \nScanOut99[4] , \nScanOut99[3] , 
        \nScanOut99[2] , \nScanOut99[1] , \nScanOut99[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut6_2[7] , \nOut6_2[6] , \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , 
        \nOut6_2[2] , \nOut6_2[1] , \nOut6_2[0] }), .SouthIn({\nOut6_4[7] , 
        \nOut6_4[6] , \nOut6_4[5] , \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , 
        \nOut6_4[1] , \nOut6_4[0] }), .EastIn({\nOut7_3[7] , \nOut7_3[6] , 
        \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , 
        \nOut7_3[0] }), .WestIn({\nOut5_3[7] , \nOut5_3[6] , \nOut5_3[5] , 
        \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , \nOut5_3[0] }), 
        .Out({\nOut6_3[7] , \nOut6_3[6] , \nOut6_3[5] , \nOut6_3[4] , 
        \nOut6_3[3] , \nOut6_3[2] , \nOut6_3[1] , \nOut6_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_138 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut139[7] , \nScanOut139[6] , 
        \nScanOut139[5] , \nScanOut139[4] , \nScanOut139[3] , \nScanOut139[2] , 
        \nScanOut139[1] , \nScanOut139[0] }), .ScanOut({\nScanOut138[7] , 
        \nScanOut138[6] , \nScanOut138[5] , \nScanOut138[4] , \nScanOut138[3] , 
        \nScanOut138[2] , \nScanOut138[1] , \nScanOut138[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_9[7] , \nOut8_9[6] , \nOut8_9[5] , \nOut8_9[4] , \nOut8_9[3] , 
        \nOut8_9[2] , \nOut8_9[1] , \nOut8_9[0] }), .SouthIn({\nOut8_11[7] , 
        \nOut8_11[6] , \nOut8_11[5] , \nOut8_11[4] , \nOut8_11[3] , 
        \nOut8_11[2] , \nOut8_11[1] , \nOut8_11[0] }), .EastIn({\nOut9_10[7] , 
        \nOut9_10[6] , \nOut9_10[5] , \nOut9_10[4] , \nOut9_10[3] , 
        \nOut9_10[2] , \nOut9_10[1] , \nOut9_10[0] }), .WestIn({\nOut7_10[7] , 
        \nOut7_10[6] , \nOut7_10[5] , \nOut7_10[4] , \nOut7_10[3] , 
        \nOut7_10[2] , \nOut7_10[1] , \nOut7_10[0] }), .Out({\nOut8_10[7] , 
        \nOut8_10[6] , \nOut8_10[5] , \nOut8_10[4] , \nOut8_10[3] , 
        \nOut8_10[2] , \nOut8_10[1] , \nOut8_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_208 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut209[7] , \nScanOut209[6] , 
        \nScanOut209[5] , \nScanOut209[4] , \nScanOut209[3] , \nScanOut209[2] , 
        \nScanOut209[1] , \nScanOut209[0] }), .ScanOut({\nScanOut208[7] , 
        \nScanOut208[6] , \nScanOut208[5] , \nScanOut208[4] , \nScanOut208[3] , 
        \nScanOut208[2] , \nScanOut208[1] , \nScanOut208[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut13_0[7] , \nOut13_0[6] , 
        \nOut13_0[5] , \nOut13_0[4] , \nOut13_0[3] , \nOut13_0[2] , 
        \nOut13_0[1] , \nOut13_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_186 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut187[7] , \nScanOut187[6] , 
        \nScanOut187[5] , \nScanOut187[4] , \nScanOut187[3] , \nScanOut187[2] , 
        \nScanOut187[1] , \nScanOut187[0] }), .ScanOut({\nScanOut186[7] , 
        \nScanOut186[6] , \nScanOut186[5] , \nScanOut186[4] , \nScanOut186[3] , 
        \nScanOut186[2] , \nScanOut186[1] , \nScanOut186[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , \nOut11_9[4] , 
        \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , \nOut11_9[0] }), 
        .SouthIn({\nOut11_11[7] , \nOut11_11[6] , \nOut11_11[5] , 
        \nOut11_11[4] , \nOut11_11[3] , \nOut11_11[2] , \nOut11_11[1] , 
        \nOut11_11[0] }), .EastIn({\nOut12_10[7] , \nOut12_10[6] , 
        \nOut12_10[5] , \nOut12_10[4] , \nOut12_10[3] , \nOut12_10[2] , 
        \nOut12_10[1] , \nOut12_10[0] }), .WestIn({\nOut10_10[7] , 
        \nOut10_10[6] , \nOut10_10[5] , \nOut10_10[4] , \nOut10_10[3] , 
        \nOut10_10[2] , \nOut10_10[1] , \nOut10_10[0] }), .Out({\nOut11_10[7] , 
        \nOut11_10[6] , \nOut11_10[5] , \nOut11_10[4] , \nOut11_10[3] , 
        \nOut11_10[2] , \nOut11_10[1] , \nOut11_10[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_35 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut36[7] , \nScanOut36[6] , 
        \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , 
        \nScanOut36[1] , \nScanOut36[0] }), .ScanOut({\nScanOut35[7] , 
        \nScanOut35[6] , \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , 
        \nScanOut35[2] , \nScanOut35[1] , \nScanOut35[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , 
        \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), .SouthIn({\nOut2_4[7] , 
        \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , 
        \nOut2_4[1] , \nOut2_4[0] }), .EastIn({\nOut3_3[7] , \nOut3_3[6] , 
        \nOut3_3[5] , \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , 
        \nOut3_3[0] }), .WestIn({\nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , 
        \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), 
        .Out({\nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , 
        \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_40 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut41[7] , \nScanOut41[6] , 
        \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , 
        \nScanOut41[1] , \nScanOut41[0] }), .ScanOut({\nScanOut40[7] , 
        \nScanOut40[6] , \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , 
        \nScanOut40[2] , \nScanOut40[1] , \nScanOut40[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , 
        \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), .SouthIn({\nOut2_9[7] , 
        \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , 
        \nOut2_9[1] , \nOut2_9[0] }), .EastIn({\nOut3_8[7] , \nOut3_8[6] , 
        \nOut3_8[5] , \nOut3_8[4] , \nOut3_8[3] , \nOut3_8[2] , \nOut3_8[1] , 
        \nOut3_8[0] }), .WestIn({\nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , 
        \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), 
        .Out({\nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , 
        \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_67 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut68[7] , \nScanOut68[6] , 
        \nScanOut68[5] , \nScanOut68[4] , \nScanOut68[3] , \nScanOut68[2] , 
        \nScanOut68[1] , \nScanOut68[0] }), .ScanOut({\nScanOut67[7] , 
        \nScanOut67[6] , \nScanOut67[5] , \nScanOut67[4] , \nScanOut67[3] , 
        \nScanOut67[2] , \nScanOut67[1] , \nScanOut67[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , \nOut4_2[4] , \nOut4_2[3] , 
        \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }), .SouthIn({\nOut4_4[7] , 
        \nOut4_4[6] , \nOut4_4[5] , \nOut4_4[4] , \nOut4_4[3] , \nOut4_4[2] , 
        \nOut4_4[1] , \nOut4_4[0] }), .EastIn({\nOut5_3[7] , \nOut5_3[6] , 
        \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , \nOut5_3[1] , 
        \nOut5_3[0] }), .WestIn({\nOut3_3[7] , \nOut3_3[6] , \nOut3_3[5] , 
        \nOut3_3[4] , \nOut3_3[3] , \nOut3_3[2] , \nOut3_3[1] , \nOut3_3[0] }), 
        .Out({\nOut4_3[7] , \nOut4_3[6] , \nOut4_3[5] , \nOut4_3[4] , 
        \nOut4_3[3] , \nOut4_3[2] , \nOut4_3[1] , \nOut4_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_144 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut145[7] , \nScanOut145[6] , 
        \nScanOut145[5] , \nScanOut145[4] , \nScanOut145[3] , \nScanOut145[2] , 
        \nScanOut145[1] , \nScanOut145[0] }), .ScanOut({\nScanOut144[7] , 
        \nScanOut144[6] , \nScanOut144[5] , \nScanOut144[4] , \nScanOut144[3] , 
        \nScanOut144[2] , \nScanOut144[1] , \nScanOut144[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut9_0[7] , \nOut9_0[6] , 
        \nOut9_0[5] , \nOut9_0[4] , \nOut9_0[3] , \nOut9_0[2] , \nOut9_0[1] , 
        \nOut9_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_163 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut164[7] , \nScanOut164[6] , 
        \nScanOut164[5] , \nScanOut164[4] , \nScanOut164[3] , \nScanOut164[2] , 
        \nScanOut164[1] , \nScanOut164[0] }), .ScanOut({\nScanOut163[7] , 
        \nScanOut163[6] , \nScanOut163[5] , \nScanOut163[4] , \nScanOut163[3] , 
        \nScanOut163[2] , \nScanOut163[1] , \nScanOut163[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), 
        .SouthIn({\nOut10_4[7] , \nOut10_4[6] , \nOut10_4[5] , \nOut10_4[4] , 
        \nOut10_4[3] , \nOut10_4[2] , \nOut10_4[1] , \nOut10_4[0] }), .EastIn(
        {\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .WestIn(
        {\nOut9_3[7] , \nOut9_3[6] , \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , 
        \nOut9_3[2] , \nOut9_3[1] , \nOut9_3[0] }), .Out({\nOut10_3[7] , 
        \nOut10_3[6] , \nOut10_3[5] , \nOut10_3[4] , \nOut10_3[3] , 
        \nOut10_3[2] , \nOut10_3[1] , \nOut10_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_178 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut179[7] , \nScanOut179[6] , 
        \nScanOut179[5] , \nScanOut179[4] , \nScanOut179[3] , \nScanOut179[2] , 
        \nScanOut179[1] , \nScanOut179[0] }), .ScanOut({\nScanOut178[7] , 
        \nScanOut178[6] , \nScanOut178[5] , \nScanOut178[4] , \nScanOut178[3] , 
        \nScanOut178[2] , \nScanOut178[1] , \nScanOut178[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut11_1[7] , \nOut11_1[6] , \nOut11_1[5] , \nOut11_1[4] , 
        \nOut11_1[3] , \nOut11_1[2] , \nOut11_1[1] , \nOut11_1[0] }), 
        .SouthIn({\nOut11_3[7] , \nOut11_3[6] , \nOut11_3[5] , \nOut11_3[4] , 
        \nOut11_3[3] , \nOut11_3[2] , \nOut11_3[1] , \nOut11_3[0] }), .EastIn(
        {\nOut12_2[7] , \nOut12_2[6] , \nOut12_2[5] , \nOut12_2[4] , 
        \nOut12_2[3] , \nOut12_2[2] , \nOut12_2[1] , \nOut12_2[0] }), .WestIn(
        {\nOut10_2[7] , \nOut10_2[6] , \nOut10_2[5] , \nOut10_2[4] , 
        \nOut10_2[3] , \nOut10_2[2] , \nOut10_2[1] , \nOut10_2[0] }), .Out({
        \nOut11_2[7] , \nOut11_2[6] , \nOut11_2[5] , \nOut11_2[4] , 
        \nOut11_2[3] , \nOut11_2[2] , \nOut11_2[1] , \nOut11_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_248 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut249[7] , \nScanOut249[6] , 
        \nScanOut249[5] , \nScanOut249[4] , \nScanOut249[3] , \nScanOut249[2] , 
        \nScanOut249[1] , \nScanOut249[0] }), .ScanOut({\nScanOut248[7] , 
        \nScanOut248[6] , \nScanOut248[5] , \nScanOut248[4] , \nScanOut248[3] , 
        \nScanOut248[2] , \nScanOut248[1] , \nScanOut248[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_8[7] , \nOut15_8[6] , 
        \nOut15_8[5] , \nOut15_8[4] , \nOut15_8[3] , \nOut15_8[2] , 
        \nOut15_8[1] , \nOut15_8[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_253 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut254[7] , \nScanOut254[6] , 
        \nScanOut254[5] , \nScanOut254[4] , \nScanOut254[3] , \nScanOut254[2] , 
        \nScanOut254[1] , \nScanOut254[0] }), .ScanOut({\nScanOut253[7] , 
        \nScanOut253[6] , \nScanOut253[5] , \nScanOut253[4] , \nScanOut253[3] , 
        \nScanOut253[2] , \nScanOut253[1] , \nScanOut253[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut15_13[7] , \nOut15_13[6] , 
        \nOut15_13[5] , \nOut15_13[4] , \nOut15_13[3] , \nOut15_13[2] , 
        \nOut15_13[1] , \nOut15_13[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_82 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut83[7] , \nScanOut83[6] , 
        \nScanOut83[5] , \nScanOut83[4] , \nScanOut83[3] , \nScanOut83[2] , 
        \nScanOut83[1] , \nScanOut83[0] }), .ScanOut({\nScanOut82[7] , 
        \nScanOut82[6] , \nScanOut82[5] , \nScanOut82[4] , \nScanOut82[3] , 
        \nScanOut82[2] , \nScanOut82[1] , \nScanOut82[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut5_1[7] , \nOut5_1[6] , \nOut5_1[5] , \nOut5_1[4] , \nOut5_1[3] , 
        \nOut5_1[2] , \nOut5_1[1] , \nOut5_1[0] }), .SouthIn({\nOut5_3[7] , 
        \nOut5_3[6] , \nOut5_3[5] , \nOut5_3[4] , \nOut5_3[3] , \nOut5_3[2] , 
        \nOut5_3[1] , \nOut5_3[0] }), .EastIn({\nOut6_2[7] , \nOut6_2[6] , 
        \nOut6_2[5] , \nOut6_2[4] , \nOut6_2[3] , \nOut6_2[2] , \nOut6_2[1] , 
        \nOut6_2[0] }), .WestIn({\nOut4_2[7] , \nOut4_2[6] , \nOut4_2[5] , 
        \nOut4_2[4] , \nOut4_2[3] , \nOut4_2[2] , \nOut4_2[1] , \nOut4_2[0] }), 
        .Out({\nOut5_2[7] , \nOut5_2[6] , \nOut5_2[5] , \nOut5_2[4] , 
        \nOut5_2[3] , \nOut5_2[2] , \nOut5_2[1] , \nOut5_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_116 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut117[7] , \nScanOut117[6] , 
        \nScanOut117[5] , \nScanOut117[4] , \nScanOut117[3] , \nScanOut117[2] , 
        \nScanOut117[1] , \nScanOut117[0] }), .ScanOut({\nScanOut116[7] , 
        \nScanOut116[6] , \nScanOut116[5] , \nScanOut116[4] , \nScanOut116[3] , 
        \nScanOut116[2] , \nScanOut116[1] , \nScanOut116[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , \nOut7_3[4] , \nOut7_3[3] , 
        \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }), .SouthIn({\nOut7_5[7] , 
        \nOut7_5[6] , \nOut7_5[5] , \nOut7_5[4] , \nOut7_5[3] , \nOut7_5[2] , 
        \nOut7_5[1] , \nOut7_5[0] }), .EastIn({\nOut8_4[7] , \nOut8_4[6] , 
        \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , \nOut8_4[1] , 
        \nOut8_4[0] }), .WestIn({\nOut6_4[7] , \nOut6_4[6] , \nOut6_4[5] , 
        \nOut6_4[4] , \nOut6_4[3] , \nOut6_4[2] , \nOut6_4[1] , \nOut6_4[0] }), 
        .Out({\nOut7_4[7] , \nOut7_4[6] , \nOut7_4[5] , \nOut7_4[4] , 
        \nOut7_4[3] , \nOut7_4[2] , \nOut7_4[1] , \nOut7_4[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_131 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut132[7] , \nScanOut132[6] , 
        \nScanOut132[5] , \nScanOut132[4] , \nScanOut132[3] , \nScanOut132[2] , 
        \nScanOut132[1] , \nScanOut132[0] }), .ScanOut({\nScanOut131[7] , 
        \nScanOut131[6] , \nScanOut131[5] , \nScanOut131[4] , \nScanOut131[3] , 
        \nScanOut131[2] , \nScanOut131[1] , \nScanOut131[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut8_2[7] , \nOut8_2[6] , \nOut8_2[5] , \nOut8_2[4] , \nOut8_2[3] , 
        \nOut8_2[2] , \nOut8_2[1] , \nOut8_2[0] }), .SouthIn({\nOut8_4[7] , 
        \nOut8_4[6] , \nOut8_4[5] , \nOut8_4[4] , \nOut8_4[3] , \nOut8_4[2] , 
        \nOut8_4[1] , \nOut8_4[0] }), .EastIn({\nOut9_3[7] , \nOut9_3[6] , 
        \nOut9_3[5] , \nOut9_3[4] , \nOut9_3[3] , \nOut9_3[2] , \nOut9_3[1] , 
        \nOut9_3[0] }), .WestIn({\nOut7_3[7] , \nOut7_3[6] , \nOut7_3[5] , 
        \nOut7_3[4] , \nOut7_3[3] , \nOut7_3[2] , \nOut7_3[1] , \nOut7_3[0] }), 
        .Out({\nOut8_3[7] , \nOut8_3[6] , \nOut8_3[5] , \nOut8_3[4] , 
        \nOut8_3[3] , \nOut8_3[2] , \nOut8_3[1] , \nOut8_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_201 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut202[7] , \nScanOut202[6] , 
        \nScanOut202[5] , \nScanOut202[4] , \nScanOut202[3] , \nScanOut202[2] , 
        \nScanOut202[1] , \nScanOut202[0] }), .ScanOut({\nScanOut201[7] , 
        \nScanOut201[6] , \nScanOut201[5] , \nScanOut201[4] , \nScanOut201[3] , 
        \nScanOut201[2] , \nScanOut201[1] , \nScanOut201[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut12_8[7] , \nOut12_8[6] , \nOut12_8[5] , \nOut12_8[4] , 
        \nOut12_8[3] , \nOut12_8[2] , \nOut12_8[1] , \nOut12_8[0] }), 
        .SouthIn({\nOut12_10[7] , \nOut12_10[6] , \nOut12_10[5] , 
        \nOut12_10[4] , \nOut12_10[3] , \nOut12_10[2] , \nOut12_10[1] , 
        \nOut12_10[0] }), .EastIn({\nOut13_9[7] , \nOut13_9[6] , \nOut13_9[5] , 
        \nOut13_9[4] , \nOut13_9[3] , \nOut13_9[2] , \nOut13_9[1] , 
        \nOut13_9[0] }), .WestIn({\nOut11_9[7] , \nOut11_9[6] , \nOut11_9[5] , 
        \nOut11_9[4] , \nOut11_9[3] , \nOut11_9[2] , \nOut11_9[1] , 
        \nOut11_9[0] }), .Out({\nOut12_9[7] , \nOut12_9[6] , \nOut12_9[5] , 
        \nOut12_9[4] , \nOut12_9[3] , \nOut12_9[2] , \nOut12_9[1] , 
        \nOut12_9[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_226 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut227[7] , \nScanOut227[6] , 
        \nScanOut227[5] , \nScanOut227[4] , \nScanOut227[3] , \nScanOut227[2] , 
        \nScanOut227[1] , \nScanOut227[0] }), .ScanOut({\nScanOut226[7] , 
        \nScanOut226[6] , \nScanOut226[5] , \nScanOut226[4] , \nScanOut226[3] , 
        \nScanOut226[2] , \nScanOut226[1] , \nScanOut226[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut14_1[7] , \nOut14_1[6] , \nOut14_1[5] , \nOut14_1[4] , 
        \nOut14_1[3] , \nOut14_1[2] , \nOut14_1[1] , \nOut14_1[0] }), 
        .SouthIn({\nOut14_3[7] , \nOut14_3[6] , \nOut14_3[5] , \nOut14_3[4] , 
        \nOut14_3[3] , \nOut14_3[2] , \nOut14_3[1] , \nOut14_3[0] }), .EastIn(
        {\nOut15_2[7] , \nOut15_2[6] , \nOut15_2[5] , \nOut15_2[4] , 
        \nOut15_2[3] , \nOut15_2[2] , \nOut15_2[1] , \nOut15_2[0] }), .WestIn(
        {\nOut13_2[7] , \nOut13_2[6] , \nOut13_2[5] , \nOut13_2[4] , 
        \nOut13_2[3] , \nOut13_2[2] , \nOut13_2[1] , \nOut13_2[0] }), .Out({
        \nOut14_2[7] , \nOut14_2[6] , \nOut14_2[5] , \nOut14_2[4] , 
        \nOut14_2[3] , \nOut14_2[2] , \nOut14_2[1] , \nOut14_2[0] }) );
endmodule

