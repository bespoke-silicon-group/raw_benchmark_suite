
module BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, 
        n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, 
        n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, 
        n94, n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, 
        n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, 
        n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, 
        n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n110) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n107), .D(n102), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[25]), .Z(n101) );
    VMW_INV U92 ( .A(A[28]), .Z(n103) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(B[25]), .Z(n98) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[24]), .Z(n90) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BubbleSort_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, 
    AIn, BIn, HiOut, LoOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] LoOut;
input  [31:0] AIn;
input  [31:0] BIn;
output [31:0] HiOut;
input  Clk, Reset, RD, WR;
    wire n159, a58;
    VMW_PULLDOWN U21 ( .Z(n159) );
    VMW_MUX2 U54 ( .A(BIn[9]), .B(AIn[9]), .S(a58), .Z(HiOut[9]) );
    VMW_MUX2 U73 ( .A(BIn[20]), .B(AIn[20]), .S(a58), .Z(HiOut[20]) );
    VMW_MUX2 U22 ( .A(AIn[9]), .B(BIn[9]), .S(a58), .Z(LoOut[9]) );
    VMW_MUX2 U26 ( .A(AIn[5]), .B(BIn[5]), .S(a58), .Z(LoOut[5]) );
    VMW_MUX2 U28 ( .A(AIn[3]), .B(BIn[3]), .S(a58), .Z(LoOut[3]) );
    VMW_MUX2 U33 ( .A(AIn[28]), .B(BIn[28]), .S(a58), .Z(LoOut[28]) );
    VMW_MUX2 U68 ( .A(BIn[25]), .B(AIn[25]), .S(a58), .Z(HiOut[25]) );
    VMW_MUX2 U34 ( .A(AIn[27]), .B(BIn[27]), .S(a58), .Z(LoOut[27]) );
    VMW_MUX2 U41 ( .A(AIn[20]), .B(BIn[20]), .S(a58), .Z(LoOut[20]) );
    VMW_MUX2 U46 ( .A(AIn[16]), .B(BIn[16]), .S(a58), .Z(LoOut[16]) );
    VMW_MUX2 U61 ( .A(BIn[31]), .B(AIn[31]), .S(a58), .Z(HiOut[31]) );
    VMW_MUX2 U84 ( .A(BIn[10]), .B(AIn[10]), .S(a58), .Z(HiOut[10]) );
    VMW_MUX2 U66 ( .A(BIn[27]), .B(AIn[27]), .S(a58), .Z(HiOut[27]) );
    VMW_MUX2 U83 ( .A(BIn[11]), .B(AIn[11]), .S(a58), .Z(HiOut[11]) );
    VMW_MUX2 U48 ( .A(AIn[14]), .B(BIn[14]), .S(a58), .Z(LoOut[14]) );
    VMW_MUX2 U27 ( .A(AIn[4]), .B(BIn[4]), .S(a58), .Z(LoOut[4]) );
    VMW_MUX2 U35 ( .A(AIn[26]), .B(BIn[26]), .S(a58), .Z(LoOut[26]) );
    VMW_MUX2 U53 ( .A(AIn[0]), .B(BIn[0]), .S(a58), .Z(LoOut[0]) );
    VMW_MUX2 U74 ( .A(BIn[1]), .B(AIn[1]), .S(a58), .Z(HiOut[1]) );
    VMW_MUX2 U40 ( .A(AIn[21]), .B(BIn[21]), .S(a58), .Z(LoOut[21]) );
    VMW_MUX2 U82 ( .A(BIn[12]), .B(AIn[12]), .S(a58), .Z(HiOut[12]) );
    VMW_MUX2 U52 ( .A(AIn[10]), .B(BIn[10]), .S(a58), .Z(LoOut[10]) );
    VMW_MUX2 U67 ( .A(BIn[26]), .B(AIn[26]), .S(a58), .Z(HiOut[26]) );
    VMW_MUX2 U75 ( .A(BIn[19]), .B(AIn[19]), .S(a58), .Z(HiOut[19]) );
    VMW_MUX2 U29 ( .A(AIn[31]), .B(BIn[31]), .S(a58), .Z(LoOut[31]) );
    VMW_MUX2 U47 ( .A(AIn[15]), .B(BIn[15]), .S(a58), .Z(LoOut[15]) );
    VMW_MUX2 U49 ( .A(AIn[13]), .B(BIn[13]), .S(a58), .Z(LoOut[13]) );
    VMW_MUX2 U55 ( .A(BIn[8]), .B(AIn[8]), .S(a58), .Z(HiOut[8]) );
    VMW_MUX2 U69 ( .A(BIn[24]), .B(AIn[24]), .S(a58), .Z(HiOut[24]) );
    VMW_MUX2 U72 ( .A(BIn[21]), .B(AIn[21]), .S(a58), .Z(HiOut[21]) );
    VMW_MUX2 U60 ( .A(BIn[3]), .B(AIn[3]), .S(a58), .Z(HiOut[3]) );
    VMW_MUX2 U32 ( .A(AIn[29]), .B(BIn[29]), .S(a58), .Z(LoOut[29]) );
    VMW_MUX2 U85 ( .A(BIn[0]), .B(AIn[0]), .S(a58), .Z(HiOut[0]) );
    VMW_MUX2 U39 ( .A(AIn[22]), .B(BIn[22]), .S(a58), .Z(LoOut[22]) );
    VMW_MUX2 U57 ( .A(BIn[6]), .B(AIn[6]), .S(a58), .Z(HiOut[6]) );
    VMW_MUX2 U70 ( .A(BIn[23]), .B(AIn[23]), .S(a58), .Z(HiOut[23]) );
    VMW_MUX2 U23 ( .A(AIn[8]), .B(BIn[8]), .S(a58), .Z(LoOut[8]) );
    VMW_MUX2 U24 ( .A(AIn[7]), .B(BIn[7]), .S(a58), .Z(LoOut[7]) );
    VMW_MUX2 U25 ( .A(AIn[6]), .B(BIn[6]), .S(a58), .Z(LoOut[6]) );
    VMW_MUX2 U30 ( .A(AIn[30]), .B(BIn[30]), .S(a58), .Z(LoOut[30]) );
    VMW_MUX2 U79 ( .A(BIn[15]), .B(AIn[15]), .S(a58), .Z(HiOut[15]) );
    BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 gt_41 ( .A(BIn), .B(AIn), .LEQ(n159
        ), .TC(n159), .LT_LE(a58) );
    VMW_MUX2 U37 ( .A(AIn[24]), .B(BIn[24]), .S(a58), .Z(LoOut[24]) );
    VMW_MUX2 U42 ( .A(AIn[1]), .B(BIn[1]), .S(a58), .Z(LoOut[1]) );
    VMW_MUX2 U45 ( .A(AIn[17]), .B(BIn[17]), .S(a58), .Z(LoOut[17]) );
    VMW_MUX2 U62 ( .A(BIn[30]), .B(AIn[30]), .S(a58), .Z(HiOut[30]) );
    VMW_MUX2 U65 ( .A(BIn[28]), .B(AIn[28]), .S(a58), .Z(HiOut[28]) );
    VMW_MUX2 U80 ( .A(BIn[14]), .B(AIn[14]), .S(a58), .Z(HiOut[14]) );
    VMW_MUX2 U59 ( .A(BIn[4]), .B(AIn[4]), .S(a58), .Z(HiOut[4]) );
    VMW_MUX2 U36 ( .A(AIn[25]), .B(BIn[25]), .S(a58), .Z(LoOut[25]) );
    VMW_MUX2 U50 ( .A(AIn[12]), .B(BIn[12]), .S(a58), .Z(LoOut[12]) );
    VMW_MUX2 U77 ( .A(BIn[17]), .B(AIn[17]), .S(a58), .Z(HiOut[17]) );
    VMW_MUX2 U58 ( .A(BIn[5]), .B(AIn[5]), .S(a58), .Z(HiOut[5]) );
    VMW_MUX2 U43 ( .A(AIn[19]), .B(BIn[19]), .S(a58), .Z(LoOut[19]) );
    VMW_MUX2 U64 ( .A(BIn[29]), .B(AIn[29]), .S(a58), .Z(HiOut[29]) );
    VMW_MUX2 U81 ( .A(BIn[13]), .B(AIn[13]), .S(a58), .Z(HiOut[13]) );
    VMW_MUX2 U51 ( .A(AIn[11]), .B(BIn[11]), .S(a58), .Z(LoOut[11]) );
    VMW_MUX2 U76 ( .A(BIn[18]), .B(AIn[18]), .S(a58), .Z(HiOut[18]) );
    VMW_MUX2 U31 ( .A(AIn[2]), .B(BIn[2]), .S(a58), .Z(LoOut[2]) );
    VMW_MUX2 U38 ( .A(AIn[23]), .B(BIn[23]), .S(a58), .Z(LoOut[23]) );
    VMW_MUX2 U44 ( .A(AIn[18]), .B(BIn[18]), .S(a58), .Z(LoOut[18]) );
    VMW_MUX2 U56 ( .A(BIn[7]), .B(AIn[7]), .S(a58), .Z(HiOut[7]) );
    VMW_MUX2 U71 ( .A(BIn[22]), .B(AIn[22]), .S(a58), .Z(HiOut[22]) );
    VMW_MUX2 U63 ( .A(BIn[2]), .B(AIn[2]), .S(a58), .Z(HiOut[2]) );
    VMW_MUX2 U78 ( .A(BIn[16]), .B(AIn[16]), .S(a58), .Z(HiOut[16]) );
endmodule


module BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, In, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[31] , \ScanOut[5]1 , \ScanOut[4]1 , n245, n262, n217, n230, 
        n222, n199, n205, n257, n239, \ScanOut[23]1 , \ScanOut[8]1 , n202, 
        n250, n219, n225, n259, n210, n237, \ScanOut[10]1 , \ScanOut[22]1 , 
        \ScanOut[11]1 , n242, \ScanOut[9]1 , n197, n203, n224, n251, n206, 
        \ScanOut[19]1 , n196, n218, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , \ScanOut[0]1 , n258, n243, \ScanOut[15]1 , n211, n236, 
        n216, n231, \ScanOut[27]1 , n244, \ScanOut[14]1 , n256, n238, n223, 
        n198, n204, n233, n228, n261, n246, n214, \ScanOut[28]1 , n221, 
        \ScanOut[3]1 , \ScanOut[30]1 , \ScanOut[29]1 , \ScanOut[2]1 , n254, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, 
        \ScanOut[16]1 , n226, n201, n213, n234, n241, n194, n208, 
        \ScanOut[6]1 , n200, n227, n249, \ScanOut[7]1 , n252, n195, n209, n212, 
        n240, n235, n215, n260, n232, n247, \ScanOut[21]1 , n229, 
        \ScanOut[13]1 , \ScanOut[12]1 , n255, \ScanOut[20]1 , n207, n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U54 ( .A(\ScanOut[25]1 ), .B(n194), .C(n220), .Z(n237) );
    VMW_AO22 U73 ( .A(ScanIn[30]), .B(n230), .C(In[30]), .D(n228), .Z(n225) );
    VMW_AO22 U68 ( .A(ScanIn[6]), .B(n230), .C(In[6]), .D(n228), .Z(n201) );
    VMW_AO22 U96 ( .A(ScanIn[0]), .B(n230), .C(In[0]), .D(n228), .Z(n195) );
    VMW_AO21 U33 ( .A(\ScanOut[4]1 ), .B(n194), .C(n199), .Z(n258) );
    VMW_AO21 U34 ( .A(\ScanOut[5]1 ), .B(n194), .C(n200), .Z(n257) );
    VMW_AO21 U41 ( .A(\ScanOut[12]1 ), .B(n194), .C(n207), .Z(n250) );
    VMW_AO21 U46 ( .A(\ScanOut[17]1 ), .B(n194), .C(n212), .Z(n245) );
    VMW_NOR2 U61 ( .A(Reset), .B(n194), .Z(n227) );
    VMW_AO22 U84 ( .A(ScanIn[20]), .B(n230), .C(In[20]), .D(n228), .Z(n215) );
    VMW_AO22 U66 ( .A(ScanIn[8]), .B(n230), .C(In[8]), .D(n228), .Z(n203) );
    VMW_AO22 U83 ( .A(ScanIn[21]), .B(n230), .C(In[21]), .D(n228), .Z(n216) );
    VMW_AO21 U35 ( .A(\ScanOut[6]1 ), .B(n194), .C(n201), .Z(n256) );
    VMW_AO21 U48 ( .A(\ScanOut[19]1 ), .B(n194), .C(n214), .Z(n243) );
    VMW_AO21 U53 ( .A(\ScanOut[24]1 ), .B(n194), .C(n219), .Z(n238) );
    VMW_AO22 U91 ( .A(ScanIn[14]), .B(n230), .C(In[14]), .D(n228), .Z(n209) );
    VMW_AO22 U74 ( .A(ScanIn[2]), .B(n230), .C(In[2]), .D(n228), .Z(n197) );
    VMW_FD \Out_reg[25]  ( .D(n237), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n246), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_AO21 U29 ( .A(\ScanOut[0]1 ), .B(n194), .C(n195), .Z(n262) );
    VMW_AO21 U40 ( .A(\ScanOut[11]1 ), .B(n194), .C(n206), .Z(n251) );
    VMW_AO22 U82 ( .A(ScanIn[22]), .B(n230), .C(In[22]), .D(n228), .Z(n217) );
    VMW_FD \Out_reg[5]  ( .D(n257), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO21 U47 ( .A(\ScanOut[18]1 ), .B(n194), .C(n213), .Z(n244) );
    VMW_AO21 U49 ( .A(\ScanOut[20]1 ), .B(n194), .C(n215), .Z(n242) );
    VMW_AO21 U52 ( .A(\ScanOut[23]1 ), .B(n194), .C(n218), .Z(n239) );
    VMW_AO22 U67 ( .A(ScanIn[7]), .B(n230), .C(In[7]), .D(n228), .Z(n202) );
    VMW_AO22 U75 ( .A(ScanIn[29]), .B(n230), .C(In[29]), .D(n228), .Z(n224) );
    VMW_FD \Out_reg[12]  ( .D(n250), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(ScanIn[15]), .B(n230), .C(In[15]), .D(n228), .Z(n210) );
    VMW_FD \Out_reg[21]  ( .D(n241), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_FD \Out_reg[31]  ( .D(n231), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n234), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n254), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n261), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO21 U55 ( .A(\ScanOut[26]1 ), .B(n194), .C(n221), .Z(n236) );
    VMW_AO22 U69 ( .A(ScanIn[5]), .B(n230), .C(In[5]), .D(n228), .Z(n200) );
    VMW_FD \Out_reg[19]  ( .D(n243), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(ScanIn[31]), .B(n230), .C(In[31]), .D(n228), .Z(n226) );
    VMW_INV U97 ( .A(n227), .Z(n229) );
    VMW_FD \Out_reg[3]  ( .D(n259), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[23]  ( .D(n239), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n252), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_AO21 U60 ( .A(\ScanOut[31] ), .B(n194), .C(n226), .Z(n231) );
    VMW_FD \Out_reg[7]  ( .D(n255), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO21 U32 ( .A(\ScanOut[3]1 ), .B(n194), .C(n198), .Z(n259) );
    VMW_AO22 U85 ( .A(ScanIn[1]), .B(n230), .C(In[1]), .D(n228), .Z(n196) );
    VMW_FD \Out_reg[27]  ( .D(n235), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n248), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_AO21 U30 ( .A(\ScanOut[1]1 ), .B(n194), .C(n196), .Z(n261) );
    VMW_AO21 U39 ( .A(\ScanOut[10]1 ), .B(n194), .C(n205), .Z(n252) );
    VMW_AO21 U57 ( .A(\ScanOut[28]1 ), .B(n194), .C(n223), .Z(n234) );
    VMW_FD \Out_reg[6]  ( .D(n256), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(ScanIn[4]), .B(n230), .C(In[4]), .D(n228), .Z(n199) );
    VMW_AO22 U79 ( .A(ScanIn[25]), .B(n230), .C(In[25]), .D(n228), .Z(n220) );
    VMW_AO22 U95 ( .A(ScanIn[10]), .B(n230), .C(In[10]), .D(n228), .Z(n205) );
    VMW_FD \Out_reg[26]  ( .D(n236), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n247), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n244), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO21 U31 ( .A(\ScanOut[2]1 ), .B(n194), .C(n197), .Z(n260) );
    VMW_AO21 U36 ( .A(\ScanOut[7]1 ), .B(n194), .C(n202), .Z(n255) );
    VMW_AO21 U37 ( .A(\ScanOut[8]1 ), .B(n194), .C(n203), .Z(n254) );
    VMW_AO21 U42 ( .A(\ScanOut[13]1 ), .B(n194), .C(n208), .Z(n249) );
    VMW_AO21 U45 ( .A(\ScanOut[16]1 ), .B(n194), .C(n211), .Z(n246) );
    VMW_AO22 U87 ( .A(ScanIn[18]), .B(n230), .C(In[18]), .D(n228), .Z(n213) );
    VMW_FD \Out_reg[2]  ( .D(n260), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[11]  ( .D(n251), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_NOR2 U62 ( .A(n229), .B(ScanEnable), .Z(n228) );
    VMW_FD \Out_reg[22]  ( .D(n240), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_AO22 U65 ( .A(ScanIn[9]), .B(n230), .C(In[9]), .D(n228), .Z(n204) );
    VMW_FD \Out_reg[20]  ( .D(n242), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n249), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(ScanIn[24]), .B(n230), .C(In[24]), .D(n228), .Z(n219) );
    VMW_FD \Out_reg[9]  ( .D(n253), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_AO21 U50 ( .A(\ScanOut[21]1 ), .B(n194), .C(n216), .Z(n241) );
    VMW_AO21 U59 ( .A(\ScanOut[30]1 ), .B(n194), .C(n225), .Z(n232) );
    VMW_FD \Out_reg[30]  ( .D(n232), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n262), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n233), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(ScanIn[27]), .B(n230), .C(In[27]), .D(n228), .Z(n222) );
    VMW_AO22 U89 ( .A(ScanIn[16]), .B(n230), .C(In[16]), .D(n228), .Z(n211) );
    VMW_AO22 U92 ( .A(ScanIn[13]), .B(n230), .C(In[13]), .D(n228), .Z(n208) );
    VMW_FD \Out_reg[24]  ( .D(n238), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n245), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n258), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_AO21 U58 ( .A(\ScanOut[29]1 ), .B(n194), .C(n224), .Z(n233) );
    VMW_AO21 U38 ( .A(\ScanOut[9]1 ), .B(n194), .C(n204), .Z(n253) );
    VMW_AO21 U43 ( .A(\ScanOut[14]1 ), .B(n194), .C(n209), .Z(n248) );
    VMW_NOR3 U64 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n194) );
    VMW_AO22 U81 ( .A(ScanIn[23]), .B(n230), .C(In[23]), .D(n228), .Z(n218) );
    VMW_AO21 U51 ( .A(\ScanOut[22]1 ), .B(n194), .C(n217), .Z(n240) );
    VMW_AO22 U76 ( .A(ScanIn[28]), .B(n230), .C(In[28]), .D(n228), .Z(n223) );
    VMW_AO22 U88 ( .A(ScanIn[17]), .B(n230), .C(In[17]), .D(n228), .Z(n212) );
    VMW_AO22 U93 ( .A(ScanIn[12]), .B(n230), .C(In[12]), .D(n228), .Z(n207) );
    VMW_AO21 U44 ( .A(\ScanOut[15]1 ), .B(n194), .C(n210), .Z(n247) );
    VMW_AO21 U56 ( .A(\ScanOut[27]1 ), .B(n194), .C(n222), .Z(n235) );
    VMW_AO22 U94 ( .A(ScanIn[11]), .B(n230), .C(In[11]), .D(n228), .Z(n206) );
    VMW_AO22 U71 ( .A(ScanIn[3]), .B(n230), .C(In[3]), .D(n228), .Z(n198) );
    VMW_AND2 U63 ( .A(ScanEnable), .B(n227), .Z(n230) );
    VMW_AO22 U86 ( .A(ScanIn[19]), .B(n230), .C(In[19]), .D(n228), .Z(n214) );
    VMW_AO22 U78 ( .A(ScanIn[26]), .B(n230), .C(In[26]), .D(n228), .Z(n221) );
endmodule


module BubbleSort_Control_CWIDTH8_IDWIDTH1_WIDTH32_SCAN1_DW01_dec_8_0 ( A, SUM
     );
input  [7:0] A;
output [7:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n11, n10;
    VMW_AO21 U3 ( .A(n5), .B(A[5]), .C(n6), .Z(SUM[5]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n7), .Z(SUM[1]) );
    VMW_OAI21 U6 ( .A(n10), .B(n11), .C(n5), .Z(SUM[4]) );
    VMW_NOR2 U14 ( .A(n5), .B(A[5]), .Z(n6) );
    VMW_INV U7 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO21 U8 ( .A(n9), .B(A[3]), .C(n10), .Z(SUM[3]) );
    VMW_NAND2 U13 ( .A(n10), .B(n11), .Z(n5) );
    VMW_NOR2 U9 ( .A(A[6]), .B(n13), .Z(n12) );
    VMW_NOR2 U12 ( .A(n9), .B(A[3]), .Z(n10) );
    VMW_XOR2 U15 ( .A(A[7]), .B(n12), .Z(SUM[7]) );
    VMW_INV U17 ( .A(A[2]), .Z(n8) );
    VMW_NOR2 U10 ( .A(A[0]), .B(A[1]), .Z(n7) );
    VMW_NAND2 U11 ( .A(n7), .B(n8), .Z(n9) );
    VMW_INV U19 ( .A(n6), .Z(n13) );
    VMW_OAI21 U4 ( .A(n7), .B(n8), .C(n9), .Z(SUM[2]) );
    VMW_INV U18 ( .A(A[4]), .Z(n11) );
    VMW_MUX2I U16 ( .A(n13), .B(n6), .S(A[6]), .Z(SUM[6]) );
endmodule


module BubbleSort_Control_CWIDTH8_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, 
    Addr, DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n317, n330, \count[2] , n362, n345, \count[6] , n339, n357, n322, 
        n325, n350, n319, \count[4] , n342, \count[0] , n359, n356, n337, n318, 
        n351, \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , \count260[3] , n324, 
        \ScanReg[18] , n336, n358, \count260[7] , n343, \ScanReg[22] , 
        \ScanReg[11] , \ScanReg[6] , n363, \ScanReg[20] , \ScanReg[13] , 
        \ScanReg[4] , \count260[5] , n344, n316, \count260[1] , \ScanReg[29] , 
        \ScanReg[30] , n331, n323, \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , 
        \ScanReg[9] , n338, n314, \count260[0] , n333, \ScanReg[16] , 
        \ScanReg[25] , n361, n346, \ScanReg[1] , \ScanReg[8] , \ScanReg[7] , 
        n328, \ScanReg[5] , \count260[4] , \ScanReg[21] , \ScanReg[12] , n354, 
        \ScanReg[28] , \ScanReg[31] , n321, n326, \ScanReg[19] , n348, 
        \count260[6] , n353, \ScanReg[10] , \ScanReg[23] , n341, \ScanReg[14] , 
        \ScanReg[27] , n313, \ScanReg[3] , \count260[2] , n334, \count[1] , 
        n352, n349, n327, n335, n360, n340, \count[5] , \count[7] , n347, n329, 
        n332, n315, \count[3] , n320, n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U73 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_AND2 U113 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_INV U134 ( .A(n313), .Z(Enable) );
    VMW_AND2 U68 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AND2 U96 ( .A(\ScanReg[28] ), .B(n317), .Z(n338) );
    VMW_AND2 U108 ( .A(\ScanReg[19] ), .B(n317), .Z(n323) );
    VMW_BUFIZ U141 ( .A(n329), .E(n328), .Z(\arr[4] ) );
    VMW_BUFIZ U166 ( .A(n354), .E(n328), .Z(\arr[1] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n357), .CP(Clk), .Q(\count[6] ) );
    VMW_AND2 U53 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U61 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U84 ( .A(\ScanReg[8] ), .B(n317), .Z(n355) );
    VMW_BUFIZ U148 ( .A(n336), .E(n328), .Z(\arr[31] ) );
    VMW_BUFIZ U153 ( .A(n341), .E(n328), .Z(\arr[30] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \count_reg[2]  ( .D(n361), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U66 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U101 ( .A(\ScanReg[25] ), .B(n317), .Z(n332) );
    VMW_AND2 U106 ( .A(\ScanReg[23] ), .B(n317), .Z(n325) );
    VMW_OAI21 U121 ( .A(RD), .B(WR), .C(n322), .Z(n321) );
    VMW_AO22 U126 ( .A(\count[3] ), .B(n318), .C(\ScanReg[3] ), .D(n317), .Z(
        n344) );
    VMW_AO22 U83 ( .A(ScanOut[7]), .B(n315), .C(\count260[7] ), .D(n316), .Z(
        n356) );
    VMW_FD \count_reg[0]  ( .D(n363), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U91 ( .A(\ScanReg[24] ), .B(n317), .Z(n345) );
    VMW_AND2 U98 ( .A(\ScanReg[31] ), .B(n317), .Z(n336) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(\count[1] ), .B(n318), .C(\ScanReg[1] ), .D(n317), .Z(
        n354) );
    VMW_BUFIZ U154 ( .A(n342), .E(n328), .Z(\arr[29] ) );
    VMW_FD \count_reg[4]  ( .D(n359), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n334), .E(n328), .Z(\arr[12] ) );
    VMW_BUFIZ U161 ( .A(n349), .E(n328), .Z(\arr[26] ) );
    VMW_AND2 U74 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_AND2 U114 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_XNOR2 U133 ( .A(Addr[0]), .B(ScanId), .Z(n322) );
    VMW_AND2 U99 ( .A(\ScanReg[12] ), .B(n317), .Z(n334) );
    VMW_BUFIZ U155 ( .A(n343), .E(n328), .Z(\arr[20] ) );
    VMW_AND2 U52 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U67 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AO22 U82 ( .A(ScanOut[6]), .B(n315), .C(\count260[6] ), .D(n316), .Z(
        n357) );
    VMW_AO21 U107 ( .A(RD), .B(ScanEnable), .C(n318), .Z(n328) );
    VMW_AND2 U120 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U55 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U69 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U75 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U115 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_INV U132 ( .A(n318), .Z(n317) );
    VMW_AND2 U90 ( .A(\ScanReg[17] ), .B(n317), .Z(n346) );
    VMW_XNOR2 U109 ( .A(Addr[0]), .B(Id), .Z(n318) );
    VMW_AO22 U129 ( .A(\count[0] ), .B(n318), .C(\ScanReg[0] ), .D(n317), .Z(
        n324) );
    VMW_BUFIZ U147 ( .A(n335), .E(n328), .Z(\arr[6] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n348), .E(n328), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U97 ( .A(\ScanReg[21] ), .B(n317), .Z(n337) );
    VMW_BUFIZ U140 ( .A(n327), .E(n328), .Z(\arr[9] ) );
    VMW_BUFIZ U167 ( .A(n355), .E(n328), .Z(\arr[8] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AND2 U112 ( .A(n319), .B(n318), .Z(n315) );
    VMW_INV U135 ( .A(n321), .Z(ScanEnable) );
    BubbleSort_Control_CWIDTH8_IDWIDTH1_WIDTH32_SCAN1_DW01_dec_8_0 sub_202 ( 
        .A({\count[7] , \count[6] , \count[5] , \count[4] , \count[3] , 
        \count[2] , \count[1] , \count[0] }), .SUM({\count260[7] , 
        \count260[6] , \count260[5] , \count260[4] , \count260[3] , 
        \count260[2] , \count260[1] , \count260[0] }) );
    VMW_AND2 U60 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U85 ( .A(\ScanReg[11] ), .B(n317), .Z(n353) );
    VMW_AND2 U100 ( .A(\ScanReg[16] ), .B(n317), .Z(n333) );
    VMW_AO22 U127 ( .A(\count[2] ), .B(n318), .C(\ScanReg[2] ), .D(n317), .Z(
        n339) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n337), .E(n328), .Z(\arr[21] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n340), .E(n328), .Z(\arr[13] ) );
    VMW_NOR5 U51 ( .A(\count[0] ), .B(\count[1] ), .C(\count[6] ), .D(
        \count[3] ), .E(n314), .Z(n313) );
    VMW_AND2 U57 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_BUFIZ U137 ( .A(n324), .E(n328), .Z(\arr[0] ) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U58 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U62 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U70 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AO22 U79 ( .A(ScanOut[3]), .B(n315), .C(\count260[3] ), .D(n316), .Z(
        n360) );
    VMW_AND2 U95 ( .A(\ScanReg[13] ), .B(n317), .Z(n340) );
    VMW_AOI21 U110 ( .A(n320), .B(n313), .C(Reset), .Z(n319) );
    VMW_BUFIZ U159 ( .A(n347), .E(n328), .Z(\arr[7] ) );
    VMW_AND2 U119 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_BUFIZ U142 ( .A(n330), .E(n328), .Z(\arr[27] ) );
    VMW_BUFIZ U165 ( .A(n353), .E(n328), .Z(\arr[11] ) );
    VMW_AND2 U87 ( .A(\ScanReg[18] ), .B(n317), .Z(n351) );
    VMW_BUFIZ U150 ( .A(n338), .E(n328), .Z(\arr[28] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(\count[4] ), .B(n318), .C(\ScanReg[4] ), .D(n317), .Z(
        n329) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U65 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U102 ( .A(\ScanReg[14] ), .B(n317), .Z(n331) );
    VMW_AND2 U105 ( .A(\ScanReg[10] ), .B(n317), .Z(n326) );
    VMW_AO22 U80 ( .A(ScanOut[4]), .B(n315), .C(\count260[4] ), .D(n316), .Z(
        n359) );
    VMW_AO22 U122 ( .A(\count[7] ), .B(n318), .C(\ScanReg[7] ), .D(n317), .Z(
        n347) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_BUFIZ U139 ( .A(n326), .E(n328), .Z(\arr[10] ) );
    VMW_BUFIZ U157 ( .A(n345), .E(n328), .Z(\arr[24] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO22 U77 ( .A(ScanOut[1]), .B(n315), .C(\count260[1] ), .D(n316), .Z(
        n362) );
    VMW_AND2 U89 ( .A(\ScanReg[26] ), .B(n317), .Z(n349) );
    VMW_AND2 U92 ( .A(\ScanReg[20] ), .B(n317), .Z(n343) );
    VMW_BUFIZ U145 ( .A(n333), .E(n328), .Z(\arr[16] ) );
    VMW_BUFIZ U162 ( .A(n350), .E(n328), .Z(\arr[15] ) );
    VMW_AND2 U117 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_OR4 U130 ( .A(\count[4] ), .B(\count[5] ), .C(\count[2] ), .D(
        \count[7] ), .Z(n314) );
    VMW_BUFIZ U138 ( .A(n325), .E(n328), .Z(\arr[23] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n358), .CP(Clk), .Q(\count[5] ) );
    VMW_AND2 U64 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AO22 U81 ( .A(ScanOut[5]), .B(n315), .C(\count260[5] ), .D(n316), .Z(
        n358) );
    VMW_BUFIZ U156 ( .A(n344), .E(n328), .Z(\arr[3] ) );
    VMW_AND2 U104 ( .A(\ScanReg[9] ), .B(n317), .Z(n327) );
    VMW_AO22 U76 ( .A(ScanOut[0]), .B(n315), .C(\count260[0] ), .D(n316), .Z(
        n363) );
    VMW_AND2 U116 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AO22 U123 ( .A(\count[6] ), .B(n318), .C(\ScanReg[6] ), .D(n317), .Z(
        n335) );
    VMW_AND2 U56 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U88 ( .A(\ScanReg[15] ), .B(n317), .Z(n350) );
    VMW_AND2 U93 ( .A(\ScanReg[29] ), .B(n317), .Z(n342) );
    VMW_NAND2 U131 ( .A(n318), .B(WR), .Z(n320) );
    VMW_FD \count_reg[1]  ( .D(n362), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[30] ), .B(n317), .Z(n341) );
    VMW_BUFIZ U143 ( .A(n331), .E(n328), .Z(\arr[14] ) );
    VMW_BUFIZ U144 ( .A(n332), .E(n328), .Z(\arr[25] ) );
    VMW_BUFIZ U163 ( .A(n351), .E(n328), .Z(\arr[18] ) );
    VMW_BUFIZ U158 ( .A(n346), .E(n328), .Z(\arr[17] ) );
    VMW_BUFIZ U164 ( .A(n352), .E(n328), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_FD \count_reg[3]  ( .D(n360), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n323), .E(n328), .Z(\arr[19] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U63 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U71 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_AND2 U111 ( .A(n319), .B(n320), .Z(n316) );
    VMW_AO22 U124 ( .A(\count[5] ), .B(n318), .C(\ScanReg[5] ), .D(n317), .Z(
        n348) );
    VMW_AO22 U78 ( .A(ScanOut[2]), .B(n315), .C(\count260[2] ), .D(n316), .Z(
        n361) );
    VMW_AND2 U86 ( .A(\ScanReg[22] ), .B(n317), .Z(n352) );
    VMW_AND2 U103 ( .A(\ScanReg[27] ), .B(n317), .Z(n330) );
    VMW_AND2 U118 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U151 ( .A(n339), .E(n328), .Z(\arr[2] ) );
    VMW_FD \count_reg[7]  ( .D(n356), .CP(Clk), .Q(\count[7] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wRegInA0[9] , \wAMid11[23] , \wAMid64[13] , \wBIn108[25] , 
        \wRegInB70[9] , \wRegInB30[28] , \wRegInB45[18] , \wRegInB66[30] , 
        \ScanLink213[0] , \wAMid27[26] , \wBIn28[21] , \wAIn29[19] , 
        \wAMid32[12] , \wAMid47[22] , \wRegInB13[19] , \wRegInB30[31] , 
        \wBIn48[25] , \wRegInB66[29] , \wAIn38[9] , \wAMid52[16] , 
        \ScanLink173[5] , \wBIn40[5] , \wAMid71[27] , \wAIn1[3] , \wAIn2[0] , 
        \wBMid9[13] , \wAIn25[6] , \wBMid38[18] , \ScanLink72[19] , 
        \ScanLink51[31] , \ScanLink51[28] , \ScanLink50[8] , \ScanLink24[18] , 
        \wBIn92[3] , \wBIn118[2] , \ScanLink219[19] , \wAMid65[2] , 
        \wAMid66[1] , \wBMid95[18] , \wRegInB120[13] , \wRegInB2[12] , 
        \wRegInA4[17] , \wRegInB103[22] , \ScanLink89[18] , \wRegInB116[16] , 
        \wAMid8[18] , \wBMid9[20] , \wAIn26[5] , \wBIn43[6] , \wAIn84[19] , 
        \wBIn90[15] , \wBIn91[0] , \ScanLink210[3] , \ScanLink0[13] , 
        \wBMid117[14] , \wBIn85[21] , \wBMid102[20] , \wBMid121[11] , 
        \ScanLink170[6] , \wBMid75[9] , \wAIn117[31] , \wAIn117[28] , 
        \wRegInB107[5] , \wRegInA69[7] , \wAMid27[15] , \wBIn28[12] , 
        \wAIn41[2] , \wAIn108[9] , \wAMid52[25] , \wAMid71[14] , 
        \wRegInA80[31] , \ScanLink29[3] , \wBIn0[27] , \wBIn0[9] , 
        \wRegInA0[26] , \wRegInA0[15] , \wAIn3[21] , \wAIn3[12] , \wBMid2[9] , 
        \wAMid3[27] , \wAMid3[14] , \wAIn7[10] , \wAMid11[10] , 
        \wRegInA80[28] , \wBIn24[1] , \wAMid32[21] , \wAMid64[20] , 
        \wBMid68[6] , \wBIn108[16] , \wAIn93[4] , \wRegInA74[8] , \wAIn115[6] , 
        \wBIn27[2] , \wAMid47[11] , \wBIn48[16] , \wBIn85[12] , \wBMid102[13] , 
        \ScanLink117[1] , \wAIn90[7] , \wBMid121[22] , \wRegInB119[9] , 
        \wRegInA58[18] , \wAIn116[5] , \ScanLink114[2] , \wBMid26[13] , 
        \wAIn42[1] , \wBIn90[26] , \ScanLink0[20] , \wBMid117[27] , 
        \wRegInA4[24] , \wRegInB104[6] , \wRegInB116[25] , \ScanLink171[30] , 
        \ScanLink152[18] , \wBMid53[23] , \wBMid70[12] , \wRegInB2[21] , 
        \wRegInB120[20] , \ScanLink127[28] , \wRegInB103[11] , 
        \ScanLink171[29] , \ScanLink127[31] , \ScanLink104[19] , 
        \wRegInB76[7] , \ScanLink212[26] , \ScanLink84[0] , \ScanLink19[22] , 
        \ScanLink244[27] , \wRegInA6[7] , \ScanLink231[17] , \ScanLink194[10] , 
        \ScanLink251[13] , \wBMid33[27] , \wBMid46[17] , \wRegInA110[18] , 
        \ScanLink224[23] , \ScanLink181[24] , \wAIn109[10] , \ScanLink79[26] , 
        \wAIn7[23] , \wBMid10[16] , \wBMid65[26] , \wBIn103[3] , \wBIn89[2] , 
        \wRegInA16[2] , \ScanLink207[12] , \wAIn14[23] , \wAIn37[12] , 
        \wAIn42[22] , \wRegInB78[22] , \wAMid59[29] , \ScanLink56[6] , 
        \wAIn14[10] , \wBIn15[31] , \wBIn15[28] , \wBMid14[0] , \wBMid17[3] , 
        \wAMid59[30] , \wAIn61[13] , \ScanLink208[1] , \wAIn22[26] , 
        \wAIn23[8] , \wAIn74[27] , \wAMid121[2] , \wAIn57[16] , 
        \wRegInB18[26] , \ScanLink168[4] , \wBIn58[7] , \wAMid81[19] , 
        \wAMid122[1] , \wRegInA26[24] , \wRegInA53[14] , \wRegInA70[25] , 
        \wRegInA46[20] , \wRegInB83[23] , \ScanLink55[5] , \wRegInA10[21] , 
        \wRegInA33[10] , \wRegInB96[17] , \wRegInA65[11] , \wBIn43[30] , 
        \wBIn45[8] , \wBIn100[0] , \wRegInB75[4] , \ScanLink97[13] , 
        \ScanLink9[6] , \ScanLink139[10] , \ScanLink87[3] , \wRegInA15[1] , 
        \ScanLink159[14] , \wBIn60[18] , \wBIn103[29] , \wRegInA5[4] , 
        \ScanLink176[8] , \ScanLink82[27] , \wAIn74[14] , \wBIn36[19] , 
        \wBIn43[29] , \wAIn57[25] , \wBIn103[30] , \wBIn120[18] , 
        \wRegInB18[15] , \ScanLink32[2] , \wAIn22[15] , \wAIn37[21] , 
        \wAIn42[11] , \wAIn88[5] , \wAIn61[20] , \wRegInB78[11] , 
        \wBMid33[14] , \wBMid73[7] , \ScanLink224[10] , \ScanLink181[17] , 
        \wRegInB12[3] , \ScanLink251[20] , \ScanLink79[15] , \wBMid10[25] , 
        \wBMid46[24] , \ScanLink207[21] , \wBMid65[15] , \wAIn109[23] , 
        \wBIn18[5] , \wAMid19[4] , \wBMid26[20] , \wBMid70[21] , 
        \wRegInA72[6] , \ScanLink212[15] , \wAIn113[8] , \wBMid53[10] , 
        \ScanLink231[24] , \ScanLink194[23] , \ScanLink19[11] , \wRegInB11[0] , 
        \ScanLink244[14] , \ScanLink159[27] , \ScanLink82[14] , \wAIn59[0] , 
        \ScanLink97[20] , \wAIn60[9] , \wBMid70[4] , \wAIn96[9] , 
        \ScanLink139[23] , \wAMid105[30] , \wAMid105[29] , \wRegInA33[23] , 
        \wRegInA71[5] , \wRegInB96[24] , \wAMid126[18] , \wRegInA10[12] , 
        \wRegInA46[13] , \ScanLink31[1] , \wRegInB102[8] , \wRegInA65[22] , 
        \wBMid86[4] , \wRegInA26[17] , \wRegInA70[16] , \wRegInA53[27] , 
        \wRegInB83[10] , \wRegInA55[3] , \ScanLink128[26] , \ScanLink86[25] , 
        \wRegInB35[6] , \ScanLink93[11] , \wRegInA42[22] , \ScanLink148[22] , 
        \wBMid118[30] , \wRegInA87[5] , \wBMid54[2] , \wAMid101[18] , 
        \wRegInA37[12] , \wRegInB92[15] , \wBMid118[29] , \wAMid122[30] , 
        \wRegInA61[13] , \wAMid122[29] , \wRegInA14[23] , \wBIn8[1] , 
        \wBIn11[19] , \wRegInA22[26] , \wRegInB28[9] , \wRegInA74[27] , 
        \wRegInA57[16] , \wRegInB87[21] , \ScanLink15[7] , \wAIn26[24] , 
        \wBIn32[31] , \wBMid57[1] , \wAIn70[25] , \wBMid98[8] , \wBIn124[30] , 
        \wBIn107[18] , \wBIn64[29] , \wRegInB69[14] , \wRegInA84[6] , 
        \wBIn32[28] , \wBIn124[29] , \ScanLink128[6] , \wAIn10[21] , 
        \wAIn33[10] , \wBIn47[18] , \wAIn53[14] , \wBIn64[30] , \wAIn46[20] , 
        \ScanLink16[4] , \wAIn65[11] , \ScanLink248[3] , \wAMid7[16] , 
        \wBMid37[25] , \wBMid42[15] , \ScanLink255[11] , \wBMid85[7] , 
        \ScanLink220[21] , \ScanLink185[26] , \wRegInA99[9] , \wBMid14[14] , 
        \wBMid61[24] , \wRegInA56[0] , \ScanLink203[10] , \ScanLink135[9] , 
        \wAIn19[2] , \wBMid22[11] , \wBMid57[21] , \wBMid74[10] , 
        \wAIn118[26] , \ScanLink216[24] , \wRegInB36[5] , \ScanLink240[25] , 
        \ScanLink68[10] , \wBMid30[6] , \wAMid44[9] , \ScanLink235[15] , 
        \ScanLink190[12] , \wAMid85[28] , \wRegInA74[14] , \wAMid59[6] , 
        \wAMid85[31] , \wAMid106[7] , \wRegInA22[15] , \wRegInB87[12] , 
        \wRegInA14[10] , \wRegInA37[21] , \wRegInA57[25] , \wRegInB92[26] , 
        \ScanLink180[8] , \wRegInA42[11] , \ScanLink71[3] , \wRegInA61[20] , 
        \wRegInB83[4] , \wRegInB119[18] , \ScanLink93[22] , \wBMid22[22] , 
        \wBMid74[23] , \wBIn124[6] , \wRegInA31[7] , \wBIn127[5] , 
        \wRegInA32[4] , \wRegInB51[2] , \wRegInA113[8] , \ScanLink148[11] , 
        \ScanLink128[15] , \ScanLink86[16] , \ScanLink216[17] , \wAIn118[15] , 
        \ScanLink68[23] , \wBMid37[16] , \wBMid57[12] , \ScanLink235[26] , 
        \ScanLink190[21] , \wRegInB52[1] , \ScanLink240[16] , 
        \ScanLink220[12] , \ScanLink185[15] , \wRegInA114[29] , 
        \ScanLink231[8] , \wAMid7[25] , \wBMid14[27] , \wBMid42[26] , 
        \ScanLink255[22] , \ScanLink203[23] , \wBMid61[17] , \wRegInA114[30] , 
        \wAIn10[12] , \wAMid28[28] , \wAIn33[23] , \wAIn46[13] , \wAMid105[4] , 
        \wBMid33[5] , \wAIn65[22] , \wAMid88[3] , \wAIn26[17] , \wAMid28[31] , 
        \wAIn53[27] , \wAIn70[16] , \wRegInB80[7] , \wRegInB69[27] , 
        \ScanLink72[0] , \wBIn81[23] , \wBIn94[17] , \wBMid106[22] , 
        \wBMid113[16] , \wBMid125[13] , \wRegInA29[19] , \wRegInB33[8] , 
        \ScanLink130[4] , \ScanLink250[1] , \ScanLink4[11] , \wBMid4[7] , 
        \wAMid26[3] , \wAIn66[7] , \wBMid116[1] , \wRegInB112[14] , 
        \wRegInB6[10] , \wRegInB124[11] , \ScanLink100[31] , \ScanLink123[19] , 
        \wRegInB107[20] , \ScanLink156[29] , \ScanLink100[28] , 
        \ScanLink13[9] , \wBMid7[4] , \wAMid25[0] , \wAIn65[4] , 
        \wRegInB120[0] , \ScanLink175[18] , \ScanLink156[30] , \wAIn113[19] , 
        \wRegInA82[8] , \wBMid115[2] , \wRegInB123[3] , \wAMid15[21] , 
        \wAMid23[24] , \wAMid56[14] , \wBIn59[13] , \ScanLink133[7] , 
        \wAMid60[11] , \wAMid75[25] , \wBMid83[9] , \wBIn119[13] , 
        \wRegInA84[19] , \ScanLink253[2] , \wAMid36[10] , \wAMid43[20] , 
        \wBMid36[8] , \wBIn39[17] , \wAMid42[7] , \wBMid91[29] , \wAMid100[9] , 
        \wRegInB6[23] , \wRegInB124[22] , \ScanLink186[6] , \wRegInB107[13] , 
        \wBMid91[30] , \wAIn2[18] , \wBIn5[4] , \wAMid5[0] , \wBIn67[0] , 
        \wAIn80[31] , \wRegInA108[9] , \wRegInB112[27] , \wBIn122[8] , 
        \wRegInA37[9] , \wRegInB99[19] , \ScanLink154[0] , \wAIn80[28] , 
        \wAMid90[1] , \wBIn81[10] , \wBIn94[24] , \wBMid113[25] , 
        \ScanLink4[22] , \wBMid106[11] , \wRegInB98[5] , \wAMid6[3] , 
        \wAMid15[12] , \wAMid93[2] , \wBMid125[20] , \wRegInA115[6] , 
        \ScanLink234[5] , \wRegInB41[29] , \wAMid23[17] , \wBMid28[4] , 
        \wRegInB17[31] , \wRegInB34[19] , \wAMid36[23] , \wAMid60[22] , 
        \wRegInB41[30] , \wRegInB62[18] , \wBIn39[24] , \wAMid43[13] , 
        \wBIn64[3] , \wRegInB17[28] , \wAIn58[18] , \ScanLink157[3] , 
        \wAMid56[27] , \wBIn59[20] , \wRegInA116[5] , \wAMid75[16] , 
        \ScanLink69[1] , \wBIn119[20] , \ScanLink237[6] , \wBMid7[17] , 
        \wBIn10[20] , \wAIn11[18] , \wAMid41[4] , \wBMid49[19] , \wAMid57[0] , 
        \wRegInB9[0] , \wRegInA29[5] , \ScanLink76[28] , \ScanLink20[30] , 
        \wRegInB49[0] , \wRegInB86[9] , \ScanLink185[5] , \ScanLink20[29] , 
        \ScanLink76[31] , \ScanLink55[19] , \wAIn64[28] , \wBIn70[24] , 
        \wAMid98[9] , \wBIn113[15] , \wAIn17[4] , \wAIn32[30] , \wAIn47[19] , 
        \wBIn53[15] , \wAIn64[31] , \wBIn26[25] , \wAMid29[22] , \wAIn32[29] , 
        \ScanLink193[1] , \wBIn33[11] , \wBIn46[21] , \wBIn125[10] , 
        \wAMid49[26] , \wBIn65[10] , \wBIn106[21] , \wBMid23[31] , 
        \wBMid23[28] , \wBMid56[18] , \wBMid75[30] , \wAMid85[6] , 
        \wRegInA100[17] , \ScanLink69[29] , \wRegInA123[26] , \wBMid75[29] , 
        \wAMid108[1] , \ScanLink69[30] , \wAIn14[7] , \wBIn71[4] , \wBIn72[7] , 
        \wRegInA100[1] , \ScanLink202[29] , \ScanLink141[7] , \wRegInA115[23] , 
        \ScanLink254[31] , \ScanLink221[18] , \ScanLink202[30] , 
        \ScanLink254[28] , \ScanLink221[2] , \ScanLink142[4] , 
        \ScanLink92[31] , \wAMid86[5] , \wRegInB1[8] , \wRegInB41[8] , 
        \wRegInB118[12] , \ScanLink92[28] , \wRegInA103[2] , \ScanLink222[1] , 
        \wAMid54[3] , \wAMid115[15] , \wRegInB86[18] , \ScanLink190[2] , 
        \wAMid84[22] , \wAMid91[16] , \wBMid119[10] , \wAMid123[10] , 
        \wAMid100[21] , \wRegInA89[3] , \ScanLink61[9] , \ScanLink125[3] , 
        \wBIn16[3] , \wAIn127[4] , \wBIn4[25] , \wBIn6[7] , \wBMid7[24] , 
        \wRegInA100[24] , \wRegInA115[10] , \ScanLink245[6] , 
        \ScanLink191[18] , \wBIn10[13] , \wBIn33[22] , \wAIn73[0] , 
        \wRegInA123[15] , \wBIn46[12] , \wBIn125[23] , \wAMid49[15] , 
        \wBIn15[0] , \wBIn26[16] , \wAMid29[11] , \wAMid33[4] , \wBIn65[23] , 
        \wBMid88[2] , \wBIn106[12] , \wBIn70[17] , \wBMid103[6] , 
        \wBIn113[26] , \wAMid30[7] , \wBIn53[26] , \wRegInA43[31] , 
        \wRegInA60[19] , \wBMid44[8] , \wAMid91[25] , \wBMid119[23] , 
        \wBMid100[5] , \wRegInA15[29] , \wBMid59[7] , \wAIn70[3] , 
        \wAMid123[23] , \wRegInA43[28] , \wRegInA58[6] , \wAMid84[11] , 
        \wAMid100[12] , \wRegInA15[30] , \wRegInA36[18] , \wAMid115[26] , 
        \wRegInB38[3] , \wRegInA45[9] , \wAIn124[7] , \ScanLink126[0] , 
        \wAIn9[14] , \wBIn69[6] , \wAIn107[14] , \wRegInB118[21] , 
        \ScanLink246[5] , \ScanLink149[31] , \ScanLink149[28] , 
        \ScanLink18[2] , \wAMid113[0] , \ScanLink21[23] , \ScanLink209[16] , 
        \ScanLink54[13] , \wAIn12[9] , \wAMid14[18] , \wBMid25[1] , 
        \wBMid48[13] , \wAIn124[25] , \wBMid28[17] , \wRegInB96[3] , 
        \ScanLink77[22] , \ScanLink62[16] , \ScanLink17[26] , \wAMid37[30] , 
        \wAMid37[29] , \wAIn112[20] , \ScanLink34[17] , \wRegInA24[0] , 
        \wRegInB63[12] , \ScanLink64[4] , \ScanLink41[27] , \wAMid42[19] , 
        \wAIn59[12] , \wAMid61[31] , \wBIn74[9] , \wRegInB16[22] , 
        \ScanLink188[0] , \ScanLink147[9] , \wRegInB40[23] , \wBMid26[2] , 
        \wAIn39[16] , \wAMid61[28] , \wAMid83[8] , \wRegInB4[5] , 
        \wRegInB35[13] , \wRegInA90[14] , \wRegInB20[27] , \wRegInB44[5] , 
        \wRegInB55[17] , \wRegInA85[20] , \wAIn81[22] , \wRegInB7[6] , 
        \wRegInB76[26] , \ScanLink5[28] , \wAIn94[16] , \wRegInA27[3] , 
        \wRegInA48[24] , \wRegInA28[20] , \wRegInB98[13] , \ScanLink5[31] , 
        \wRegInB7[30] , \wRegInB47[6] , \wRegInB106[19] , \ScanLink174[21] , 
        \wRegInB125[31] , \ScanLink101[11] , \ScanLink157[10] , \wBMid85[17] , 
        \wBMid90[23] , \wAMid110[3] , \wRegInB125[28] , \ScanLink159[5] , 
        \ScanLink122[20] , \wRegInB7[29] , \wRegInA118[3] , \ScanLink142[24] , 
        \ScanLink67[7] , \ScanLink137[14] , \wBIn4[16] , \wAMid8[5] , 
        \wRegInB95[0] , \ScanLink99[17] , \ScanLink161[15] , \wAIn9[27] , 
        \wAMid28[5] , \wBIn118[19] , \ScanLink239[0] , \ScanLink114[25] , 
        \wRegInB20[14] , \wRegInA85[13] , \wBMid28[24] , \wAIn39[25] , 
        \wBIn58[19] , \wAIn68[1] , \wBMid93[3] , \wBMid118[7] , 
        \wRegInB55[24] , \wRegInA40[4] , \wAIn59[21] , \wRegInB16[11] , 
        \wRegInB76[15] , \wRegInB20[1] , \wRegInB35[20] , \wRegInB63[21] , 
        \wRegInA90[27] , \wRegInB40[10] , \ScanLink243[8] , \ScanLink62[25] , 
        \wBMid41[5] , \ScanLink17[15] , \wBMid105[8] , \wAIn107[27] , 
        \wAIn112[13] , \wRegInA92[2] , \ScanLink41[14] , \ScanLink34[24] , 
        \ScanLink209[25] , \ScanLink54[20] , \wAIn124[16] , \ScanLink77[11] , 
        \ScanLink21[10] , \wAMid36[9] , \wBMid48[20] , \wBMid85[24] , 
        \wRegInA91[1] , \ScanLink142[17] , \ScanLink137[27] , \wBMid42[6] , 
        \ScanLink114[16] , \ScanLink99[24] , \wBIn80[30] , \wBMid90[10] , 
        \ScanLink174[12] , \ScanLink161[26] , \ScanLink101[22] , 
        \ScanLink122[13] , \wBMid107[31] , \wAIn122[9] , \wRegInA28[13] , 
        \wRegInA43[7] , \ScanLink157[23] , \wBMid124[19] , \wBMid9[2] , 
        \wBIn80[29] , \wBMid107[28] , \wBMid90[0] , \wAIn94[25] , \wAIn81[11] , 
        \wRegInB23[2] , \wBMid81[15] , \wRegInA48[17] , \wRegInB98[20] , 
        \ScanLink146[26] , \ScanLink27[5] , \ScanLink133[16] , \wBIn0[14] , 
        \wAMid9[12] , \wAIn28[20] , \wBIn29[18] , \wBIn37[8] , \wBMid66[0] , 
        \ScanLink170[23] , \ScanLink165[17] , \ScanLink110[27] , 
        \ScanLink105[13] , \ScanLink88[21] , \wBIn84[18] , \wAIn90[14] , 
        \wBMid94[21] , \ScanLink153[12] , \ScanLink126[22] , \ScanLink119[7] , 
        \wBMid120[28] , \wRegInA59[12] , \wRegInB89[25] , \wRegInB109[3] , 
        \wBMid120[31] , \wAIn85[20] , \wBMid103[19] , \wRegInA39[16] , 
        \wRegInA67[1] , \ScanLink104[8] , \wRegInB24[25] , \wRegInB51[15] , 
        \wRegInA81[22] , \wAIn48[24] , \wRegInB72[24] , \wRegInA64[2] , 
        \ScanLink39[9] , \wRegInB67[10] , \wAIn51[8] , \wBMid59[25] , 
        \wRegInB12[20] , \wRegInB31[11] , \wRegInB44[21] , \wRegInA94[16] , 
        \ScanLink13[24] , \wAIn103[16] , \wAIn116[22] , \wRegInB19[8] , 
        \ScanLink66[14] , \ScanLink30[15] , \ScanLink218[20] , 
        \ScanLink45[25] , \ScanLink24[6] , \ScanLink25[21] , \wBIn29[4] , 
        \wAIn118[3] , \wBMid39[21] , \wBMid65[3] , \wAIn120[27] , 
        \ScanLink50[11] , \wBMid81[26] , \wAIn85[13] , \wRegInB63[0] , 
        \ScanLink73[20] , \ScanLink200[9] , \wAIn90[27] , \wBIn116[4] , 
        \wRegInA39[25] , \ScanLink1[19] , \ScanLink91[7] , \wRegInA59[21] , 
        \wRegInB89[16] , \wBMid94[12] , \wRegInB3[18] , \wRegInB102[31] , 
        \wRegInB102[28] , \ScanLink105[20] , \wRegInB121[19] , 
        \ScanLink170[10] , \ScanLink88[12] , \ScanLink126[11] , 
        \ScanLink153[21] , \ScanLink43[1] , \ScanLink146[15] , 
        \ScanLink133[25] , \ScanLink110[14] , \wBMid3[15] , \wAIn6[30] , 
        \wBMid8[19] , \wAMid9[21] , \wAIn103[25] , \ScanLink165[24] , 
        \ScanLink50[22] , \ScanLink40[2] , \wBMid39[12] , \ScanLink25[12] , 
        \wBMid59[16] , \wAMid75[8] , \wAIn120[14] , \ScanLink73[13] , 
        \ScanLink66[27] , \ScanLink13[17] , \wBIn108[8] , \ScanLink218[13] , 
        \ScanLink45[16] , \wAMid10[30] , \wAIn28[13] , \wAMid46[28] , 
        \wBIn82[9] , \ScanLink30[26] , \wAIn116[11] , \wRegInB12[13] , 
        \wRegInA122[9] , \wRegInB67[23] , \wAMid10[29] , \wAMid33[18] , 
        \wAMid46[31] , \wRegInB31[22] , \wRegInA94[25] , \ScanLink92[4] , 
        \wRegInB60[3] , \wAMid65[19] , \wRegInB44[12] , \wAMid14[1] , 
        \wAIn28[3] , \wAMid68[7] , \wRegInB24[16] , \wRegInA81[11] , 
        \wRegInB51[26] , \wAIn48[17] , \wAIn54[5] , \wAMid95[14] , 
        \wBIn115[7] , \wRegInA11[18] , \wRegInB72[17] , \wRegInB112[2] , 
        \wRegInA32[30] , \wRegInA64[28] , \wAMid104[23] , \wRegInA32[29] , 
        \wRegInA47[19] , \wRegInA64[31] , \wAMid111[17] , \wBIn31[6] , 
        \wAMid80[20] , \wAIn86[3] , \wBMid108[26] , \wBMid124[3] , 
        \wRegInB8[14] , \wRegInB109[24] , \wAIn100[1] , \ScanLink138[29] , 
        \ScanLink102[6] , \ScanLink138[30] , \wAIn6[29] , \wAIn108[29] , 
        \wRegInA111[21] , \wAIn85[0] , \wAIn108[30] , \wRegInA104[15] , 
        \wRegInA127[24] , \ScanLink195[29] , \wAIn103[2] , \ScanLink195[30] , 
        \wBIn14[22] , \wBIn32[5] , \wBIn37[13] , \wBIn42[23] , \wBIn121[12] , 
        \ScanLink101[5] , \wAMid38[14] , \wBIn61[12] , \wBIn102[23] , 
        \ScanLink22[8] , \wRegInB111[1] , \wAMid17[2] , \wBIn74[26] , 
        \wBMid19[5] , \wBIn22[27] , \wAIn57[6] , \wBIn57[17] , \wAMid58[10] , 
        \wBIn117[17] , \wRegInA127[4] , \ScanLink206[7] , \ScanLink97[9] , 
        \ScanLink96[19] , \ScanLink58[0] , \wBIn55[2] , \wRegInB109[17] , 
        \wAMid80[13] , \wAMid111[24] , \wRegInB8[27] , \ScanLink166[2] , 
        \wRegInB82[29] , \wBIn0[0] , \wBIn3[3] , \wBMid3[26] , \wBIn14[11] , 
        \wAIn15[30] , \wAIn15[29] , \wAIn30[1] , \wAMid70[5] , \wBMid108[15] , 
        \wRegInB78[1] , \wRegInB82[30] , \ScanLink4[3] , \wAMid95[27] , 
        \wRegInA8[1] , \wRegInA18[4] , \wBIn87[4] , \wAMid104[10] , 
        \ScanLink7[0] , \wBIn22[14] , \wAIn36[18] , \wAIn43[31] , \wAIn60[19] , 
        \wRegInB79[31] , \wBIn74[15] , \wBIn117[24] , \wAIn33[2] , 
        \wAIn43[28] , \wBIn57[24] , \wAMid58[23] , \wRegInB79[28] , 
        \ScanLink89[5] , \wBIn37[20] , \wAMid38[27] , \wBIn42[10] , 
        \wBIn84[7] , \wBIn121[21] , \wAMid73[6] , \wBMid27[19] , \wBMid52[29] , 
        \wBIn61[21] , \wBIn102[10] , \wRegInA104[26] , \ScanLink18[28] , 
        \wBMid52[30] , \ScanLink205[4] , \wRegInA124[7] , \ScanLink18[31] , 
        \wAMid14[22] , \wAMid37[13] , \wAMid42[23] , \wBIn56[1] , 
        \wBMid71[18] , \wBIn99[8] , \wBIn113[9] , \wRegInA127[17] , 
        \ScanLink225[30] , \ScanLink206[18] , \ScanLink165[1] , \wAIn59[28] , 
        \wRegInB16[18] , \wRegInB35[30] , \wRegInA111[12] , \ScanLink250[19] , 
        \ScanLink225[29] , \wRegInB63[28] , \wBIn38[14] , \wAIn59[31] , 
        \wRegInB20[8] , \wRegInB35[29] , \wAMid61[12] , \wRegInB40[19] , 
        \wRegInB63[31] , \ScanLink243[1] , \wAMid22[27] , \wAMid57[17] , 
        \wBIn58[10] , \wAMid74[26] , \wBIn118[10] , \wAIn68[8] , 
        \ScanLink123[4] , \wBIn10[4] , \wBIn13[7] , \wAMid35[3] , 
        \wBMid48[30] , \wAIn121[3] , \ScanLink54[29] , \ScanLink21[19] , 
        \wBMid48[29] , \ScanLink77[18] , \ScanLink54[30] , \wAMid36[0] , 
        \wAIn75[7] , \wBMid105[1] , \wAIn76[4] , \wBMid90[19] , \wRegInB7[13] , 
        \wRegInB106[23] , \wRegInB125[12] , \wRegInA91[8] , \wRegInA1[16] , 
        \wAIn81[18] , \wBIn95[14] , \wBMid106[2] , \wRegInB113[17] , 
        \wBMid112[15] , \wRegInB98[30] , \ScanLink240[2] , \ScanLink5[12] , 
        \wRegInB98[29] , \wAIn122[0] , \wBMid124[10] , \ScanLink120[7] , 
        \wRegInA0[0] , \wBIn1[24] , \wAIn2[22] , \wAIn2[11] , \wAMid6[15] , 
        \wAIn11[3] , \wBIn80[20] , \wBMid90[9] , \wBMid107[21] , \wAIn112[30] , 
        \wAIn112[29] , \wRegInB59[3] , \wAMid113[9] , \wRegInA39[6] , 
        \wAIn12[0] , \wAMid14[11] , \wAMid22[14] , \wBMid25[8] , \wAMid51[7] , 
        \ScanLink195[6] , \wAMid74[15] , \wBIn118[23] , \wRegInA85[29] , 
        \ScanLink227[5] , \wAMid37[20] , \wAMid57[24] , \wBIn58[23] , 
        \wRegInA106[6] , \wRegInA24[9] , \wRegInA85[30] , \ScanLink79[2] , 
        \wBIn38[27] , \wAMid42[10] , \wBIn74[0] , \ScanLink188[9] , 
        \ScanLink147[0] , \wBMid38[7] , \wAMid83[1] , \wAMid52[4] , 
        \wAMid61[21] , \wBIn77[3] , \wBIn80[13] , \wBMid124[23] , 
        \wRegInA105[5] , \wRegInA28[29] , \wAMid80[2] , \wBMid107[12] , 
        \wRegInA28[30] , \wRegInB88[6] , \ScanLink224[6] , \wBIn95[27] , 
        \wBMid112[26] , \ScanLink144[3] , \ScanLink5[21] , \wRegInA1[25] , 
        \wRegInB95[9] , \wRegInB113[24] , \ScanLink239[9] , \ScanLink174[28] , 
        \wRegInB106[10] , \ScanLink122[30] , \ScanLink101[18] , 
        \ScanLink174[31] , \wBMid23[12] , \wBMid56[22] , \wRegInB7[20] , 
        \wRegInB125[21] , \ScanLink157[19] , \ScanLink196[5] , 
        \ScanLink122[29] , \wRegInB26[6] , \ScanLink241[26] , \ScanLink69[13] , 
        \wBMid75[13] , \ScanLink234[16] , \ScanLink191[11] , \wAIn119[25] , 
        \ScanLink217[27] , \wBMid15[17] , \wBMid60[27] , \wRegInA46[3] , 
        \ScanLink202[13] , \wAMid6[26] , \wBIn10[30] , \wAIn11[22] , 
        \wBMid36[26] , \wBMid43[16] , \ScanLink254[12] , \wBMid95[4] , 
        \wRegInA115[19] , \ScanLink221[22] , \ScanLink184[25] , \wBIn15[9] , 
        \wAIn27[27] , \wAMid29[18] , \wAIn64[12] , \wAIn32[13] , \wAIn47[23] , 
        \wAIn73[9] , \wRegInA94[5] , \wRegInB68[17] , \wBMid44[1] , 
        \wBMid47[2] , \wAIn52[17] , \ScanLink138[5] , \wAIn71[26] , 
        \wAMid84[18] , \wRegInA23[25] , \wRegInA56[15] , \wRegInB86[22] , 
        \wRegInA60[10] , \wRegInA75[24] , \wBMid96[7] , \wRegInA15[20] , 
        \wRegInB25[5] , \wRegInA36[11] , \wRegInA43[21] , \wRegInA97[6] , 
        \wRegInB93[16] , \wRegInB118[31] , \ScanLink149[21] , \ScanLink92[12] , 
        \wRegInB118[28] , \ScanLink87[26] , \wRegInA45[0] , \ScanLink129[25] , 
        \wAIn27[14] , \wBIn33[18] , \wBIn46[28] , \wAIn52[24] , \wBIn106[31] , 
        \ScanLink126[9] , \wBIn125[19] , \wRegInB68[24] , \ScanLink62[3] , 
        \wBIn10[29] , \wBIn46[31] , \wBIn65[19] , \wBIn106[28] , 
        \wRegInB90[4] , \wAIn71[15] , \wAIn11[11] , \wBMid23[6] , \wAMid57[9] , 
        \wAIn64[21] , \wAMid98[0] , \wBMid15[24] , \wAIn32[20] , \wAIn47[10] , 
        \wAMid115[7] , \ScanLink202[20] , \ScanLink193[8] , \wBMid60[14] , 
        \wRegInA100[8] , \wBMid36[15] , \wRegInB42[2] , \ScanLink221[11] , 
        \ScanLink184[16] , \wAMid2[24] , \wAMid2[17] , \wBIn14[18] , 
        \wBMid20[5] , \wBMid23[21] , \wBMid43[25] , \ScanLink254[21] , 
        \ScanLink69[20] , \wAMid49[5] , \wBMid56[11] , \wRegInB2[2] , 
        \ScanLink234[25] , \ScanLink191[22] , \wBMid75[20] , \wAMid108[8] , 
        \wRegInA22[7] , \ScanLink241[15] , \ScanLink217[14] , \wAIn119[16] , 
        \wRegInB1[1] , \wRegInA21[4] , \wRegInB41[1] , \ScanLink222[8] , 
        \ScanLink129[16] , \ScanLink87[15] , \ScanLink149[12] , \wAMid100[31] , 
        \wAMid123[19] , \wRegInA15[13] , \ScanLink92[21] , \wRegInB93[7] , 
        \wAMid100[28] , \wBMid119[19] , \wRegInA60[23] , \wRegInA36[22] , 
        \wRegInB93[25] , \wAMid116[4] , \wRegInA43[12] , \wEnable[0] , 
        \ScanLink61[0] , \wRegInA23[16] , \wRegInB86[11] , \wRegInA56[26] , 
        \wRegInA75[17] , \wAIn23[25] , \wAIn30[8] , \wBIn110[3] , 
        \ScanLink83[24] , \wRegInA8[8] , \wRegInA64[12] , \wRegInB65[7] , 
        \ScanLink158[17] , \ScanLink138[13] , \ScanLink97[0] , \ScanLink58[9] , 
        \ScanLink96[10] , \wRegInA11[22] , \wRegInA47[23] , \wBIn48[4] , 
        \wAMid104[19] , \wRegInA32[13] , \wRegInB97[14] , \wRegInA27[27] , 
        \wRegInA52[17] , \wRegInB82[20] , \wRegInA71[26] , \wRegInB78[8] , 
        \ScanLink45[6] , \wBIn37[29] , \wBIn42[19] , \wBIn121[28] , 
        \wRegInB19[25] , \ScanLink178[7] , \wAIn56[15] , \wBIn61[31] , 
        \wAIn15[20] , \wBIn37[30] , \wBIn61[28] , \wAIn75[24] , \wBIn102[19] , 
        \wBIn121[31] , \wAIn36[11] , \wAIn60[10] , \ScanLink7[9] , 
        \ScanLink218[2] , \wAIn43[21] , \wRegInB79[21] , \wAIn108[13] , 
        \ScanLink46[5] , \wAIn6[13] , \wBMid11[15] , \wBMid64[25] , 
        \wBIn113[0] , \wBIn99[1] , \ScanLink206[11] , \ScanLink165[8] , 
        \wBIn56[8] , \ScanLink250[10] , \wAIn9[2] , \wBMid47[14] , 
        \ScanLink225[20] , \ScanLink180[27] , \wBMid11[26] , \wAMid14[8] , 
        \wBMid27[10] , \wBMid32[24] , \wBMid52[20] , \wRegInB66[4] , 
        \ScanLink78[25] , \ScanLink18[21] , \ScanLink245[24] , \wBMid71[11] , 
        \ScanLink230[14] , \ScanLink195[13] , \wAMid80[30] , \wRegInA27[14] , 
        \wRegInB82[13] , \ScanLink213[25] , \ScanLink94[3] , \wRegInA52[24] , 
        \wBMid27[23] , \wAIn49[3] , \wBMid60[7] , \wAMid80[29] , 
        \wRegInA11[11] , \wRegInA71[15] , \wRegInA32[20] , \wRegInA64[21] , 
        \wRegInA47[10] , \wRegInB97[27] , \ScanLink21[2] , \wAIn100[8] , 
        \wRegInA61[6] , \ScanLink138[20] , \ScanLink158[24] , \ScanLink96[23] , 
        \ScanLink83[17] , \wBMid52[13] , \ScanLink230[27] , \ScanLink195[20] , 
        \ScanLink18[12] , \wBMid71[22] , \wAIn85[9] , \wRegInA62[5] , 
        \ScanLink245[17] , \ScanLink213[16] , \wRegInA111[31] , 
        \ScanLink206[22] , \wBMid64[16] , \wAIn108[20] , \wBMid2[25] , 
        \wBMid2[16] , \wAIn6[20] , \wBMid32[17] , \ScanLink225[13] , 
        \ScanLink180[14] , \wRegInA111[28] , \ScanLink78[16] , 
        \ScanLink250[23] , \wBMid8[23] , \wBMid8[10] , \wAIn15[13] , 
        \wBMid47[27] , \wAIn60[23] , \wAIn23[16] , \wAIn36[22] , \wAIn43[12] , 
        \wAMid58[19] , \wBMid63[4] , \wAIn98[6] , \wAIn56[26] , 
        \wRegInB19[16] , \wRegInB79[12] , \ScanLink22[1] , \wAIn35[5] , 
        \wAIn36[6] , \wBIn53[5] , \wAIn75[17] , \wRegInB111[8] , 
        \wBMid120[12] , \wBIn84[22] , \wBMid103[23] , \wRegInA59[28] , 
        \ScanLink160[5] , \wBIn91[16] , \wRegInA59[31] , \wRegInB63[9] , 
        \ScanLink200[0] , \ScanLink1[10] , \wBMid116[17] , \wRegInA121[3] , 
        \wAMid75[1] , \wAMid76[2] , \wBIn81[3] , \wRegInA5[14] , 
        \wRegInB3[11] , \wRegInB102[21] , \wRegInB117[15] , \wRegInB121[10] , 
        \ScanLink170[19] , \ScanLink153[31] , \ScanLink105[29] , 
        \ScanLink2[4] , \ScanLink126[18] , \ScanLink105[30] , 
        \ScanLink153[28] , \ScanLink43[8] , \wBIn82[0] , \wBIn108[1] , 
        \wAMid9[31] , \wAMid9[28] , \wAIn116[18] , \ScanLink1[7] , 
        \wAMid10[20] , \wAMid26[25] , \wBIn29[22] , \wAMid53[15] , 
        \wAMid70[24] , \wRegInA81[18] , \ScanLink163[6] , \wAMid33[11] , 
        \wAMid46[21] , \wBIn50[6] , \wRegInA122[0] , \wBIn49[26] , 
        \wAMid65[10] , \wBIn109[26] , \ScanLink203[3] , \wAMid10[13] , 
        \wAMid12[6] , \wAIn28[29] , \wBIn37[1] , \wAIn52[2] , \wBMid66[9] , 
        \wBMid122[4] , \wRegInB102[12] , \ScanLink88[28] , \wBMid94[31] , 
        \wAIn80[4] , \wAIn85[30] , \wAIn85[29] , \wBMid94[28] , 
        \wRegInB121[23] , \ScanLink88[31] , \wRegInB3[22] , \wRegInA5[27] , 
        \wRegInB114[5] , \wRegInB117[26] , \wBIn91[25] , \ScanLink1[23] , 
        \wBMid116[24] , \wRegInA67[8] , \wAIn106[6] , \ScanLink104[1] , 
        \wAIn83[7] , \wBIn84[11] , \wBMid103[10] , \wBMid120[21] , 
        \wRegInB44[31] , \wRegInB67[19] , \wAMid33[22] , \wBIn34[2] , 
        \wAIn105[5] , \wRegInB12[29] , \wAMid46[12] , \wBIn49[15] , 
        \wRegInB44[28] , \ScanLink107[2] , \wAMid11[5] , \wAMid26[16] , 
        \wAIn28[30] , \wBIn29[11] , \wAMid65[23] , \wBMid78[5] , 
        \wRegInB12[30] , \wBIn109[15] , \wRegInB31[18] , \wAMid70[17] , 
        \wBMid39[31] , \wAIn51[1] , \wAMid53[26] , \wRegInA79[4] , 
        \ScanLink39[0] , \ScanLink73[30] , \ScanLink50[18] , \ScanLink25[28] , 
        \wBMid39[28] , \wBMid121[7] , \ScanLink25[31] , \ScanLink73[29] , 
        \wRegInB19[1] , \wRegInB117[6] , \ScanLink218[30] , \wAIn14[19] , 
        \wBIn23[24] , \wAIn42[18] , \ScanLink218[29] , \wAIn47[5] , 
        \wBIn56[14] , \wAMid59[13] , \wAIn61[30] , \wAIn37[28] , \wAIn61[29] , 
        \wBIn75[25] , \wRegInB78[18] , \wBIn116[14] , \wBIn15[21] , 
        \wAIn37[31] , \wBIn60[11] , \wBIn103[20] , \wRegInB101[2] , 
        \wBMid26[30] , \wBIn36[10] , \wBIn43[20] , \wBIn120[11] , 
        \wAMid39[17] , \wAIn95[3] , \wRegInA126[27] , \wAIn113[1] , 
        \wAIn7[19] , \wBIn21[5] , \wBIn22[6] , \wBMid70[28] , \wBMid26[29] , 
        \ScanLink111[6] , \wBMid53[19] , \wBMid70[31] , \wRegInA105[16] , 
        \wAIn59[9] , \wRegInA110[22] , \ScanLink224[19] , \ScanLink19[18] , 
        \ScanLink207[31] , \ScanLink251[30] , \ScanLink251[29] , 
        \ScanLink207[28] , \ScanLink97[29] , \wAIn96[0] , \wAIn110[2] , 
        \ScanLink112[5] , \ScanLink97[30] , \wAIn44[6] , \wAMid81[23] , 
        \wRegInB9[17] , \wRegInB11[9] , \wRegInB108[27] , \wBMid109[25] , 
        \wAMid110[14] , \wAMid94[17] , \wAMid105[20] , \wRegInB83[19] , 
        \wAMid126[11] , \wRegInB102[1] , \ScanLink31[8] , \wBIn46[2] , 
        \wAIn109[19] , \wRegInA110[11] , \ScanLink175[2] , \wAIn4[7] , 
        \wBIn15[12] , \wAMid63[5] , \wRegInA105[25] , \wRegInA126[14] , 
        \ScanLink84[9] , \ScanLink215[7] , \ScanLink194[19] , \wBIn103[13] , 
        \wAIn7[4] , \wBMid14[9] , \wAIn20[2] , \wAIn23[1] , \wBIn60[22] , 
        \wBIn23[17] , \wBIn36[23] , \wAMid39[24] , \wBIn43[13] , \wBIn94[4] , 
        \wBIn120[22] , \wBIn56[27] , \wAMid59[20] , \wBIn75[16] , 
        \ScanLink99[6] , \wBIn116[27] , \wRegInA46[29] , \ScanLink208[8] , 
        \wAMid60[6] , \wBIn97[7] , \wAMid122[8] , \wRegInA10[31] , 
        \wRegInA33[19] , \wAMid105[13] , \wRegInA46[30] , \wRegInA65[18] , 
        \wAMid94[24] , \wAMid126[22] , \wRegInA10[28] , \wAMid8[11] , 
        \wBMid38[22] , \wBIn45[1] , \wAMid81[10] , \wBIn100[9] , 
        \wBMid109[16] , \wAMid110[27] , \wRegInB68[2] , \wRegInA15[8] , 
        \wBMid75[0] , \wAIn121[24] , \wRegInB9[24] , \wRegInB108[14] , 
        \ScanLink176[1] , \ScanLink216[4] , \ScanLink139[19] , \ScanLink48[3] , 
        \wAIn102[15] , \ScanLink72[23] , \ScanLink24[22] , \wBMid9[30] , 
        \wBMid9[29] , \wBIn39[7] , \wAIn108[0] , \ScanLink51[12] , 
        \wBMid58[26] , \wAIn117[21] , \ScanLink31[16] , \ScanLink219[23] , 
        \ScanLink44[26] , \ScanLink34[5] , \ScanLink12[27] , \wAMid11[19] , 
        \wAMid32[31] , \wRegInB45[22] , \ScanLink67[17] , \wBIn24[8] , 
        \wAIn29[23] , \wAMid32[28] , \wAMid64[29] , \wRegInB30[12] , 
        \wRegInA95[15] , \wRegInB66[13] , \wRegInA74[1] , \wAIn42[8] , 
        \wAMid47[18] , \wAMid64[30] , \wRegInB13[23] , \ScanLink117[8] , 
        \wAIn49[27] , \wRegInB73[27] , \wAIn84[23] , \wRegInB14[4] , 
        \wRegInB25[26] , \wRegInB50[16] , \wRegInA80[21] , \wRegInA38[15] , 
        \wRegInA77[2] , \ScanLink0[30] , \ScanLink0[29] , \wAIn91[17] , 
        \wRegInB17[7] , \wRegInA58[11] , \wRegInB119[0] , \wRegInB88[26] , 
        \wBMid76[3] , \wBMid95[22] , \wRegInB2[28] , \wRegInB120[29] , 
        \ScanLink152[11] , \ScanLink127[21] , \ScanLink109[4] , \wRegInB2[31] , 
        \wRegInB103[18] , \ScanLink171[20] , \ScanLink104[10] , 
        \ScanLink89[22] , \wRegInB120[30] , \wBIn28[28] , \wAIn38[0] , 
        \wBMid80[16] , \ScanLink164[14] , \ScanLink147[25] , \ScanLink111[24] , 
        \ScanLink37[6] , \ScanLink132[15] , \wAIn49[14] , \wBIn105[4] , 
        \wRegInA10[5] , \wRegInB73[14] , \wBIn1[17] , \wAIn2[9] , \wBIn28[31] , 
        \wAMid78[4] , \wRegInB25[15] , \wRegInA80[12] , \wAIn29[10] , 
        \wRegInB13[10] , \wRegInB30[21] , \wRegInB50[25] , \wRegInB70[0] , 
        \wRegInB45[11] , \wRegInA95[26] , \ScanLink213[9] , \wRegInB66[20] , 
        \wAIn117[12] , \ScanLink219[10] , \ScanLink82[7] , \ScanLink44[15] , 
        \ScanLink31[25] , \ScanLink67[24] , \wAMid8[22] , \wBMid11[4] , 
        \wBMid58[15] , \ScanLink12[14] , \wBMid38[11] , \wAIn102[26] , 
        \wAIn121[17] , \ScanLink72[10] , \ScanLink51[21] , \ScanLink50[1] , 
        \wBMid12[7] , \wAMid66[8] , \ScanLink24[11] , \ScanLink111[17] , 
        \wBIn5[26] , \wBMid80[25] , \ScanLink164[27] , \wAIn84[10] , 
        \wBIn85[31] , \wBIn85[28] , \wBIn91[9] , \wAMid124[6] , 
        \ScanLink147[16] , \ScanLink132[26] , \wBMid95[11] , \ScanLink127[12] , 
        \wRegInA3[3] , \ScanLink171[13] , \ScanLink152[22] , \ScanLink104[23] , 
        \ScanLink53[2] , \ScanLink89[11] , \wAIn91[24] , \wBMid102[29] , 
        \wBIn106[7] , \wRegInA13[6] , \wRegInB88[15] , \wBMid102[30] , 
        \wBMid121[18] , \wRegInA38[26] , \wRegInA58[22] , \wRegInB73[3] , 
        \ScanLink81[4] , \wAMid5[9] , \wBMid36[1] , \wBMid84[14] , 
        \wRegInB85[3] , \ScanLink98[14] , \wRegInA108[0] , \ScanLink229[3] , 
        \ScanLink160[16] , \ScanLink115[26] , \ScanLink143[27] , 
        \ScanLink77[4] , \wBMid91[20] , \wAMid100[0] , \ScanLink156[13] , 
        \ScanLink136[17] , \ScanLink149[6] , \ScanLink123[23] , 
        \ScanLink175[22] , \ScanLink100[12] , \wBIn81[19] , \wAIn95[15] , 
        \wBMid125[30] , \wBMid106[18] , \wRegInB57[5] , \wAIn8[17] , 
        \wBMid29[14] , \wAIn38[15] , \wBIn67[9] , \wBIn122[1] , \wBMid125[29] , 
        \wRegInA29[23] , \wRegInA37[0] , \wRegInA49[27] , \wRegInB99[10] , 
        \ScanLink154[9] , \wAIn80[21] , \wAMid90[8] , \wAIn58[11] , 
        \wBIn59[30] , \wBIn59[29] , \wRegInB77[25] , \wBIn119[30] , 
        \ScanLink69[8] , \wRegInB54[14] , \wRegInB54[6] , \wBIn119[29] , 
        \wRegInA84[23] , \wBIn121[2] , \wRegInB21[24] , \wRegInA34[3] , 
        \wRegInB34[10] , \wRegInB41[20] , \wRegInB62[11] , \wRegInA91[17] , 
        \wRegInB17[21] , \ScanLink198[3] , \wAIn113[23] , \ScanLink35[14] , 
        \wRegInB49[9] , \wRegInB86[0] , \ScanLink74[7] , \ScanLink40[24] , 
        \ScanLink16[25] , \ScanLink63[15] , \wBMid35[2] , \wBMid49[10] , 
        \wAIn125[26] , \wRegInB9[9] , \wBIn79[5] , \wAMid103[3] , 
        \wAIn106[17] , \ScanLink76[21] , \ScanLink20[20] , \ScanLink208[15] , 
        \wAIn80[12] , \wRegInB33[1] , \wRegInA49[14] , \wRegInB99[23] , 
        \ScanLink55[10] , \ScanLink250[8] , \wBMid80[3] , \wAIn95[26] , 
        \ScanLink4[18] , \wBMid91[13] , \wRegInA29[10] , \wRegInA53[4] , 
        \wRegInB107[30] , \wRegInB124[18] , \ScanLink123[10] , \wRegInB6[19] , 
        \ScanLink156[20] , \wAMid0[4] , \wAIn3[28] , \wAMid3[7] , \wBIn5[15] , 
        \wBMid52[5] , \wRegInB107[29] , \ScanLink13[0] , \wRegInB120[9] , 
        \ScanLink100[21] , \ScanLink175[11] , \ScanLink115[15] , \wBMid116[8] , 
        \ScanLink98[27] , \wAIn8[24] , \wBMid84[27] , \ScanLink160[25] , 
        \wAIn125[15] , \wRegInA81[2] , \ScanLink143[14] , \ScanLink136[24] , 
        \ScanLink76[12] , \wAMid15[31] , \wAMid15[28] , \wAMid25[9] , 
        \wBMid29[27] , \wBMid49[23] , \wAIn106[24] , \ScanLink208[26] , 
        \ScanLink55[23] , \ScanLink10[3] , \wAIn113[10] , \wRegInA82[1] , 
        \ScanLink20[13] , \ScanLink40[17] , \ScanLink35[27] , \ScanLink63[26] , 
        \wAMid43[30] , \wBMid51[6] , \ScanLink16[16] , \wRegInB30[2] , 
        \wRegInB34[23] , \wRegInA91[24] , \wAMid60[18] , \wRegInB41[13] , 
        \wAMid43[29] , \wRegInB17[12] , \wAIn58[22] , \wRegInB62[22] , 
        \wAMid36[19] , \wAIn38[26] , \wAIn78[2] , \wRegInA50[7] , \wAMid38[6] , 
        \wRegInB21[17] , \wRegInB77[16] , \wRegInA84[10] , \wAMid44[0] , 
        \wBMid83[0] , \wAMid90[15] , \wAMid101[22] , \wBMid108[4] , 
        \wRegInB54[27] , \wRegInA37[28] , \wBMid118[13] , \wAMid122[13] , 
        \wRegInA14[19] , \wRegInA42[18] , \wRegInA61[30] , \wRegInA37[31] , 
        \wRegInA61[29] , \wAMid85[21] , \wAMid114[16] , \wRegInA113[1] , 
        \ScanLink180[1] , \wBIn61[7] , \wAMid96[6] , \ScanLink232[2] , 
        \wRegInB119[11] , \ScanLink152[7] , \ScanLink148[18] , \wRegInB52[8] , 
        \wRegInA114[20] , \ScanLink231[1] , \wBMid1[3] , \wAIn3[31] , 
        \wRegInA110[2] , \wBMid2[0] , \wBMid6[14] , \wAMid118[2] , 
        \wRegInA122[25] , \ScanLink190[31] , \wBIn11[23] , \wBIn62[4] , 
        \wBIn64[13] , \wAMid95[5] , \wRegInA101[14] , \ScanLink151[4] , 
        \wBIn107[22] , \ScanLink190[28] , \wBIn27[26] , \wAMid28[21] , 
        \wBIn32[12] , \wBIn47[22] , \wBIn124[13] , \wAMid48[25] , 
        \ScanLink72[9] , \wBIn52[16] , \wAMid47[3] , \ScanLink183[2] , 
        \wBMid49[4] , \wBIn71[27] , \wBIn112[16] , \wRegInB119[22] , 
        \ScanLink256[6] , \ScanLink93[18] , \ScanLink136[3] , \wAIn10[31] , 
        \wAMid20[4] , \wAIn60[0] , \wAMid85[12] , \wAMid114[25] , 
        \wRegInB28[0] , \wRegInB87[31] , \wRegInB126[7] , \wRegInA48[5] , 
        \wRegInB87[28] , \wAMid101[11] , \wAMid28[12] , \wAIn33[19] , 
        \wAMid90[26] , \wBMid118[20] , \wBMid110[6] , \wAMid122[20] , 
        \wAIn10[28] , \wBIn27[15] , \wAIn46[29] , \wBIn52[25] , 
        \wRegInB125[4] , \wAMid2[30] , \wBMid3[11] , \wBMid6[27] , \wBIn8[8] , 
        \wBIn11[10] , \wAIn46[30] , \wAIn65[18] , \wBIn71[14] , \wBIn112[25] , 
        \wAMid23[7] , \wBIn32[21] , \wBMid57[8] , \wBIn64[20] , \wBMid98[1] , 
        \wBIn107[11] , \wBMid113[5] , \wAIn63[3] , \wBIn47[11] , \wBIn124[20] , 
        \wAMid48[16] , \wBMid57[31] , \wBMid74[19] , \wBIn14[26] , 
        \wAMid17[6] , \wBIn22[23] , \wBMid22[18] , \wBMid57[28] , 
        \wRegInA122[16] , \wRegInA101[27] , \wAIn57[2] , \wBIn57[13] , 
        \wRegInA56[9] , \wRegInA99[0] , \wRegInA114[13] , \ScanLink255[18] , 
        \ScanLink255[5] , \ScanLink68[19] , \ScanLink220[28] , 
        \ScanLink220[31] , \ScanLink203[19] , \ScanLink135[0] , \wAMid58[14] , 
        \wBIn61[16] , \wBMid63[9] , \wBIn74[22] , \wBIn117[13] , \wBIn102[27] , 
        \wRegInB111[5] , \wBIn37[17] , \wAMid38[10] , \wBIn42[27] , 
        \wBIn121[16] , \wAIn85[4] , \wRegInA127[20] , \wRegInA62[8] , 
        \wBIn32[1] , \wAIn103[6] , \wRegInA104[11] , \ScanLink101[1] , 
        \wRegInA111[25] , \ScanLink180[19] , \wAMid2[29] , \wBMid3[22] , 
        \wBMid11[18] , \wAMid14[5] , \wBIn31[2] , \wAIn86[7] , \wAIn100[5] , 
        \ScanLink102[2] , \wRegInB8[10] , \wRegInB109[20] , \ScanLink158[29] , 
        \ScanLink158[30] , \wBMid32[30] , \wBMid32[29] , \wBMid47[19] , 
        \wAIn54[1] , \wAMid80[24] , \wBMid108[22] , \wAMid111[13] , 
        \wBMid124[7] , \wRegInA52[30] , \wRegInA71[18] , \wBMid64[31] , 
        \wAMid95[10] , \wAMid104[27] , \wRegInA27[19] , \wRegInA52[29] , 
        \wRegInB112[6] , \wBMid64[28] , \wRegInA111[16] , \ScanLink78[28] , 
        \ScanLink165[5] , \wBIn56[5] , \ScanLink78[31] , \wBIn14[15] , 
        \wRegInB66[9] , \wRegInA124[3] , \wRegInA127[13] , \ScanLink245[30] , 
        \ScanLink213[28] , \wRegInA104[22] , \ScanLink245[29] , 
        \ScanLink230[19] , \ScanLink205[0] , \ScanLink213[31] , \wBIn22[10] , 
        \wAIn23[31] , \wAIn23[28] , \wAIn33[6] , \wBIn61[25] , \wAMid73[2] , 
        \wBIn102[14] , \wRegInB19[31] , \wAIn75[29] , \wBIn37[24] , 
        \wAMid38[23] , \wBIn42[14] , \wAIn56[18] , \wBIn84[3] , \wBIn121[25] , 
        \wRegInB19[28] , \wAIn75[30] , \wAIn30[5] , \wBIn57[20] , 
        \wAMid58[27] , \wBIn74[11] , \ScanLink89[1] , \ScanLink46[8] , 
        \ScanLink7[4] , \wBIn117[20] , \wRegInA18[0] , \wBIn48[9] , 
        \wRegInB97[19] , \wAMid70[1] , \wBIn87[0] , \wAMid104[14] , 
        \wAMid80[17] , \wAMid95[23] , \wRegInA8[5] , \wBMid108[11] , 
        \wBIn0[23] , \wAMid9[16] , \wAMid11[8] , \wBMid19[1] , \wBIn55[6] , 
        \wAMid111[20] , \wRegInB78[5] , \ScanLink4[7] , \ScanLink83[30] , 
        \wRegInB8[23] , \ScanLink166[6] , \ScanLink83[29] , \wAIn120[23] , 
        \wRegInB109[13] , \wRegInA127[0] , \ScanLink206[3] , \ScanLink58[4] , 
        \wBMid39[25] , \wBMid65[7] , \ScanLink73[24] , \wAIn103[12] , 
        \wRegInA79[9] , \ScanLink25[25] , \wAIn28[24] , \wBIn29[0] , 
        \wAIn118[7] , \wBMid59[21] , \wAIn116[26] , \ScanLink50[15] , 
        \ScanLink30[11] , \ScanLink218[24] , \ScanLink45[21] , \ScanLink24[2] , 
        \wBMid78[8] , \wRegInB44[25] , \ScanLink66[10] , \ScanLink13[20] , 
        \wBIn109[18] , \wRegInA94[12] , \wRegInB31[15] , \wRegInA64[6] , 
        \wRegInB67[14] , \wAIn48[20] , \wBIn49[18] , \wAIn105[8] , 
        \wRegInB12[24] , \wRegInB72[20] , \wBMid66[4] , \wAIn80[9] , 
        \wRegInB24[21] , \wRegInB51[11] , \wRegInA81[26] , \wAIn85[24] , 
        \wBIn91[31] , \wBMid116[30] , \wRegInA67[5] , \wBIn91[28] , 
        \wBMid116[29] , \wRegInA39[12] , \wAIn90[10] , \wBMid94[25] , 
        \wRegInA59[16] , \wRegInB109[7] , \wRegInB89[21] , \ScanLink153[16] , 
        \ScanLink126[26] , \ScanLink119[3] , \ScanLink170[27] , 
        \ScanLink105[17] , \ScanLink88[25] , \wBMid122[9] , \wBIn0[10] , 
        \wAMid9[25] , \wAMid26[31] , \wAMid26[28] , \wAIn28[7] , \wBMid81[11] , 
        \wRegInB114[8] , \ScanLink165[13] , \ScanLink146[22] , 
        \ScanLink110[23] , \ScanLink27[1] , \ScanLink133[12] , \wAIn48[13] , 
        \wAMid53[18] , \wAMid70[30] , \wBIn115[3] , \wAMid68[3] , 
        \wAMid70[29] , \wRegInB72[13] , \wRegInB24[12] , \wRegInA81[15] , 
        \wAIn28[17] , \wRegInB12[17] , \wRegInB31[26] , \wRegInB51[22] , 
        \wRegInB60[7] , \wRegInA94[21] , \wRegInB44[16] , \wRegInB67[27] , 
        \wAIn35[8] , \ScanLink92[0] , \ScanLink45[12] , \wBMid39[16] , 
        \wBMid59[12] , \wAIn116[15] , \ScanLink218[17] , \ScanLink30[22] , 
        \ScanLink66[23] , \ScanLink73[17] , \ScanLink13[13] , \wAIn103[21] , 
        \wAIn120[10] , \ScanLink50[26] , \ScanLink40[6] , \wRegInA5[19] , 
        \ScanLink25[16] , \wRegInB117[18] , \ScanLink110[10] , \wRegInA0[22] , 
        \wRegInA0[11] , \wBIn4[21] , \wBIn53[8] , \wBMid81[22] , 
        \ScanLink165[20] , \wAIn90[23] , \wBMid94[16] , \ScanLink146[11] , 
        \ScanLink133[21] , \ScanLink126[15] , \ScanLink170[14] , 
        \ScanLink153[25] , \ScanLink105[24] , \ScanLink43[5] , \ScanLink2[9] , 
        \ScanLink88[16] , \wBIn116[0] , \wRegInB89[12] , \wAIn85[17] , 
        \wRegInA39[21] , \wRegInA59[25] , \ScanLink160[8] , \wRegInB63[4] , 
        \ScanLink91[3] , \wBIn4[12] , \wAMid8[1] , \wRegInB95[4] , 
        \ScanLink161[11] , \ScanLink99[13] , \wAIn9[10] , \wAMid22[19] , 
        \wBMid26[6] , \wAMid52[9] , \wBMid85[13] , \wRegInA1[31] , 
        \wRegInA1[28] , \wRegInB113[29] , \ScanLink239[4] , \ScanLink114[21] , 
        \wRegInA118[7] , \ScanLink142[20] , \ScanLink67[3] , \wBMid90[27] , 
        \wAMid110[7] , \wRegInB113[30] , \ScanLink137[10] , \ScanLink157[14] , 
        \ScanLink196[8] , \ScanLink159[1] , \ScanLink122[24] , 
        \ScanLink174[25] , \ScanLink101[15] , \wAIn39[12] , \wAIn81[26] , 
        \wAIn94[12] , \wRegInB7[2] , \wRegInA27[7] , \wRegInA28[24] , 
        \wRegInB47[2] , \wRegInA105[8] , \wRegInA48[20] , \wRegInB98[17] , 
        \wBMid28[13] , \wAMid57[30] , \wAMid57[29] , \wRegInB76[22] , 
        \wRegInB44[1] , \wRegInB55[13] , \ScanLink227[8] , \wAIn59[16] , 
        \wAMid74[18] , \wRegInB4[1] , \wRegInB20[23] , \wRegInB40[27] , 
        \wRegInA85[24] , \wRegInB16[26] , \wRegInA24[4] , \wRegInB35[17] , 
        \wRegInA90[10] , \wRegInB63[16] , \ScanLink188[4] , \wAIn112[24] , 
        \ScanLink34[13] , \wRegInB96[7] , \ScanLink64[0] , \ScanLink41[23] , 
        \ScanLink17[22] , \ScanLink62[12] , \wBMid9[6] , \wBMid25[5] , 
        \wBMid48[17] , \wAIn124[21] , \wBIn69[2] , \wAIn107[10] , 
        \ScanLink77[26] , \wAMid113[4] , \ScanLink21[27] , \ScanLink209[12] , 
        \wRegInA48[13] , \wRegInB98[24] , \ScanLink54[17] , \wBMid42[2] , 
        \wAIn81[15] , \wRegInB23[6] , \wBMid90[14] , \wBMid90[4] , 
        \wAIn94[21] , \wBIn95[19] , \wBMid112[18] , \wRegInA28[17] , 
        \wRegInA43[3] , \ScanLink122[17] , \ScanLink174[16] , 
        \ScanLink157[27] , \ScanLink101[26] , \ScanLink114[12] , 
        \ScanLink99[20] , \wBIn5[0] , \wBIn6[3] , \wBMid7[13] , \wAIn9[23] , 
        \wAIn76[9] , \wBMid85[20] , \ScanLink161[22] , \ScanLink137[23] , 
        \wAIn124[12] , \wRegInA91[5] , \ScanLink142[13] , \ScanLink77[15] , 
        \wBIn10[9] , \wBMid28[20] , \wBMid48[24] , \wAIn107[23] , 
        \ScanLink209[21] , \ScanLink54[24] , \wAIn112[17] , \wRegInA92[6] , 
        \ScanLink21[14] , \ScanLink41[10] , \ScanLink34[20] , \wBIn38[19] , 
        \wBMid41[1] , \ScanLink62[21] , \ScanLink17[11] , \wAIn59[25] , 
        \wRegInB16[15] , \wRegInB20[5] , \wRegInB35[24] , \wRegInA90[23] , 
        \wRegInB40[14] , \wRegInB63[25] , \wAIn39[21] , \wAIn68[5] , 
        \wRegInA40[0] , \ScanLink123[9] , \wRegInB76[11] , \wAIn14[3] , 
        \wBMid20[8] , \wAMid28[1] , \wRegInB20[10] , \wRegInA85[17] , 
        \wAMid54[7] , \wAMid91[12] , \wBMid93[7] , \wAMid100[25] , 
        \wBMid118[3] , \wRegInB55[20] , \wRegInB93[28] , \wAMid123[14] , 
        \wRegInB93[31] , \wBMid119[14] , \wAMid84[26] , \wAMid115[11] , 
        \wAMid116[9] , \wBMid15[30] , \wAMid49[8] , \wAMid86[1] , 
        \wRegInA103[6] , \ScanLink190[6] , \ScanLink222[5] , \ScanLink87[18] , 
        \wRegInB118[16] , \wBIn71[0] , \wRegInA21[9] , \ScanLink142[0] , 
        \wRegInA115[27] , \wBMid15[29] , \wBMid36[18] , \wBMid43[28] , 
        \ScanLink221[6] , \wBMid43[31] , \wRegInA100[5] , \wBMid60[19] , 
        \wAMid108[5] , \wRegInA123[22] , \ScanLink234[31] , \ScanLink217[19] , 
        \wBIn10[24] , \wAIn52[30] , \wBIn65[14] , \wAIn71[18] , \wBIn72[3] , 
        \wAMid85[2] , \wRegInA100[13] , \ScanLink141[3] , \wBIn106[25] , 
        \ScanLink241[18] , \ScanLink234[28] , \wRegInB90[9] , \wRegInB68[30] , 
        \wBIn15[4] , \wAIn17[0] , \wAIn27[19] , \wBIn46[25] , \wAMid49[22] , 
        \wBIn125[14] , \wAIn52[29] , \wRegInB68[29] , \wBIn33[15] , 
        \wBIn53[11] , \wBIn26[21] , \wAMid29[26] , \wAMid57[4] , \wBIn70[20] , 
        \ScanLink193[5] , \wBIn113[11] , \wRegInB25[8] , \wRegInB118[25] , 
        \ScanLink246[1] , \ScanLink18[6] , \wAIn124[3] , \ScanLink129[28] , 
        \ScanLink126[4] , \wAMid6[18] , \wBMid7[20] , \wBIn10[17] , 
        \wBIn26[12] , \wAMid30[3] , \wBMid59[3] , \wAIn70[7] , \wAMid84[15] , 
        \ScanLink129[31] , \wAMid115[22] , \wRegInA23[31] , \wRegInB38[7] , 
        \wRegInA75[29] , \wRegInA56[18] , \wRegInA75[30] , \wRegInA23[28] , 
        \wRegInA58[2] , \wAMid100[16] , \wAMid91[21] , \wBMid100[1] , 
        \wBMid119[27] , \wAMid123[27] , \wAMid29[15] , \wAMid33[0] , 
        \wBIn53[22] , \wBIn70[13] , \wBIn113[22] , \wBIn33[26] , \wBIn65[27] , 
        \wBMid88[6] , \wBIn106[16] , \wAIn73[4] , \wBMid103[2] , 
        \wRegInA94[8] , \wBIn46[16] , \wAMid49[11] , \wBIn125[27] , 
        \ScanLink138[8] , \wBMid95[9] , \wAIn119[31] , \wAIn119[28] , 
        \wRegInA123[11] , \wRegInA100[20] , \ScanLink245[2] , 
        \ScanLink184[28] , \wRegInA89[7] , \wRegInA115[14] , \ScanLink184[31] , 
        \ScanLink125[7] , \wBMid4[3] , \wAIn8[30] , \wAMid15[25] , \wBIn16[7] , 
        \wAMid36[14] , \wBIn39[13] , \wAMid43[24] , \wAIn127[0] , 
        \wRegInA91[30] , \wAMid60[15] , \wRegInA91[29] , \ScanLink253[6] , 
        \wAMid23[20] , \wAMid56[10] , \wAMid75[21] , \wBMid108[9] , 
        \wBIn119[17] , \wBIn59[17] , \ScanLink133[3] , \wAIn8[29] , 
        \wBMid7[0] , \wAIn106[29] , \wRegInB123[7] , \wAMid25[4] , 
        \wAIn106[30] , \wAIn125[18] , \wAIn65[0] , \wBMid115[6] , 
        \wRegInB107[24] , \wAIn66[3] , \wRegInB6[14] , \wRegInB120[4] , 
        \wRegInB124[15] , \ScanLink160[31] , \ScanLink136[29] , 
        \ScanLink143[19] , \wBIn5[18] , \wAMid26[7] , \wRegInB112[10] , 
        \ScanLink136[30] , \ScanLink115[18] , \wAMid5[4] , \wAMid6[7] , 
        \wBMid29[19] , \wBMid52[8] , \wBMid116[5] , \wBIn81[27] , \wBIn94[13] , 
        \wBMid113[12] , \ScanLink250[5] , \ScanLink160[28] , \ScanLink4[15] , 
        \wBMid125[17] , \wRegInA49[19] , \wRegInA53[9] , \ScanLink130[0] , 
        \wBMid106[26] , \wRegInB49[4] , \ScanLink16[28] , \ScanLink63[18] , 
        \wAMid41[0] , \wBIn79[8] , \wRegInA29[1] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink35[19] , \ScanLink16[31] , 
        \ScanLink208[18] , \ScanLink185[1] , \wAMid75[12] , \wRegInB9[4] , 
        \wRegInB54[19] , \wRegInB77[31] , \wBIn119[24] , \ScanLink237[2] , 
        \wRegInB21[29] , \wAMid15[16] , \wAMid23[13] , \wAMid36[27] , 
        \wAIn38[18] , \wBIn39[20] , \wAMid56[23] , \wRegInB77[28] , 
        \wRegInA116[1] , \wBIn59[24] , \wRegInB21[30] , \ScanLink69[5] , 
        \wAMid43[17] , \wBIn64[7] , \ScanLink157[7] , \wBMid28[0] , 
        \wAMid93[6] , \wAMid60[26] , \wBIn81[14] , \wBMid125[24] , 
        \wRegInA115[2] , \wAIn95[18] , \wBMid106[15] , \wRegInB57[8] , 
        \wRegInB98[1] , \wBIn67[4] , \wAMid90[5] , \ScanLink234[1] , 
        \wBIn94[20] , \wBMid113[21] , \ScanLink4[26] , \ScanLink154[4] , 
        \wBMid84[19] , \ScanLink98[19] , \ScanLink77[9] , \wAMid0[9] , 
        \wAIn3[25] , \wAIn3[16] , \wAMid7[12] , \wBMid22[15] , \wAMid42[3] , 
        \wRegInB112[23] , \wBMid57[25] , \wRegInB6[27] , \wRegInB107[17] , 
        \wRegInB124[26] , \ScanLink186[2] , \wRegInB36[1] , \ScanLink240[21] , 
        \wBMid74[14] , \ScanLink255[8] , \ScanLink68[14] , \ScanLink235[11] , 
        \ScanLink190[16] , \wAIn118[22] , \ScanLink216[20] , \wBMid14[10] , 
        \wBMid61[20] , \wRegInA56[4] , \ScanLink203[14] , \ScanLink255[15] , 
        \wAMid7[21] , \wBIn8[5] , \wAIn10[25] , \wBMid37[21] , \wBMid42[11] , 
        \wBMid85[3] , \ScanLink220[25] , \ScanLink185[22] , \wRegInB125[9] , 
        \wAIn26[20] , \wBIn27[18] , \wBIn52[31] , \wBIn71[19] , \wAIn65[15] , 
        \wBIn112[28] , \ScanLink248[7] , \wAIn33[14] , \wAIn46[24] , 
        \wBIn52[28] , \wBIn112[31] , \ScanLink16[0] , \wRegInB69[10] , 
        \wRegInA84[2] , \ScanLink128[2] , \wAIn10[16] , \wBIn18[1] , 
        \wAMid20[9] , \wAIn53[10] , \wBMid57[5] , \wAIn70[21] , \wBMid113[8] , 
        \wAMid114[31] , \wAMid114[28] , \wRegInA57[12] , \wRegInA22[22] , 
        \wRegInA74[23] , \wRegInB87[25] , \ScanLink15[3] , \wBMid54[6] , 
        \wRegInA14[27] , \wRegInA61[17] , \wRegInA42[26] , \wRegInA48[8] , 
        \wRegInA87[1] , \ScanEnable[0] , \wAIn26[13] , \wAMid48[28] , 
        \wBMid49[9] , \wRegInB35[2] , \wRegInA37[16] , \wRegInB92[11] , 
        \ScanLink148[26] , \ScanLink93[15] , \ScanLink86[21] , \wAIn53[23] , 
        \wBMid86[0] , \wRegInA55[7] , \ScanLink128[22] , \wRegInB69[23] , 
        \ScanLink72[4] , \wAMid48[31] , \wAIn70[12] , \wRegInB80[3] , 
        \wAIn65[26] , \wAMid88[7] , \wBMid14[23] , \wAIn33[27] , \wBMid33[1] , 
        \wAIn46[17] , \wAMid105[0] , \ScanLink203[27] , \wBMid61[13] , 
        \wBMid37[12] , \ScanLink220[16] , \ScanLink185[11] , \wRegInB52[5] , 
        \ScanLink255[26] , \wAIn1[7] , \wBMid2[31] , \wAMid3[10] , \wAIn7[9] , 
        \wBMid6[19] , \wBMid22[26] , \wBMid42[22] , \wRegInA101[19] , 
        \wBMid57[16] , \wAMid95[8] , \wRegInA122[31] , \ScanLink235[22] , 
        \ScanLink68[27] , \ScanLink190[25] , \wBIn62[9] , \wBIn127[1] , 
        \wRegInA32[0] , \ScanLink240[12] , \wRegInA122[28] , \ScanLink216[13] , 
        \wBMid74[27] , \wBMid14[4] , \wAIn19[6] , \wAIn118[11] , 
        \ScanLink151[9] , \wRegInB51[6] , \ScanLink128[11] , \ScanLink86[12] , 
        \wBMid30[2] , \wAMid59[2] , \wBIn124[2] , \wRegInA31[3] , 
        \ScanLink148[15] , \wAMid90[18] , \wRegInA14[14] , \ScanLink93[26] , 
        \wRegInA61[24] , \wRegInB83[0] , \wAMid106[3] , \wRegInA37[25] , 
        \wRegInB92[22] , \wRegInA42[15] , \ScanLink71[7] , \wRegInA22[11] , 
        \wRegInA57[21] , \wRegInB87[16] , \wAMid94[29] , \wBIn100[4] , 
        \wRegInA5[0] , \wRegInA74[10] , \wRegInB9[30] , \wRegInB108[19] , 
        \ScanLink82[23] , \wRegInB9[29] , \wRegInA15[5] , \ScanLink159[10] , 
        \wRegInA65[15] , \wRegInB75[0] , \ScanLink139[14] , \ScanLink87[7] , 
        \ScanLink97[17] , \ScanLink216[9] , \ScanLink9[2] , \wRegInA10[25] , 
        \wAIn14[27] , \wBMid17[7] , \wAIn22[22] , \wBIn58[3] , \wAMid94[30] , 
        \wAMid122[5] , \wRegInA46[24] , \wAMid121[6] , \wRegInA26[20] , 
        \wRegInA33[14] , \wRegInB96[13] , \wRegInA53[10] , \wRegInA70[21] , 
        \wRegInB83[27] , \ScanLink55[1] , \wAMid39[30] , \wAMid39[29] , 
        \wAIn57[12] , \wBIn94[9] , \wRegInB18[22] , \ScanLink168[0] , 
        \wAMid63[8] , \wAIn74[23] , \wAIn37[16] , \wAIn61[17] , 
        \ScanLink208[5] , \wAIn42[26] , \wRegInB78[26] , \wBIn103[7] , 
        \wAIn109[14] , \ScanLink56[2] , \wAIn7[14] , \wBMid10[12] , 
        \wBMid65[22] , \wRegInA16[6] , \wBIn89[6] , \ScanLink207[16] , 
        \wRegInA6[3] , \wBMid33[23] , \wBMid46[13] , \ScanLink251[17] , 
        \ScanLink224[27] , \ScanLink181[20] , \ScanLink79[22] , \wBMid2[28] , 
        \wBMid26[17] , \wBMid53[27] , \wRegInB76[3] , \ScanLink19[26] , 
        \ScanLink244[23] , \wRegInA105[28] , \ScanLink231[13] , 
        \ScanLink194[14] , \wAMid3[23] , \wBMid10[21] , \wAMid19[0] , 
        \wBIn21[8] , \wAIn59[4] , \wBMid70[16] , \wBMid70[0] , \wBMid109[31] , 
        \wAMid110[19] , \wRegInA105[31] , \wRegInA126[19] , \ScanLink212[22] , 
        \ScanLink84[4] , \wRegInA26[13] , \wRegInB83[14] , \wBMid109[28] , 
        \wRegInA53[23] , \wRegInA70[12] , \wRegInA10[16] , \wRegInA33[27] , 
        \wRegInA65[26] , \wRegInB96[20] , \wRegInA46[17] , \ScanLink31[5] , 
        \wRegInA71[1] , \ScanLink139[27] , \ScanLink112[8] , \wBMid26[24] , 
        \wRegInB11[4] , \ScanLink97[24] , \ScanLink159[23] , \ScanLink82[10] , 
        \wBMid53[14] , \ScanLink231[20] , \ScanLink194[27] , \wBMid70[25] , 
        \wRegInA72[2] , \ScanLink244[10] , \ScanLink19[15] , \ScanLink212[11] , 
        \ScanLink207[25] , \wBMid65[11] , \wAIn109[27] , \wAIn7[27] , 
        \wBMid33[10] , \wRegInB12[7] , \ScanLink224[14] , \ScanLink181[13] , 
        \ScanLink79[11] , \wAIn14[14] , \wBIn23[30] , \wBMid46[20] , 
        \ScanLink251[24] , \wAIn61[24] , \wBIn75[28] , \wBIn116[19] , 
        \wBMid73[3] , \wAIn22[11] , \wBIn23[29] , \wAIn37[25] , \wAIn42[15] , 
        \wBIn56[19] , \wBIn75[31] , \wAIn47[8] , \wAIn88[1] , \wAIn57[21] , 
        \wRegInB18[11] , \wRegInB78[15] , \ScanLink32[6] , \wAIn26[1] , 
        \wBIn43[2] , \wAIn74[10] , \wAIn91[30] , \wRegInB88[18] , 
        \wBMid80[28] , \wBIn85[25] , \wAIn91[29] , \wBMid121[15] , 
        \ScanLink170[2] , \wBMid102[24] , \wBIn90[11] , \ScanLink210[7] , 
        \wBMid117[10] , \ScanLink81[9] , \ScanLink0[17] , \wAMid66[5] , 
        \wBIn91[4] , \wRegInA4[13] , \wBMid80[31] , \wRegInB116[12] , 
        \wAIn2[4] , \wBMid58[18] , \wAMid65[6] , \wRegInB2[16] , 
        \wRegInB103[26] , \wRegInB120[17] , \ScanLink67[29] , \ScanLink12[19] , 
        \ScanLink31[31] , \wBMid9[17] , \wBMid11[9] , \wAIn25[2] , \wBIn92[7] , 
        \wBIn118[6] , \ScanLink67[30] , \ScanLink44[18] , \wAMid71[23] , 
        \ScanLink31[28] , \wAMid78[9] , \wRegInB25[18] , \wBIn1[30] , 
        \wAMid11[27] , \wAMid27[22] , \wAIn49[19] , \wAMid52[12] , 
        \wRegInB50[28] , \wBIn105[9] , \wRegInA10[8] , \ScanLink173[1] , 
        \wBIn28[25] , \wAMid32[16] , \wBIn40[1] , \wAMid47[26] , \wBIn48[21] , 
        \wRegInB50[31] , \wRegInB73[19] , \wAMid64[17] , \wBIn108[21] , 
        \ScanLink213[4] , \wAIn42[5] , \wRegInB103[15] , \wRegInB2[25] , 
        \wRegInB120[24] , \ScanLink109[9] , \wBIn1[29] , \wRegInB104[2] , 
        \ScanLink147[28] , \ScanLink132[18] , \ScanLink111[30] , \wAMid11[14] , 
        \wBIn24[5] , \wBIn27[6] , \wAIn90[3] , \wBIn90[22] , \wRegInA4[20] , 
        \ScanLink164[19] , \ScanLink147[31] , \wRegInB116[21] , 
        \ScanLink111[29] , \wBMid117[23] , \ScanLink0[24] , \wAIn116[1] , 
        \wRegInA38[18] , \ScanLink114[6] , \wAMid32[25] , \wBIn85[16] , 
        \wBMid102[17] , \wBMid121[26] , \wAIn93[0] , \wAIn115[2] , 
        \wAMid47[15] , \wBIn48[12] , \ScanLink117[5] , \wAMid64[24] , 
        \wBMid68[2] , \wBIn108[12] , \wRegInA95[18] , \wAMid71[10] , 
        \wRegInB14[9] , \wRegInA0[18] , \wAMid0[0] , \wBMid6[10] , 
        \wBMid9[24] , \wAMid27[11] , \wBIn28[16] , \wAIn41[6] , \wAMid52[21] , 
        \wAIn102[18] , \wAIn121[30] , \wRegInA69[3] , \ScanLink29[7] , 
        \wAIn121[29] , \wRegInB107[1] , \wBIn11[27] , \wBIn27[22] , 
        \wBMid33[8] , \wAMid47[7] , \wBIn71[23] , \ScanLink34[8] , 
        \wBIn112[12] , \wBIn52[12] , \wAMid105[9] , \wAMid28[25] , 
        \wBIn32[16] , \wBIn47[26] , \wAMid48[21] , \wBIn124[17] , 
        \ScanLink183[6] , \wBIn64[17] , \wBIn107[26] , \wAMid95[1] , 
        \wRegInA101[10] , \wAMid118[6] , \wBIn127[8] , \wRegInA32[9] , 
        \wRegInA122[21] , \wAMid7[28] , \wBIn62[0] , \wAIn118[18] , 
        \wRegInA110[6] , \ScanLink151[0] , \wRegInA114[24] , \ScanLink185[18] , 
        \ScanLink231[5] , \wBMid1[7] , \wAMid3[3] , \wAMid7[31] , \wBIn61[3] , 
        \ScanLink152[3] , \wAMid96[2] , \wRegInB119[15] , \wBMid6[23] , 
        \wBMid14[19] , \wBMid37[31] , \wAMid44[4] , \wAMid114[12] , 
        \wRegInA113[5] , \ScanLink232[6] , \ScanLink128[18] , \wRegInA22[18] , 
        \wRegInA57[28] , \ScanLink180[5] , \wBMid61[29] , \wAMid85[25] , 
        \wAMid90[11] , \wAMid122[17] , \wRegInA57[31] , \wRegInA74[19] , 
        \wRegInB83[9] , \wAMid101[26] , \wBMid118[17] , \wRegInA99[4] , 
        \ScanLink135[4] , \wBMid37[28] , \wBMid42[18] , \wBMid61[30] , 
        \wRegInB36[8] , \wRegInA114[17] , \wRegInA101[23] , \ScanLink240[28] , 
        \ScanLink255[1] , \ScanLink235[18] , \ScanLink216[30] , \wBIn11[14] , 
        \wAMid23[3] , \wAIn26[29] , \wBIn32[25] , \wAIn63[7] , \wRegInB69[19] , 
        \wRegInA122[12] , \ScanLink240[31] , \ScanLink216[29] , \wBIn47[15] , 
        \wAMid48[12] , \wAIn53[19] , \wBIn124[24] , \wAIn70[31] , \wAIn26[30] , 
        \wBIn64[24] , \wBMid98[5] , \wBIn107[15] , \wAIn70[28] , \wBMid113[1] , 
        \wRegInB125[0] , \wBMid2[4] , \wBIn18[8] , \wAMid20[0] , \wBIn27[11] , 
        \wBIn71[10] , \wBIn112[21] , \wAMid28[16] , \wBIn52[21] , 
        \ScanLink16[9] , \wAIn60[4] , \wAMid90[22] , \wBMid110[2] , 
        \wBMid118[24] , \wAMid122[24] , \wRegInA48[1] , \wRegInA87[8] , 
        \wRegInB92[18] , \wAMid101[15] , \wAMid114[21] , \wBIn5[22] , 
        \wAIn8[13] , \wBMid49[0] , \wAMid85[16] , \wRegInB28[4] , 
        \wRegInB126[3] , \ScanLink86[28] , \wBIn79[1] , \wBMid86[9] , 
        \wAMid103[7] , \wAIn106[13] , \wRegInB119[26] , \ScanLink256[2] , 
        \ScanLink136[7] , \ScanLink86[31] , \wRegInA29[8] , \ScanLink20[24] , 
        \ScanLink208[11] , \ScanLink185[8] , \ScanLink55[14] , \wBMid28[9] , 
        \wBMid29[10] , \wBMid35[6] , \wAMid41[9] , \wBMid49[14] , 
        \wAIn125[22] , \wRegInB86[4] , \ScanLink76[25] , \ScanLink16[21] , 
        \wBIn39[30] , \wBIn39[29] , \wAIn113[27] , \ScanLink63[11] , 
        \ScanLink35[10] , \wBIn121[6] , \wRegInA34[7] , \wRegInB62[15] , 
        \ScanLink74[3] , \ScanLink40[20] , \wAIn58[15] , \wRegInB17[25] , 
        \ScanLink198[7] , \wRegInB41[24] , \wRegInB34[14] , \wRegInA91[13] , 
        \wBMid36[5] , \wAIn38[11] , \wRegInB21[20] , \wRegInB54[10] , 
        \wRegInB54[2] , \wRegInA84[27] , \wAIn80[25] , \wBIn94[29] , 
        \wRegInB77[21] , \wRegInA116[8] , \wBMid113[28] , \wBIn94[30] , 
        \wRegInA49[23] , \wAIn95[11] , \wBMid113[31] , \wBIn122[5] , 
        \wRegInA37[4] , \wRegInA29[27] , \wRegInB99[14] , \wRegInB57[1] , 
        \wRegInB98[8] , \ScanLink234[8] , \ScanLink175[26] , \ScanLink100[16] , 
        \wBMid84[10] , \wBMid91[24] , \wAMid100[4] , \ScanLink156[17] , 
        \ScanLink149[2] , \ScanLink123[27] , \wRegInA108[4] , 
        \ScanLink143[23] , \ScanLink77[0] , \ScanLink136[13] , \wAIn8[20] , 
        \wBMid7[9] , \wAMid23[30] , \wAMid38[2] , \wAMid75[28] , 
        \wRegInB85[7] , \ScanLink160[12] , \ScanLink98[10] , \ScanLink229[7] , 
        \ScanLink115[22] , \wRegInB21[13] , \wRegInA84[14] , \wAMid23[29] , 
        \wAMid56[19] , \wAMid75[31] , \wBMid83[4] , \wBMid108[0] , 
        \wRegInB54[23] , \wAIn78[6] , \wRegInA50[3] , \wBMid29[23] , 
        \wAIn38[22] , \wAIn58[26] , \wRegInB17[16] , \wRegInB77[12] , 
        \wRegInB30[6] , \wRegInB34[27] , \wRegInB62[26] , \wRegInA91[20] , 
        \wRegInB41[17] , \wBMid51[2] , \ScanLink63[22] , \ScanLink16[12] , 
        \wAIn65[9] , \wRegInA82[5] , \wAIn106[20] , \wAIn113[14] , 
        \ScanLink40[13] , \ScanLink35[23] , \ScanLink208[22] , 
        \ScanLink55[27] , \ScanLink20[17] , \ScanLink10[7] , \wAIn125[11] , 
        \ScanLink76[16] , \wBMid49[27] , \wBMid84[23] , \wRegInA81[6] , 
        \ScanLink136[20] , \ScanLink143[10] , \wBIn1[20] , \wBIn5[11] , 
        \wBMid52[1] , \wRegInB112[19] , \ScanLink115[11] , \ScanLink98[23] , 
        \wAIn80[16] , \wBMid80[7] , \wBMid91[17] , \ScanLink175[15] , 
        \ScanLink160[21] , \ScanLink100[25] , \ScanLink123[14] , \wAIn95[22] , 
        \wRegInA29[14] , \wRegInA53[0] , \ScanLink156[24] , \ScanLink13[4] , 
        \ScanLink130[9] , \wRegInB33[5] , \wBMid80[12] , \wRegInA4[30] , 
        \wRegInA49[10] , \wRegInB99[27] , \ScanLink147[21] , \ScanLink37[2] , 
        \wRegInB116[31] , \ScanLink132[11] , \wAMid52[31] , \wBMid76[7] , 
        \wRegInA4[29] , \ScanLink164[10] , \wRegInB116[28] , \ScanLink171[24] , 
        \ScanLink111[20] , \ScanLink104[14] , \ScanLink89[26] , \wAIn84[27] , 
        \wAIn91[13] , \wBMid95[26] , \ScanLink152[15] , \ScanLink127[25] , 
        \ScanLink109[0] , \wRegInB17[3] , \wRegInA58[15] , \wRegInB88[22] , 
        \wRegInB119[4] , \wAIn116[8] , \wRegInA38[11] , \wRegInA77[6] , 
        \wRegInB14[0] , \wRegInB50[12] , \wAMid71[19] , \wBIn0[19] , 
        \wRegInA0[4] , \wBIn1[13] , \wAMid8[15] , \wAMid27[18] , 
        \wRegInB25[22] , \wRegInA80[25] , \wAIn29[27] , \wAIn49[23] , 
        \wAMid52[28] , \wRegInB73[23] , \wAIn93[9] , \wRegInA74[5] , 
        \wRegInB66[17] , \wBMid58[22] , \wRegInB13[27] , \wRegInB30[16] , 
        \wRegInB45[26] , \wRegInA95[11] , \wAIn102[11] , \wAIn117[25] , 
        \wRegInB107[8] , \ScanLink12[23] , \ScanLink67[13] , \ScanLink31[12] , 
        \ScanLink219[27] , \ScanLink44[22] , \ScanLink34[1] , \ScanLink24[26] , 
        \wBMid12[3] , \wAIn26[8] , \wBIn39[3] , \wAIn108[4] , \wBMid38[26] , 
        \wBMid75[4] , \wAIn121[20] , \ScanLink51[16] , \ScanLink72[27] , 
        \wBMid80[21] , \wAIn84[14] , \wRegInB73[7] , \wBIn90[18] , 
        \wBMid117[19] , \wAIn91[20] , \wBIn106[3] , \wRegInA38[22] , 
        \ScanLink81[0] , \wRegInA3[7] , \wRegInA13[2] , \wRegInA58[26] , 
        \wRegInB88[11] , \wBMid95[15] , \ScanLink171[17] , \ScanLink104[27] , 
        \ScanLink127[16] , \ScanLink89[15] , \ScanLink152[26] , 
        \ScanLink53[6] , \wAMid124[2] , \ScanLink147[12] , \ScanLink132[22] , 
        \ScanLink111[13] , \wAMid8[26] , \wAIn102[22] , \ScanLink164[23] , 
        \ScanLink51[25] , \ScanLink50[5] , \wBMid11[0] , \wBMid38[15] , 
        \ScanLink72[14] , \ScanLink24[15] , \wBMid58[11] , \wAIn121[13] , 
        \ScanLink67[20] , \ScanLink12[10] , \wAIn29[14] , \wBIn48[28] , 
        \wBIn108[31] , \wAIn117[16] , \ScanLink219[14] , \ScanLink44[11] , 
        \ScanLink31[21] , \wRegInB13[14] , \wRegInB66[24] , \wBIn48[31] , 
        \wBIn108[28] , \ScanLink82[3] , \wRegInB30[25] , \wRegInB70[4] , 
        \wRegInA95[22] , \wRegInB45[15] , \wBMid2[21] , \wBMid2[12] , 
        \wBMid10[31] , \wBMid10[28] , \wAMid19[9] , \wBIn21[1] , \wAIn38[4] , 
        \wAMid78[0] , \wRegInB25[11] , \wRegInA80[16] , \wRegInB50[21] , 
        \wBIn40[8] , \wAIn49[10] , \wBIn105[0] , \wRegInA10[1] , 
        \wRegInB73[10] , \ScanLink173[8] , \wAIn44[2] , \wAMid94[13] , 
        \wAMid126[15] , \wRegInB96[30] , \wRegInB102[5] , \wAMid105[24] , 
        \wRegInB96[29] , \wBMid70[9] , \wAMid81[27] , \wBMid109[21] , 
        \wAMid110[10] , \wAIn96[4] , \wRegInB9[13] , \wRegInB108[23] , 
        \ScanLink82[19] , \wRegInA71[8] , \wAIn110[6] , \ScanLink112[1] , 
        \wBMid46[30] , \wBMid65[18] , \wBMid33[19] , \wRegInA110[26] , 
        \wBMid46[29] , \ScanLink79[18] , \wAIn95[7] , \wRegInA105[12] , 
        \wRegInA126[23] , \ScanLink244[19] , \ScanLink231[29] , 
        \ScanLink231[30] , \ScanLink212[18] , \wAIn4[3] , \wAIn7[0] , 
        \wBIn15[25] , \wAIn22[18] , \wBIn22[2] , \wAIn113[5] , \wBIn43[24] , 
        \wBIn120[15] , \wRegInB18[18] , \ScanLink111[2] , \wAIn57[28] , 
        \wBIn36[14] , \wAMid39[13] , \wAIn57[31] , \wAIn74[19] , \wBIn103[24] , 
        \wRegInB101[6] , \wBIn60[15] , \wBIn23[20] , \wAIn47[1] , \wBIn56[10] , 
        \wBIn75[21] , \wAIn88[8] , \wBIn116[10] , \wAMid59[17] , \wBIn45[5] , 
        \wRegInA5[9] , \wRegInB75[9] , \ScanLink48[7] , \ScanLink216[0] , 
        \wRegInB108[10] , \ScanLink159[19] , \wAMid60[2] , \wAMid81[14] , 
        \wBMid109[12] , \wAMid110[23] , \wRegInB9[20] , \wRegInA53[19] , 
        \ScanLink176[5] , \wRegInA70[31] , \wRegInA26[29] , \ScanLink55[8] , 
        \wRegInA26[30] , \wRegInB68[6] , \wRegInA70[28] , \wAMid94[20] , 
        \wAMid126[26] , \wBIn15[16] , \wAIn20[6] , \wAIn23[5] , \wBIn23[13] , 
        \wBIn75[12] , \wBIn97[3] , \wAMid105[17] , \wBIn116[23] , \wBIn56[23] , 
        \wAMid59[24] , \ScanLink99[2] , \wBIn36[27] , \wAMid39[20] , 
        \wBIn43[17] , \wBIn94[0] , \wBIn120[26] , \ScanLink168[9] , 
        \wAMid63[1] , \wBIn103[17] , \wBIn60[26] , \wRegInA105[21] , 
        \ScanLink215[3] , \wAMid3[19] , \wRegInA126[10] , \wBMid8[14] , 
        \wAMid10[24] , \wBIn46[6] , \ScanLink181[30] , \ScanLink175[6] , 
        \wAMid65[14] , \wBIn109[22] , \wRegInA110[15] , \ScanLink181[29] , 
        \wRegInA94[28] , \ScanLink203[7] , \wAMid26[21] , \wAMid33[15] , 
        \wAMid46[25] , \wBIn49[22] , \wRegInA94[31] , \wRegInA122[4] , 
        \ScanLink92[9] , \wAMid53[11] , \ScanLink163[2] , \wBIn29[26] , 
        \wAIn35[1] , \wBIn50[2] , \wAMid70[20] , \wAIn103[31] , \ScanLink1[3] , 
        \wAIn103[28] , \wAIn120[19] , \wBIn82[4] , \wBIn108[5] , \wAMid75[5] , 
        \wAMid76[6] , \wRegInB3[15] , \wRegInB121[14] , \wRegInA5[10] , 
        \wRegInB102[25] , \ScanLink2[0] , \wRegInB117[11] , \ScanLink133[31] , 
        \ScanLink110[19] , \wAMid2[13] , \wAIn6[17] , \wBMid8[27] , 
        \wAIn36[2] , \ScanLink165[29] , \ScanLink133[28] , \wBIn53[1] , 
        \wBIn81[7] , \ScanLink165[30] , \wBIn84[26] , \wBIn91[12] , 
        \wRegInA39[31] , \wRegInA39[28] , \ScanLink146[18] , \wRegInA121[7] , 
        \ScanLink200[4] , \wBMid103[27] , \wBMid116[13] , \ScanLink1[14] , 
        \wBIn116[9] , \wBMid120[16] , \ScanLink160[1] , \wAMid10[17] , 
        \wAMid11[1] , \wBMid59[31] , \ScanLink30[18] , \ScanLink13[30] , 
        \wBMid59[28] , \ScanLink45[28] , \ScanLink13[29] , \wRegInB19[5] , 
        \wRegInB117[2] , \ScanLink66[19] , \ScanLink45[31] , \wAMid26[12] , 
        \wBIn29[9] , \wAIn51[5] , \wBMid121[3] , \wRegInA79[0] , \wBIn29[15] , 
        \wAIn48[30] , \wAIn48[29] , \wRegInB72[29] , \wAMid53[22] , 
        \wAMid70[13] , \wRegInB24[31] , \ScanLink39[4] , \wRegInB51[18] , 
        \wRegInB72[30] , \wRegInB24[28] , \wAMid12[2] , \wAMid33[26] , 
        \wAMid65[27] , \wBMid78[1] , \wBIn109[11] , \wAIn83[3] , \wBIn34[6] , 
        \wAIn105[1] , \wBIn37[5] , \wAMid46[16] , \wBIn49[11] , \wAIn80[0] , 
        \wBIn84[15] , \wBMid103[14] , \ScanLink107[6] , \wAIn90[19] , 
        \wBMid120[25] , \wRegInB89[31] , \wRegInB89[28] , \wAIn106[2] , 
        \ScanLink104[5] , \wAIn52[6] , \wBMid81[18] , \wBIn91[21] , 
        \wBMid116[20] , \wRegInA5[23] , \wRegInB114[1] , \ScanLink1[27] , 
        \wRegInB117[22] , \ScanLink27[8] , \wRegInB3[26] , \wRegInB121[27] , 
        \wBMid27[14] , \wBMid52[24] , \wBMid71[15] , \wBMid122[0] , 
        \wRegInB102[16] , \ScanLink213[21] , \ScanLink94[7] , \wRegInB66[0] , 
        \ScanLink18[25] , \ScanLink245[20] , \ScanLink230[10] , 
        \ScanLink195[17] , \ScanLink205[9] , \wAIn9[6] , \wBMid47[10] , 
        \ScanLink250[14] , \ScanLink225[24] , \ScanLink180[23] , \wBMid32[20] , 
        \ScanLink78[21] , \wAIn108[17] , \wBIn113[4] , \wBMid11[11] , 
        \wBMid64[21] , \wBIn99[5] , \ScanLink206[15] , \wAIn15[24] , 
        \wBIn22[19] , \wAIn36[15] , \wAIn43[25] , \wRegInB79[25] , 
        \wBIn57[29] , \ScanLink46[1] , \wBIn117[30] , \ScanLink89[8] , 
        \wAIn23[21] , \wBIn57[30] , \wAIn60[14] , \wBIn74[18] , \wAIn75[20] , 
        \wBIn117[29] , \ScanLink218[6] , \wAIn56[11] , \wRegInB19[21] , 
        \ScanLink178[3] , \wBIn0[31] , \wBIn0[28] , \wBIn0[4] , \wAIn2[26] , 
        \wAIn2[15] , \wAMid2[20] , \wAIn6[24] , \wAIn15[17] , \wBMid19[8] , 
        \wBIn48[0] , \wBMid108[18] , \wAMid111[30] , \wRegInA71[22] , 
        \wAMid111[29] , \wRegInA52[13] , \wRegInA18[9] , \wRegInA27[23] , 
        \wRegInB82[24] , \ScanLink45[2] , \wRegInA47[27] , \wAMid70[8] , 
        \wBIn87[9] , \wRegInA32[17] , \wRegInB97[10] , \wBIn110[7] , 
        \wRegInA11[26] , \wRegInA64[16] , \wRegInB65[3] , \ScanLink96[14] , 
        \wRegInA127[9] , \ScanLink138[17] , \ScanLink97[4] , \ScanLink158[13] , 
        \ScanLink83[20] , \wAIn23[12] , \wAMid38[19] , \wAIn56[22] , 
        \wAIn75[13] , \wRegInB19[12] , \ScanLink22[5] , \wAIn36[26] , 
        \wAIn43[16] , \wAIn98[2] , \wAIn60[27] , \wRegInB79[16] , \wBMid63[0] , 
        \wBMid32[13] , \ScanLink225[17] , \ScanLink180[10] , \ScanLink78[12] , 
        \wBMid11[22] , \wBMid47[23] , \ScanLink250[27] , \ScanLink206[26] , 
        \wBMid64[12] , \wAIn108[24] , \wBMid3[18] , \wBIn32[8] , 
        \wRegInA62[1] , \wRegInA127[29] , \ScanLink213[12] , \wAIn11[26] , 
        \wAIn27[23] , \wBMid27[27] , \wBMid71[26] , \wRegInA104[18] , 
        \ScanLink101[8] , \wRegInA127[30] , \wAMid33[9] , \wBMid44[5] , 
        \wAIn49[7] , \wBMid52[17] , \ScanLink230[23] , \ScanLink195[24] , 
        \wRegInB8[19] , \wRegInB109[30] , \ScanLink245[13] , \ScanLink18[16] , 
        \wRegInB109[29] , \ScanLink158[20] , \ScanLink96[27] , 
        \ScanLink83[13] , \wAIn54[8] , \wBMid60[3] , \wAMid95[19] , 
        \wRegInA11[15] , \wRegInA32[24] , \wRegInA61[2] , \ScanLink138[24] , 
        \wRegInA47[14] , \wRegInB97[23] , \ScanLink21[6] , \wRegInA64[25] , 
        \wRegInA71[11] , \wAMid91[31] , \wBMid96[3] , \wRegInA27[10] , 
        \wRegInB82[17] , \wRegInA45[4] , \wRegInA52[20] , \ScanLink129[21] , 
        \ScanLink87[22] , \wRegInB25[1] , \ScanLink92[16] , \wRegInA43[25] , 
        \ScanLink246[8] , \ScanLink149[25] , \wRegInA97[2] , \wAMid91[28] , 
        \wRegInA36[15] , \wRegInA60[14] , \wRegInB93[12] , \wRegInA15[24] , 
        \wBMid100[8] , \wRegInA23[21] , \wRegInA56[11] , \wRegInA75[20] , 
        \wRegInB86[26] , \wBMid47[6] , \wAIn71[22] , \wRegInB68[13] , 
        \wRegInA94[1] , \wAIn32[17] , \wAMid49[18] , \ScanLink138[1] , 
        \wAIn52[13] , \wAIn47[27] , \wAIn64[16] , \ScanLink254[16] , 
        \wBIn5[9] , \wAMid6[11] , \wBMid36[22] , \wBMid43[12] , \wBMid95[0] , 
        \ScanLink221[26] , \ScanLink184[21] , \wBMid60[23] , \wRegInA46[7] , 
        \wBMid7[30] , \wBMid7[29] , \wBMid15[13] , \wAIn127[9] , 
        \ScanLink202[17] , \wBMid75[17] , \wAIn119[21] , \wRegInA100[30] , 
        \wRegInA123[18] , \ScanLink217[23] , \wBMid20[1] , \wBMid23[16] , 
        \wBMid56[26] , \wRegInB26[2] , \ScanLink241[22] , \wRegInA100[29] , 
        \ScanLink69[17] , \ScanLink234[12] , \ScanLink191[15] , \wBMid23[25] , 
        \wAMid49[1] , \wAMid86[8] , \wAMid115[18] , \wRegInA75[13] , 
        \wAMid116[0] , \wRegInA15[17] , \wRegInA23[12] , \wRegInB86[15] , 
        \wRegInA36[26] , \wRegInA56[22] , \wRegInA43[16] , \wRegInB93[21] , 
        \ScanLink61[4] , \wRegInA60[27] , \wRegInB93[3] , \wRegInB1[5] , 
        \wBIn71[9] , \wRegInA21[0] , \ScanLink92[25] , \ScanLink142[9] , 
        \wBMid75[24] , \wRegInA22[3] , \wRegInB41[5] , \ScanLink149[16] , 
        \ScanLink129[12] , \ScanLink87[11] , \ScanLink217[10] , \wAIn119[12] , 
        \wBMid36[11] , \wBMid56[15] , \wRegInB2[6] , \ScanLink234[21] , 
        \ScanLink191[26] , \ScanLink69[24] , \ScanLink241[11] , 
        \ScanLink221[15] , \ScanLink184[12] , \wRegInB42[6] , 
        \ScanLink254[25] , \wAMid6[22] , \wBMid15[20] , \wBMid43[21] , 
        \ScanLink202[24] , \wBMid60[10] , \wAIn11[15] , \wAIn17[9] , 
        \wAIn47[14] , \wBIn53[18] , \wBIn70[30] , \wBIn26[28] , \wAIn32[24] , 
        \wAMid115[3] , \wAIn64[25] , \wBIn70[29] , \wAMid98[4] , \wBIn113[18] , 
        \wBIn13[3] , \wBMid23[2] , \wBIn26[31] , \wAIn27[10] , \wAIn52[20] , 
        \wAIn71[11] , \wRegInB90[0] , \wRegInB68[20] , \ScanLink62[7] , 
        \wBIn80[24] , \wAIn94[28] , \wBMid107[25] , \wBMid124[14] , 
        \wAIn94[31] , \wAIn122[4] , \ScanLink120[3] , \wBIn3[7] , 
        \wBMid28[30] , \wAMid36[4] , \wBMid85[30] , \wBIn95[10] , 
        \wBMid112[11] , \ScanLink240[6] , \ScanLink5[16] , \wRegInA1[12] , 
        \wAIn75[3] , \wAIn76[0] , \wBMid85[29] , \wBMid106[6] , 
        \wRegInB113[13] , \ScanLink99[29] , \wRegInB7[17] , \wRegInB125[16] , 
        \ScanLink99[30] , \wRegInB106[27] , \ScanLink41[19] , \ScanLink62[31] , 
        \wBMid28[29] , \ScanLink62[28] , \ScanLink34[29] , \wAMid35[7] , 
        \wAIn39[28] , \wBMid41[8] , \wBMid105[5] , \ScanLink34[30] , 
        \ScanLink17[18] , \wAMid57[13] , \ScanLink209[31] , \ScanLink209[28] , 
        \wBIn58[14] , \wRegInA40[9] , \ScanLink123[0] , \wBIn4[31] , 
        \wBIn4[28] , \wBIn10[0] , \wAMid22[23] , \wRegInB55[30] , \wAIn12[4] , 
        \wAMid14[26] , \wAMid28[8] , \wAMid74[22] , \wAIn121[7] , 
        \wRegInB76[18] , \wAIn39[31] , \wBIn118[14] , \wRegInB20[19] , 
        \wAMid61[16] , \wRegInB55[29] , \ScanLink243[5] , \wAMid37[17] , 
        \wBIn38[10] , \wAMid42[27] , \wAMid52[0] , \wRegInB7[24] , 
        \wRegInB125[25] , \ScanLink159[8] , \ScanLink196[1] , \wRegInB106[14] , 
        \wAMid8[8] , \wRegInA1[21] , \ScanLink161[18] , \ScanLink142[30] , 
        \wRegInB113[20] , \ScanLink114[28] , \wAIn9[19] , \wAMid14[15] , 
        \wBIn77[7] , \wRegInA48[29] , \ScanLink142[29] , \ScanLink137[19] , 
        \ScanLink114[31] , \ScanLink144[7] , \wBIn80[17] , \wAMid80[6] , 
        \wBIn95[23] , \wBMid112[22] , \wRegInA48[30] , \ScanLink5[25] , 
        \wAMid83[5] , \wBMid107[16] , \wBMid124[27] , \wRegInB88[2] , 
        \wRegInA105[1] , \ScanLink224[2] , \wAMid22[10] , \wAMid37[24] , 
        \wBIn38[23] , \wBMid38[3] , \wRegInB4[8] , \wAMid61[25] , 
        \wRegInA90[19] , \wAMid42[14] , \wBIn74[4] , \ScanLink147[4] , 
        \wAMid51[3] , \wAMid57[20] , \wRegInA106[2] , \wBIn58[27] , 
        \wAMid74[11] , \wRegInB44[8] , \ScanLink79[6] , \wBIn118[27] , 
        \ScanLink227[1] , \wAIn124[28] , \wBMid8[16] , \wAIn11[7] , 
        \wAIn107[19] , \wAIn124[31] , \wRegInA39[2] , \wAIn36[0] , \wBIn53[3] , 
        \wBIn84[24] , \wRegInB59[7] , \ScanLink195[2] , \ScanLink64[9] , 
        \wAIn90[31] , \wAIn90[28] , \wBMid103[25] , \wBMid120[14] , 
        \wAMid76[4] , \wBMid81[30] , \wBIn91[10] , \wBMid116[11] , 
        \wRegInB89[19] , \ScanLink160[3] , \wRegInA121[5] , \ScanLink91[8] , 
        \ScanLink200[6] , \ScanLink1[16] , \wBIn81[5] , \wRegInA5[12] , 
        \wRegInB117[13] , \wBMid81[29] , \wRegInB3[17] , \wRegInB121[16] , 
        \wRegInB102[27] , \ScanLink30[29] , \ScanLink2[2] , \wAMid10[26] , 
        \wAMid26[23] , \wBIn29[24] , \wAIn35[3] , \wBIn82[6] , 
        \ScanLink66[31] , \ScanLink45[19] , \wBMid59[19] , \wBIn108[7] , 
        \ScanLink30[30] , \wAMid75[7] , \ScanLink66[28] , \ScanLink13[18] , 
        \ScanLink1[1] , \wAIn48[18] , \wBIn50[0] , \wRegInB72[18] , 
        \ScanLink163[0] , \wRegInB51[30] , \wAMid53[13] , \wAMid68[8] , 
        \wAMid70[22] , \wBIn115[8] , \wRegInB51[29] , \wRegInB24[19] , 
        \wAMid12[0] , \wAMid33[17] , \wAMid65[16] , \wBIn109[20] , 
        \ScanLink203[5] , \wAMid46[27] , \wRegInA122[6] , \wBIn49[20] , 
        \wAIn52[4] , \wRegInB3[24] , \wRegInB121[25] , \ScanLink119[8] , 
        \wBMid122[2] , \wRegInB102[14] , \wRegInA5[21] , \wRegInB117[20] , 
        \ScanLink110[28] , \wRegInB114[3] , \ScanLink165[18] , 
        \ScanLink146[30] , \ScanLink133[19] , \ScanLink110[31] , \wBIn0[6] , 
        \wAIn2[24] , \wAIn2[17] , \wAMid2[22] , \wAMid2[11] , \wAIn6[15] , 
        \wAIn9[4] , \wBMid8[25] , \wAMid10[15] , \wBIn37[7] , \wRegInA39[19] , 
        \ScanLink146[29] , \ScanLink104[7] , \wAMid65[25] , \wBMid78[3] , 
        \wAIn80[2] , \wAIn106[0] , \wBIn84[17] , \wBIn91[23] , \wBMid116[22] , 
        \ScanLink1[25] , \wBMid103[16] , \wBMid120[27] , \wBIn109[13] , 
        \wRegInA94[19] , \wAMid11[3] , \wAMid26[10] , \wBIn29[17] , 
        \wAMid33[24] , \wBIn34[4] , \wAMid46[14] , \wAIn105[3] , 
        \ScanLink107[4] , \wBIn49[13] , \wAIn83[1] , \wAMid53[20] , 
        \ScanLink39[6] , \wAMid70[11] , \wAIn120[28] , \wBMid121[1] , 
        \wAIn51[7] , \wAIn103[19] , \wAIn120[31] , \wRegInA79[2] , 
        \ScanLink24[9] , \wAIn15[26] , \wAIn23[23] , \wAMid38[31] , 
        \wBIn48[2] , \wBIn110[5] , \wRegInB8[28] , \wRegInB19[7] , 
        \wRegInB117[0] , \ScanLink158[11] , \wRegInB8[31] , \wRegInB109[18] , 
        \wRegInA32[15] , \wRegInB65[1] , \ScanLink206[8] , \ScanLink83[22] , 
        \ScanLink96[16] , \wRegInB97[12] , \ScanLink138[15] , \ScanLink97[6] , 
        \wAIn75[22] , \wAMid95[31] , \wRegInA47[25] , \wAMid95[28] , 
        \wRegInA11[24] , \wRegInA64[14] , \wRegInA27[21] , \wRegInA71[20] , 
        \ScanLink45[0] , \wRegInA52[11] , \wRegInB82[26] , \wAMid38[28] , 
        \wAIn56[13] , \wAMid73[9] , \wBIn84[8] , \wRegInB19[23] , 
        \ScanLink178[1] , \wAIn36[17] , \wAIn43[27] , \ScanLink46[3] , 
        \wAIn60[16] , \wRegInB79[27] , \ScanLink218[4] , \wBMid32[22] , 
        \ScanLink225[26] , \ScanLink180[21] , \ScanLink250[16] , 
        \ScanLink78[23] , \wBMid11[13] , \wBMid47[12] , \wBIn99[7] , 
        \ScanLink206[17] , \wBMid64[23] , \wAIn108[15] , \wBMid3[30] , 
        \wBMid3[29] , \wBIn113[6] , \wRegInA104[30] , \wRegInA127[18] , 
        \ScanLink213[23] , \ScanLink94[5] , \wBMid27[16] , \wBMid71[17] , 
        \wRegInA104[29] , \wRegInA124[8] , \wBMid52[26] , \wRegInB66[2] , 
        \ScanLink230[12] , \ScanLink195[15] , \ScanLink18[27] , \wAIn6[26] , 
        \wBMid27[25] , \wBIn31[9] , \wBMid60[1] , \wBMid108[29] , 
        \ScanLink245[22] , \wBMid108[30] , \wRegInA71[13] , \wAMid111[18] , 
        \wRegInA52[22] , \wRegInA11[17] , \wRegInA27[12] , \wRegInA32[26] , 
        \wRegInA47[16] , \wRegInB82[15] , \wRegInB97[21] , \ScanLink21[4] , 
        \wRegInA64[27] , \ScanLink102[9] , \ScanLink96[25] , \wAIn49[5] , 
        \wBMid52[15] , \wBMid71[24] , \wRegInA61[0] , \ScanLink138[26] , 
        \ScanLink158[22] , \ScanLink83[11] , \wRegInA62[3] , \ScanLink213[10] , 
        \ScanLink18[14] , \ScanLink245[11] , \ScanLink250[25] , 
        \ScanLink230[21] , \ScanLink195[26] , \wBMid32[11] , \wBMid47[21] , 
        \ScanLink225[15] , \ScanLink180[12] , \wAIn108[26] , \ScanLink78[10] , 
        \wBMid11[20] , \wBMid64[10] , \ScanLink206[24] , \wAIn15[15] , 
        \wBIn22[28] , \wAIn36[24] , \wAIn43[14] , \wAIn98[0] , \wRegInB79[14] , 
        \wAIn57[9] , \wBIn57[18] , \wBIn74[30] , \wBIn22[31] , \wAIn23[10] , 
        \wAIn60[25] , \wBMid63[2] , \wBIn74[29] , \wAIn75[11] , \wBIn117[18] , 
        \wBMid23[14] , \wAIn56[20] , \wRegInB19[10] , \ScanLink22[7] , 
        \wBMid75[15] , \ScanLink217[21] , \wAIn119[23] , \ScanLink69[15] , 
        \wBMid36[20] , \wBMid56[24] , \ScanLink245[9] , \ScanLink234[10] , 
        \ScanLink191[17] , \wBMid95[2] , \wRegInB26[0] , \ScanLink241[20] , 
        \ScanLink221[24] , \ScanLink184[23] , \wBIn6[8] , \wAMid6[13] , 
        \wBMid15[11] , \wBMid43[10] , \ScanLink254[14] , \ScanLink202[15] , 
        \wBMid60[21] , \wRegInA46[5] , \wAIn11[24] , \wBIn26[19] , 
        \wAIn32[15] , \wAIn47[25] , \wBIn53[29] , \wBIn113[30] , \wBIn53[30] , 
        \wAIn64[14] , \wBIn70[18] , \wBIn113[29] , \wAIn27[21] , \wBMid47[4] , 
        \wAIn71[20] , \wBMid103[9] , \wAIn52[11] , \ScanLink138[3] , 
        \wRegInB68[11] , \wRegInA94[3] , \wAMid30[8] , \wBMid44[7] , 
        \wAMid115[30] , \wAMid115[29] , \wRegInA75[22] , \wRegInA23[23] , 
        \wRegInA36[17] , \wRegInA56[13] , \wRegInB86[24] , \wRegInB93[10] , 
        \wRegInA43[27] , \wRegInA58[9] , \wRegInA97[0] , \wRegInA15[26] , 
        \wRegInA60[16] , \wAIn124[8] , \wRegInB25[3] , \ScanLink92[14] , 
        \ScanLink149[27] , \ScanLink129[23] , \wAIn11[17] , \wBMid23[0] , 
        \wAIn27[12] , \wAMid49[30] , \wBMid59[8] , \wRegInA45[6] , 
        \wAIn71[13] , \wBMid96[1] , \wRegInB90[2] , \ScanLink87[20] , 
        \wRegInB68[22] , \wAIn32[26] , \wAMid49[29] , \ScanLink62[5] , 
        \wAIn52[22] , \wAIn47[16] , \wAMid115[1] , \wAIn64[27] , \wAMid98[6] , 
        \wBIn3[5] , \wAMid6[20] , \wBMid36[13] , \wBMid43[23] , 
        \ScanLink254[27] , \wRegInB42[4] , \ScanLink221[17] , 
        \ScanLink184[10] , \wBMid7[18] , \wBMid15[22] , \wBMid60[12] , 
        \ScanLink202[26] , \wBMid75[26] , \wAIn14[8] , \wBMid20[3] , 
        \wBMid23[27] , \wBMid56[17] , \wBIn72[8] , \wAIn119[10] , 
        \wRegInA22[1] , \wRegInA123[29] , \ScanLink141[8] , \ScanLink217[12] , 
        \wRegInA123[30] , \ScanLink241[13] , \ScanLink69[26] , \wAMid49[3] , 
        \wAMid85[9] , \wRegInA100[18] , \wRegInB1[7] , \wRegInB2[4] , 
        \wRegInB41[7] , \ScanLink234[23] , \ScanLink191[24] , 
        \ScanLink129[10] , \ScanLink87[13] , \ScanLink92[27] , \wAMid91[19] , 
        \wRegInA21[2] , \ScanLink149[14] , \wRegInA36[24] , \wRegInA43[14] , 
        \wRegInB93[23] , \ScanLink61[6] , \wRegInA60[25] , \wRegInA15[15] , 
        \wRegInA75[11] , \wRegInB93[1] , \wAMid116[2] , \wRegInA56[20] , 
        \wAMid14[24] , \wRegInA23[10] , \wRegInB86[17] , \wAMid22[21] , 
        \wAMid37[15] , \wAMid61[14] , \wRegInA90[28] , \ScanLink243[7] , 
        \wBIn38[12] , \wAMid42[25] , \wRegInA90[31] , \wBIn4[19] , \wAIn9[31] , 
        \wAIn9[28] , \wBIn10[2] , \wAIn121[5] , \ScanLink123[2] , 
        \wAMid57[11] , \wBIn58[16] , \wAMid74[20] , \wBMid118[8] , 
        \wAIn107[31] , \wBIn118[16] , \wAIn124[19] , \wAIn107[28] , 
        \wAMid35[5] , \wAIn75[1] , \wBMid105[7] , \wBMid42[9] , \wRegInB7[15] , 
        \wRegInB125[14] , \wRegInB106[25] , \wBMid106[4] , \wBIn13[1] , 
        \wAMid36[6] , \ScanLink161[29] , \wAIn76[2] , \wRegInA1[10] , 
        \wRegInB113[11] , \ScanLink114[19] , \ScanLink161[30] , 
        \ScanLink142[18] , \ScanLink137[31] , \ScanLink137[28] , \wBIn80[26] , 
        \wBIn95[12] , \wRegInA48[18] , \ScanLink240[4] , \wBMid107[27] , 
        \wBMid112[13] , \ScanLink5[14] , \wAIn122[6] , \wBMid124[16] , 
        \wRegInA0[30] , \wAMid0[2] , \wAMid3[1] , \wAIn11[5] , \wBMid28[18] , 
        \wRegInA43[8] , \ScanLink120[1] , \ScanLink41[31] , \ScanLink41[28] , 
        \ScanLink34[18] , \ScanLink17[30] , \wAMid51[1] , \wRegInB59[5] , 
        \ScanLink62[19] , \ScanLink17[29] , \wBIn69[9] , \ScanLink209[19] , 
        \ScanLink195[0] , \wRegInA39[0] , \wAIn12[6] , \wAMid14[17] , 
        \wAMid22[12] , \wAIn39[19] , \wAMid57[22] , \wBIn58[25] , 
        \wRegInB20[31] , \ScanLink79[4] , \wBMid38[1] , \wAMid74[13] , 
        \wRegInB76[29] , \wRegInA106[0] , \ScanLink227[3] , \wBIn118[25] , 
        \wRegInB20[28] , \wRegInB55[18] , \wRegInB76[30] , \wAMid61[27] , 
        \wAMid37[26] , \wAMid42[16] , \wBIn74[6] , \wAMid83[7] , 
        \ScanLink147[6] , \wBIn38[21] , \wBIn77[5] , \wBIn80[15] , 
        \wAIn94[19] , \ScanLink224[0] , \wBMid107[14] , \wRegInB47[9] , 
        \wBMid124[25] , \wRegInB88[0] , \wRegInA105[3] , \ScanLink144[5] , 
        \wAMid80[4] , \wBMid85[18] , \wBIn95[21] , \wRegInB7[9] , 
        \wBMid112[20] , \wRegInA1[23] , \ScanLink5[27] , \wRegInB113[22] , 
        \ScanLink99[18] , \ScanLink67[8] , \wRegInB7[26] , \wRegInB125[27] , 
        \ScanLink196[3] , \wBMid30[9] , \wAMid52[2] , \wRegInB106[16] , 
        \wAMid85[27] , \wAMid90[13] , \wBMid118[15] , \wAMid101[24] , 
        \wAMid122[15] , \wRegInB92[30] , \wRegInB92[29] , \wAMid106[8] , 
        \wAMid114[10] , \ScanLink180[7] , \wAMid44[6] , \wBMid14[28] , 
        \wBMid42[30] , \wAMid59[9] , \wBIn61[1] , \wRegInA113[7] , 
        \ScanLink232[4] , \ScanLink86[19] , \ScanLink152[1] , \wAMid96[0] , 
        \wBIn124[9] , \wRegInA31[8] , \wBMid61[18] , \wRegInB119[17] , 
        \wRegInA110[4] , \ScanLink231[7] , \wBMid1[5] , \wBMid2[6] , 
        \wBMid6[12] , \wBMid14[31] , \wBMid37[19] , \wBMid42[29] , \wBIn62[2] , 
        \wAMid95[3] , \wRegInA101[12] , \wRegInA114[26] , \ScanLink240[19] , 
        \ScanLink235[29] , \wBIn11[25] , \wAIn26[18] , \wBIn32[14] , 
        \wAMid118[4] , \wRegInA122[23] , \ScanLink151[2] , \wRegInB69[28] , 
        \ScanLink235[30] , \ScanLink216[18] , \wBIn47[24] , \wAIn53[28] , 
        \wBIn124[15] , \wAMid48[23] , \wRegInB69[31] , \wBIn27[20] , 
        \wAMid28[27] , \wAMid47[5] , \wAIn53[31] , \wBIn107[24] , 
        \wRegInB80[8] , \wBIn64[15] , \wAIn70[19] , \wBIn71[21] , 
        \wBIn112[10] , \ScanLink183[4] , \wBMid49[2] , \wBIn52[10] , 
        \wRegInB35[9] , \wRegInB119[24] , \ScanLink256[0] , \ScanLink128[30] , 
        \wAMid85[14] , \wAMid114[23] , \ScanLink136[5] , \ScanLink128[29] , 
        \wRegInA22[30] , \wRegInA22[29] , \wRegInA57[19] , \wRegInA74[31] , 
        \ScanLink15[8] , \wAMid20[2] , \wBMid110[0] , \wRegInB28[6] , 
        \wRegInA74[28] , \wRegInB126[1] , \wAMid122[26] , \wAIn60[6] , 
        \wAMid90[20] , \wBMid118[26] , \wAMid101[17] , \wRegInA48[3] , 
        \wBIn71[12] , \wBIn112[23] , \wRegInB125[2] , \wBMid6[21] , 
        \wBIn11[16] , \wBIn27[13] , \wAMid28[14] , \wBIn52[23] , \wBIn32[27] , 
        \wBIn47[17] , \wBIn124[26] , \ScanLink128[9] , \wAMid48[10] , 
        \wAIn63[5] , \wRegInA84[9] , \wBIn64[26] , \wBMid98[7] , \wBIn107[17] , 
        \wBMid113[3] , \wAMid23[1] , \wAIn118[30] , \wRegInA101[21] , 
        \ScanLink255[3] , \wRegInA122[10] , \wAMid7[19] , \wAIn118[29] , 
        \wRegInA99[6] , \ScanLink185[30] , \ScanLink135[6] , \wBMid84[12] , 
        \wBMid85[8] , \ScanLink185[29] , \wRegInA114[15] , \ScanLink77[2] , 
        \wRegInA0[29] , \wRegInA108[6] , \wRegInB112[31] , \ScanLink136[11] , 
        \ScanLink143[21] , \wRegInA0[6] , \wBIn1[22] , \wBIn5[20] , 
        \wRegInB112[28] , \ScanLink229[5] , \ScanLink115[20] , 
        \ScanLink98[12] , \wBIn5[13] , \wBMid4[8] , \wAIn8[11] , \wAMid23[18] , 
        \wBMid36[7] , \wRegInB85[5] , \ScanLink160[10] , \ScanLink100[14] , 
        \wAMid42[8] , \ScanLink175[24] , \wAMid56[31] , \wAMid75[19] , 
        \wAIn80[27] , \wBMid91[26] , \ScanLink149[0] , \ScanLink123[25] , 
        \wAIn95[13] , \wAMid100[6] , \ScanLink186[9] , \wRegInA29[25] , 
        \ScanLink156[15] , \wRegInB57[3] , \wRegInA115[9] , \wBIn122[7] , 
        \wRegInA49[21] , \wRegInB99[16] , \wRegInA37[6] , \ScanLink237[9] , 
        \wAMid56[28] , \wRegInB21[22] , \wRegInB54[12] , \wRegInB54[0] , 
        \wRegInA84[25] , \wBMid29[12] , \wAIn38[13] , \wAIn58[17] , 
        \wRegInB17[27] , \wRegInB77[23] , \ScanLink198[5] , \wBIn121[4] , 
        \wRegInA34[5] , \wRegInB34[16] , \wRegInB62[17] , \wRegInA91[11] , 
        \wRegInB41[26] , \ScanLink63[13] , \wBMid35[4] , \wBIn79[3] , 
        \wAIn113[25] , \wRegInB86[6] , \ScanLink74[1] , \ScanLink40[22] , 
        \ScanLink16[23] , \ScanLink35[12] , \wAMid103[5] , \wAIn106[11] , 
        \ScanLink208[13] , \ScanLink55[16] , \ScanLink20[26] , \wAIn125[20] , 
        \ScanLink76[27] , \wBMid49[16] , \wAIn80[14] , \wBIn94[18] , 
        \wBMid113[19] , \wBMid80[5] , \wAIn95[20] , \wRegInA29[16] , 
        \wRegInB33[7] , \wRegInA49[12] , \wRegInA53[2] , \wRegInB99[25] , 
        \ScanLink175[17] , \ScanLink100[27] , \wAIn66[8] , \wBMid84[21] , 
        \wBMid91[15] , \ScanLink156[26] , \ScanLink123[16] , \ScanLink13[6] , 
        \ScanLink143[12] , \wRegInA81[4] , \ScanLink136[22] , \wAIn8[22] , 
        \wBMid52[3] , \wAIn106[22] , \ScanLink160[23] , \ScanLink98[21] , 
        \ScanLink115[13] , \ScanLink10[5] , \ScanLink208[20] , 
        \ScanLink20[15] , \ScanLink55[25] , \wAMid8[17] , \wBMid29[21] , 
        \wBMid49[25] , \wAIn125[13] , \wBMid51[0] , \ScanLink76[14] , 
        \ScanLink16[10] , \ScanLink63[20] , \wAIn38[20] , \wAMid38[0] , 
        \wBIn39[18] , \wAIn113[16] , \ScanLink35[21] , \wRegInB62[24] , 
        \wRegInA82[7] , \ScanLink40[11] , \wAIn58[24] , \wRegInB17[14] , 
        \wBMid83[6] , \wRegInB30[4] , \wRegInB41[15] , \wRegInB34[25] , 
        \wRegInA91[22] , \wBMid108[2] , \wRegInB54[21] , \wRegInB21[11] , 
        \wRegInA84[16] , \wBIn39[1] , \wAIn78[4] , \wRegInB77[10] , 
        \ScanLink133[8] , \wRegInA50[1] , \wAIn102[13] , \wAIn108[6] , 
        \wRegInA69[8] , \ScanLink51[14] , \wAIn29[25] , \wBMid38[24] , 
        \wBMid75[6] , \ScanLink24[24] , \wBIn48[19] , \wBMid58[20] , 
        \wAIn121[22] , \ScanLink72[25] , \ScanLink67[11] , \ScanLink12[21] , 
        \wAIn115[9] , \wAIn117[27] , \ScanLink219[25] , \ScanLink44[20] , 
        \ScanLink34[3] , \ScanLink31[10] , \wRegInB13[25] , \wRegInB66[15] , 
        \wRegInA74[7] , \wAIn49[21] , \wBMid68[9] , \wBIn108[19] , 
        \wRegInA95[13] , \wRegInB30[14] , \wRegInB14[2] , \wRegInB25[20] , 
        \wRegInB45[24] , \wRegInB50[10] , \wRegInA80[27] , \wBMid76[5] , 
        \wAIn84[25] , \wRegInB73[21] , \wAIn90[8] , \wBIn90[30] , \wBIn90[29] , 
        \wBMid117[28] , \wRegInA38[13] , \wBMid117[31] , \wAIn91[11] , 
        \wRegInA58[17] , \wRegInA77[4] , \wRegInB88[20] , \wRegInB17[1] , 
        \wRegInB119[6] , \ScanLink104[16] , \wBMid80[10] , \wBMid95[24] , 
        \ScanLink171[26] , \ScanLink127[27] , \ScanLink89[24] , 
        \ScanLink109[2] , \ScanLink152[17] , \wRegInB104[9] , 
        \ScanLink147[23] , \ScanLink132[13] , \ScanLink37[0] , 
        \ScanLink111[22] , \wAMid27[30] , \ScanLink164[12] , \wAMid71[28] , 
        \wRegInB50[23] , \wAMid78[2] , \wRegInB25[13] , \wRegInA80[14] , 
        \wAMid27[29] , \wAIn38[6] , \wAIn49[12] , \wAMid52[19] , 
        \wRegInB73[12] , \wAMid71[31] , \wBIn105[2] , \wRegInA10[3] , 
        \wRegInA0[20] , \wRegInA0[13] , \wBIn1[11] , \wAMid8[24] , 
        \wBMid11[2] , \wAIn29[16] , \wRegInB66[26] , \ScanLink82[1] , 
        \wBMid58[13] , \wRegInB13[16] , \wRegInB30[27] , \wRegInB45[17] , 
        \wRegInB70[6] , \wRegInA95[20] , \ScanLink12[12] , \wAIn25[9] , 
        \wAIn117[14] , \ScanLink67[22] , \ScanLink31[23] , \wAIn102[20] , 
        \ScanLink219[16] , \ScanLink44[13] , \ScanLink50[7] , \ScanLink24[17] , 
        \wBMid38[17] , \wAIn121[11] , \ScanLink51[27] , \wBMid80[23] , 
        \ScanLink147[10] , \ScanLink72[16] , \wAMid124[0] , \ScanLink132[20] , 
        \wBMid2[23] , \wBMid2[10] , \wBMid12[1] , \wBIn15[27] , \wBIn23[22] , 
        \wBIn43[9] , \wBMid95[17] , \wRegInA4[18] , \ScanLink164[21] , 
        \wRegInB116[19] , \ScanLink111[11] , \ScanLink171[15] , 
        \ScanLink152[24] , \ScanLink104[25] , \ScanLink89[17] , 
        \ScanLink127[14] , \ScanLink53[4] , \wBMid73[8] , \wAIn84[16] , 
        \wAIn91[22] , \wBIn106[1] , \wRegInA13[0] , \wRegInA58[24] , 
        \ScanLink170[9] , \wRegInB88[13] , \wRegInA3[5] , \wRegInA38[20] , 
        \wRegInB73[5] , \ScanLink81[2] , \wBIn75[23] , \wBIn116[12] , 
        \wBIn36[16] , \wAIn47[3] , \wBIn56[12] , \wAMid59[15] , \wAMid39[11] , 
        \wBIn43[26] , \wBIn120[17] , \wBIn22[0] , \wBIn60[17] , \wBIn103[26] , 
        \wRegInB101[4] , \wRegInA105[10] , \wAIn113[7] , \wAMid3[31] , 
        \wAMid3[28] , \wAIn95[5] , \ScanLink111[0] , \wRegInA72[9] , 
        \wRegInA126[21] , \wBMid10[19] , \wBIn21[3] , \wRegInA110[24] , 
        \ScanLink181[18] , \ScanLink112[3] , \wAIn44[0] , \wAIn96[6] , 
        \wAIn110[4] , \wAMid110[12] , \wRegInB9[11] , \wRegInB108[21] , 
        \ScanLink159[31] , \ScanLink159[28] , \wRegInA53[28] , \wAMid81[25] , 
        \wRegInA26[18] , \wAMid94[11] , \wBMid109[23] , \wRegInA53[31] , 
        \wRegInA70[19] , \wAMid105[26] , \wAMid126[17] , \wRegInB102[7] , 
        \ScanLink175[4] , \wBMid33[31] , \wBIn46[4] , \ScanLink79[30] , 
        \wBMid33[28] , \wBMid65[29] , \wRegInA110[17] , \ScanLink79[29] , 
        \wBMid46[18] , \wRegInA6[8] , \wBMid65[30] , \wRegInB76[8] , 
        \wRegInA105[23] , \ScanLink231[18] , \ScanLink212[30] , 
        \ScanLink215[1] , \wRegInA126[12] , \ScanLink244[28] , 
        \ScanLink212[29] , \wAIn4[1] , \wAIn22[29] , \wAIn23[7] , \wBIn43[15] , 
        \wAIn74[31] , \wBIn94[2] , \wBIn120[24] , \wRegInB18[29] , 
        \ScanLink244[31] , \wAIn57[19] , \wBIn36[25] , \wAMid39[22] , 
        \wAIn7[2] , \wBIn15[14] , \wAIn22[30] , \wBIn60[24] , \wAIn74[28] , 
        \wBIn103[15] , \wRegInB18[30] , \wAMid63[3] , \wBIn23[11] , 
        \wBIn56[21] , \wAMid59[26] , \wBIn75[10] , \wBIn116[21] , 
        \ScanLink56[9] , \ScanLink99[0] , \wAIn20[4] , \wBIn58[8] , 
        \wAMid60[0] , \wAMid126[24] , \wAMid94[22] , \wBIn97[1] , 
        \wAMid105[15] , \wRegInB96[18] , \wAMid26[5] , \wBIn45[7] , 
        \wAMid81[16] , \wAMid110[21] , \wBMid109[10] , \wRegInB68[4] , 
        \wRegInB108[12] , \ScanLink82[28] , \wAIn66[1] , \wBIn81[25] , 
        \wAIn95[30] , \wRegInB9[22] , \ScanLink216[2] , \ScanLink176[7] , 
        \ScanLink82[31] , \ScanLink48[5] , \ScanLink9[9] , \wBMid106[24] , 
        \wBMid125[15] , \ScanLink130[2] , \wBMid84[28] , \wBIn94[11] , 
        \wAIn95[29] , \ScanLink250[7] , \wBMid113[10] , \ScanLink98[31] , 
        \ScanLink4[17] , \wBMid116[7] , \ScanLink98[28] , \wBMid84[31] , 
        \wBIn5[30] , \wBMid4[1] , \wRegInB112[12] , \wBMid7[2] , \wAMid25[6] , 
        \wBMid29[28] , \wBMid51[9] , \wRegInB6[16] , \wRegInB107[26] , 
        \wRegInB120[6] , \wRegInB124[17] , \ScanLink35[31] , \ScanLink16[19] , 
        \wBMid115[4] , \ScanLink63[29] , \wBMid29[31] , \ScanLink35[28] , 
        \wAIn65[2] , \ScanLink63[30] , \wRegInB123[5] , \ScanLink208[29] , 
        \ScanLink40[18] , \ScanLink208[30] , \wAMid15[27] , \wAMid23[22] , 
        \wAIn38[30] , \wAMid38[9] , \wAMid75[23] , \wRegInB54[28] , 
        \wBIn119[15] , \wRegInB21[18] , \wAMid36[16] , \wAIn38[29] , 
        \ScanLink133[1] , \wAMid56[12] , \wBIn59[15] , \wRegInB54[31] , 
        \wRegInB77[19] , \wRegInA50[8] , \wBIn39[11] , \wAMid43[26] , 
        \wAMid42[1] , \wAMid60[17] , \ScanLink253[4] , \wRegInB107[15] , 
        \wRegInB6[25] , \wRegInB124[24] , \ScanLink186[0] , \ScanLink149[9] , 
        \ScanLink136[18] , \ScanLink115[30] , \ScanLink143[28] , \wAIn3[27] , 
        \wAIn3[14] , \wBIn5[29] , \wRegInB112[21] , \ScanLink115[29] , 
        \wAMid5[6] , \wBIn67[6] , \wAMid90[7] , \ScanLink160[19] , 
        \ScanLink143[31] , \wBIn94[22] , \wRegInA49[31] , \wBMid113[23] , 
        \ScanLink154[6] , \ScanLink4[24] , \wBMid125[26] , \wRegInA49[28] , 
        \wRegInA115[0] , \wAMid6[5] , \wAMid15[14] , \wBMid28[2] , 
        \wAMid36[25] , \wAMid43[15] , \wBIn64[5] , \wBIn81[16] , 
        \wBMid106[17] , \ScanLink234[3] , \wRegInB98[3] , \ScanLink157[5] , 
        \wBIn39[22] , \wRegInA91[18] , \wAMid60[24] , \wAMid93[4] , 
        \wAMid75[10] , \ScanLink237[0] , \wAMid7[10] , \wAIn8[18] , 
        \wAMid23[11] , \wAMid56[21] , \wBIn59[26] , \wBIn119[26] , 
        \wRegInB54[9] , \ScanLink69[7] , \wAIn106[18] , \wRegInA116[3] , 
        \ScanLink185[3] , \wAIn125[30] , \wRegInA29[3] , \wBIn8[7] , 
        \wBIn18[3] , \wAMid41[2] , \wBMid54[4] , \wBMid86[2] , \wAIn125[29] , 
        \wRegInB9[6] , \wRegInB49[6] , \ScanLink74[8] , \wBMid110[9] , 
        \wRegInB35[0] , \wRegInA55[5] , \ScanLink128[20] , \ScanLink86[23] , 
        \ScanLink256[9] , \ScanLink148[24] , \ScanLink93[17] , \wAMid90[29] , 
        \wRegInA14[25] , \wRegInA61[15] , \wRegInA37[14] , \wRegInB92[13] , 
        \wAMid90[30] , \wRegInA42[24] , \wRegInA22[20] , \wRegInA87[3] , 
        \wRegInB87[27] , \ScanLink15[1] , \wRegInA57[10] , \wRegInA74[21] , 
        \wRegInB126[8] , \wAIn10[27] , \wAMid23[8] , \wAIn26[22] , 
        \wAMid48[19] , \wAIn53[12] , \ScanLink128[0] , \wRegInB69[12] , 
        \wRegInA84[0] , \wBMid57[7] , \wAIn70[23] , \wAIn65[17] , 
        \ScanLink248[5] , \wBMid14[12] , \wAIn33[16] , \wAIn46[26] , 
        \ScanLink16[2] , \ScanLink203[16] , \wBMid61[22] , \wRegInA56[6] , 
        \wBMid37[23] , \wBMid85[1] , \ScanLink220[27] , \ScanLink185[20] , 
        \wAMid3[8] , \wBMid6[31] , \wBMid22[17] , \wBMid42[13] , 
        \ScanLink255[17] , \wRegInA101[28] , \ScanLink68[16] , \wBMid57[27] , 
        \ScanLink235[13] , \ScanLink190[14] , \wRegInB36[3] , \wBMid6[28] , 
        \wBMid74[16] , \wRegInA101[31] , \ScanLink240[23] , \wRegInA122[19] , 
        \ScanLink216[22] , \wAIn19[4] , \wBMid30[0] , \wAMid106[1] , 
        \wAIn118[20] , \wRegInA57[23] , \wAMid114[19] , \wRegInA22[13] , 
        \wRegInB87[14] , \wRegInA74[12] , \wBIn61[8] , \wRegInA14[16] , 
        \wRegInA61[26] , \wRegInA37[27] , \wRegInA42[17] , \wRegInB83[2] , 
        \ScanLink71[5] , \wRegInB92[20] , \ScanLink152[8] , \ScanLink148[17] , 
        \wAMid59[0] , \wAMid96[9] , \wBIn124[0] , \wRegInA31[1] , 
        \ScanLink93[24] , \wAMid7[23] , \wBMid22[24] , \wBMid57[14] , 
        \wRegInB51[4] , \ScanLink86[10] , \ScanLink128[13] , \ScanLink240[10] , 
        \ScanLink68[25] , \wBMid74[25] , \ScanLink235[20] , \ScanLink190[27] , 
        \wAIn118[13] , \wBIn127[3] , \wRegInA32[2] , \ScanLink216[11] , 
        \wBMid14[21] , \wBMid61[11] , \ScanLink203[25] , \wBMid2[19] , 
        \wAMid3[21] , \wAMid3[12] , \wAIn10[14] , \wBIn27[30] , \wBMid33[3] , 
        \wBMid37[10] , \wBMid42[20] , \ScanLink255[24] , \wRegInB52[7] , 
        \ScanLink220[14] , \ScanLink185[13] , \wBMid10[10] , \wAIn26[11] , 
        \wBIn27[29] , \wAIn65[24] , \wBIn71[28] , \wAMid88[5] , \wBIn112[19] , 
        \wAIn33[25] , \wAIn46[15] , \wBIn71[31] , \wBIn52[19] , \wAMid105[2] , 
        \wRegInB69[21] , \wBMid26[15] , \wAIn53[21] , \ScanLink72[6] , 
        \wAIn70[10] , \wRegInB80[1] , \wBMid53[25] , \wRegInB76[1] , 
        \ScanLink231[11] , \ScanLink215[8] , \ScanLink194[16] , 
        \ScanLink19[24] , \wBMid70[14] , \ScanLink244[21] , \ScanLink212[20] , 
        \ScanLink84[6] , \wBIn89[4] , \ScanLink207[14] , \wBMid65[20] , 
        \wAIn109[16] , \wRegInA16[4] , \wAIn4[8] , \wAIn7[16] , \wBMid33[21] , 
        \wBIn103[5] , \ScanLink224[25] , \ScanLink181[22] , \ScanLink251[15] , 
        \ScanLink79[20] , \wAIn14[25] , \wBMid46[11] , \wRegInA6[1] , 
        \wBIn56[31] , \wAIn61[15] , \wBIn75[19] , \wBIn116[28] , 
        \ScanLink208[7] , \wAIn22[20] , \wBIn23[18] , \wAIn37[14] , 
        \wAIn42[24] , \wBIn56[28] , \ScanLink56[0] , \wBIn116[31] , 
        \ScanLink99[9] , \wAIn57[10] , \wRegInB18[20] , \wRegInB78[24] , 
        \ScanLink168[2] , \wAMid121[4] , \wAIn14[16] , \wBMid14[6] , 
        \wBMid17[5] , \wAIn74[21] , \wBMid109[19] , \wAMid110[31] , 
        \wAMid110[28] , \wRegInA26[22] , \wRegInB83[25] , \ScanLink55[3] , 
        \wRegInA53[12] , \wRegInA10[27] , \wRegInA70[23] , \wAIn22[13] , 
        \wBIn58[1] , \wAMid60[9] , \wRegInA65[17] , \wRegInA33[16] , 
        \wRegInB96[11] , \wBIn97[8] , \wBIn100[6] , \wAMid122[7] , 
        \wRegInA46[26] , \wRegInA5[2] , \wRegInB75[2] , \ScanLink139[16] , 
        \ScanLink87[5] , \ScanLink97[15] , \ScanLink9[0] , \ScanLink82[21] , 
        \wRegInA15[7] , \ScanLink159[12] , \wAMid39[18] , \wAIn57[23] , 
        \wRegInB18[13] , \ScanLink32[4] , \wAIn74[12] , \wAIn37[27] , 
        \wAIn61[26] , \wBMid73[1] , \wAIn42[17] , \wAIn88[3] , \wRegInB78[17] , 
        \wAIn109[25] , \wAIn7[25] , \wBMid10[23] , \wBMid65[13] , 
        \ScanLink207[27] , \ScanLink251[26] , \wBMid26[26] , \wBMid33[12] , 
        \wBMid46[22] , \ScanLink224[16] , \ScanLink181[11] , \wBMid53[16] , 
        \wRegInB12[5] , \ScanLink79[13] , \ScanLink19[17] , \ScanLink244[12] , 
        \wRegInA105[19] , \wRegInA126[31] , \ScanLink231[22] , 
        \ScanLink194[25] , \wAMid11[25] , \wAMid19[2] , \wBIn22[9] , 
        \wBMid70[27] , \wAIn59[6] , \wRegInB9[18] , \wRegInB11[6] , 
        \wRegInA72[0] , \wRegInA126[28] , \ScanLink111[9] , \ScanLink212[13] , 
        \ScanLink82[12] , \wRegInB108[31] , \wRegInB108[28] , 
        \ScanLink159[21] , \wRegInA71[3] , \ScanLink139[25] , \ScanLink97[26] , 
        \wAMid32[14] , \wAIn44[9] , \wAMid94[18] , \wRegInA65[24] , 
        \wRegInA10[14] , \wRegInA33[25] , \wRegInA46[15] , \ScanLink31[7] , 
        \wRegInA53[21] , \wRegInB96[22] , \wBMid70[2] , \wRegInA26[11] , 
        \wRegInB83[16] , \wRegInA70[10] , \wAMid47[24] , \wRegInA95[30] , 
        \ScanLink82[8] , \wBIn48[23] , \wAMid64[15] , \wBIn108[23] , 
        \ScanLink213[6] , \wRegInA95[29] , \wAMid71[21] , \wAIn1[5] , 
        \wBIn1[18] , \wAIn2[6] , \wAMid27[20] , \wBIn28[27] , \wBIn40[3] , 
        \ScanLink173[3] , \wAMid52[10] , \wAIn102[30] , \wAIn102[29] , 
        \wAIn121[18] , \wBMid9[15] , \wAMid65[4] , \wBMid12[8] , \wAIn25[0] , 
        \wBIn92[5] , \wAIn26[3] , \wBIn91[6] , \wBIn118[4] , \wRegInB2[14] , 
        \wRegInB103[24] , \wRegInB120[15] , \ScanLink147[19] , \wAMid124[9] , 
        \ScanLink164[31] , \ScanLink132[29] , \wBMid9[26] , \wBIn43[0] , 
        \wAMid66[7] , \ScanLink164[28] , \wBIn90[13] , \wBMid117[12] , 
        \wRegInA4[11] , \wRegInB116[10] , \ScanLink210[5] , \ScanLink132[30] , 
        \ScanLink111[18] , \ScanLink0[15] , \wBMid121[17] , \wRegInA38[30] , 
        \wRegInA38[29] , \wBMid58[30] , \wBMid58[29] , \wBIn85[27] , 
        \wBIn106[8] , \ScanLink170[0] , \wRegInA13[9] , \wBMid102[26] , 
        \ScanLink67[18] , \ScanLink44[30] , \wRegInB107[3] , \ScanLink12[28] , 
        \ScanLink44[29] , \ScanLink31[19] , \ScanLink12[31] , \wBIn39[8] , 
        \wAIn41[4] , \wRegInA69[1] , \wAIn49[31] , \wAMid71[12] , \wBMid3[13] , 
        \wAMid11[16] , \wBIn24[7] , \wAMid27[13] , \wBIn28[14] , \wAIn49[28] , 
        \wAMid52[23] , \wRegInB25[29] , \wRegInB50[19] , \wRegInB73[31] , 
        \wRegInB25[30] , \ScanLink29[5] , \wRegInB73[28] , \wAMid32[27] , 
        \wAMid47[17] , \wAIn115[0] , \ScanLink117[7] , \wBIn48[10] , 
        \wAIn93[2] , \wAMid64[26] , \wBMid68[0] , \wBIn108[10] , \wBMid11[30] , 
        \wAMid14[7] , \wBIn27[4] , \wBIn85[14] , \wAIn91[18] , \wBMid121[24] , 
        \wRegInB88[29] , \wRegInB17[8] , \wRegInB88[30] , \wBIn90[20] , 
        \wBMid102[15] , \wBMid117[21] , \ScanLink0[26] , \ScanLink114[4] , 
        \wAIn42[7] , \wBMid80[19] , \wAIn90[1] , \wAIn116[3] , \ScanLink37[9] , 
        \wRegInB2[27] , \wRegInA4[22] , \wRegInB103[17] , \wRegInB104[0] , 
        \wRegInB116[23] , \wRegInB120[26] , \wBMid60[8] , \wAMid80[26] , 
        \wAMid95[12] , \wAMid104[25] , \wRegInB97[28] , \wRegInB97[31] , 
        \wRegInB112[4] , \wBMid108[20] , \wBMid124[5] , \wBIn31[0] , 
        \wAIn54[3] , \wAMid111[11] , \wRegInB8[12] , \wRegInB109[22] , 
        \ScanLink83[18] , \ScanLink102[0] , \wBMid32[18] , \wBMid47[28] , 
        \wAIn86[5] , \wAIn100[7] , \wRegInA61[9] , \ScanLink78[19] , 
        \wRegInA111[27] , \wBMid11[29] , \wBMid47[31] , \wBMid64[19] , 
        \wBIn32[3] , \wAIn103[4] , \wBIn14[24] , \wAIn85[6] , \ScanLink101[3] , 
        \wRegInA104[13] , \wRegInA127[22] , \ScanLink245[18] , 
        \ScanLink230[31] , \ScanLink213[19] , \ScanLink230[28] , \wAMid17[4] , 
        \wBIn22[21] , \wAIn23[19] , \wBIn37[15] , \wAIn56[30] , \wBIn61[14] , 
        \wBIn102[25] , \wAIn75[18] , \wRegInB111[7] , \wAMid38[12] , 
        \wBIn42[25] , \wAIn56[29] , \wBIn121[14] , \wRegInB19[19] , 
        \wAIn57[0] , \wBIn57[11] , \wAMid58[16] , \wAIn98[9] , \wBIn74[20] , 
        \wBMid19[3] , \wBIn55[4] , \wBIn117[11] , \wRegInB65[8] , 
        \ScanLink206[1] , \wRegInA127[2] , \ScanLink58[6] , \wRegInB8[21] , 
        \ScanLink166[4] , \ScanLink158[18] , \wRegInA27[31] , \wRegInB109[11] , 
        \wBIn0[21] , \wAMid2[18] , \wBMid3[20] , \wBIn14[17] , \wBIn22[12] , 
        \wAIn30[7] , \wAMid80[15] , \wBIn87[2] , \wAMid104[16] , 
        \wBMid108[13] , \wAMid111[22] , \wRegInA71[29] , \wRegInB78[7] , 
        \ScanLink4[5] , \wRegInA27[28] , \wRegInA52[18] , \wRegInA71[30] , 
        \ScanLink45[9] , \wRegInA18[2] , \wBIn57[22] , \wAMid58[25] , 
        \wAMid70[3] , \wAMid95[21] , \wRegInA8[7] , \ScanLink89[3] , 
        \wBIn61[27] , \wBIn74[13] , \wBIn102[16] , \wBIn117[22] , 
        \ScanLink7[6] , \wAMid73[0] , \wAIn33[4] , \wBIn42[16] , \wBIn84[1] , 
        \wBIn121[27] , \ScanLink178[8] , \wBIn37[26] , \wAMid38[21] , 
        \wRegInA124[1] , \wRegInA127[11] , \wBIn56[7] , \wRegInA104[20] , 
        \wRegInA111[14] , \ScanLink205[2] , \ScanLink180[28] , 
        \ScanLink180[31] , \ScanLink165[7] , \wRegInA5[28] , \wRegInB117[29] , 
        \ScanLink110[21] , \wBIn0[12] , \wAMid9[14] , \wAMid12[9] , 
        \wBMid66[6] , \wBMid81[13] , \ScanLink165[11] , \wBMid94[27] , 
        \wRegInA5[31] , \wRegInB117[30] , \ScanLink27[3] , \ScanLink146[20] , 
        \ScanLink133[10] , \ScanLink126[24] , \ScanLink119[1] , 
        \ScanLink153[14] , \ScanLink105[15] , \ScanLink170[25] , \wAMid26[19] , 
        \wAIn48[22] , \wAIn85[26] , \wAIn90[12] , \wRegInB109[5] , 
        \ScanLink88[27] , \wAIn106[9] , \wRegInA39[10] , \wRegInA59[14] , 
        \wRegInB89[23] , \wRegInA67[7] , \wAMid53[29] , \wAIn28[26] , 
        \wAMid53[30] , \wAMid70[18] , \wRegInB72[22] , \wAIn83[8] , 
        \wRegInB12[26] , \wRegInB24[23] , \wRegInA81[24] , \wRegInB31[17] , 
        \wRegInB51[13] , \wRegInB44[27] , \wRegInA94[10] , \wRegInA64[4] , 
        \wRegInB67[16] , \wBIn29[2] , \wBMid39[27] , \wBMid59[23] , 
        \wAIn116[24] , \ScanLink218[26] , \ScanLink45[23] , \ScanLink30[13] , 
        \ScanLink24[0] , \ScanLink66[12] , \ScanLink13[22] , \wBMid65[5] , 
        \wBMid121[8] , \wRegInB117[9] , \wAIn120[21] , \ScanLink73[26] , 
        \wAIn103[10] , \wAIn118[5] , \ScanLink50[17] , \wAIn85[15] , 
        \wBIn91[19] , \wRegInA39[23] , \ScanLink91[1] , \ScanLink25[27] , 
        \wBMid116[18] , \wAIn90[21] , \wRegInB63[6] , \wBMid94[14] , 
        \wBIn116[2] , \wRegInA59[27] , \wRegInB89[10] , \ScanLink153[27] , 
        \ScanLink126[17] , \ScanLink43[7] , \ScanLink170[16] , 
        \ScanLink105[26] , \ScanLink88[14] , \wRegInA0[2] , \wAIn1[8] , 
        \wBIn1[26] , \wBMid2[27] , \wBMid2[14] , \wBIn4[23] , \wAMid8[3] , 
        \wAIn9[12] , \wAMid9[27] , \wAIn36[9] , \wBMid81[20] , 
        \ScanLink165[22] , \ScanLink146[13] , \ScanLink110[12] , 
        \ScanLink133[23] , \wBMid39[14] , \wAIn120[12] , \ScanLink1[8] , 
        \wAIn103[23] , \ScanLink73[15] , \ScanLink40[4] , \ScanLink25[14] , 
        \wBMid25[7] , \wAIn28[15] , \wBIn49[30] , \wBMid59[10] , \wAIn116[17] , 
        \ScanLink50[24] , \ScanLink30[20] , \ScanLink218[15] , 
        \ScanLink45[10] , \ScanLink13[11] , \wBIn109[29] , \wRegInB44[14] , 
        \ScanLink66[21] , \wRegInB31[24] , \wRegInB60[5] , \wRegInA94[23] , 
        \wRegInB67[25] , \ScanLink92[2] , \wAIn28[5] , \wAIn48[11] , 
        \wBIn49[29] , \wBIn109[30] , \wRegInB12[15] , \wBIn50[9] , 
        \ScanLink163[9] , \wRegInB72[11] , \wAMid68[1] , \wBIn115[1] , 
        \wRegInB51[20] , \wRegInB24[10] , \wRegInA81[17] , \wAMid51[8] , 
        \wAIn124[23] , \ScanLink77[24] , \wBMid26[4] , \wBMid28[11] , 
        \wBMid48[15] , \wBIn69[0] , \wAIn107[12] , \wRegInA39[9] , 
        \ScanLink209[10] , \ScanLink195[9] , \ScanLink54[15] , \wAIn112[26] , 
        \wAMid113[6] , \ScanLink64[2] , \ScanLink41[21] , \ScanLink21[25] , 
        \ScanLink34[11] , \ScanLink62[10] , \wBIn38[31] , \wBMid38[8] , 
        \wRegInB96[5] , \ScanLink17[20] , \wRegInB4[3] , \wRegInB35[15] , 
        \wRegInB40[25] , \wRegInA90[12] , \wBIn38[28] , \wAIn59[14] , 
        \wRegInB16[24] , \ScanLink188[6] , \wRegInA24[6] , \wRegInB63[14] , 
        \wAIn39[10] , \wAIn81[24] , \wBIn95[31] , \wBMid112[30] , 
        \wRegInB20[21] , \wRegInB76[20] , \wRegInA85[26] , \wRegInA106[9] , 
        \wRegInA27[5] , \wRegInB44[3] , \wRegInA48[22] , \wRegInB55[11] , 
        \wRegInB98[15] , \wRegInB7[0] , \wBMid90[25] , \wAIn94[10] , 
        \wBIn95[28] , \wBMid112[29] , \wRegInB47[0] , \ScanLink224[9] , 
        \wRegInA28[26] , \wRegInB88[9] , \ScanLink159[3] , \ScanLink122[26] , 
        \wAMid110[5] , \ScanLink157[16] , \ScanLink101[17] , \ScanLink174[27] , 
        \ScanLink239[6] , \ScanLink114[23] , \ScanLink99[11] , \wBIn4[10] , 
        \wAIn9[21] , \wAMid22[31] , \wAMid22[28] , \wAIn39[23] , \wBMid85[11] , 
        \wRegInB95[6] , \ScanLink161[13] , \wRegInA118[5] , \ScanLink137[12] , 
        \ScanLink67[1] , \ScanLink142[22] , \wAMid57[18] , \wRegInB76[13] , 
        \wAIn68[7] , \wAMid74[30] , \wBMid93[5] , \wRegInA40[2] , \wAMid28[3] , 
        \wAMid74[29] , \wBMid118[1] , \wRegInB55[22] , \wBMid28[22] , 
        \wBMid41[3] , \wAIn59[27] , \wRegInB16[17] , \wRegInB20[12] , 
        \wRegInA85[15] , \wRegInB20[7] , \wRegInB35[26] , \wRegInB40[16] , 
        \wRegInA90[21] , \wRegInB63[27] , \wAIn75[8] , \wAIn112[15] , 
        \ScanLink34[22] , \wRegInA92[4] , \ScanLink41[12] , \ScanLink17[13] , 
        \ScanLink62[23] , \wBMid48[26] , \wAIn124[10] , \wAIn107[21] , 
        \ScanLink77[17] , \ScanLink209[23] , \ScanLink21[16] , 
        \ScanLink54[26] , \wBIn5[2] , \wAMid6[30] , \wBMid7[11] , \wBIn10[26] , 
        \wBMid9[4] , \wBIn13[8] , \wBMid42[0] , \wBMid85[22] , \wRegInA1[19] , 
        \ScanLink161[20] , \ScanLink99[22] , \wRegInB113[18] , 
        \ScanLink142[11] , \ScanLink114[10] , \wBMid90[16] , \wRegInA91[7] , 
        \ScanLink157[25] , \ScanLink137[21] , \ScanLink122[15] , \wBMid90[6] , 
        \wAIn94[23] , \ScanLink174[14] , \ScanLink101[24] , \wAIn81[17] , 
        \wRegInA28[15] , \wRegInA43[1] , \ScanLink120[8] , \wRegInA48[11] , 
        \wRegInB98[26] , \wAIn17[2] , \wBIn26[23] , \wAMid29[24] , 
        \wRegInB23[4] , \ScanLink193[7] , \wBIn53[13] , \wBMid23[9] , 
        \wAMid115[8] , \wAMid57[6] , \wBIn70[22] , \wBIn113[13] , \wBIn33[17] , 
        \wBIn65[16] , \wBIn106[27] , \wBIn46[27] , \wBIn125[16] , 
        \wAMid49[20] , \wBIn72[1] , \wAMid85[0] , \wAMid108[7] , \wAIn119[19] , 
        \ScanLink141[1] , \wRegInA22[8] , \wRegInA123[20] , \wRegInA100[11] , 
        \ScanLink221[4] , \wAMid6[29] , \wRegInA115[25] , \ScanLink184[19] , 
        \wAIn14[1] , \wAMid54[5] , \wBIn71[2] , \wAMid86[3] , \wRegInA100[7] , 
        \wRegInB118[14] , \ScanLink142[2] , \wAMid84[24] , \wRegInA103[4] , 
        \ScanLink129[19] , \ScanLink222[7] , \wRegInA56[30] , \wRegInA75[18] , 
        \wRegInA56[29] , \ScanLink190[4] , \wBMid36[29] , \wAMid91[10] , 
        \wAMid100[27] , \wAMid115[13] , \wRegInA23[19] , \wBMid119[16] , 
        \wAMid123[16] , \wRegInB93[8] , \wRegInA115[16] , \wBMid43[19] , 
        \wBMid60[31] , \wBIn6[1] , \wBMid7[22] , \wBIn16[5] , \wBMid15[18] , 
        \wAIn127[2] , \ScanLink125[5] , \wBMid36[30] , \wBMid60[28] , 
        \wRegInA89[5] , \wRegInA123[13] , \ScanLink217[28] , \wBIn10[15] , 
        \wBIn65[25] , \wAIn71[29] , \wBMid88[4] , \wBIn106[14] , 
        \wRegInB26[9] , \wRegInA100[22] , \ScanLink241[30] , \ScanLink245[0] , 
        \ScanLink217[31] , \ScanLink234[19] , \ScanLink241[29] , \wBMid103[0] , 
        \wBIn15[6] , \wBIn26[10] , \wAIn27[31] , \wAMid33[2] , \wAIn27[28] , 
        \wBIn46[14] , \wBIn125[25] , \wAMid49[13] , \wAIn52[18] , \wAIn71[30] , 
        \wAIn73[6] , \wRegInB68[18] , \wAMid29[17] , \wBIn33[24] , 
        \wBIn53[20] , \wAMid30[1] , \wAIn70[5] , \wBIn70[11] , \wAMid100[14] , 
        \wBIn113[20] , \wRegInB93[19] , \wRegInA58[0] , \wRegInA97[9] , 
        \wBMid100[3] , \wAMid123[25] , \wAMid84[17] , \wAMid91[23] , 
        \wBMid119[25] , \wAMid115[20] , \wRegInB38[5] , \wAIn124[1] , 
        \wAIn7[31] , \wAIn7[28] , \wBIn21[7] , \wAIn44[4] , \wBMid59[1] , 
        \ScanLink126[6] , \ScanLink87[30] , \wAMid81[21] , \wAMid94[15] , 
        \wBMid96[8] , \wAMid105[22] , \wRegInA33[28] , \wRegInA46[18] , 
        \wRegInA65[30] , \wRegInB118[27] , \ScanLink246[3] , \ScanLink87[29] , 
        \ScanLink18[4] , \wRegInA65[29] , \wBMid109[27] , \wAMid126[13] , 
        \wRegInA10[19] , \wRegInA33[31] , \wRegInB102[3] , \wAMid110[16] , 
        \wRegInB9[15] , \wRegInB108[25] , \ScanLink139[31] , \ScanLink112[7] , 
        \wAIn96[2] , \wAIn110[0] , \ScanLink139[28] , \wAIn109[31] , 
        \wAIn109[28] , \wRegInB12[8] , \wRegInA110[20] , \wBIn22[4] , 
        \wAIn4[5] , \wAIn7[6] , \wBIn15[23] , \wAIn95[1] , \wAIn113[3] , 
        \ScanLink111[4] , \wRegInA105[14] , \wRegInA126[25] , 
        \ScanLink194[31] , \ScanLink194[28] , \wAIn20[0] , \wBIn23[26] , 
        \wBIn36[12] , \wAMid39[15] , \wBIn60[13] , \wBIn103[22] , 
        \wRegInB101[0] , \ScanLink32[9] , \wBIn43[22] , \wBIn120[13] , 
        \wBIn45[3] , \wAIn47[7] , \wBIn56[16] , \wAMid59[11] , \wBIn75[27] , 
        \wBIn116[16] , \ScanLink216[6] , \ScanLink97[18] , \ScanLink87[8] , 
        \ScanLink48[1] , \wAMid81[12] , \wBMid109[14] , \wRegInB9[26] , 
        \wRegInB83[31] , \wRegInB108[16] , \ScanLink176[3] , \wBIn97[5] , 
        \wAMid105[11] , \wAMid110[25] , \wRegInB68[0] , \wRegInB83[28] , 
        \wAIn14[31] , \wAIn42[29] , \wAMid60[4] , \wAMid126[20] , 
        \wAMid94[26] , \wBIn56[25] , \wAMid59[22] , \ScanLink99[4] , 
        \wAIn14[28] , \wBIn23[15] , \wAIn37[19] , \wAIn42[30] , 
        \wRegInB78[29] , \wAIn61[18] , \wBIn75[14] , \wBIn116[25] , 
        \wRegInB78[30] , \wBIn15[10] , \wBMid17[8] , \wBIn103[11] , 
        \wBIn60[20] , \wAIn23[3] , \wBIn43[11] , \wAMid63[7] , \wBIn94[6] , 
        \wBIn120[20] , \wAMid121[9] , \wBIn36[21] , \wAMid39[26] , 
        \wRegInA126[16] , \wBMid26[18] , \wBMid53[31] , \wBMid70[19] , 
        \ScanLink19[30] , \wBIn46[0] , \wBMid53[28] , \wRegInA105[27] , 
        \ScanLink215[5] , \ScanLink19[29] , \wBIn89[9] , \wRegInA110[13] , 
        \ScanLink224[28] , \ScanLink251[18] , \ScanLink224[31] , 
        \ScanLink207[19] , \ScanLink175[0] , \wBIn103[8] , \wRegInA16[9] , 
        \ScanLink111[26] , \wBIn1[15] , \wAMid8[13] , \wBIn27[9] , 
        \wBMid76[1] , \wBMid80[14] , \ScanLink164[16] , \wBMid95[20] , 
        \ScanLink147[27] , \ScanLink132[17] , \ScanLink37[4] , 
        \ScanLink127[23] , \ScanLink109[6] , \ScanLink152[13] , 
        \ScanLink104[12] , \wBIn85[19] , \wBMid102[18] , \ScanLink171[22] , 
        \ScanLink89[20] , \wAIn91[15] , \wBMid121[30] , \wRegInB119[2] , 
        \wBMid121[29] , \wRegInB17[5] , \wRegInB88[24] , \wRegInA38[17] , 
        \wRegInA58[13] , \ScanLink114[9] , \wBIn28[19] , \wAIn49[25] , 
        \wAIn84[21] , \wRegInA77[0] , \ScanLink29[8] , \wAIn29[21] , 
        \wRegInB13[21] , \wRegInB14[6] , \wRegInB25[24] , \wRegInB73[25] , 
        \wRegInB50[14] , \wRegInA80[23] , \wRegInB30[10] , \wRegInA95[17] , 
        \wRegInB45[20] , \wRegInB66[11] , \wRegInA74[3] , \wBIn39[5] , 
        \wBMid38[20] , \wBMid58[24] , \wAIn117[23] , \ScanLink219[21] , 
        \ScanLink44[24] , \ScanLink34[7] , \ScanLink31[14] , \ScanLink67[15] , 
        \wBMid75[2] , \ScanLink12[25] , \ScanLink72[21] , \wAIn121[26] , 
        \wAIn102[17] , \wAIn108[2] , \ScanLink51[10] , \wAIn41[9] , 
        \ScanLink24[20] , \wAIn84[12] , \wRegInA38[24] , \ScanLink81[6] , 
        \ScanLink210[8] , \ScanLink0[18] , \wAIn91[26] , \wRegInB73[1] , 
        \wBMid95[13] , \wBIn106[5] , \wRegInA3[1] , \wRegInA13[4] , 
        \wRegInA58[20] , \wRegInB88[17] , \wRegInB103[30] , \ScanLink152[20] , 
        \ScanLink53[0] , \wRegInB120[18] , \ScanLink127[10] , \wRegInB2[19] , 
        \wRegInB103[29] , \ScanLink171[11] , \ScanLink89[13] , 
        \ScanLink104[21] , \wBMid12[5] , \ScanLink164[25] , \wAMid8[20] , 
        \wBMid38[13] , \wBMid80[27] , \ScanLink147[14] , \ScanLink111[15] , 
        \wAIn121[15] , \wAMid124[4] , \ScanLink132[24] , \ScanLink72[12] , 
        \wAIn102[24] , \ScanLink50[3] , \ScanLink24[13] , \wBMid9[18] , 
        \wBIn92[8] , \ScanLink51[23] , \ScanLink31[27] , \wAMid11[31] , 
        \wAMid11[28] , \wBMid11[6] , \wBMid58[17] , \wAIn117[10] , 
        \wBIn118[9] , \ScanLink44[17] , \ScanLink219[12] , \ScanLink12[16] , 
        \wAMid65[9] , \ScanLink67[26] , \wRegInB45[13] , \wAIn29[12] , 
        \wAMid32[19] , \wAMid47[30] , \wAMid64[18] , \wRegInB30[23] , 
        \wRegInA95[24] , \wRegInB70[2] , \wRegInB66[22] , \ScanLink82[5] , 
        \wAIn38[2] , \wAMid47[29] , \wRegInB13[12] , \wAIn49[16] , 
        \wRegInB73[16] , \wBIn105[6] , \wRegInA10[7] , \wRegInB50[27] , 
        \wBIn5[24] , \wAMid6[8] , \wAIn8[15] , \wBMid35[0] , \wAMid78[6] , 
        \wRegInB25[17] , \wRegInA80[10] , \wAIn125[24] , \ScanLink76[23] , 
        \wAMid15[19] , \wBMid29[16] , \wBMid49[12] , \wBIn79[7] , 
        \wAMid103[1] , \wAIn106[15] , \ScanLink208[17] , \ScanLink55[12] , 
        \wAIn113[21] , \ScanLink74[5] , \ScanLink40[26] , \ScanLink20[22] , 
        \ScanLink35[16] , \wAMid60[29] , \wRegInB34[12] , \wRegInB86[2] , 
        \ScanLink63[17] , \wRegInA91[15] , \ScanLink16[27] , \wRegInB41[22] , 
        \wAMid36[31] , \wAMid93[9] , \wAMid36[28] , \wAMid43[18] , \wBIn64[8] , 
        \wRegInB17[23] , \ScanLink198[1] , \wAIn58[13] , \wAMid60[30] , 
        \ScanLink157[8] , \wBIn121[0] , \wRegInA34[1] , \wRegInB62[13] , 
        \wAIn38[17] , \wRegInB21[26] , \wRegInB77[27] , \wBMid36[3] , 
        \wAIn80[23] , \wBIn122[3] , \wRegInA49[25] , \wRegInB54[16] , 
        \wRegInB54[4] , \wRegInA84[21] , \wRegInB99[12] , \wRegInA37[2] , 
        \ScanLink4[30] , \wBMid91[22] , \wAIn95[17] , \wRegInB57[7] , 
        \ScanLink4[29] , \wRegInB6[28] , \wRegInA29[21] , \wRegInB124[29] , 
        \ScanLink149[4] , \ScanLink123[21] , \wAMid100[2] , \wRegInB107[18] , 
        \wRegInB124[30] , \ScanLink156[11] , \ScanLink100[10] , \wRegInB6[31] , 
        \ScanLink229[1] , \ScanLink175[20] , \ScanLink115[24] , 
        \ScanLink98[16] , \wBIn5[17] , \wAIn8[26] , \wBMid29[25] , 
        \wAIn38[24] , \wBMid84[16] , \wRegInB85[1] , \ScanLink160[14] , 
        \wRegInA108[2] , \ScanLink136[15] , \ScanLink77[6] , \ScanLink143[25] , 
        \wAMid38[4] , \wBIn59[18] , \wRegInB77[14] , \wAIn78[0] , \wBMid83[2] , 
        \wRegInA50[5] , \wBMid108[6] , \wRegInB54[25] , \wBMid51[4] , 
        \wAIn58[20] , \wBIn119[18] , \wRegInB17[10] , \wRegInB21[15] , 
        \wRegInB30[0] , \wRegInB34[21] , \wRegInB41[11] , \wRegInA84[12] , 
        \wRegInA91[26] , \ScanLink253[9] , \wRegInB62[20] , \wAIn113[12] , 
        \ScanLink35[25] , \wBMid115[9] , \wRegInA82[3] , \ScanLink40[15] , 
        \ScanLink16[14] , \ScanLink63[24] , \wBMid49[21] , \wAIn125[17] , 
        \wAIn106[26] , \wRegInB123[8] , \ScanLink76[10] , \ScanLink208[24] , 
        \ScanLink20[11] , \ScanLink10[1] , \ScanLink55[21] , \wAMid26[8] , 
        \wBMid52[7] , \ScanLink98[25] , \ScanLink160[27] , \wBMid84[25] , 
        \ScanLink143[16] , \ScanLink115[17] , \wRegInA81[0] , 
        \ScanLink136[26] , \ScanLink156[22] , \ScanLink13[2] , \wBIn0[25] , 
        \wBIn0[2] , \wAMid0[6] , \wBMid6[16] , \wAIn10[19] , \wBIn27[24] , 
        \wAIn33[28] , \wAIn80[10] , \wBIn81[31] , \wBIn81[28] , \wBMid91[11] , 
        \ScanLink123[12] , \wAIn95[24] , \ScanLink175[13] , \ScanLink100[23] , 
        \wBMid80[1] , \wBMid106[29] , \wBMid125[18] , \wBMid106[30] , 
        \wRegInA29[12] , \wRegInA53[6] , \wRegInA49[16] , \wRegInB99[21] , 
        \wRegInB33[3] , \ScanLink183[0] , \wAMid28[23] , \wAIn33[31] , 
        \wAIn46[18] , \wBIn52[14] , \wAIn65[30] , \wBIn11[21] , \wAMid47[1] , 
        \wAIn65[29] , \wBIn71[25] , \wAMid88[8] , \wBIn112[14] , \wBIn32[10] , 
        \wBIn64[11] , \wBIn107[20] , \wBIn47[20] , \wAMid48[27] , 
        \wBIn124[11] , \wBIn62[6] , \wBMid74[28] , \wBMid22[30] , 
        \ScanLink151[6] , \ScanLink68[31] , \wBMid22[29] , \wBMid57[19] , 
        \wAMid118[0] , \wRegInA122[27] , \wBMid74[31] , \wRegInA101[16] , 
        \ScanLink68[28] , \wAMid95[7] , \ScanLink255[29] , \ScanLink231[3] , 
        \wBMid1[1] , \wAIn3[19] , \wAMid3[5] , \wAIn19[9] , \wBIn61[5] , 
        \wAMid96[4] , \wRegInA110[0] , \wRegInA114[22] , \ScanLink220[19] , 
        \ScanLink203[31] , \ScanLink255[30] , \ScanLink203[28] , 
        \ScanLink93[29] , \wRegInB119[13] , \ScanLink152[5] , \ScanLink93[30] , 
        \wRegInA113[3] , \wAMid44[2] , \wAMid85[23] , \wRegInB51[9] , 
        \ScanLink232[0] , \wAMid90[17] , \wAMid101[20] , \wAMid114[14] , 
        \ScanLink180[3] , \wRegInB87[19] , \ScanLink71[8] , \wBMid118[11] , 
        \wAMid122[11] , \wRegInA114[11] , \wBMid6[25] , \wRegInA99[2] , 
        \ScanLink135[2] , \wRegInA122[14] , \wBIn11[12] , \wAMid23[5] , 
        \wBIn64[22] , \wBMid98[3] , \wRegInA101[25] , \ScanLink255[7] , 
        \ScanLink190[19] , \wBIn107[13] , \wBMid113[7] , \wBIn27[17] , 
        \wBIn32[23] , \wBIn47[13] , \wAMid48[14] , \wBIn124[22] , \wAIn63[1] , 
        \wBIn52[27] , \wAMid28[10] , \wBIn71[16] , \wBIn112[27] , 
        \wRegInB125[6] , \ScanLink248[8] , \wBMid2[2] , \wAMid20[6] , 
        \wBMid54[9] , \wAIn60[2] , \wAMid101[13] , \wRegInA14[31] , 
        \wRegInA37[19] , \wRegInA42[29] , \wRegInA48[7] , \wBMid110[4] , 
        \wAMid122[22] , \wRegInA14[28] , \wRegInA42[30] , \wAMid85[10] , 
        \wAMid90[24] , \wRegInA61[18] , \wBMid118[22] , \wBIn13[5] , 
        \wBMid49[6] , \wAMid114[27] , \wRegInB28[2] , \wRegInB126[5] , 
        \wRegInA55[8] , \ScanLink136[1] , \wAIn122[2] , \wRegInB119[20] , 
        \ScanLink256[4] , \ScanLink148[30] , \ScanLink148[29] , \wBMid124[12] , 
        \wAIn2[30] , \wAIn2[20] , \wAIn2[13] , \wBIn3[1] , \wBMid9[9] , 
        \wBIn80[22] , \wBMid107[23] , \wRegInA28[18] , \ScanLink120[5] , 
        \wBIn95[16] , \ScanLink240[0] , \ScanLink5[10] , \wBMid112[17] , 
        \wAMid35[1] , \wAMid36[2] , \wAIn76[6] , \wRegInB23[9] , \wBMid106[0] , 
        \wBMid105[3] , \wRegInA1[14] , \wRegInB7[11] , \wRegInB106[21] , 
        \wRegInB113[15] , \ScanLink174[19] , \ScanLink157[31] , 
        \wRegInB125[10] , \ScanLink157[28] , \ScanLink101[29] , 
        \ScanLink122[18] , \ScanLink101[30] , \wAMid74[24] , \wAIn75[5] , 
        \wAIn112[18] , \wBMid93[8] , \wRegInA92[9] , \wBIn118[12] , 
        \wRegInA85[18] , \wAMid6[17] , \wBIn10[18] , \wBIn10[6] , 
        \wAMid22[25] , \wAIn121[1] , \ScanLink123[6] , \wAIn11[1] , 
        \wAIn12[2] , \wAMid14[20] , \wAMid37[11] , \wBIn38[16] , \wAMid57[15] , 
        \wBIn58[12] , \wAMid42[21] , \wBMid26[9] , \wAMid61[10] , 
        \ScanLink243[3] , \wBMid90[31] , \wRegInB106[12] , \wAMid52[6] , 
        \wBMid90[28] , \wRegInB125[23] , \wRegInB7[22] , \ScanLink196[7] , 
        \wAMid14[13] , \wAMid37[22] , \wBIn38[25] , \wAMid42[12] , 
        \wAIn59[19] , \wBIn74[2] , \wBIn77[1] , \wAMid80[0] , \wAMid110[8] , 
        \wRegInA1[27] , \wRegInA118[8] , \wRegInB113[26] , \wAIn81[29] , 
        \wBIn95[25] , \ScanLink5[23] , \wBMid112[24] , \wRegInB98[18] , 
        \ScanLink144[1] , \wBIn80[11] , \wAIn81[30] , \wRegInA27[8] , 
        \wBMid107[10] , \wBMid124[21] , \wRegInA105[7] , \ScanLink224[4] , 
        \wRegInB88[4] , \wRegInB16[29] , \ScanLink147[2] , \wRegInB40[31] , 
        \wRegInB63[19] , \wBMid38[5] , \wAMid61[23] , \wRegInB16[30] , 
        \wRegInB35[18] , \wAMid83[3] , \wRegInB40[28] , \wAMid22[16] , 
        \wAMid57[26] , \wAMid74[17] , \ScanLink227[7] , \wBIn118[21] , 
        \wBIn58[21] , \ScanLink79[0] , \wRegInA39[4] , \wRegInA106[4] , 
        \ScanLink195[4] , \ScanLink77[30] , \ScanLink54[18] , \ScanLink21[28] , 
        \wAIn27[25] , \wBIn33[29] , \wBMid44[3] , \wBMid48[18] , \wAMid51[5] , 
        \ScanLink77[29] , \ScanLink21[31] , \wBMid96[5] , \wRegInB59[1] , 
        \wRegInB96[8] , \wRegInA15[22] , \wRegInB25[7] , \wRegInA45[2] , 
        \ScanLink129[27] , \ScanLink87[24] , \ScanLink149[23] , 
        \ScanLink18[9] , \ScanLink92[10] , \wBIn46[19] , \wAIn52[15] , 
        \wAIn70[8] , \wAMid100[19] , \wBMid119[28] , \wAMid123[28] , 
        \wRegInA60[12] , \wAMid123[31] , \wRegInA36[13] , \wRegInB93[14] , 
        \wBMid119[31] , \wRegInA43[23] , \wBIn125[28] , \wRegInA23[27] , 
        \wRegInA97[4] , \wRegInB38[8] , \wRegInA56[17] , \wRegInB86[20] , 
        \wRegInA75[26] , \ScanLink138[7] , \wBIn65[31] , \wRegInB68[15] , 
        \wRegInA94[7] , \wBIn33[30] , \wBMid47[0] , \wBIn65[28] , \wBMid88[9] , 
        \wBIn106[19] , \wBIn125[31] , \wAIn71[24] , \wAIn11[20] , \wAIn64[10] , 
        \wBIn16[8] , \wAIn32[11] , \wAIn47[21] , \ScanLink202[11] , 
        \ScanLink125[8] , \wBMid15[15] , \wBMid60[25] , \wRegInA89[8] , 
        \wRegInA46[1] , \wBMid36[24] , \wBMid95[6] , \ScanLink221[20] , 
        \ScanLink184[27] , \ScanLink254[10] , \wAMid6[24] , \wBMid20[7] , 
        \wBMid23[10] , \wBMid43[14] , \wBMid56[20] , \wRegInB26[4] , 
        \ScanLink234[14] , \ScanLink69[11] , \ScanLink191[13] , \wBMid75[11] , 
        \ScanLink241[24] , \ScanLink217[25] , \wAMid84[30] , \wAIn119[27] , 
        \wAMid84[29] , \wAMid116[6] , \wRegInA56[24] , \ScanLink190[9] , 
        \wRegInA23[14] , \wRegInB86[13] , \wBMid23[23] , \wAMid49[7] , 
        \wAMid54[8] , \wRegInA75[15] , \wRegInB1[3] , \wRegInA15[11] , 
        \wRegInA60[21] , \wRegInA21[6] , \wRegInA36[20] , \wRegInA43[10] , 
        \wRegInB93[5] , \wRegInB93[27] , \ScanLink61[2] , \ScanLink149[10] , 
        \ScanLink92[23] , \wRegInB118[19] , \wBMid56[13] , \wRegInB41[3] , 
        \ScanLink87[17] , \wRegInA103[9] , \ScanLink129[14] , 
        \ScanLink241[17] , \wBMid75[22] , \wRegInB2[0] , \ScanLink69[22] , 
        \ScanLink234[27] , \ScanLink191[20] , \wAIn119[14] , \wRegInA22[5] , 
        \ScanLink217[16] , \wBMid15[26] , \wBMid60[16] , \wRegInA115[31] , 
        \ScanLink202[22] , \ScanLink254[23] , \ScanLink221[9] , \wAMid2[26] , 
        \wAMid2[15] , \wAIn11[13] , \wBMid36[17] , \wBMid43[27] , 
        \wRegInA115[28] , \ScanLink221[13] , \ScanLink184[14] , \wRegInB42[0] , 
        \wBMid11[17] , \wBMid23[4] , \wAMid29[30] , \wAIn27[16] , 
        \wAMid29[29] , \wAIn64[23] , \wAMid98[2] , \wAIn32[22] , \wAIn47[12] , 
        \wAMid115[5] , \wRegInB68[26] , \wBMid27[12] , \wAIn52[26] , 
        \ScanLink62[1] , \wAIn71[17] , \wRegInB90[6] , \wBMid52[22] , 
        \ScanLink230[16] , \ScanLink195[11] , \wBMid71[13] , \wRegInB66[6] , 
        \ScanLink18[23] , \ScanLink245[26] , \ScanLink213[27] , 
        \ScanLink94[1] , \wBIn99[3] , \ScanLink206[13] , \wBMid64[27] , 
        \wAIn108[11] , \wBIn113[2] , \wAIn6[11] , \wAIn9[0] , \wBMid32[26] , 
        \ScanLink225[22] , \ScanLink180[25] , \ScanLink78[27] , 
        \wRegInA111[19] , \wBIn14[30] , \wAIn15[22] , \wBMid47[16] , 
        \ScanLink250[12] , \wAMid58[31] , \wAIn60[12] , \ScanLink218[0] , 
        \wAIn23[27] , \wAIn33[9] , \wAIn36[13] , \wAIn43[23] , \wAMid58[28] , 
        \ScanLink46[7] , \wAIn56[17] , \wRegInB19[27] , \wRegInB79[23] , 
        \ScanLink178[5] , \wAIn23[14] , \wBIn48[6] , \wAIn75[26] , 
        \wAMid80[18] , \wRegInA27[25] , \ScanLink45[4] , \wRegInA52[15] , 
        \wRegInB82[22] , \wRegInA11[20] , \wRegInA71[24] , \ScanLink4[8] , 
        \wRegInA32[11] , \wRegInA64[10] , \wRegInB97[16] , \wBIn55[9] , 
        \wRegInA47[21] , \wRegInB65[5] , \ScanLink138[11] , \ScanLink97[2] , 
        \ScanLink96[12] , \ScanLink83[26] , \wBIn110[1] , \ScanLink166[9] , 
        \ScanLink158[15] , \wBIn14[29] , \wBIn37[18] , \wBIn42[28] , 
        \wBIn102[31] , \wBIn121[19] , \wRegInB19[14] , \ScanLink22[3] , 
        \wAIn56[24] , \wAIn15[11] , \wBIn42[31] , \wAIn75[15] , \wBIn102[28] , 
        \wBIn61[19] , \wBMid63[6] , \wAMid17[9] , \wAIn36[20] , \wAIn60[21] , 
        \wAIn43[10] , \wAIn98[4] , \wRegInB79[10] , \wAIn108[22] , \wAIn6[22] , 
        \wBMid11[24] , \wBMid64[14] , \ScanLink206[20] , \wBMid8[21] , 
        \wBMid8[12] , \wAMid10[22] , \wAIn28[18] , \wBMid27[21] , 
        \wBMid32[15] , \wBMid47[25] , \ScanLink250[21] , \ScanLink225[11] , 
        \ScanLink180[16] , \ScanLink78[14] , \wBMid52[11] , \ScanLink245[15] , 
        \ScanLink18[10] , \wAIn49[1] , \wBMid71[20] , \wAIn103[9] , 
        \ScanLink230[25] , \ScanLink195[22] , \wRegInA62[7] , 
        \ScanLink213[14] , \ScanLink158[26] , \ScanLink83[15] , \wBMid60[5] , 
        \wAIn86[8] , \wAMid104[31] , \wRegInA11[13] , \wRegInA61[4] , 
        \wRegInA64[23] , \ScanLink138[22] , \ScanLink96[21] , \wRegInB112[9] , 
        \wAMid104[28] , \wRegInA32[22] , \wRegInA47[12] , \wRegInB97[25] , 
        \ScanLink21[0] , \wBMid124[8] , \wRegInA27[16] , \wRegInA52[26] , 
        \wRegInA71[17] , \wRegInB82[11] , \wRegInB67[28] , \wAMid33[13] , 
        \wAMid46[23] , \wBIn49[24] , \wRegInB12[18] , \wRegInA122[2] , 
        \wRegInB31[30] , \wRegInB44[19] , \wRegInB67[31] , \wAMid26[27] , 
        \wAMid65[12] , \wBIn109[24] , \wRegInB60[8] , \ScanLink203[1] , 
        \wRegInB31[29] , \wAMid70[26] , \wAIn28[8] , \wBIn29[20] , \wBIn50[4] , 
        \ScanLink163[4] , \wBMid39[19] , \wAMid53[17] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink40[9] , \ScanLink25[19] , \ScanLink1[5] , 
        \wAMid75[3] , \ScanLink73[18] , \wAIn35[7] , \wBIn82[2] , \wAIn36[4] , 
        \wBIn81[1] , \wBMid94[19] , \wBIn108[3] , \ScanLink218[18] , 
        \wRegInB3[13] , \wRegInB102[23] , \ScanLink88[19] , \wRegInB121[12] , 
        \ScanLink2[6] , \wBIn53[7] , \wAMid76[0] , \wAIn85[18] , 
        \wRegInA5[16] , \wRegInB117[17] , \ScanLink200[2] , \wBIn91[14] , 
        \wBMid116[15] , \wRegInA121[1] , \ScanLink1[12] , \wBIn84[20] , 
        \wBMid120[10] , \ScanLink160[7] , \wBMid103[21] , \wAIn116[30] , 
        \wRegInB19[3] , \wRegInB117[4] , \wAMid9[19] , \wAIn51[3] , 
        \wAIn116[29] , \wAIn118[8] , \wRegInA79[6] , \wAMid10[11] , 
        \wAMid11[7] , \wBMid65[8] , \wBMid121[5] , \wAMid26[14] , 
        \wAMid53[24] , \wAMid70[15] , \wRegInA81[29] , \wRegInA81[30] , 
        \ScanLink39[2] , \wBIn29[13] , \wAMid33[20] , \wBIn34[0] , 
        \wAMid46[10] , \wBIn49[17] , \wAIn105[7] , \ScanLink107[0] , 
        \wAIn83[5] , \wRegInA64[9] , \wAMid65[21] , \wBMid78[7] , 
        \wBIn109[17] , \wAMid12[4] , \wBIn37[3] , \wBIn84[13] , \wBMid120[23] , 
        \wRegInA59[19] , \wRegInB109[8] , \wBIn91[27] , \wBMid103[12] , 
        \wBMid116[26] , \ScanLink104[3] , \ScanLink1[21] , \wAIn80[6] , 
        \wAIn106[4] , \wBMid122[6] , \wRegInA5[25] , \wRegInB102[10] , 
        \wRegInB114[7] , \wRegInB117[24] , \ScanLink105[18] , 
        \ScanLink126[30] , \ScanLink170[28] , \wAIn14[5] , \wAIn52[0] , 
        \wRegInB3[20] , \wRegInB121[21] , \ScanLink126[29] , \wAMid91[14] , 
        \wRegInA60[28] , \ScanLink170[31] , \ScanLink153[19] , \wAMid100[23] , 
        \wBMid119[12] , \wAMid123[12] , \wRegInA15[18] , \wRegInA36[30] , 
        \wRegInA36[29] , \wRegInA43[19] , \wRegInA60[31] , \wAMid115[17] , 
        \ScanLink190[0] , \wAMid54[1] , \wAMid84[20] , \wBIn71[6] , 
        \wRegInA103[0] , \ScanLink222[3] , \ScanLink142[6] , \wAMid86[7] , 
        \ScanLink149[19] , \wRegInB118[10] , \wAIn2[29] , \wRegInA100[3] , 
        \wBIn3[8] , \wBIn4[27] , \wBIn5[6] , \wBIn6[5] , \wBMid7[15] , 
        \wBIn72[5] , \wAMid85[4] , \wRegInB42[9] , \ScanLink221[0] , 
        \wRegInA100[15] , \wRegInA115[21] , \ScanLink191[29] , \wRegInB2[9] , 
        \wBIn10[22] , \wBIn33[13] , \wAMid108[3] , \wRegInA123[24] , 
        \ScanLink141[5] , \ScanLink191[30] , \wBIn46[23] , \wAMid49[24] , 
        \wBIn125[12] , \ScanLink62[8] , \wBIn15[2] , \wAIn17[6] , \wBIn26[27] , 
        \wAMid57[2] , \wBIn65[12] , \wBIn106[23] , \wBIn70[26] , \wBIn113[17] , 
        \ScanLink193[3] , \wAMid29[20] , \wBIn53[17] , \wBMid59[5] , 
        \wRegInB118[23] , \ScanLink246[7] , \ScanLink18[0] , \ScanLink92[19] , 
        \wAIn124[5] , \wBMid7[26] , \wBIn10[11] , \wAIn11[30] , \wAIn11[29] , 
        \wAMid30[5] , \wAMid84[13] , \wAMid115[24] , \ScanLink126[2] , 
        \wRegInB86[30] , \wRegInB86[29] , \wBMid100[7] , \wRegInB38[1] , 
        \wAMid123[21] , \wAIn47[31] , \wAIn70[1] , \wAMid91[27] , 
        \wAMid100[10] , \wBMid119[21] , \wRegInA58[4] , \wBIn70[15] , 
        \wAIn64[19] , \wBIn113[24] , \wBIn26[14] , \wAIn47[28] , \wBIn53[24] , 
        \wAMid29[13] , \wAIn32[18] , \wBIn33[20] , \wBIn46[10] , \wAMid49[17] , 
        \wBIn125[21] , \wAIn73[2] , \wAMid33[6] , \wBMid47[9] , \wBMid88[0] , 
        \wBIn106[10] , \wBIn65[21] , \wBMid103[4] , \wBMid23[19] , 
        \ScanLink69[18] , \wBMid56[29] , \wRegInA100[26] , \ScanLink245[4] , 
        \wBMid75[18] , \wRegInA123[17] , \wBMid56[30] , \ScanLink221[30] , 
        \wAMid8[7] , \wBIn16[1] , \wAIn127[6] , \ScanLink202[18] , 
        \ScanLink125[1] , \wBMid85[15] , \wRegInA46[8] , \wRegInA89[1] , 
        \wRegInA115[12] , \ScanLink221[29] , \ScanLink254[19] , 
        \wRegInA118[1] , \ScanLink137[16] , \ScanLink67[5] , \ScanLink142[26] , 
        \ScanLink239[2] , \ScanLink114[27] , \ScanLink99[15] , \wBIn4[14] , 
        \wAIn9[16] , \wAIn11[8] , \wBMid26[0] , \wRegInB95[2] , 
        \ScanLink161[17] , \ScanLink101[13] , \wBMid28[15] , \wAIn39[14] , 
        \wBIn58[31] , \wBIn77[8] , \wBIn80[18] , \wBMid90[21] , 
        \ScanLink174[23] , \ScanLink159[7] , \ScanLink122[22] , \wAMid110[1] , 
        \wBMid124[28] , \wRegInA28[22] , \ScanLink157[12] , \wAMid80[9] , 
        \wAIn94[14] , \wBMid107[19] , \wRegInB47[4] , \wBMid124[31] , 
        \wAIn81[20] , \wRegInB7[4] , \wRegInB98[11] , \ScanLink144[8] , 
        \wRegInA27[1] , \wRegInA48[26] , \wBIn58[28] , \wBIn118[28] , 
        \wRegInA85[22] , \wRegInB20[25] , \wRegInB44[7] , \wRegInB55[15] , 
        \wBIn118[31] , \ScanLink79[9] , \wAIn59[10] , \wRegInB16[20] , 
        \wRegInB76[24] , \ScanLink188[2] , \wRegInB4[7] , \wRegInA24[2] , 
        \wRegInB35[11] , \wRegInB63[10] , \wRegInB40[21] , \wRegInA90[16] , 
        \wBIn69[4] , \wAIn112[22] , \wRegInB59[8] , \wRegInB96[1] , 
        \ScanLink62[14] , \ScanLink17[24] , \ScanLink64[6] , \ScanLink41[25] , 
        \ScanLink34[15] , \wAIn107[16] , \ScanLink209[14] , \ScanLink54[11] , 
        \wAMid113[2] , \wBMid25[3] , \ScanLink21[21] , \wAIn124[27] , 
        \ScanLink77[20] , \wBMid9[0] , \wBMid48[11] , \wAIn81[13] , 
        \ScanLink240[9] , \ScanLink5[19] , \wBMid85[26] , \wBMid90[12] , 
        \wBMid90[2] , \wAIn94[27] , \wRegInB23[0] , \wRegInA28[11] , 
        \wRegInA43[5] , \wRegInA48[15] , \wRegInB98[22] , \wRegInB7[18] , 
        \wRegInB106[31] , \wRegInB106[28] , \ScanLink174[10] , 
        \ScanLink101[20] , \ScanLink157[21] , \wRegInB125[19] , 
        \ScanLink122[11] , \ScanLink142[15] , \wRegInA91[3] , 
        \ScanLink137[25] , \wAIn9[25] , \wBMid42[4] , \wBMid106[9] , 
        \ScanLink99[26] , \wAIn107[25] , \ScanLink161[24] , \ScanLink114[14] , 
        \ScanLink209[27] , \ScanLink21[12] , \ScanLink54[22] , \wAMid14[30] , 
        \wBMid28[26] , \wBMid41[7] , \wBMid48[22] , \wAIn124[14] , 
        \ScanLink77[13] , \ScanLink17[17] , \wAMid35[8] , \ScanLink62[27] , 
        \wAMid37[18] , \wAIn112[11] , \ScanLink34[26] , \wRegInB63[23] , 
        \wRegInA92[0] , \ScanLink41[16] , \wAMid14[29] , \wAMid42[28] , 
        \wAIn59[23] , \wRegInB16[13] , \wRegInB40[12] , \wAMid28[7] , 
        \wAMid42[31] , \wAMid61[19] , \wRegInB20[3] , \wRegInB35[22] , 
        \wRegInA90[25] , \wBMid93[1] , \wBMid118[5] , \wRegInB55[26] , 
        \wAIn39[27] , \wRegInB20[16] , \wRegInA85[11] , \wBMid8[31] , 
        \wAMid9[10] , \wBIn29[6] , \wAIn68[3] , \wAIn121[8] , \wRegInB76[17] , 
        \wRegInA40[6] , \wAIn103[14] , \wAIn118[1] , \ScanLink50[13] , 
        \wBMid39[23] , \wBMid65[1] , \ScanLink25[23] , \ScanLink73[22] , 
        \wAIn120[25] , \ScanLink66[16] , \wBMid8[28] , \wBMid59[27] , 
        \ScanLink218[22] , \ScanLink45[27] , \ScanLink13[26] , 
        \ScanLink30[17] , \ScanLink24[4] , \wAMid10[18] , \wAIn28[22] , 
        \wBIn34[9] , \wAIn116[20] , \wRegInB12[22] , \wAMid46[19] , 
        \wAMid65[31] , \wRegInA64[0] , \wRegInB67[12] , \ScanLink107[9] , 
        \wAMid33[29] , \wAMid65[28] , \wRegInB31[13] , \wRegInA94[14] , 
        \wRegInB44[23] , \wAMid33[30] , \wAIn48[26] , \wRegInB24[27] , 
        \wRegInA81[20] , \wRegInB51[17] , \wAIn52[9] , \wBMid66[2] , 
        \wAIn85[22] , \wRegInB72[26] , \wAIn90[16] , \wRegInA39[14] , 
        \ScanLink1[28] , \wRegInA59[10] , \wRegInA67[3] , \ScanLink1[31] , 
        \wRegInB89[27] , \wRegInB102[19] , \wRegInB109[1] , \wRegInB121[31] , 
        \ScanLink105[11] , \wBMid94[23] , \wRegInB3[30] , \wRegInB121[28] , 
        \ScanLink170[21] , \ScanLink126[20] , \ScanLink119[5] , 
        \ScanLink88[23] , \wRegInB3[29] , \ScanLink153[10] , \wBMid81[17] , 
        \ScanLink146[24] , \ScanLink133[14] , \ScanLink27[7] , 
        \ScanLink110[25] , \wBIn0[16] , \wAMid9[23] , \wAIn28[11] , 
        \wAIn28[1] , \wBIn29[30] , \ScanLink165[15] , \wBIn29[29] , 
        \wAMid68[5] , \wRegInB51[24] , \wRegInB24[14] , \wRegInA81[13] , 
        \wAIn48[15] , \wRegInB72[15] , \wBIn115[5] , \wRegInB67[21] , 
        \ScanLink92[6] , \wBMid59[14] , \wRegInB12[11] , \wRegInB31[20] , 
        \wRegInB44[10] , \wRegInB60[1] , \ScanLink203[8] , \wRegInA94[27] , 
        \wAIn103[27] , \wAIn116[13] , \ScanLink66[25] , \ScanLink13[15] , 
        \ScanLink30[24] , \ScanLink218[11] , \ScanLink45[14] , \ScanLink40[0] , 
        \ScanLink25[10] , \wBMid39[10] , \wAIn120[16] , \ScanLink50[20] , 
        \ScanLink73[11] , \wBIn81[8] , \wBMid81[24] , \ScanLink146[17] , 
        \ScanLink133[27] , \wBMid3[24] , \wBMid3[17] , \wBIn14[20] , 
        \wAIn15[18] , \wAIn36[30] , \wAMid76[9] , \ScanLink165[26] , 
        \wBIn84[30] , \wBMid94[10] , \ScanLink170[12] , \ScanLink110[16] , 
        \ScanLink153[23] , \ScanLink105[22] , \ScanLink88[10] , 
        \ScanLink126[13] , \ScanLink43[3] , \wBMid103[31] , \wBMid120[19] , 
        \wBIn84[29] , \wAIn90[25] , \wBIn116[6] , \wRegInA59[23] , 
        \wRegInB89[14] , \wBMid103[28] , \wAIn85[11] , \wRegInA39[27] , 
        \wRegInB63[2] , \ScanLink91[5] , \wRegInA121[8] , \wAMid17[0] , 
        \wAIn60[28] , \wBIn22[25] , \wAIn36[29] , \wBIn74[24] , \wBIn117[15] , 
        \wBIn37[11] , \wAMid38[16] , \wAIn43[19] , \wBIn57[15] , 
        \wRegInB79[19] , \wAMid58[12] , \wAIn60[31] , \wAIn57[4] , 
        \wBIn42[21] , \wBIn121[10] , \wBMid27[28] , \wBMid52[18] , 
        \wBIn61[10] , \wBIn102[21] , \wRegInB111[3] , \ScanLink18[19] , 
        \wBMid71[30] , \wRegInA104[17] , \wBIn32[7] , \wAIn6[18] , \wAIn9[9] , 
        \wAMid14[3] , \wBMid27[31] , \wBMid71[29] , \wAIn85[2] , \wAIn103[0] , 
        \ScanLink101[7] , \wRegInA127[26] , \wBIn31[4] , \wRegInA111[23] , 
        \ScanLink250[31] , \ScanLink250[28] , \ScanLink206[29] , 
        \ScanLink225[18] , \ScanLink206[30] , \ScanLink102[4] , 
        \ScanLink96[31] , \wAIn49[8] , \wAIn100[3] , \wAIn54[7] , \wAIn86[1] , 
        \wAMid111[15] , \wRegInB8[16] , \wRegInB109[26] , \ScanLink96[28] , 
        \wAMid80[22] , \wBMid108[24] , \wRegInB82[18] , \wBMid124[1] , 
        \wBIn56[3] , \wAMid95[16] , \wAMid104[21] , \wRegInB112[0] , 
        \ScanLink21[9] , \ScanLink165[3] , \wAIn108[18] , \wRegInA111[10] , 
        \wRegInA104[24] , \wRegInA127[15] , \ScanLink205[6] , 
        \ScanLink195[18] , \ScanLink94[8] , \wBIn14[13] , \wAIn33[0] , 
        \wBIn42[12] , \wBIn84[5] , \wBIn121[23] , \wRegInA124[5] , 
        \wBIn37[22] , \wAMid38[25] , \wBIn61[23] , \wBIn102[12] , \wBIn22[16] , 
        \wBIn57[26] , \wAMid73[4] , \wBIn74[17] , \wBIn117[26] , 
        \ScanLink218[9] , \ScanLink7[2] , \wAMid58[21] , \ScanLink89[7] , 
        \wAIn30[3] , \wAMid70[7] , \wRegInA11[29] , \wRegInA47[31] , 
        \wBIn87[6] , \wAMid95[25] , \wRegInA8[3] , \wRegInA64[19] , 
        \wAMid104[12] , \wRegInA11[30] , \wRegInA32[18] , \wRegInA18[6] , 
        \wRegInA47[28] , \wBMid108[17] , \wAMid111[26] , \wAIn1[1] , 
        \wBMid19[7] , \wAMid80[11] , \wRegInB78[3] , \ScanLink4[1] , 
        \wBIn43[4] , \wBIn55[0] , \wRegInB109[15] , \wBIn85[23] , \wBIn110[8] , 
        \wRegInB8[25] , \ScanLink166[0] , \wRegInA127[6] , \ScanLink138[18] , 
        \ScanLink58[2] , \ScanLink206[5] , \wBMid102[22] , \wRegInA3[8] , 
        \wRegInA58[30] , \wBIn90[17] , \wBMid117[16] , \wBMid121[13] , 
        \wRegInA58[29] , \ScanLink210[1] , \ScanLink170[4] , \wRegInB73[8] , 
        \ScanLink0[11] , \wAIn2[2] , \wBMid9[11] , \wAIn26[7] , \wAMid66[3] , 
        \wBIn91[2] , \wRegInA4[15] , \wRegInB116[14] , \wRegInB2[10] , 
        \wRegInB120[11] , \ScanLink152[29] , \ScanLink53[9] , 
        \ScanLink127[19] , \ScanLink104[31] , \wRegInB103[20] , 
        \ScanLink171[18] , \ScanLink152[30] , \ScanLink104[28] , \wAIn25[4] , 
        \wBIn92[1] , \wAIn117[19] , \wBIn118[0] , \wAMid8[30] , \wAMid65[0] , 
        \wAMid8[29] , \wAMid27[24] , \wBIn28[23] , \wBIn40[7] , 
        \ScanLink173[7] , \wAMid52[14] , \wAMid71[25] , \wRegInA80[19] , 
        \wAMid11[21] , \wAMid11[12] , \wBIn27[0] , \wAMid32[10] , 
        \wAMid64[11] , \wBIn108[27] , \ScanLink213[2] , \wAIn42[3] , 
        \wAMid47[20] , \wBIn48[27] , \wBMid95[29] , \wRegInB2[23] , 
        \wRegInB120[22] , \wBMid76[8] , \wBMid95[30] , \wRegInB103[13] , 
        \ScanLink89[30] , \wRegInA4[26] , \ScanLink89[29] , \wRegInB104[4] , 
        \wRegInB116[27] , \ScanLink114[0] , \wAMid64[22] , \wBMid68[4] , 
        \wAIn84[31] , \wAIn90[5] , \wAIn116[7] , \wRegInA77[9] , \wAIn84[28] , 
        \wBIn90[24] , \wBMid117[25] , \ScanLink0[22] , \wBIn85[10] , 
        \wBMid102[11] , \wBIn108[14] , \wBMid121[20] , \wRegInB30[19] , 
        \wRegInB13[31] , \wRegInB45[29] , \wBIn24[3] , \wAIn29[31] , 
        \wAMid27[17] , \wAIn29[28] , \wAMid32[23] , \wAMid47[13] , 
        \wBIn48[14] , \wAIn115[4] , \wRegInB13[28] , \ScanLink117[3] , 
        \wAIn93[6] , \wRegInB45[30] , \wRegInB66[18] , \wAMid52[27] , 
        \ScanLink29[1] , \wBIn28[10] , \wAMid71[16] , \wRegInA0[24] , 
        \wRegInA0[17] , \wBMid1[8] , \wAIn3[10] , \wAMid3[25] , \wAMid3[16] , 
        \wAIn7[12] , \wBMid9[22] , \wBMid38[30] , \wBMid38[29] , 
        \ScanLink72[28] , \ScanLink24[30] , \wAIn41[0] , \wRegInA69[5] , 
        \ScanLink72[31] , \ScanLink51[19] , \ScanLink219[28] , 
        \ScanLink24[29] , \wAIn14[21] , \wBIn15[19] , \wBMid14[2] , 
        \wAIn20[9] , \wBIn58[5] , \wBIn100[2] , \wRegInA15[3] , 
        \wRegInB107[7] , \ScanLink219[31] , \ScanLink159[16] , \wRegInA5[6] , 
        \ScanLink82[25] , \wRegInA33[12] , \wRegInB75[6] , \ScanLink97[11] , 
        \ScanLink139[12] , \ScanLink87[1] , \ScanLink9[4] , \ScanLink48[8] , 
        \wRegInB96[15] , \wAMid105[18] , \wAMid126[30] , \wRegInA46[22] , 
        \wAMid122[3] , \wBMid17[1] , \wBIn60[29] , \wBIn103[18] , 
        \wAMid126[29] , \wRegInA10[23] , \wRegInA26[26] , \wRegInA65[13] , 
        \wRegInB68[9] , \wRegInA70[27] , \wRegInB83[21] , \ScanLink55[7] , 
        \wRegInA53[16] , \wBIn120[30] , \wAIn74[25] , \wBIn36[31] , 
        \wAIn22[24] , \wBIn36[28] , \wBIn43[18] , \wAIn57[14] , \wBIn60[30] , 
        \wBIn120[29] , \wRegInB18[24] , \ScanLink168[6] , \wAMid121[0] , 
        \wAIn37[10] , \wAIn42[20] , \ScanLink56[4] , \wAIn61[11] , 
        \wRegInB78[20] , \ScanLink208[3] , \wBMid33[25] , \ScanLink224[21] , 
        \ScanLink181[26] , \ScanLink79[24] , \wBMid10[14] , \wBIn46[9] , 
        \wBMid46[15] , \wRegInA6[5] , \ScanLink251[11] , \wBIn89[0] , 
        \ScanLink207[10] , \ScanLink175[9] , \wBMid65[24] , \wAIn109[12] , 
        \wRegInA16[0] , \wBIn103[1] , \wAIn7[21] , \wAMid19[6] , \wBMid26[11] , 
        \wBMid70[10] , \ScanLink212[24] , \ScanLink84[2] , \wBMid53[21] , 
        \ScanLink231[15] , \ScanLink194[12] , \wBMid70[6] , \wAMid81[28] , 
        \wRegInB76[5] , \ScanLink19[20] , \ScanLink244[25] , \wRegInA70[14] , 
        \wAMid81[31] , \wRegInA10[10] , \wRegInA26[15] , \wRegInA53[25] , 
        \wRegInB83[12] , \wRegInA33[21] , \wRegInA46[11] , \ScanLink31[3] , 
        \wRegInA65[20] , \wRegInB96[26] , \ScanLink97[22] , \wBMid26[22] , 
        \wBMid53[12] , \wAIn59[2] , \wAIn110[9] , \wBMid70[23] , 
        \wRegInB11[2] , \wRegInA71[7] , \ScanLink159[25] , \ScanLink139[21] , 
        \ScanLink82[16] , \wAIn95[8] , \wRegInA72[4] , \ScanLink212[17] , 
        \ScanLink244[16] , \ScanLink19[13] , \ScanLink231[26] , 
        \ScanLink194[21] , \wBMid33[16] , \wBMid46[26] , \ScanLink251[22] , 
        \wRegInB12[1] , \wRegInA110[29] , \ScanLink224[12] , \ScanLink181[15] , 
        \ScanLink79[17] , \wAIn109[21] , \wBMid10[27] , \wBMid65[17] , 
        \ScanLink207[23] , \wAIn14[12] , \wAIn37[23] , \wRegInA110[30] , 
        \wAIn42[13] , \wAIn88[7] , \wRegInB78[13] , \wAMid59[18] , 
        \wBMid73[5] , \wAIn22[17] , \wAIn61[22] , \wAIn74[16] , 
        \wRegInB101[9] , \wBMid22[13] , \wAIn57[27] , \wRegInB18[17] , 
        \ScanLink32[0] , \wBMid74[12] , \ScanLink216[26] , \wAIn118[24] , 
        \wBMid37[27] , \wBMid57[23] , \wRegInB36[7] , \ScanLink235[17] , 
        \ScanLink190[10] , \ScanLink68[12] , \wBMid85[5] , \ScanLink240[27] , 
        \ScanLink220[23] , \ScanLink185[24] , \wRegInA114[18] , 
        \ScanLink255[13] , \wAMid7[14] , \wBMid14[16] , \wBMid42[17] , 
        \ScanLink203[12] , \wBMid61[26] , \wRegInA56[2] , \wAIn10[23] , 
        \wAMid28[19] , \wAIn33[12] , \wAIn46[22] , \ScanLink16[6] , 
        \wAIn65[13] , \ScanLink248[1] , \wAIn3[23] , \wBIn8[3] , \wBMid57[3] , 
        \wAIn70[27] , \wAIn10[10] , \wBIn11[31] , \wBIn11[28] , \wBIn18[7] , 
        \wAIn26[26] , \wAIn53[16] , \ScanLink128[4] , \wAIn63[8] , 
        \wRegInB69[16] , \wRegInA84[4] , \wAMid85[19] , \wRegInA22[24] , 
        \wRegInA74[25] , \wRegInB87[23] , \ScanLink15[5] , \wRegInA37[10] , 
        \wRegInA57[14] , \wRegInB92[17] , \wBMid54[0] , \wRegInA14[21] , 
        \wRegInA42[20] , \wRegInA87[7] , \wBMid86[6] , \wRegInB35[4] , 
        \wRegInA61[11] , \wRegInB119[29] , \ScanLink93[13] , \wRegInA55[1] , 
        \wRegInB119[30] , \ScanLink148[20] , \ScanLink136[8] , 
        \ScanLink128[24] , \ScanLink86[27] , \wBIn47[30] , \wBIn107[29] , 
        \wRegInB80[5] , \wBIn64[18] , \wAIn70[14] , \wRegInB69[25] , 
        \wAIn26[15] , \wBIn32[19] , \ScanLink72[2] , \wAIn33[21] , 
        \wBIn47[29] , \wBIn107[30] , \wBIn124[18] , \wAIn53[25] , 
        \ScanLink183[9] , \wAIn46[11] , \wAMid105[6] , \wBMid33[7] , 
        \wAMid47[8] , \wAIn65[20] , \wAMid88[1] , \ScanLink255[20] , 
        \wBMid4[5] , \wAMid7[27] , \wBMid37[14] , \wBMid42[24] , 
        \ScanLink220[10] , \ScanLink185[17] , \wRegInB52[3] , \wBMid7[6] , 
        \wBMid14[25] , \wBMid61[15] , \wRegInA110[9] , \ScanLink203[21] , 
        \wAMid15[23] , \wAIn19[0] , \wBMid22[20] , \wBMid57[10] , 
        \wBMid74[21] , \wAIn118[17] , \wAMid118[9] , \wBIn127[7] , 
        \wRegInA32[6] , \ScanLink216[15] , \ScanLink240[14] , \wAMid59[4] , 
        \wRegInB51[0] , \ScanLink235[24] , \ScanLink190[23] , \ScanLink68[21] , 
        \ScanLink232[9] , \ScanLink128[17] , \ScanLink86[14] , 
        \ScanLink93[20] , \ScanLink148[13] , \wBMid30[4] , \wAMid101[30] , 
        \wAMid101[29] , \wBIn124[4] , \wRegInA31[5] , \wRegInA37[23] , 
        \wRegInA42[13] , \ScanLink71[1] , \wRegInB92[24] , \wBMid118[18] , 
        \wRegInA61[22] , \wRegInA14[12] , \wAMid122[18] , \wRegInB83[6] , 
        \wAMid106[5] , \wRegInA57[27] , \wRegInA74[16] , \wRegInA22[17] , 
        \wRegInB87[10] , \wRegInB41[18] , \wRegInB62[30] , \wAMid23[26] , 
        \wAMid36[12] , \wBIn39[15] , \wAIn58[30] , \wRegInB30[9] , 
        \wRegInB34[28] , \ScanLink253[0] , \wAMid60[13] , \wRegInB62[29] , 
        \wAMid43[22] , \wRegInB17[19] , \wRegInB34[31] , \wAIn58[29] , 
        \wBMid49[28] , \wAMid56[16] , \wAIn78[9] , \ScanLink133[5] , 
        \wBIn59[11] , \wAMid75[27] , \wBIn119[11] , \wRegInB123[1] , 
        \wAMid25[2] , \wBMid49[31] , \ScanLink76[19] , \ScanLink55[31] , 
        \ScanLink10[8] , \wAIn65[6] , \ScanLink55[28] , \ScanLink20[18] , 
        \wBMid115[0] , \wBMid91[18] , \wRegInB124[13] , \wRegInB6[12] , 
        \wAMid26[1] , \wBMid116[3] , \wRegInB107[22] , \wRegInB120[2] , 
        \wAMid5[2] , \wAMid6[1] , \wAMid23[15] , \wBMid35[9] , \wAIn66[5] , 
        \wRegInA81[9] , \wRegInB112[16] , \wAIn80[19] , \wRegInB99[28] , 
        \ScanLink250[3] , \wBIn81[21] , \wBIn94[15] , \ScanLink4[13] , 
        \wBMid106[20] , \wBMid113[14] , \wRegInB99[31] , \wBMid80[8] , 
        \wAIn113[31] , \wAIn113[28] , \wBMid125[11] , \ScanLink130[6] , 
        \wRegInB49[2] , \wAMid41[6] , \wAMid56[25] , \wAMid103[8] , 
        \wRegInB9[2] , \wRegInA29[7] , \ScanLink185[7] , \wBIn59[22] , 
        \wRegInA84[31] , \ScanLink69[3] , \wAMid75[14] , \wRegInA116[7] , 
        \ScanLink237[4] , \wAMid15[10] , \wBMid28[6] , \wBIn119[22] , 
        \wRegInA84[28] , \wAMid60[20] , \wAMid36[21] , \wBIn39[26] , 
        \wAMid43[11] , \wBIn64[1] , \wAMid93[0] , \ScanLink198[8] , 
        \ScanLink157[1] , \wBIn121[9] , \wRegInA34[8] , \wBIn67[2] , 
        \wBIn81[12] , \wBMid106[13] , \wRegInA29[31] , \ScanLink234[7] , 
        \wBMid125[22] , \wRegInA29[28] , \wRegInB98[7] , \wRegInA115[4] , 
        \ScanLink154[2] , \wAMid90[3] , \wBIn94[26] , \ScanLink4[20] , 
        \wBMid113[27] , \wAIn1[25] , \wBMid0[31] , \wBMid0[28] , \wBMid0[5] , 
        \wAMid42[5] , \wRegInB6[21] , \wRegInB85[8] , \wRegInB112[25] , 
        \ScanLink229[8] , \wRegInB124[20] , \ScanLink123[28] , 
        \ScanLink186[4] , \wRegInB107[11] , \ScanLink175[30] , 
        \ScanLink156[18] , \ScanLink175[29] , \ScanLink123[31] , 
        \ScanLink100[19] , \wRegInA6[20] , \wRegInB114[21] , \ScanLink113[29] , 
        \wAMid1[23] , \wAMid1[2] , \wBIn3[30] , \wBIn3[29] , \wRegInB124[2] , 
        \ScanLink166[19] , \ScanLink145[31] , \ScanLink145[28] , 
        \ScanLink130[18] , \ScanLink113[30] , \wBMid3[6] , \wAMid13[14] , 
        \wAMid22[1] , \wAIn62[5] , \wRegInB0[25] , \wRegInB122[24] , 
        \ScanLink129[9] , \wBMid99[7] , \wBMid112[3] , \wRegInA85[9] , 
        \wRegInB101[15] , \wAMid25[11] , \wAMid50[21] , \wBMid84[8] , 
        \wBIn87[16] , \wBMid100[17] , \ScanLink254[3] , \wAMid88[11] , 
        \wAMid119[26] , \wBMid123[26] , \wRegInA19[30] , \wRegInA19[29] , 
        \wRegInA98[6] , \ScanLink134[6] , \wBIn92[22] , \wBMid115[23] , 
        \ScanLink2[24] , \wBMid48[2] , \wAMid66[24] , \wAMid73[10] , 
        \wRegInB34[9] , \wBIn69[23] , \wRegInA97[18] , \wAMid30[25] , 
        \wAMid45[15] , \ScanLink137[5] , \wRegInB127[1] , \wRegInB29[6] , 
        \ScanLink14[8] , \wAMid21[2] , \wBMid111[0] , \wRegInA119[10] , 
        \wAIn61[6] , \wAIn123[29] , \wBIn92[11] , \wAIn100[18] , \wAIn123[30] , 
        \wRegInA49[3] , \wRegInA111[4] , \wBMid115[10] , \ScanLink2[17] , 
        \wAMid2[1] , \wAMid13[27] , \wBMid31[9] , \wAMid46[5] , \wBIn63[2] , 
        \wBIn87[25] , \wAIn93[29] , \ScanLink230[7] , \wBMid100[24] , 
        \wAMid88[22] , \wAMid94[3] , \ScanLink150[2] , \wAIn93[30] , 
        \wAMid119[15] , \wAMid119[4] , \wBMid123[15] , \wRegInB0[16] , 
        \wRegInA6[13] , \wRegInB81[8] , \wRegInB122[17] , \wRegInB101[26] , 
        \wRegInB114[12] , \wBMid79[29] , \wBMid82[31] , \wBMid82[28] , 
        \ScanLink182[4] , \wRegInA119[23] , \ScanLink181[7] , \wAMid107[8] , 
        \ScanLink46[18] , \ScanLink33[28] , \ScanLink65[30] , \wAMid45[6] , 
        \wBMid79[30] , \ScanLink10[19] , \ScanLink33[31] , \ScanLink233[4] , 
        \ScanLink65[29] , \wAIn5[27] , \wBIn8[16] , \wAMid25[22] , 
        \wAMid30[16] , \wAMid66[17] , \wBIn69[10] , \wAMid45[26] , \wBIn60[1] , 
        \wRegInA112[7] , \wRegInB52[31] , \wRegInB71[19] , \ScanLink153[1] , 
        \wAMid50[12] , \wAIn68[31] , \wBIn125[9] , \wRegInA30[8] , 
        \wBMid50[0] , \wAMid58[9] , \wRegInB52[28] , \wAIn68[28] , 
        \wRegInB27[18] , \wAMid73[23] , \wAMid97[0] , \wRegInA12[16] , 
        \wRegInA31[27] , \wRegInA44[17] , \ScanLink11[5] , \wRegInA67[26] , 
        \wRegInB94[20] , \wRegInA72[12] , \wAIn98[25] , \wBMid109[2] , 
        \wAMid112[19] , \wRegInA24[13] , \wRegInA51[23] , \wRegInB81[14] , 
        \wRegInB31[4] , \wRegInA83[7] , \ScanLink178[12] , \ScanLink80[10] , 
        \wAMid39[0] , \wBMid82[6] , \ScanLink95[24] , \wBMid44[20] , 
        \wAIn79[4] , \wBMid89[24] , \wRegInA51[1] , \ScanLink132[8] , 
        \ScanLink118[16] , \wBMid31[10] , \wRegInB32[7] , \ScanLink253[24] , 
        \wBMid67[11] , \ScanLink226[14] , \ScanLink183[13] , \wBMid5[8] , 
        \wBMid12[21] , \wBMid24[24] , \wBMid51[14] , \wBMid72[25] , 
        \ScanLink205[25] , \ScanLink58[20] , \ScanLink38[24] , \wBMid81[5] , 
        \wRegInA52[2] , \ScanLink210[11] , \ScanLink246[10] , 
        \ScanLink233[20] , \ScanLink196[27] , \wAIn76[10] , \wRegInB39[20] , 
        \wBIn8[25] , \wAIn16[14] , \wAIn20[11] , \ScanLink12[6] , \wBIn21[30] , 
        \wBIn21[29] , \wAIn35[25] , \wAIn55[21] , \wAIn40[15] , \wBIn54[19] , 
        \wAIn67[8] , \wRegInA80[4] , \wBIn77[31] , \wBMid53[3] , 
        \wRegInB59[24] , \wAIn63[24] , \wBIn114[19] , \wRegInA89[13] , 
        \wBIn77[28] , \wRegInB55[0] , \ScanLink236[9] , \ScanLink118[25] , 
        \ScanLink95[17] , \wAIn16[27] , \wAIn35[16] , \wBMid34[4] , 
        \wBIn78[3] , \wBMid89[17] , \wAIn98[16] , \wBIn120[4] , 
        \ScanLink199[5] , \wRegInA35[5] , \wRegInA72[21] , \ScanLink178[21] , 
        \ScanLink80[23] , \wRegInA24[20] , \wRegInB81[27] , \wRegInB87[6] , 
        \wRegInA51[10] , \ScanLink75[1] , \wAMid96[30] , \wAMid102[5] , 
        \wRegInA31[14] , \wRegInB94[13] , \wRegInA44[24] , \ScanLink9[31] , 
        \wAIn40[26] , \wAMid96[29] , \wRegInA12[25] , \wRegInA67[15] , 
        \ScanLink9[28] , \wRegInA109[6] , \ScanLink76[2] , \wAIn63[17] , 
        \wRegInA89[20] , \ScanLink228[5] , \wRegInB59[17] , \wRegInB84[5] , 
        \wAMid18[18] , \wBMid37[7] , \wAIn76[23] , \wRegInB39[13] , 
        \wAIn20[22] , \wAMid43[8] , \wAIn55[12] , \ScanLink187[9] , 
        \ScanLink148[0] , \wBMid72[16] , \wAMid101[6] , \wRegInA107[31] , 
        \wRegInA124[19] , \ScanLink210[22] , \wRegInA114[9] , \ScanLink38[17] , 
        \wBMid24[17] , \ScanLink233[13] , \ScanLink196[14] , \wRegInA107[28] , 
        \ScanLink246[23] , \wAMid1[10] , \wAIn5[14] , \wBMid31[23] , 
        \wBMid51[27] , \wRegInB56[3] , \wBMid44[13] , \ScanLink226[27] , 
        \ScanLink183[20] , \wBMid12[12] , \ScanLink253[17] , \wBIn123[7] , 
        \ScanLink205[16] , \ScanLink58[13] , \wBMid4[19] , \wAIn12[16] , 
        \wAIn31[27] , \wBMid67[22] , \wRegInA36[6] , \wAIn44[17] , 
        \wAMid125[0] , \wBMid13[1] , \wAIn24[13] , \wAIn67[26] , 
        \wRegInB28[16] , \wAMid69[19] , \wRegInB48[12] , \wAIn72[12] , 
        \wRegInA98[25] , \ScanLink52[4] , \wBIn42[9] , \wAIn51[23] , 
        \ScanLink171[9] , \wBMid20[26] , \wBMid55[16] , \wBMid76[27] , 
        \wBIn107[1] , \wRegInA12[0] , \ScanLink214[13] , \ScanLink49[16] , 
        \wRegInA120[28] , \ScanLink242[12] , \wRegInA2[5] , \ScanLink237[22] , 
        \ScanLink192[25] , \wRegInA103[19] , \wBMid40[22] , \wRegInA120[31] , 
        \wAIn1[16] , \wAMid5[21] , \wBMid35[12] , \wBMid63[13] , 
        \wRegInB72[5] , \ScanLink222[16] , \ScanLink187[11] , \ScanLink29[12] , 
        \wBMid10[2] , \wBMid16[23] , \ScanLink80[2] , \wAIn39[6] , 
        \wAMid79[2] , \ScanLink201[27] , \ScanLink169[24] , \ScanLink91[26] , 
        \wBIn104[2] , \wRegInA1[6] , \wRegInA11[3] , \wBMid98[12] , 
        \ScanLink83[1] , \wRegInB71[6] , \ScanLink84[12] , \ScanLink109[20] , 
        \wAIn24[9] , \wRegInA20[11] , \wRegInA55[21] , \wRegInA76[10] , 
        \wRegInB85[16] , \wBMid35[21] , \wAIn89[13] , \wAMid92[18] , 
        \wAMid126[3] , \wRegInA35[25] , \wRegInA40[15] , \ScanLink51[7] , 
        \wRegInB90[22] , \wRegInA16[14] , \wRegInA63[24] , \wBMid40[11] , 
        \ScanLink222[25] , \ScanLink187[22] , \wAIn5[1] , \wAMid5[12] , 
        \wBMid16[10] , \ScanLink201[14] , \wAIn6[2] , \wAIn12[25] , 
        \wBMid20[15] , \wBMid63[20] , \wBMid76[14] , \wAIn91[8] , 
        \wRegInA76[4] , \ScanLink214[20] , \ScanLink29[21] , \ScanLink49[25] , 
        \ScanLink237[11] , \ScanLink192[16] , \wAIn24[20] , \wAIn51[10] , 
        \wBMid55[25] , \wRegInB16[1] , \ScanLink242[21] , \wRegInB118[6] , 
        \wAIn72[21] , \wBMid77[5] , \wRegInB48[21] , \wRegInA98[16] , 
        \ScanLink108[2] , \wBIn25[18] , \wAIn44[24] , \wBIn110[31] , 
        \wBIn50[28] , \ScanLink36[0] , \wAIn31[14] , \wBIn50[31] , 
        \wBIn73[19] , \wBIn110[28] , \wRegInB28[25] , \wAIn67[15] , 
        \wRegInB105[9] , \wBIn38[1] , \wBMid69[9] , \wBMid74[6] , \wAIn109[6] , 
        \wRegInA16[27] , \wRegInA35[16] , \wRegInA40[26] , \wRegInA68[8] , 
        \wRegInB90[11] , \wBIn88[18] , \wAIn89[20] , \wAMid116[31] , 
        \wRegInA63[17] , \wRegInA76[23] , \wBMid98[21] , \wAMid116[28] , 
        \wRegInA20[22] , \wRegInB85[25] , \ScanLink35[3] , \wRegInA55[12] , 
        \wAIn114[9] , \wRegInA75[7] , \ScanLink109[13] , \wRegInB15[2] , 
        \ScanLink169[17] , \ScanLink84[21] , \ScanLink91[15] , \wAMid17[16] , 
        \wAIn21[4] , \wBIn59[8] , \wAMid61[0] , \ScanLink229[29] , \wBIn96[1] , 
        \ScanLink229[30] , \wAMid62[26] , \wRegInB69[4] , \wRegInA108[26] , 
        \ScanLink61[18] , \ScanLink42[29] , \ScanLink37[19] , \ScanLink14[31] , 
        \ScanLink42[30] , \ScanLink14[28] , \wBIn18[11] , \wAIn19[30] , 
        \wAMid21[13] , \wAMid34[27] , \wAMid41[17] , \wBIn44[7] , 
        \ScanLink177[7] , \wAMid54[23] , \wRegInB23[30] , \ScanLink49[5] , 
        \wRegInB75[28] , \wAIn19[29] , \wAMid77[12] , \wBIn78[15] , 
        \wRegInB23[29] , \wRegInB56[19] , \wRegInB75[31] , \ScanLink217[2] , 
        \ScanLink8[9] , \wAIn22[7] , \wBIn47[4] , \wAMid108[10] , \wBIn83[14] , 
        \wBIn96[20] , \wAMid99[27] , \ScanLink174[4] , \ScanLink6[26] , 
        \wBMid111[21] , \wRegInA7[8] , \ScanLink214[1] , \wBIn95[2] , 
        \wAIn97[18] , \wBMid104[15] , \wRegInB77[8] , \wRegInB4[27] , 
        \wRegInB126[26] , \wAMid17[25] , \wBIn20[3] , \wAMid62[3] , 
        \wRegInB105[17] , \wBMid86[19] , \wRegInA2[22] , \wRegInB110[23] , 
        \ScanLink98[0] , \ScanLink57[9] , \wAMid21[20] , \wAIn111[4] , 
        \ScanLink113[3] , \wAMid54[10] , \wAIn97[6] , \wAMid77[21] , 
        \wBIn78[26] , \wBIn18[22] , \wAMid34[14] , \wAMid62[15] , 
        \wRegInA93[29] , \wAMid41[24] , \wAIn45[0] , \wRegInA93[30] , 
        \ScanLink199[30] , \wAIn104[30] , \wRegInA108[15] , \ScanLink199[29] , 
        \wAIn104[29] , \wAIn127[18] , \wRegInB103[7] , \wAMid4[18] , 
        \wBIn7[18] , \ScanLink162[28] , \wAMid10[3] , \wBIn23[0] , \wAIn46[3] , 
        \wBMid72[8] , \wRegInA2[11] , \wRegInB110[10] , \ScanLink134[30] , 
        \ScanLink117[18] , \ScanLink162[31] , \ScanLink141[19] , \wBIn83[27] , 
        \wRegInB4[14] , \ScanLink134[29] , \wRegInB100[4] , \wRegInB126[15] , 
        \wRegInB105[24] , \wBMid104[26] , \ScanLink110[0] , \wBIn35[4] , 
        \wBMid79[3] , \wAIn94[5] , \wAIn112[7] , \wBIn96[13] , \wAMid99[14] , 
        \wAMid108[23] , \wRegInA68[31] , \wRegInA73[9] , \ScanLink6[15] , 
        \wBMid111[12] , \wRegInA68[28] , \ScanLink108[19] , \ScanLink106[4] , 
        \wAIn82[1] , \wAIn104[3] , \wAMid93[21] , \wBMid120[1] , 
        \wAMid121[27] , \wRegInA8[24] , \ScanLink38[6] , \wBIn12[17] , 
        \wAMid13[0] , \wBIn31[26] , \wBIn44[16] , \wAIn50[7] , \wAMid102[16] , 
        \wAMid86[15] , \wAMid117[22] , \wRegInA21[28] , \wRegInA78[2] , 
        \ScanLink25[9] , \wRegInB18[7] , \wRegInA21[31] , \wRegInA54[18] , 
        \wRegInA77[30] , \wRegInA77[29] , \wRegInB116[0] , \wBIn89[12] , 
        \wBIn127[27] , \ScanLink118[8] , \wAIn53[4] , \wBIn67[27] , 
        \wAMid68[20] , \wBIn104[16] , \wBMid123[2] , \wBIn24[12] , 
        \wBIn51[22] , \wBIn72[13] , \wBIn111[22] , \wRegInB115[3] , 
        \wBIn36[7] , \wAIn81[2] , \wAIn107[0] , \ScanLink186[31] , 
        \ScanLink105[7] , \wBIn6[21] , \wBIn6[12] , \wBMid5[20] , 
        \wRegInA102[20] , \wRegInA117[14] , \ScanLink186[28] , 
        \wRegInA121[11] , \wBMid5[13] , \wAIn34[3] , \wBIn83[6] , \wBIn109[7] , 
        \wBIn51[0] , \wAMid74[7] , \wAMid86[26] , \wAMid117[11] , \wBIn89[21] , 
        \wAIn88[19] , \wAMid93[12] , \wAMid102[25] , \wAMid121[14] , 
        \wRegInB91[31] , \ScanLink0[1] , \wRegInB91[28] , \wAMid69[8] , 
        \wBIn114[8] , \ScanLink162[0] , \wBMid99[18] , \wRegInA8[17] , 
        \ScanLink202[5] , \ScanLink85[18] , \wRegInA102[13] , \wRegInA123[6] , 
        \ScanLink243[18] , \ScanLink236[28] , \ScanLink161[3] , \wBIn12[24] , 
        \wBMid17[30] , \wBMid17[29] , \wBMid41[31] , \wBIn52[3] , 
        \wRegInA121[22] , \ScanLink236[31] , \ScanLink215[19] , \wBMid62[19] , 
        \ScanLink28[18] , \ScanLink90[8] , \wBMid41[28] , \wRegInA120[5] , 
        \wRegInA117[27] , \ScanLink201[6] , \wBIn24[21] , \wBMid34[18] , 
        \wBIn72[20] , \wBIn111[11] , \wAMid77[4] , \wBIn80[5] , \wAIn25[19] , 
        \wAIn37[0] , \wBIn51[11] , \wBIn31[15] , \wBIn44[25] , \wAIn50[29] , 
        \wBIn127[14] , \wAIn50[30] , \wBIn67[14] , \wAIn73[18] , 
        \wRegInB49[18] , \ScanLink3[2] , \wAIn56[9] , \wAMid68[13] , 
        \wAIn83[15] , \wAIn96[21] , \wBIn104[25] , \wRegInA63[3] , 
        \wBIn97[19] , \wAMid109[30] , \wBMid110[18] , \wRegInA69[22] , 
        \wAMid109[29] , \ScanLink140[13] , \ScanLink135[23] , \wBMid62[2] , 
        \wBMid87[20] , \wAIn99[0] , \ScanLink163[22] , \wAIn18[10] , 
        \wBMid61[1] , \wBMid92[14] , \ScanLink176[16] , \ScanLink116[12] , 
        \ScanLink155[27] , \ScanLink103[26] , \ScanLink23[7] , 
        \ScanLink120[17] , \wBMid69[15] , \wAIn110[17] , \ScanLink248[14] , 
        \ScanLink198[23] , \ScanLink15[11] , \ScanLink60[21] , 
        \ScanLink43[10] , \ScanLink36[20] , \wAIn105[23] , \ScanLink23[14] , 
        \wAIn126[12] , \ScanLink56[24] , \ScanLink20[4] , \wRegInB57[20] , 
        \ScanLink228[10] , \ScanLink75[15] , \wBIn19[31] , \wBIn30[9] , 
        \wRegInB22[10] , \wRegInA87[17] , \wRegInB74[11] , \wAIn48[5] , 
        \wRegInA60[0] , \ScanLink103[9] , \wBIn19[28] , \wRegInB14[15] , 
        \wRegInB61[25] , \wAMid72[9] , \wAIn78[14] , \wRegInB42[14] , 
        \wRegInB37[24] , \wRegInA92[23] , \ScanLink103[15] , \wBIn85[8] , 
        \wBMid92[27] , \ScanLink176[25] , \wBMid87[13] , \wRegInA3[31] , 
        \wRegInB111[30] , \ScanLink179[1] , \ScanLink120[24] , 
        \ScanLink155[14] , \ScanLink135[10] , \ScanLink47[3] , \wRegInA3[28] , 
        \wRegInB111[29] , \ScanLink219[4] , \ScanLink140[20] , 
        \ScanLink116[21] , \ScanLink163[11] , \wAIn8[4] , \wAIn83[26] , 
        \wBIn98[7] , \wRegInA69[11] , \wAIn18[23] , \wAMid55[30] , 
        \wAIn78[27] , \wAIn96[12] , \wBIn112[6] , \wRegInA125[8] , 
        \ScanLink95[5] , \wBIn111[5] , \wRegInB14[26] , \wRegInB67[2] , 
        \wRegInB61[16] , \wRegInB22[23] , \wRegInB37[17] , \wRegInB42[27] , 
        \wRegInA92[10] , \wRegInA87[24] , \wAMid76[18] , \ScanLink207[8] , 
        \wRegInB57[13] , \wRegInB64[1] , \wAMid20[19] , \wAMid55[29] , 
        \wRegInB74[22] , \ScanLink96[6] , \wAMid24[31] , \wBIn49[2] , 
        \ScanLink56[17] , \wBMid69[26] , \wAIn105[10] , \ScanLink23[27] , 
        \wAIn110[24] , \wAIn126[21] , \ScanLink228[23] , \ScanLink75[26] , 
        \ScanLink248[27] , \ScanLink198[10] , \ScanLink60[12] , 
        \ScanLink44[0] , \ScanLink15[22] , \ScanLink43[23] , \wRegInB10[17] , 
        \wRegInB65[27] , \ScanLink36[13] , \wRegInB33[26] , \wRegInB46[16] , 
        \wRegInB40[7] , \wRegInA96[21] , \wRegInB53[22] , \wAMid24[28] , 
        \wAMid48[3] , \wRegInB26[12] , \wRegInA83[15] , \wAIn69[22] , 
        \wAMid72[29] , \wRegInB0[7] , \wRegInB70[13] , \wAMid72[30] , 
        \wRegInA20[2] , \wBIn2[10] , \wAIn15[8] , \wBMid18[27] , \wAMid51[18] , 
        \wAIn101[21] , \ScanLink60[6] , \ScanLink27[16] , \wBMid21[3] , 
        \wAIn122[10] , \wRegInA118[30] , \ScanLink52[26] , \wRegInB92[1] , 
        \wRegInA118[29] , \ScanLink71[17] , \ScanLink189[15] , \wBMid78[23] , 
        \wAIn114[15] , \ScanLink239[26] , \ScanLink11[13] , \ScanLink64[23] , 
        \ScanLink32[22] , \wAMid117[2] , \ScanLink47[12] , \wBMid22[0] , 
        \wBMid83[22] , \wBMid96[16] , \wRegInB91[2] , \ScanLink172[14] , 
        \ScanLink107[24] , \ScanLink151[25] , \ScanLink63[5] , \wAMid114[1] , 
        \ScanLink144[11] , \ScanLink124[15] , \ScanLink131[21] , 
        \ScanLink167[20] , \wBMid18[14] , \wBIn73[8] , \wAIn87[17] , 
        \wAMid99[6] , \wRegInB115[18] , \ScanLink112[10] , \wRegInA7[19] , 
        \wAMid89[31] , \wRegInA18[10] , \wRegInB43[4] , \ScanLink140[8] , 
        \wBMid78[10] , \wAMid84[9] , \wAMid89[28] , \wRegInA23[1] , 
        \wRegInA78[14] , \wAIn92[23] , \wAIn114[26] , \wRegInB3[4] , 
        \ScanLink239[15] , \ScanLink64[10] , \ScanLink47[21] , 
        \ScanLink11[20] , \ScanLink32[11] , \wAMid31[8] , \wBMid45[7] , 
        \wAIn101[12] , \wRegInA96[0] , \ScanLink52[15] , \ScanLink27[25] , 
        \wRegInA59[9] , \ScanLink189[26] , \ScanLink71[24] , \wAIn122[23] , 
        \wAIn69[11] , \wRegInB26[21] , \wRegInA83[26] , \wRegInB24[3] , 
        \wRegInB53[11] , \wAIn0[26] , \wAMid0[30] , \wAMid0[29] , \wBIn2[23] , 
        \wBIn7[8] , \wBIn68[30] , \wRegInB70[20] , \wBMid58[8] , \wBIn68[29] , 
        \wAIn125[8] , \wRegInB10[24] , \wRegInA44[6] , \wRegInB65[14] , 
        \wBMid97[1] , \wBMid83[11] , \wAIn87[24] , \wAIn92[10] , 
        \wRegInB27[0] , \wRegInB33[15] , \wRegInB46[25] , \wRegInA96[12] , 
        \wRegInA78[27] , \ScanLink244[9] , \wBIn93[28] , \wBMid94[2] , 
        \wBMid114[29] , \wRegInA18[23] , \wBIn93[31] , \wBMid114[30] , 
        \wRegInA47[5] , \ScanLink131[12] , \ScanLink167[13] , 
        \ScanLink144[22] , \ScanLink112[23] , \wBMid1[22] , \wBMid46[4] , 
        \wBMid96[25] , \wBMid102[9] , \ScanLink172[27] , \ScanLink107[17] , 
        \wRegInB46[9] , \wRegInB89[0] , \wRegInA95[3] , \ScanLink151[16] , 
        \ScanLink139[3] , \ScanLink124[26] , \wRegInA106[22] , 
        \ScanLink232[19] , \ScanLink225[0] , \ScanLink211[31] , 
        \ScanLink247[29] , \wRegInA125[13] , \ScanLink211[28] , 
        \ScanLink247[30] , \wAIn10[5] , \wAIn13[6] , \wBMid13[18] , 
        \wBMid30[30] , \wRegInA104[3] , \wBIn76[5] , \ScanLink59[19] , 
        \wBIn20[10] , \wBMid30[29] , \wBMid66[28] , \ScanLink145[5] , 
        \wBMid45[19] , \wBMid66[31] , \wRegInA113[16] , \wBIn55[20] , 
        \wBIn76[11] , \wAMid79[16] , \wAMid81[4] , \wBIn115[20] , 
        \wRegInB6[9] , \ScanLink66[8] , \wAIn21[28] , \wBIn35[24] , 
        \wBIn40[14] , \wAIn54[18] , \ScanLink197[3] , \wAIn77[30] , 
        \wBIn123[25] , \wBIn16[15] , \wBIn63[25] , \wAIn77[29] , \wBIn100[14] , 
        \wRegInB38[19] , \wAMid19[12] , \wAMid53[2] , \wAIn21[31] , 
        \wAMid50[1] , \wAMid82[17] , \wAMid113[20] , \wRegInB58[5] , 
        \wAMid97[23] , \wBIn98[24] , \wAMid125[25] , \ScanLink8[22] , 
        \wBIn68[9] , \wAMid106[14] , \wRegInB95[19] , \ScanLink194[0] , 
        \wBIn16[26] , \wBIn35[17] , \wBMid39[1] , \wRegInA38[0] , 
        \wRegInA107[0] , \ScanLink78[4] , \ScanLink226[3] , \wBIn75[6] , 
        \wAMid82[7] , \ScanLink81[29] , \ScanLink146[6] , \ScanLink81[30] , 
        \wBIn40[27] , \wBIn123[16] , \wAMid19[21] , \wBIn20[23] , \wAMid37[6] , 
        \wBMid43[9] , \wBIn63[16] , \wBIn100[27] , \wBMid107[4] , 
        \wBIn115[13] , \wRegInA88[19] , \wBIn76[22] , \wAMid79[25] , 
        \wBIn55[13] , \wAIn77[2] , \wBIn1[6] , \wRegInA106[11] , 
        \wRegInA113[25] , \ScanLink241[4] , \ScanLink182[19] , \wBIn2[5] , 
        \wBMid1[11] , \ScanLink121[1] , \wBIn11[2] , \wBIn12[1] , \wAIn123[6] , 
        \wAIn120[5] , \wRegInA42[8] , \wRegInA125[20] , \ScanLink242[7] , 
        \ScanLink179[18] , \wAMid4[22] , \wBIn6[31] , \wAMid34[5] , 
        \wAIn74[1] , \wAMid97[10] , \wBIn98[17] , \wBMid119[8] , 
        \ScanLink122[2] , \ScanLink8[11] , \wAMid106[27] , \wAMid125[16] , 
        \wRegInA25[19] , \wRegInA50[29] , \wAMid82[24] , \wBMid104[7] , 
        \wAMid113[13] , \wRegInA50[30] , \wRegInA73[18] , \ScanLink140[29] , 
        \ScanLink135[19] , \ScanLink116[31] , \ScanLink88[3] , \wBIn6[28] , 
        \wRegInA3[21] , \wRegInB111[20] , \ScanLink116[28] , \ScanLink163[18] , 
        \ScanLink140[30] , \ScanLink6[6] , \wAMid15[7] , \wAMid16[15] , 
        \wBMid18[3] , \wAMid20[10] , \wAIn32[4] , \wAMid72[0] , 
        \wRegInB104[14] , \wBIn85[1] , \wRegInB127[25] , \wRegInB5[24] , 
        \ScanLink179[8] , \wAMid55[20] , \wBIn57[7] , \wBIn82[17] , 
        \wBMid126[27] , \wRegInA125[1] , \ScanLink204[2] , \wBIn97[23] , 
        \wAMid98[24] , \wBMid105[16] , \ScanLink7[25] , \wBMid110[22] , 
        \wAMid109[13] , \wRegInA69[18] , \wAMid76[11] , \wBIn79[16] , 
        \ScanLink164[7] , \wRegInB64[8] , \ScanLink207[1] , \ScanLink59[6] , 
        \wRegInA126[2] , \wAMid35[24] , \wAMid40[14] , \wBIn54[4] , 
        \ScanLink167[4] , \wAMid63[25] , \wRegInA92[19] , \wAMid16[4] , 
        \wBIn19[12] , \wAIn31[7] , \wBIn86[2] , \wRegInB79[7] , 
        \wRegInA109[25] , \ScanLink198[19] , \ScanLink44[9] , \ScanLink5[5] , 
        \wBIn33[3] , \wAMid71[3] , \wAIn105[19] , \wAIn126[31] , 
        \wRegInA19[2] , \wAIn126[28] , \wRegInA9[7] , \wAIn96[31] , 
        \wBIn97[10] , \wAMid98[17] , \ScanLink7[16] , \wBMid110[11] , 
        \wAMid109[20] , \wBMid126[14] , \ScanLink100[3] , \wAIn56[0] , 
        \wBIn82[24] , \wAIn84[6] , \wAIn102[4] , \wAIn96[28] , \wBMid105[25] , 
        \wRegInB127[16] , \wRegInB5[17] , \wRegInB104[27] , \wRegInB110[7] , 
        \wBMid87[30] , \wBMid87[29] , \wAIn99[9] , \wBMid126[6] , 
        \wRegInA3[12] , \wRegInB111[13] , \wBMid61[8] , \wBMid125[5] , 
        \wRegInB113[4] , \ScanLink228[19] , \ScanLink36[30] , \ScanLink15[18] , 
        \wAMid16[26] , \wAMid35[17] , \wAIn55[3] , \wRegInA109[16] , 
        \ScanLink60[28] , \ScanLink43[19] , \ScanLink36[29] , \ScanLink60[31] , 
        \wAMid40[27] , \wAIn18[19] , \wBIn19[21] , \wAMid63[16] , 
        \wRegInB57[29] , \wAMid20[23] , \wBIn30[0] , \wAMid76[22] , 
        \wBIn79[25] , \wRegInB22[19] , \wRegInB57[30] , \wAIn101[7] , 
        \wRegInB74[18] , \ScanLink103[0] , \wAIn29[5] , \wBIn51[9] , 
        \wAMid55[13] , \wAIn87[5] , \wRegInA60[9] , \wAIn88[10] , \wBIn89[31] , 
        \wRegInA17[17] , \wRegInA62[27] , \wRegInA34[26] , \wRegInA41[16] , 
        \ScanLink41[4] , \ScanLink0[8] , \wRegInB91[21] , \wRegInA54[22] , 
        \wBIn89[28] , \wAMid117[18] , \wRegInA21[12] , \wRegInB84[15] , 
        \wRegInA77[13] , \wBMid99[11] , \wRegInB61[5] , \ScanLink85[11] , 
        \ScanLink108[23] , \ScanLink93[2] , \wBIn114[1] , \ScanLink162[9] , 
        \wBMid62[10] , \wAMid69[1] , \ScanLink168[27] , \ScanLink90[25] , 
        \ScanLink28[11] , \wBMid17[20] , \ScanLink90[1] , \wBMid41[21] , 
        \ScanLink200[24] , \ScanLink256[25] , \wAIn0[15] , \wAMid4[11] , 
        \wBMid5[30] , \wAIn13[26] , \wAIn13[15] , \wBMid21[25] , \wBMid34[11] , 
        \wBMid54[15] , \wRegInB62[6] , \ScanLink243[11] , \ScanLink223[15] , 
        \ScanLink186[12] , \ScanLink236[21] , \ScanLink193[26] , \wAIn25[10] , 
        \wBMid77[24] , \wBIn117[2] , \ScanLink215[10] , \ScanLink48[15] , 
        \ScanLink42[7] , \wAIn50[20] , \wAIn73[11] , \wRegInB49[11] , 
        \wRegInA99[26] , \wBIn24[31] , \wBIn24[28] , \wAIn30[24] , 
        \wAIn66[25] , \wBIn111[18] , \wRegInB29[15] , \wBIn72[29] , 
        \wBIn28[2] , \wAIn37[9] , \wAIn45[14] , \wBIn51[18] , \wBMid64[5] , 
        \wBIn72[30] , \wAIn82[8] , \wBMid99[22] , \ScanLink168[14] , 
        \ScanLink108[10] , \ScanLink90[16] , \ScanLink85[22] , \wRegInA65[4] , 
        \wRegInA17[24] , \wRegInA21[21] , \wRegInA54[11] , \wRegInB84[26] , 
        \ScanLink25[0] , \wRegInA77[20] , \wRegInB116[9] , \wAIn88[23] , 
        \wBMid120[8] , \wAMid93[28] , \wRegInA62[14] , \wAIn66[16] , 
        \wAMid93[31] , \wAIn119[5] , \wRegInA34[15] , \wRegInB91[12] , 
        \wRegInB29[26] , \wRegInA41[25] , \wAMid13[9] , \wAIn25[23] , 
        \wAIn30[17] , \wAIn45[27] , \ScanLink26[3] , \wAIn50[13] , 
        \wAMid68[30] , \ScanLink118[1] , \wBMid67[6] , \wAMid68[29] , 
        \wAIn73[22] , \wRegInA99[15] , \wBMid21[16] , \wRegInB49[22] , 
        \ScanLink236[12] , \ScanLink193[15] , \wRegInA102[29] , 
        \ScanLink243[22] , \wBMid5[29] , \wBMid54[26] , \wRegInB108[5] , 
        \wRegInA102[30] , \wRegInA121[18] , \ScanLink215[23] , 
        \ScanLink48[26] , \wBMid17[13] , \wBMid77[17] , \wAIn107[9] , 
        \ScanLink200[17] , \wBMid34[22] , \wBMid62[23] , \wRegInA66[7] , 
        \ScanLink28[22] , \wBMid41[12] , \ScanLink223[26] , \ScanLink186[21] , 
        \ScanLink256[16] , \wAMid0[20] , \wBMid1[18] , \wBIn12[8] , 
        \wAIn17[17] , \wBMid43[0] , \wRegInB58[27] , \wAMid19[31] , 
        \wAIn21[12] , \wAIn34[26] , \wAIn62[27] , \wRegInA88[10] , 
        \wAIn41[16] , \wRegInA90[7] , \wAMid19[28] , \wAIn54[22] , 
        \wBMid25[27] , \wBMid50[17] , \wAIn77[13] , \wBMid91[6] , 
        \wRegInB38[23] , \ScanLink247[13] , \wRegInA106[18] , 
        \ScanLink232[23] , \ScanLink197[24] , \wRegInA125[30] , 
        \ScanLink121[8] , \wBMid73[26] , \ScanLink39[27] , \wBMid66[12] , 
        \wRegInA42[1] , \ScanLink211[12] , \wRegInA125[29] , \wAMid0[13] , 
        \wAIn4[24] , \wBMid13[22] , \wBMid45[23] , \ScanLink204[26] , 
        \ScanLink59[23] , \wBIn9[15] , \wBMid8[4] , \wBMid30[13] , 
        \wRegInB22[4] , \ScanLink252[27] , \wAIn69[7] , \wBMid88[27] , 
        \wRegInA41[2] , \ScanLink227[17] , \ScanLink182[10] , \wBMid119[1] , 
        \wBMid13[11] , \wAMid29[3] , \wBMid92[5] , \ScanLink94[27] , 
        \wBMid40[3] , \wAIn74[8] , \wRegInB21[7] , \ScanLink179[11] , 
        \ScanLink119[15] , \ScanLink81[13] , \wRegInA25[10] , \wRegInA50[20] , 
        \wRegInB80[17] , \wRegInA93[4] , \wRegInA73[11] , \wAMid97[19] , 
        \wAIn99[26] , \wRegInA13[15] , \wRegInA66[25] , \ScanLink8[18] , 
        \wRegInA30[24] , \wRegInA45[14] , \wRegInB95[23] , \ScanLink204[15] , 
        \ScanLink59[10] , \wAIn4[17] , \wBMid30[20] , \wBMid66[21] , 
        \wRegInA26[5] , \wBMid45[10] , \ScanLink227[24] , \ScanLink182[23] , 
        \wRegInB6[0] , \wBIn7[1] , \wBIn9[26] , \wAMid9[3] , \wAIn21[21] , 
        \wBMid25[14] , \ScanLink252[14] , \ScanLink232[10] , \ScanLink225[9] , 
        \ScanLink197[17] , \wBMid50[24] , \wRegInB89[9] , \ScanLink247[20] , 
        \wAIn54[11] , \wBMid73[15] , \wRegInB46[0] , \ScanLink211[21] , 
        \ScanLink39[14] , \ScanLink158[3] , \wBMid27[4] , \wAIn77[20] , 
        \wAMid111[5] , \wBIn76[18] , \wBIn115[29] , \wRegInB38[10] , 
        \ScanLink238[6] , \wRegInA88[23] , \wAIn17[24] , \wBIn55[30] , 
        \wAIn62[14] , \wRegInB58[14] , \wRegInB94[6] , \wBIn20[19] , 
        \wAIn41[25] , \wBIn115[30] , \wBIn55[29] , \ScanLink66[1] , 
        \wBMid24[7] , \wAIn34[15] , \wRegInA119[5] , \wBMid39[8] , 
        \wAMid50[8] , \wRegInA13[26] , \wBIn68[0] , \wRegInA66[16] , 
        \wAIn99[15] , \wAMid112[6] , \wRegInA30[17] , \wRegInB95[10] , 
        \ScanLink194[9] , \wAMid113[30] , \wAMid113[29] , \wRegInA25[23] , 
        \wRegInA38[9] , \wRegInA45[27] , \wRegInB80[24] , \ScanLink65[2] , 
        \wRegInA50[13] , \wRegInA73[22] , \wRegInB97[5] , \wBMid88[14] , 
        \wRegInB5[3] , \wRegInA25[6] , \ScanLink189[6] , \ScanLink179[22] , 
        \ScanLink81[20] , \wRegInB45[3] , \wRegInA107[9] , \ScanLink119[26] , 
        \ScanLink94[14] , \wAMid31[1] , \wAIn71[5] , \wRegInA96[9] , 
        \wBMid101[3] , \wRegInA59[0] , \wRegInA118[13] , \wAMid44[16] , 
        \wBMid78[19] , \wRegInB39[5] , \ScanLink64[19] , \ScanLink47[31] , 
        \ScanLink47[28] , \ScanLink11[29] , \ScanLink32[18] , \ScanLink11[30] , 
        \wAMid12[17] , \wBIn14[6] , \wAIn125[1] , \ScanLink127[6] , 
        \wAMid31[26] , \wBMid58[1] , \wAMid67[27] , \wBMid97[8] , \wBIn68[20] , 
        \wAMid51[22] , \wAIn69[18] , \wAMid72[13] , \wRegInB26[28] , 
        \wRegInB26[31] , \wRegInB53[18] , \wRegInB70[30] , \ScanLink247[3] , 
        \ScanLink19[4] , \wBIn4[2] , \wBIn17[5] , \wAMid24[12] , 
        \wRegInB70[29] , \wBIn93[21] , \wBMid114[20] , \wAIn126[2] , 
        \ScanLink3[27] , \wAMid12[24] , \wAMid24[21] , \wAMid32[2] , 
        \wBIn86[15] , \wBMid101[14] , \wAMid118[25] , \wRegInA88[5] , 
        \ScanLink124[5] , \wBMid122[25] , \ScanLink244[0] , \wAMid89[12] , 
        \wBMid89[4] , \wAIn92[19] , \wBMid102[0] , \wRegInB27[9] , 
        \wRegInB100[16] , \wBIn70[2] , \wAIn72[6] , \wRegInB1[26] , 
        \wRegInB123[27] , \wAMid72[20] , \wBMid83[18] , \wRegInA7[23] , 
        \wRegInB115[22] , \wAMid87[3] , \ScanLink143[2] , \wAMid31[15] , 
        \wAMid51[11] , \wAMid44[25] , \wRegInA96[31] , \wRegInA102[4] , 
        \ScanLink223[7] , \wAIn15[1] , \wAMid55[5] , \wAMid67[14] , 
        \wBIn68[13] , \wRegInA96[28] , \ScanLink191[4] , \wAIn16[2] , 
        \wAIn101[31] , \wAIn101[28] , \wAIn122[19] , \wRegInB92[8] , 
        \wRegInA118[20] , \ScanLink192[7] , \ScanLink167[30] , 
        \ScanLink144[18] , \ScanLink131[28] , \wAMid114[8] , \wAIn0[5] , 
        \wBMid0[21] , \wAMid1[19] , \wBIn2[19] , \ScanLink167[29] , 
        \wAMid7[5] , \wBMid22[9] , \wBMid29[2] , \wAMid56[6] , \wRegInA7[10] , 
        \wRegInB115[11] , \ScanLink131[31] , \ScanLink112[19] , \wBIn65[5] , 
        \wBIn73[1] , \wRegInB1[15] , \wRegInB100[25] , \wRegInB123[14] , 
        \ScanLink140[1] , \wAMid84[0] , \wBIn86[26] , \wBMid101[27] , 
        \wAMid109[7] , \wBMid122[16] , \wAMid118[16] , \wRegInA23[8] , 
        \wAMid89[21] , \wBIn93[12] , \wBMid114[13] , \wRegInA18[19] , 
        \ScanLink220[4] , \ScanLink3[14] , \wRegInA101[7] , \ScanLink156[5] , 
        \ScanLink178[31] , \wAMid92[4] , \ScanLink178[28] , \wBIn17[16] , 
        \wAMid40[2] , \wAMid96[20] , \wBIn99[27] , \wAMid107[17] , 
        \wRegInB55[9] , \ScanLink236[0] , \wRegInA117[3] , \ScanLink68[7] , 
        \wAMid124[26] , \wRegInA28[3] , \ScanLink184[3] , \wRegInB8[6] , 
        \ScanLink9[21] , \wBIn62[26] , \wAMid83[14] , \wRegInA24[30] , 
        \wRegInB48[6] , \wRegInA72[28] , \wAMid112[23] , \wRegInA24[29] , 
        \ScanLink75[8] , \wRegInA51[19] , \wRegInA72[31] , \wBIn101[17] , 
        \wAMid18[11] , \wBIn21[13] , \wBIn34[27] , \wBIn41[17] , \wAMid43[1] , 
        \ScanLink187[0] , \wBIn122[26] , \ScanLink148[9] , \wBIn54[23] , 
        \wRegInA89[30] , \wBIn66[6] , \wBIn77[12] , \wAMid78[15] , 
        \wBIn114[23] , \wRegInA89[29] , \wAMid91[7] , \wRegInA112[15] , 
        \ScanLink183[29] , \ScanLink183[30] , \ScanLink155[6] , 
        \wRegInA124[10] , \wBMid0[12] , \wAMid4[6] , \wRegInA107[21] , 
        \wRegInA114[0] , \ScanLink235[3] , \wBMid6[2] , \wAMid24[6] , 
        \wBMid50[9] , \wBMid114[4] , \wRegInB99[3] , \wAMid83[27] , 
        \wAIn64[2] , \wAMid112[10] , \wAMid96[13] , \wBIn99[14] , 
        \wAMid107[24] , \wRegInB94[29] , \ScanLink9[12] , \wAMid39[9] , 
        \wAMid124[15] , \wRegInB94[30] , \wRegInB122[5] , \wRegInA51[8] , 
        \ScanLink132[1] , \ScanLink252[4] , \ScanLink80[19] , \ScanLink131[2] , 
        \wAMid2[8] , \wBIn3[13] , \wBMid5[1] , \wBMid12[31] , \wBMid44[29] , 
        \wRegInA107[12] , \wRegInA124[23] , \ScanLink233[30] , 
        \ScanLink210[18] , \ScanLink246[19] , \ScanLink233[29] , 
        \ScanLink251[7] , \ScanLink58[30] , \wBMid12[28] , \wBMid31[19] , 
        \wRegInA112[26] , \wBMid44[30] , \wBMid67[18] , \ScanLink58[29] , 
        \wBIn17[25] , \wBIn21[20] , \wAMid27[5] , \wBIn54[10] , \wAIn67[1] , 
        \wBIn114[10] , \wBMid117[7] , \wBIn77[21] , \wAMid78[26] , 
        \wAMid18[22] , \wAIn55[31] , \wAIn76[19] , \wRegInB121[6] , 
        \wBIn62[15] , \wAIn20[18] , \wBIn101[24] , \wRegInB39[29] , 
        \wBMid32[3] , \wBIn34[14] , \wBIn41[24] , \wAIn55[28] , \wAIn86[14] , 
        \wAIn93[20] , \wBIn122[15] , \wRegInB39[30] , \wRegInA79[17] , 
        \wBIn126[3] , \wRegInA33[2] , \wBIn92[18] , \wBMid115[19] , 
        \wRegInA19[13] , \wRegInB53[7] , \ScanLink166[23] , \wAIn18[4] , 
        \wBMid19[24] , \wBMid31[0] , \wBMid79[20] , \wBMid82[21] , 
        \wAMid89[5] , \ScanLink113[13] , \wAMid104[2] , \ScanLink145[12] , 
        \ScanLink130[22] , \wBMid97[15] , \ScanLink150[26] , \ScanLink73[6] , 
        \wAIn115[16] , \wRegInB81[1] , \ScanLink173[17] , \ScanLink125[16] , 
        \ScanLink106[27] , \ScanLink33[21] , \wAMid107[1] , \ScanLink46[11] , 
        \wAIn100[22] , \wAIn123[13] , \ScanLink238[25] , \ScanLink10[10] , 
        \ScanLink65[20] , \wRegInB82[2] , \ScanLink70[14] , \ScanLink188[16] , 
        \ScanLink70[5] , \ScanLink26[15] , \wBIn60[8] , \wRegInB71[10] , 
        \ScanLink53[25] , \wBIn125[0] , \ScanLink153[8] , \wRegInA30[1] , 
        \wAMid58[0] , \wRegInB27[11] , \wRegInB52[21] , \wRegInA82[16] , 
        \wAIn68[21] , \wAMid97[9] , \wRegInB47[15] , \wBIn3[20] , \wBIn9[7] , 
        \wBIn69[19] , \wBMid97[26] , \wRegInB11[14] , \wRegInB32[25] , 
        \wRegInB50[4] , \wRegInA97[22] , \wRegInB64[24] , \wAMid22[8] , 
        \wBMid56[7] , \wRegInA85[0] , \ScanLink150[15] , \ScanLink129[0] , 
        \ScanLink125[25] , \ScanLink106[14] , \wRegInA6[29] , \wRegInB114[28] , 
        \ScanLink173[24] , \ScanLink249[5] , \ScanLink113[20] , 
        \ScanLink166[10] , \wAIn5[8] , \wBIn7[22] , \wBIn7[11] , \wAMid18[2] , 
        \wAIn19[13] , \wBIn19[3] , \wBMid19[17] , \wAMid25[18] , \wAMid50[28] , 
        \wBMid82[12] , \wRegInA6[30] , \wRegInB114[31] , \ScanLink130[11] , 
        \ScanLink17[2] , \wBMid84[1] , \wRegInA57[6] , \ScanLink145[21] , 
        \wAIn86[27] , \wRegInA19[20] , \wBMid87[2] , \wAMid88[18] , 
        \wAIn93[13] , \wRegInB37[3] , \wRegInA79[24] , \wRegInB11[27] , 
        \wRegInB32[16] , \wRegInA97[11] , \wRegInB47[26] , \wRegInA54[5] , 
        \wRegInB64[17] , \wRegInB71[23] , \wAMid50[31] , \wRegInB27[22] , 
        \wRegInA82[25] , \wBMid55[4] , \wAIn68[12] , \wAMid73[19] , 
        \wRegInB34[0] , \wRegInB52[12] , \wRegInA119[19] , \ScanLink70[27] , 
        \wBMid111[9] , \ScanLink188[25] , \wAIn123[20] , \ScanLink53[16] , 
        \wAMid21[29] , \wAIn79[17] , \wBMid79[13] , \wAIn100[11] , 
        \wRegInA86[3] , \ScanLink26[26] , \wAIn115[25] , \ScanLink46[22] , 
        \ScanLink14[1] , \ScanLink33[12] , \wRegInB127[8] , \ScanLink238[16] , 
        \ScanLink65[13] , \wRegInB43[17] , \ScanLink10[23] , \wRegInB10[6] , 
        \wRegInB15[16] , \wRegInB36[27] , \wRegInA93[20] , \wRegInB60[26] , 
        \wRegInB75[12] , \wAMid54[19] , \wAIn58[6] , \wAMid77[31] , 
        \wRegInA70[3] , \wRegInB56[23] , \wAMid21[30] , \wRegInB23[13] , 
        \wRegInA86[14] , \wAIn45[9] , \wBMid68[16] , \wAMid77[28] , 
        \wAIn127[11] , \ScanLink229[13] , \ScanLink74[16] , \wAIn104[20] , 
        \ScanLink22[17] , \wAIn111[14] , \ScanLink57[27] , \ScanLink30[7] , 
        \ScanLink37[23] , \wBMid71[2] , \ScanLink42[13] , \wBMid72[1] , 
        \wBMid93[17] , \ScanLink249[17] , \ScanLink199[20] , \ScanLink14[12] , 
        \ScanLink154[24] , \ScanLink61[22] , \ScanLink33[4] , 
        \ScanLink177[15] , \ScanLink121[14] , \ScanLink162[21] , 
        \ScanLink102[25] , \wBMid15[6] , \wBIn23[9] , \wAIn82[16] , 
        \wBMid86[23] , \wAIn89[3] , \wRegInA2[18] , \wRegInB110[19] , 
        \ScanLink117[11] , \ScanLink141[10] , \ScanLink134[20] , \wAIn97[22] , 
        \wRegInB13[5] , \wRegInA68[21] , \ScanLink110[9] , \wAIn111[27] , 
        \wRegInA73[0] , \ScanLink54[3] , \ScanLink42[20] , \ScanLink249[24] , 
        \ScanLink199[13] , \ScanLink37[10] , \ScanLink61[11] , 
        \ScanLink74[25] , \ScanLink14[21] , \wBIn18[18] , \wAIn19[20] , 
        \wBIn59[1] , \wAMid61[9] , \ScanLink229[20] , \wBIn96[8] , 
        \wAIn127[22] , \ScanLink57[14] , \wBMid68[25] , \wAIn104[13] , 
        \wAMid123[7] , \ScanLink22[24] , \wRegInB23[20] , \wRegInB75[21] , 
        \ScanLink86[5] , \wRegInB56[10] , \wRegInA86[27] , \ScanLink8[0] , 
        \wRegInB74[2] , \wAIn79[24] , \wRegInB36[14] , \wRegInA93[13] , 
        \wAIn82[25] , \wBIn88[4] , \wAIn97[11] , \wBIn101[6] , \wRegInA4[2] , 
        \wRegInA14[7] , \wRegInB15[25] , \wRegInB43[24] , \wRegInB60[15] , 
        \ScanLink214[8] , \wAMid108[19] , \wRegInB77[1] , \ScanLink85[6] , 
        \wBIn96[30] , \wBIn96[29] , \wBIn102[5] , \wBMid111[31] , 
        \wRegInA17[4] , \wBMid111[28] , \wRegInA7[1] , \wRegInA68[12] , 
        \ScanLink209[7] , \ScanLink162[12] , \ScanLink117[22] , \wBMid16[5] , 
        \wBMid86[10] , \ScanLink134[13] , \ScanLink98[9] , \ScanLink57[0] , 
        \wBMid93[24] , \ScanLink141[23] , \wAMid120[4] , \ScanLink169[2] , 
        \ScanLink121[27] , \ScanLink154[17] , \ScanLink102[16] , \wBMid4[23] , 
        \wRegInA120[12] , \ScanLink214[29] , \ScanLink177[26] , 
        \ScanLink242[31] , \wBIn13[27] , \wBIn13[14] , \wBMid16[19] , 
        \wBIn26[4] , \wBMid35[28] , \wRegInB16[8] , \wRegInA103[23] , 
        \ScanLink237[18] , \ScanLink214[30] , \ScanLink242[28] , \wBMid40[18] , 
        \wBMid63[30] , \wRegInA116[17] , \ScanLink29[31] , \wBMid35[31] , 
        \wAIn24[30] , \wBIn25[11] , \wBIn50[21] , \wBMid63[29] , \wAIn91[1] , 
        \wAIn117[3] , \ScanLink115[4] , \ScanLink29[28] , \ScanLink36[9] , 
        \wBIn66[24] , \wBIn73[10] , \wBIn110[21] , \wRegInB105[0] , 
        \wAMid69[23] , \wAIn72[28] , \wBIn105[15] , \wAIn24[29] , \wBIn30[25] , 
        \wBIn45[15] , \wAIn51[19] , \wRegInB48[28] , \wAIn72[31] , 
        \wBIn126[24] , \wBIn25[7] , \wBIn38[8] , \wAIn43[7] , \wAMid87[16] , 
        \wRegInB48[31] , \wRegInB106[3] , \wBIn88[11] , \wAMid103[15] , 
        \wAMid116[21] , \wRegInB90[18] , \wAIn40[4] , \wAIn89[30] , 
        \wAIn89[29] , \wAMid92[22] , \wAMid120[24] , \wRegInA68[1] , 
        \wBMid98[28] , \wRegInA9[27] , \ScanLink28[5] , \ScanLink116[7] , 
        \wBMid69[0] , \wAIn92[2] , \wAIn114[0] , \ScanLink84[31] , 
        \wBMid98[31] , \ScanLink84[28] , \wBIn25[22] , \wBIn30[16] , 
        \wBIn66[17] , \wAMid69[10] , \wBIn105[26] , \wBIn45[26] , \wBIn90[6] , 
        \wBIn126[17] , \wAIn27[3] , \wAMid125[9] , \wBIn50[12] , \wBIn1[2] , 
        \wBIn2[1] , \wBMid1[26] , \wAIn3[6] , \wBMid4[10] , \wAMid5[31] , 
        \wBMid13[8] , \wAMid67[7] , \wBIn73[23] , \wBIn110[12] , \wAMid5[28] , 
        \wRegInA116[24] , \ScanLink211[5] , \ScanLink187[18] , 
        \ScanLink171[0] , \wBIn41[3] , \wBIn42[0] , \wBIn107[8] , 
        \wRegInA120[21] , \wRegInA9[14] , \wRegInA12[9] , \wRegInA103[10] , 
        \ScanLink212[6] , \ScanLink109[30] , \ScanLink83[8] , 
        \ScanLink109[29] , \wAMid87[25] , \wAMid92[11] , \wAMid103[26] , 
        \ScanLink172[3] , \wAMid120[17] , \wRegInA55[31] , \wRegInA76[19] , 
        \wAIn10[1] , \wAIn24[0] , \wAMid64[4] , \wBIn88[22] , \wBIn93[5] , 
        \wRegInA55[28] , \wAMid116[12] , \wBIn119[4] , \wRegInA20[18] , 
        \wBMid39[5] , \wBIn75[2] , \ScanLink146[2] , \wAMid82[3] , 
        \wBMid88[19] , \ScanLink226[7] , \ScanLink94[19] , \ScanLink78[0] , 
        \wAMid106[10] , \wRegInA107[4] , \ScanLink194[4] , \wAIn13[2] , 
        \wBIn16[11] , \wAMid19[16] , \wBMid27[9] , \wAMid50[5] , \wAMid97[27] , 
        \wAMid125[21] , \wRegInA38[4] , \ScanLink8[26] , \wBIn98[20] , 
        \wBIn63[21] , \wAMid82[13] , \wAIn99[18] , \wRegInB58[1] , 
        \wRegInB80[30] , \wRegInB97[8] , \wAMid113[24] , \wRegInB80[29] , 
        \wBIn100[10] , \wAMid53[6] , \wBIn35[20] , \wBIn40[10] , 
        \ScanLink197[7] , \wBIn123[21] , \wAIn17[30] , \wBIn20[14] , 
        \wAIn34[18] , \wAIn41[28] , \wBIn55[24] , \wAMid111[8] , 
        \wRegInA119[8] , \wAIn17[29] , \wAIn41[31] , \wAIn62[19] , 
        \wBIn115[24] , \wBIn76[15] , \wAMid79[12] , \wRegInB58[19] , 
        \wBMid50[30] , \wBIn76[1] , \wAMid81[0] , \wRegInA113[12] , 
        \ScanLink252[19] , \ScanLink227[29] , \wRegInA26[8] , 
        \ScanLink227[30] , \ScanLink204[18] , \ScanLink145[1] , 
        \wRegInA125[17] , \wBMid73[18] , \wRegInA104[7] , \ScanLink39[19] , 
        \wBIn9[18] , \wBMid25[19] , \wRegInA106[26] , \ScanLink225[4] , 
        \wAMid34[1] , \wBMid50[29] , \wRegInB89[4] , \wAMid82[20] , 
        \wBMid104[3] , \wAIn74[5] , \wAMid113[17] , \wBMid92[8] , 
        \wAMid97[14] , \wAMid106[23] , \wRegInA45[19] , \wRegInA93[9] , 
        \wRegInA66[31] , \wRegInA30[29] , \ScanLink8[15] , \wBIn98[13] , 
        \wAMid125[12] , \wRegInA66[28] , \wRegInA13[18] , \wRegInA30[30] , 
        \wBIn11[6] , \wAIn120[1] , \ScanLink119[18] , \ScanLink242[3] , 
        \ScanLink122[6] , \wBIn2[14] , \wBMid1[15] , \wAIn123[2] , 
        \ScanLink121[5] , \wAIn4[30] , \wAIn4[29] , \wBIn12[5] , 
        \wRegInA106[15] , \wRegInA125[24] , \ScanLink197[30] , 
        \ScanLink197[29] , \wBMid8[9] , \wRegInB22[9] , \wRegInA113[21] , 
        \ScanLink241[0] , \wBIn16[22] , \wAMid19[25] , \wBIn20[27] , 
        \wAMid37[2] , \wBIn55[17] , \wAIn77[6] , \wBIn76[26] , \wBMid107[0] , 
        \wBIn115[17] , \wAMid79[21] , \wBMid22[4] , \wBIn35[13] , \wBIn63[12] , 
        \wBIn100[23] , \wBIn40[23] , \wAIn87[13] , \wAIn92[27] , \wBIn123[12] , 
        \wRegInA78[10] , \wRegInB3[0] , \wRegInA23[5] , \wRegInA18[14] , 
        \wRegInB43[0] , \ScanLink220[9] , \ScanLink3[19] , \ScanLink167[24] , 
        \wBMid18[23] , \wBMid21[7] , \wBMid78[27] , \wBMid83[26] , 
        \wAMid99[2] , \ScanLink112[14] , \wAMid114[5] , \ScanLink144[15] , 
        \ScanLink131[25] , \wBMid96[12] , \wRegInB1[18] , \ScanLink151[21] , 
        \ScanLink63[1] , \wAIn114[11] , \wRegInB91[6] , \wRegInB100[31] , 
        \wRegInB123[19] , \ScanLink124[11] , \ScanLink172[10] , 
        \wRegInB100[28] , \ScanLink107[20] , \ScanLink191[9] , \wAMid117[6] , 
        \ScanLink32[26] , \ScanLink47[16] , \wAMid55[8] , \ScanLink11[17] , 
        \wAIn101[25] , \wAIn122[14] , \ScanLink239[22] , \ScanLink64[27] , 
        \wRegInB92[5] , \ScanLink71[13] , \ScanLink189[11] , \ScanLink27[12] , 
        \ScanLink60[2] , \ScanLink52[22] , \wRegInA20[6] , \wRegInB70[17] , 
        \wBIn2[27] , \wAMid12[30] , \wAMid12[29] , \wAMid48[7] , 
        \wRegInB26[16] , \wRegInB53[26] , \wRegInA83[11] , \wAIn69[26] , 
        \wRegInB0[3] , \wAMid44[31] , \wRegInB46[12] , \wAMid67[19] , 
        \wRegInB33[22] , \wRegInB40[3] , \wRegInA96[25] , \wAMid31[18] , 
        \wAMid44[28] , \wRegInB65[23] , \wBMid46[0] , \wBMid96[21] , 
        \wRegInB10[13] , \wRegInA102[9] , \wRegInA95[7] , \ScanLink139[7] , 
        \ScanLink124[22] , \ScanLink151[12] , \wBMid89[9] , \ScanLink107[13] , 
        \ScanLink172[23] , \ScanLink167[17] , \ScanLink112[27] , \wBIn17[8] , 
        \wBMid83[15] , \ScanLink131[16] , \ScanLink144[26] , \wBIn86[18] , 
        \wAIn87[20] , \wBMid94[6] , \wRegInA18[27] , \wRegInA47[1] , 
        \ScanLink124[8] , \wRegInA88[8] , \wAIn92[14] , \wAMid118[31] , 
        \wRegInB27[4] , \wRegInA78[23] , \wBMid122[31] , \wBMid97[5] , 
        \wBMid101[19] , \wAMid118[28] , \wBMid122[28] , \wRegInB10[20] , 
        \wRegInB33[11] , \wRegInB46[21] , \wRegInA96[16] , \wRegInA44[2] , 
        \wRegInB65[10] , \ScanLink19[9] , \wAIn0[18] , \wBIn6[25] , 
        \wBIn6[16] , \wAIn18[14] , \wBMid18[10] , \wBMid45[3] , \wAIn69[15] , 
        \wRegInB26[25] , \wRegInB70[24] , \wRegInA83[22] , \wRegInB24[7] , 
        \wRegInB53[15] , \ScanLink71[20] , \wAIn122[27] , \ScanLink189[22] , 
        \ScanLink52[11] , \wAIn48[1] , \wAIn71[8] , \wAIn78[10] , 
        \wBMid78[14] , \wAIn101[16] , \wRegInA96[4] , \ScanLink27[21] , 
        \wAIn114[22] , \ScanLink47[25] , \wRegInB39[8] , \ScanLink239[11] , 
        \ScanLink32[15] , \ScanLink64[14] , \wRegInB42[10] , \ScanLink11[24] , 
        \wBIn79[31] , \wAIn87[8] , \wRegInB14[11] , \wRegInB37[20] , 
        \wRegInB61[21] , \wRegInA92[27] , \wRegInB74[15] , \wRegInA60[4] , 
        \wRegInB57[24] , \wBMid61[5] , \wBMid69[11] , \wBIn79[28] , 
        \wRegInB22[14] , \wRegInA87[13] , \wAIn126[16] , \wRegInB113[9] , 
        \ScanLink228[14] , \ScanLink75[11] , \ScanLink23[10] , \wAIn105[27] , 
        \ScanLink20[0] , \wAIn110[13] , \ScanLink56[20] , \ScanLink43[14] , 
        \ScanLink36[24] , \wBMid62[6] , \wBMid92[10] , \wBMid125[8] , 
        \ScanLink248[10] , \ScanLink198[27] , \ScanLink15[15] , 
        \ScanLink155[23] , \ScanLink60[25] , \ScanLink23[3] , 
        \ScanLink176[12] , \ScanLink120[13] , \ScanLink163[26] , 
        \ScanLink103[22] , \wAIn8[0] , \wAMid16[18] , \wAMid16[9] , 
        \ScanLink116[16] , \wAIn18[27] , \wBIn49[6] , \wBIn82[30] , 
        \wBIn82[29] , \wAIn83[11] , \wBMid87[24] , \ScanLink140[17] , 
        \ScanLink135[27] , \wAIn99[4] , \wBMid105[28] , \wRegInA69[26] , 
        \wAIn96[25] , \wAIn102[9] , \wBMid105[31] , \wAIn110[20] , 
        \wBMid126[19] , \wRegInA63[7] , \wRegInA109[31] , \ScanLink44[4] , 
        \ScanLink43[27] , \wAIn126[25] , \wRegInA109[28] , \ScanLink198[14] , 
        \ScanLink36[17] , \ScanLink248[23] , \ScanLink60[16] , 
        \ScanLink228[27] , \ScanLink75[22] , \ScanLink15[26] , \ScanLink5[8] , 
        \ScanLink56[13] , \wBMid69[22] , \ScanLink23[23] , \wAIn105[14] , 
        \wRegInB22[27] , \wRegInB74[26] , \ScanLink96[2] , \wRegInA87[20] , 
        \wRegInB57[17] , \wRegInB64[5] , \wAMid35[30] , \wAMid63[28] , 
        \wAIn78[23] , \wRegInB37[13] , \wRegInA92[14] , \wAMid35[29] , 
        \wAMid40[19] , \wAMid63[31] , \wRegInB42[23] , \ScanLink167[9] , 
        \wBIn54[9] , \wRegInB14[22] , \wAIn96[16] , \wBIn111[1] , 
        \wRegInB61[12] , \wBIn98[3] , \wRegInB67[6] , \ScanLink95[1] , 
        \wAMid98[30] , \wBIn112[2] , \ScanLink7[31] , \wAIn83[22] , 
        \wAMid98[29] , \ScanLink7[28] , \wRegInA69[15] , \ScanLink219[0] , 
        \ScanLink116[25] , \ScanLink163[15] , \wBMid5[24] , \wAIn32[9] , 
        \wBMid87[17] , \ScanLink135[14] , \ScanLink47[7] , \wBMid92[23] , 
        \ScanLink140[24] , \wRegInB127[28] , \wRegInB5[29] , \ScanLink179[5] , 
        \ScanLink120[20] , \ScanLink155[10] , \wRegInB127[31] , \wRegInB5[30] , 
        \wRegInB104[19] , \ScanLink103[11] , \wRegInA121[15] , 
        \ScanLink176[21] , \wRegInA102[24] , \ScanLink193[18] , 
        \wRegInB108[8] , \wRegInA117[10] , \wAIn5[5] , \wBMid5[17] , 
        \wAMid10[7] , \wBIn12[13] , \wBIn24[16] , \wBIn36[3] , \wBIn51[26] , 
        \wAIn81[6] , \wAIn107[4] , \ScanLink105[3] , \wBIn67[23] , 
        \wAMid68[24] , \wBIn72[17] , \wBIn111[26] , \wRegInB115[7] , 
        \wBIn104[12] , \wBMid123[6] , \wRegInA99[18] , \wAMid13[4] , 
        \wBIn31[22] , \wBIn44[12] , \wBIn127[23] , \wAIn50[3] , \wAIn53[0] , 
        \wAMid86[11] , \wBIn89[16] , \wRegInB18[3] , \wRegInB116[4] , 
        \wAMid102[12] , \wAMid117[26] , \wAIn119[8] , \wRegInA17[30] , 
        \wRegInA34[18] , \wBMid64[8] , \wBMid120[5] , \wAMid121[23] , 
        \wRegInA41[28] , \wRegInA78[6] , \wRegInA17[29] , \wAMid93[25] , 
        \wRegInA62[19] , \wBIn12[20] , \wBIn35[0] , \wRegInA8[20] , 
        \wRegInA41[31] , \ScanLink168[19] , \ScanLink106[0] , \ScanLink38[2] , 
        \wBMid79[7] , \wAIn82[5] , \wAIn104[7] , \wRegInA65[9] , \wAIn13[18] , 
        \wBIn24[25] , \wBIn31[11] , \wBIn67[10] , \wAMid68[17] , 
        \ScanLink3[6] , \wBIn104[21] , \wBIn44[21] , \wBIn80[1] , 
        \wBIn127[10] , \wAIn30[29] , \wAIn37[4] , \wAIn45[19] , \wBIn51[15] , 
        \wAIn66[31] , \wAIn30[30] , \wAIn66[28] , \wBIn72[24] , \wAMid77[0] , 
        \wBIn111[15] , \wRegInB29[18] , \wRegInA117[23] , \ScanLink256[28] , 
        \ScanLink201[2] , \wRegInA120[1] , \ScanLink256[31] , 
        \ScanLink223[18] , \ScanLink200[30] , \ScanLink200[29] , 
        \ScanLink161[7] , \wBMid16[8] , \wBMid21[31] , \wBIn52[7] , 
        \wBMid77[29] , \wRegInA121[26] , \wBMid21[28] , \wBMid54[18] , 
        \wBMid77[30] , \ScanLink48[18] , \wAIn29[8] , \wBIn51[4] , 
        \wRegInA8[13] , \wRegInB61[8] , \wRegInA102[17] , \wRegInA123[2] , 
        \ScanLink202[1] , \ScanLink90[28] , \ScanLink162[4] , \ScanLink90[31] , 
        \wAIn34[7] , \wAMid74[3] , \wAMid86[22] , \wBIn89[25] , \wAMid93[16] , 
        \wAMid102[21] , \ScanLink41[9] , \wAMid121[10] , \ScanLink0[5] , 
        \wBIn83[2] , \wBIn109[3] , \wRegInB84[18] , \wAMid117[15] , 
        \wRegInA2[26] , \wRegInB110[27] , \ScanLink98[4] , \wBMid93[30] , 
        \wAIn6[6] , \wAMid17[12] , \wBIn18[15] , \wAMid21[17] , \wAIn22[3] , 
        \wAMid62[7] , \wRegInB105[13] , \wBMid93[29] , \wRegInB4[23] , 
        \wBIn95[6] , \wRegInB126[22] , \wAMid120[9] , \wBIn47[0] , 
        \wAIn82[28] , \wBIn83[10] , \ScanLink214[5] , \wBMid104[11] , 
        \wBIn96[24] , \wBMid111[25] , \wAMid99[23] , \ScanLink6[22] , 
        \wAMid108[14] , \wAMid54[27] , \wAMid77[16] , \wAIn82[31] , 
        \wBIn88[9] , \ScanLink174[0] , \wBIn102[8] , \wRegInA17[9] , 
        \wBIn78[11] , \ScanLink217[6] , \ScanLink49[1] , \ScanLink86[8] , 
        \wAMid34[23] , \wAMid41[13] , \wBIn44[3] , \wAIn79[30] , 
        \wRegInB15[28] , \ScanLink177[3] , \wAMid62[22] , \wAIn79[29] , 
        \wRegInB43[30] , \wRegInB60[18] , \wRegInB15[31] , \wRegInB36[19] , 
        \wAIn21[0] , \wBMid68[28] , \wBIn96[5] , \wRegInB43[29] , 
        \wRegInB69[0] , \wRegInA108[22] , \ScanLink249[29] , \ScanLink249[30] , 
        \ScanLink74[31] , \ScanLink57[19] , \ScanLink22[29] , \wBIn23[4] , 
        \wAMid61[4] , \wBMid68[31] , \ScanLink74[28] , \ScanLink22[30] , 
        \wBIn96[17] , \wBMid111[16] , \wAMid99[10] , \ScanLink6[11] , 
        \wAMid108[27] , \wRegInB13[8] , \ScanLink110[4] , \wAIn46[7] , 
        \wBIn83[23] , \wAIn94[1] , \wAIn112[3] , \wBMid104[22] , 
        \wRegInB4[10] , \wRegInB100[0] , \ScanLink177[18] , \ScanLink154[30] , 
        \wRegInB105[20] , \ScanLink102[28] , \ScanLink154[29] , 
        \ScanLink33[9] , \wRegInB126[11] , \ScanLink102[31] , 
        \ScanLink121[19] , \wRegInA2[15] , \wRegInB110[14] , \wAIn0[8] , 
        \wAIn1[21] , \wAMid5[25] , \wBMid10[6] , \wAMid17[21] , \wBIn18[26] , 
        \wAMid34[10] , \wAIn45[4] , \wAIn111[19] , \wRegInB103[3] , 
        \wRegInA108[11] , \wAMid41[20] , \wBIn20[7] , \wAMid62[11] , 
        \wAMid77[25] , \wRegInA86[19] , \wBIn78[22] , \wAMid21[24] , 
        \wAIn111[0] , \ScanLink113[7] , \wAMid54[14] , \wAIn97[2] , 
        \wAMid87[31] , \wAIn89[17] , \wBIn93[8] , \wRegInA16[10] , 
        \wRegInA63[20] , \wRegInA35[21] , \wRegInA40[11] , \ScanLink51[3] , 
        \wRegInA55[25] , \wRegInB90[26] , \wBIn119[9] , \wAMid126[7] , 
        \wRegInA20[15] , \wRegInB85[12] , \wRegInA76[14] , \wAIn39[2] , 
        \wAMid64[9] , \wAMid87[28] , \wBMid98[16] , \wRegInB71[2] , 
        \ScanLink109[24] , \ScanLink84[16] , \ScanLink83[5] , \wBIn104[6] , 
        \wRegInA11[7] , \wBMid63[17] , \wAMid79[6] , \ScanLink169[20] , 
        \ScanLink91[22] , \wRegInA1[2] , \wRegInA9[19] , \ScanLink29[16] , 
        \wBMid16[27] , \ScanLink80[6] , \wBMid40[26] , \wRegInA116[30] , 
        \ScanLink201[23] , \wBMid20[22] , \wBMid35[16] , \wRegInB72[1] , 
        \ScanLink211[8] , \wBMid55[12] , \wRegInA116[29] , \ScanLink242[16] , 
        \ScanLink222[12] , \ScanLink187[15] , \wRegInA2[1] , \ScanLink237[26] , 
        \ScanLink192[21] , \wAIn24[17] , \wBMid76[23] , \wBIn107[5] , 
        \wRegInA12[4] , \ScanLink214[17] , \ScanLink49[12] , \ScanLink52[0] , 
        \wAIn51[27] , \wAIn72[16] , \wRegInB48[16] , \wRegInA98[21] , 
        \wAIn0[1] , \wAIn1[31] , \wAIn1[12] , \wAMid5[16] , \wAIn12[21] , 
        \wAIn12[12] , \wBMid13[5] , \wAIn31[23] , \wAIn67[22] , 
        \wRegInB28[12] , \wBIn38[5] , \wAIn44[13] , \wAMid125[4] , 
        \wBMid74[2] , \wBMid98[25] , \wRegInB15[6] , \ScanLink28[8] , 
        \ScanLink169[13] , \ScanLink109[17] , \ScanLink91[11] , 
        \ScanLink84[25] , \wAMid120[29] , \wRegInA20[26] , \wRegInA75[3] , 
        \wRegInB85[21] , \wRegInA55[16] , \ScanLink35[7] , \wRegInA76[27] , 
        \wAIn89[24] , \wRegInA16[23] , \wAMid103[18] , \wRegInA63[13] , 
        \wAMid120[30] , \wAIn40[9] , \wAIn109[2] , \wRegInA35[12] , 
        \wRegInB90[15] , \wAIn67[11] , \wRegInB28[21] , \wRegInA40[22] , 
        \wBIn13[19] , \wAIn24[24] , \wAIn31[10] , \wAIn44[20] , 
        \ScanLink36[4] , \wBIn45[18] , \wAIn51[14] , \wBIn66[30] , 
        \wBIn126[29] , \ScanLink108[6] , \wBIn30[28] , \wBIn66[29] , 
        \wAIn72[25] , \wBMid77[1] , \wBIn105[18] , \wBIn126[30] , 
        \wRegInA98[12] , \wBMid16[14] , \wBMid20[11] , \wBIn30[31] , 
        \wRegInB48[25] , \ScanLink237[15] , \ScanLink192[12] , \wBMid55[21] , 
        \ScanLink242[25] , \wBMid76[10] , \wRegInB16[5] , \wRegInB118[2] , 
        \ScanLink214[24] , \ScanLink49[21] , \wBIn26[9] , \ScanLink201[10] , 
        \ScanLink115[9] , \wBMid35[25] , \wBMid63[24] , \wRegInA76[0] , 
        \ScanLink29[25] , \wBMid40[15] , \ScanLink222[21] , \ScanLink187[26] , 
        \wBMid0[1] , \wAMid1[27] , \wAIn16[10] , \wRegInB59[20] , \wBIn17[31] , 
        \wAMid27[8] , \wBMid53[7] , \wAIn63[20] , \wRegInA89[17] , 
        \wBIn34[19] , \wAIn35[21] , \wAIn40[11] , \wRegInA80[0] , 
        \ScanLink12[2] , \wBIn17[28] , \wAIn20[15] , \wBIn41[29] , 
        \wAIn55[25] , \wBIn101[30] , \wBIn122[18] , \wBMid24[20] , 
        \wBIn41[30] , \wBIn62[18] , \wBMid51[10] , \wAIn76[14] , \wBMid81[1] , 
        \wBIn101[29] , \wRegInB39[24] , \ScanLink246[14] , \ScanLink233[24] , 
        \ScanLink196[23] , \wBMid67[15] , \wBMid72[21] , \wRegInA52[6] , 
        \ScanLink210[15] , \ScanLink38[20] , \wAMid1[14] , \wAIn5[23] , 
        \wBMid12[25] , \ScanLink58[24] , \wBMid44[24] , \ScanLink205[21] , 
        \ScanLink253[20] , \wBIn8[12] , \wBMid31[14] , \wAIn79[0] , 
        \wRegInB32[3] , \wRegInA51[5] , \ScanLink226[10] , \ScanLink183[17] , 
        \wBMid89[20] , \wBMid109[6] , \wBMid12[16] , \wAMid39[4] , 
        \wBMid82[2] , \ScanLink95[20] , \wBMid50[4] , \wRegInA24[17] , 
        \wRegInB31[0] , \ScanLink252[9] , \ScanLink118[12] , \ScanLink178[16] , 
        \ScanLink80[14] , \wRegInA51[27] , \wRegInB81[10] , \wRegInA83[3] , 
        \wAIn98[21] , \wBMid114[9] , \wRegInA72[16] , \wBIn99[19] , 
        \wAMid107[30] , \wAMid124[18] , \wRegInA67[22] , \wAMid107[29] , 
        \wRegInA12[12] , \wRegInB122[8] , \wRegInA44[13] , \ScanLink11[1] , 
        \wRegInA31[23] , \wRegInB94[24] , \ScanLink58[17] , \ScanLink205[12] , 
        \wBMid3[2] , \wAIn5[10] , \wBMid31[27] , \wBMid67[26] , \wBIn123[3] , 
        \wRegInA36[2] , \wRegInA112[18] , \wBMid44[17] , \ScanLink226[23] , 
        \ScanLink183[24] , \ScanLink253[13] , \wAMid7[8] , \wAIn16[23] , 
        \wAIn20[26] , \wBMid24[13] , \ScanLink233[17] , \ScanLink196[10] , 
        \wBMid51[23] , \wRegInB56[7] , \ScanLink246[27] , \wAIn55[16] , 
        \wBMid72[12] , \ScanLink210[26] , \ScanLink38[13] , \ScanLink148[4] , 
        \wBMid37[3] , \wAMid101[2] , \wAIn63[13] , \wAIn76[27] , \wAMid78[18] , 
        \wRegInB39[17] , \wRegInA89[24] , \ScanLink228[1] , \wRegInB59[13] , 
        \wRegInB84[1] , \wAIn35[12] , \wAIn40[22] , \ScanLink76[6] , 
        \wBMid34[0] , \wRegInA12[21] , \wRegInA109[2] , \wBIn65[8] , 
        \wBIn78[7] , \wRegInA67[11] , \wAMid83[19] , \wAMid102[1] , 
        \wRegInA31[10] , \wRegInB94[17] , \wRegInA24[24] , \wRegInA44[20] , 
        \wRegInB81[23] , \wRegInA51[14] , \ScanLink75[5] , \wRegInA72[25] , 
        \wAMid92[9] , \wAIn98[12] , \wRegInB87[2] , \ScanLink199[1] , 
        \ScanLink178[25] , \ScanLink80[27] , \ScanLink156[8] , \wBMid89[13] , 
        \wBIn120[0] , \wRegInA35[1] , \wBIn8[21] , \wRegInB55[4] , 
        \ScanLink118[21] , \ScanLink95[13] , \wAMid21[6] , \wBMid55[9] , 
        \wAIn61[2] , \ScanLink188[31] , \wBMid111[4] , \wRegInA49[7] , 
        \wRegInA119[14] , \ScanLink188[28] , \wAIn115[31] , \wRegInB127[5] , 
        \wRegInB29[2] , \wAMid13[10] , \wAMid30[21] , \wAMid45[11] , 
        \wAIn115[28] , \ScanLink137[1] , \wBMid48[6] , \wAMid66[20] , 
        \wBIn69[27] , \wRegInA54[8] , \wAMid22[5] , \wAMid25[15] , 
        \wAMid50[25] , \wAMid73[14] , \wRegInA82[28] , \wRegInA82[31] , 
        \wBIn87[12] , \wAMid88[15] , \wBIn92[26] , \ScanLink2[20] , 
        \wBMid115[27] , \wAMid119[22] , \wRegInA98[2] , \ScanLink134[2] , 
        \wBMid123[22] , \wRegInA79[30] , \wRegInA79[29] , \ScanLink254[7] , 
        \wBMid100[13] , \wBMid99[3] , \wBMid112[7] , \ScanLink125[31] , 
        \wRegInB101[11] , \ScanLink106[19] , \wAIn62[1] , \wRegInB0[21] , 
        \ScanLink173[29] , \wRegInB122[20] , \ScanLink125[28] , 
        \ScanLink173[30] , \ScanLink150[18] , \wRegInA6[24] , \wRegInB114[25] , 
        \ScanLink249[8] , \wAMid1[6] , \wAMid2[5] , \wAMid13[23] , \wAIn18[9] , 
        \wAMid25[26] , \wBIn60[5] , \wAMid73[27] , \wRegInB124[6] , 
        \wAMid97[4] , \ScanLink153[5] , \wAMid50[16] , \wAMid30[12] , 
        \wAMid45[22] , \wRegInB64[29] , \wRegInB11[19] , \wRegInB32[31] , 
        \wRegInA112[3] , \ScanLink233[0] , \wRegInB64[30] , \wBMid19[30] , 
        \wBMid19[29] , \wAMid45[2] , \wAMid66[13] , \wBIn69[14] , 
        \wRegInB47[18] , \wRegInB32[28] , \wRegInB50[9] , \ScanLink238[28] , 
        \ScanLink238[31] , \ScanLink181[3] , \ScanLink70[8] , \ScanLink26[18] , 
        \wRegInA119[27] , \ScanLink70[19] , \ScanLink53[28] , \wAMid46[1] , 
        \wAMid89[8] , \ScanLink182[0] , \ScanLink53[31] , \wRegInA6[17] , 
        \wRegInB114[16] , \wBIn63[6] , \wBMid97[18] , \wRegInB101[22] , 
        \wBMid123[11] , \wRegInB0[12] , \wRegInB122[13] , \ScanLink150[6] , 
        \wBIn87[21] , \wAMid88[26] , \wAMid119[11] , \wAMid119[0] , 
        \wBMid100[20] , \wBIn92[15] , \wAMid94[7] , \ScanLink2[13] , 
        \wBMid115[14] , \wAIn3[2] , \wBMid4[27] , \wAIn12[31] , \wAIn12[28] , 
        \wBIn13[10] , \wBIn25[3] , \wBMid69[4] , \wAIn86[19] , \wRegInA111[0] , 
        \ScanLink230[3] , \ScanLink116[3] , \wBIn30[21] , \wAIn40[0] , 
        \wAIn92[6] , \wAIn114[4] , \wAMid92[26] , \wAMid120[20] , 
        \wRegInA9[23] , \ScanLink28[1] , \ScanLink91[18] , \wAMid103[11] , 
        \wBIn45[11] , \wAMid87[12] , \wBIn88[15] , \wAMid116[25] , 
        \wRegInA68[5] , \wRegInB85[28] , \wRegInB85[31] , \wRegInB106[7] , 
        \wBIn126[20] , \wAIn43[3] , \wBIn66[20] , \wAMid69[27] , \wBMid77[8] , 
        \wBIn105[11] , \wAIn44[30] , \wAIn67[18] , \wBIn110[25] , 
        \wRegInB28[28] , \wBIn73[14] , \wAIn31[19] , \wAIn44[29] , 
        \wBIn50[25] , \wRegInB28[31] , \wRegInB105[4] , \wBMid20[18] , 
        \wBIn25[15] , \wBIn26[0] , \wAIn91[5] , \wAIn117[7] , \wRegInA76[9] , 
        \ScanLink222[31] , \ScanLink201[19] , \ScanLink115[0] , 
        \wRegInA103[27] , \wRegInA116[13] , \ScanLink222[28] , 
        \ScanLink49[31] , \wBMid55[31] , \wBMid55[28] , \wRegInA120[16] , 
        \ScanLink49[28] , \wAIn24[4] , \wBMid76[19] , \wBIn93[1] , 
        \wBIn119[0] , \wBIn88[26] , \wAMid116[16] , \wBMid4[14] , \wBIn41[7] , 
        \wAMid64[0] , \wAMid87[21] , \wAMid92[15] , \wAMid103[22] , 
        \wAMid120[13] , \wRegInA63[29] , \wRegInA16[19] , \wRegInA35[31] , 
        \wRegInA40[18] , \wRegInA63[30] , \wRegInA35[28] , \ScanLink169[30] , 
        \wRegInA2[8] , \wRegInA9[10] , \ScanLink172[7] , \ScanLink169[29] , 
        \ScanLink212[2] , \wRegInA103[14] , \ScanLink192[28] , 
        \ScanLink171[4] , \wBIn42[4] , \wRegInA120[25] , \ScanLink192[31] , 
        \wAIn1[28] , \ScanLink211[1] , \wRegInB72[8] , \wRegInA116[20] , 
        \wBMid0[25] , \wBMid0[8] , \wBIn3[17] , \wBIn7[26] , \wBIn7[15] , 
        \wBIn13[23] , \wBIn25[26] , \wAMid67[3] , \wBIn110[16] , \wBIn73[27] , 
        \wBIn90[2] , \wAIn27[7] , \wBIn30[12] , \wBIn50[16] , \ScanLink52[9] , 
        \wBIn45[22] , \wBIn126[13] , \wRegInA98[31] , \wBIn66[13] , 
        \wAMid69[14] , \wBMid72[5] , \wAIn82[12] , \wAIn94[8] , \wBIn105[22] , 
        \wRegInA98[28] , \wRegInA73[4] , \wAIn97[26] , \wBMid86[27] , 
        \wAMid99[19] , \wRegInB13[1] , \wRegInA68[25] , \ScanLink6[18] , 
        \ScanLink141[14] , \ScanLink134[24] , \wAIn89[7] , \ScanLink162[25] , 
        \wBMid16[1] , \wAMid17[31] , \wAMid18[6] , \wAIn19[17] , \wBMid68[12] , 
        \wBMid71[6] , \wBMid93[13] , \wRegInB100[9] , \ScanLink177[11] , 
        \ScanLink117[15] , \wRegInB105[29] , \ScanLink154[20] , 
        \ScanLink102[21] , \ScanLink33[0] , \wRegInB4[19] , \wRegInB105[30] , 
        \wRegInB126[18] , \ScanLink121[10] , \wAIn111[10] , \wRegInA108[18] , 
        \ScanLink249[13] , \ScanLink199[24] , \ScanLink14[16] , 
        \ScanLink61[26] , \ScanLink42[17] , \ScanLink37[27] , \ScanLink22[13] , 
        \wAIn104[24] , \ScanLink30[3] , \wAIn127[15] , \ScanLink57[23] , 
        \wRegInB56[27] , \ScanLink229[17] , \ScanLink74[12] , \wRegInB23[17] , 
        \wRegInA86[10] , \wAIn58[2] , \wAIn111[9] , \wRegInA70[7] , 
        \wRegInB75[16] , \wAMid17[28] , \wAMid34[19] , \wAMid41[29] , 
        \wRegInB60[22] , \wRegInB15[12] , \wAMid41[30] , \wAIn79[13] , 
        \wRegInB43[13] , \wAMid62[18] , \wRegInB10[2] , \wRegInB36[23] , 
        \wRegInA93[24] , \wBMid86[14] , \wBMid93[20] , \ScanLink177[22] , 
        \ScanLink102[12] , \wAMid120[0] , \ScanLink169[6] , \ScanLink154[13] , 
        \ScanLink121[23] , \ScanLink134[17] , \ScanLink57[4] , 
        \ScanLink209[3] , \ScanLink141[27] , \ScanLink117[26] , 
        \ScanLink162[16] , \wBMid15[2] , \wAIn19[24] , \wBIn47[9] , 
        \wAIn82[21] , \wRegInA7[5] , \wRegInA68[16] , \wBIn78[18] , 
        \wAIn79[20] , \wBIn83[19] , \wBIn88[0] , \ScanLink174[9] , 
        \wAIn97[15] , \wBIn102[1] , \wRegInA17[0] , \ScanLink85[2] , 
        \wBMid104[18] , \wRegInB77[5] , \wBIn101[2] , \wRegInA14[3] , 
        \wRegInB15[21] , \wRegInB60[11] , \wRegInA4[6] , \wRegInB36[10] , 
        \wRegInA93[17] , \wRegInB23[24] , \wRegInB43[20] , \wRegInA86[23] , 
        \wRegInB56[14] , \wRegInB74[6] , \ScanLink8[4] , \wAIn21[9] , 
        \wBIn59[5] , \wRegInB75[25] , \ScanLink86[1] , \ScanLink49[8] , 
        \ScanLink57[10] , \ScanLink22[20] , \wBMid68[21] , \wAIn104[17] , 
        \wAMid123[3] , \ScanLink229[24] , \ScanLink74[21] , \wAIn18[0] , 
        \wAMid58[4] , \wAIn111[23] , \wAIn127[26] , \wRegInB69[9] , 
        \ScanLink199[17] , \ScanLink61[15] , \ScanLink249[20] , 
        \ScanLink54[7] , \ScanLink14[25] , \ScanLink42[24] , \wRegInB11[10] , 
        \wRegInB64[20] , \ScanLink37[14] , \wRegInB27[15] , \wRegInB32[21] , 
        \wRegInB47[11] , \ScanLink233[9] , \wRegInA97[26] , \wRegInB50[0] , 
        \wRegInB52[25] , \wRegInA82[12] , \wAIn68[25] , \wBIn125[4] , 
        \wRegInB71[14] , \wRegInA30[5] , \wBMid19[20] , \wAIn100[26] , 
        \ScanLink26[11] , \ScanLink70[1] , \ScanLink53[21] , \wBMid31[4] , 
        \wAIn123[17] , \wRegInB82[6] , \ScanLink70[10] , \ScanLink188[12] , 
        \wBMid32[7] , \wBMid79[24] , \wAIn115[12] , \ScanLink238[21] , 
        \ScanLink10[14] , \ScanLink65[24] , \wBMid82[25] , \wBMid97[11] , 
        \wAMid107[5] , \ScanLink33[25] , \wRegInB81[5] , \ScanLink173[13] , 
        \ScanLink46[15] , \ScanLink150[22] , \ScanLink106[23] , 
        \ScanLink73[2] , \wAMid104[6] , \ScanLink182[9] , \ScanLink145[16] , 
        \ScanLink125[12] , \ScanLink130[26] , \ScanLink166[27] , \wAMid13[19] , 
        \wBIn19[7] , \wBMid19[13] , \wAMid46[8] , \wAMid89[1] , 
        \ScanLink113[17] , \wBMid79[17] , \wAIn86[10] , \wBIn87[31] , 
        \wRegInA19[17] , \wRegInB53[3] , \wRegInA111[9] , \wBIn87[28] , 
        \wBMid100[30] , \wAMid119[18] , \wAMid119[9] , \wBMid123[18] , 
        \wBIn126[7] , \wRegInA33[6] , \wRegInA79[13] , \wAIn93[24] , 
        \wBMid100[29] , \wAIn115[21] , \ScanLink238[12] , \ScanLink65[17] , 
        \ScanLink46[26] , \ScanLink14[5] , \ScanLink10[27] , \ScanLink53[12] , 
        \ScanLink33[16] , \wAMid30[31] , \wAMid30[28] , \wAMid45[18] , 
        \wBMid55[0] , \wAIn100[15] , \wRegInA86[7] , \ScanLink26[22] , 
        \ScanLink188[21] , \ScanLink70[23] , \wAMid66[30] , \wAIn68[16] , 
        \wAIn123[24] , \wRegInB27[26] , \wRegInA82[21] , \wRegInB34[4] , 
        \wRegInB52[16] , \wRegInB71[27] , \ScanLink137[8] , \wRegInB11[23] , 
        \wAMid66[29] , \wRegInA54[1] , \wRegInB64[13] , \wBMid87[6] , 
        \wRegInB32[12] , \wRegInA97[15] , \wBMid82[16] , \wBMid84[5] , 
        \wAIn93[17] , \wRegInB37[7] , \wRegInB47[22] , \wRegInA79[20] , 
        \wRegInA19[24] , \wAIn86[23] , \ScanLink2[29] , \wRegInA57[2] , 
        \ScanLink130[15] , \ScanLink2[30] , \ScanLink17[6] , \ScanLink249[1] , 
        \ScanLink145[25] , \ScanLink166[14] , \ScanLink113[24] , \wBIn3[24] , 
        \wAMid4[2] , \wBIn9[3] , \wBMid56[3] , \wRegInB0[31] , \wBMid97[22] , 
        \wRegInB0[28] , \wRegInB101[18] , \ScanLink106[10] , \wRegInB122[30] , 
        \ScanLink173[20] , \wAIn62[8] , \wRegInA85[4] , \wRegInB122[29] , 
        \ScanLink129[4] , \ScanLink125[21] , \wRegInA107[25] , 
        \ScanLink235[7] , \ScanLink196[19] , \ScanLink150[11] , \wRegInB99[7] , 
        \wRegInA114[4] , \wRegInA124[14] , \wBMid0[16] , \wAIn5[19] , 
        \wBIn66[2] , \wRegInA112[11] , \ScanLink155[2] , \wBMid5[5] , 
        \wAMid7[1] , \wBIn8[31] , \wBIn17[12] , \wAMid18[15] , \wBIn21[17] , 
        \wBIn54[27] , \wBIn77[16] , \wAMid91[3] , \wBIn114[27] , 
        \ScanLink228[8] , \wAMid78[11] , \wRegInB84[8] , \wBIn34[23] , 
        \wBIn41[13] , \ScanLink187[4] , \wBIn122[22] , \wAMid43[5] , 
        \wBIn62[22] , \wBIn101[13] , \wBMid34[9] , \wAMid83[10] , 
        \wAMid112[27] , \wRegInB48[2] , \wAMid124[22] , \wAMid40[6] , 
        \wAMid96[24] , \wRegInA12[28] , \ScanLink9[25] , \wBIn99[23] , 
        \wRegInB8[2] , \wRegInA67[18] , \wAMid102[8] , \wAMid107[13] , 
        \wRegInA44[30] , \wRegInA12[31] , \wRegInA31[19] , \ScanLink184[7] , 
        \wRegInA28[7] , \wRegInA44[29] , \wRegInA117[7] , \ScanLink118[31] , 
        \ScanLink68[3] , \ScanLink118[28] , \wBIn8[28] , \ScanLink236[4] , 
        \wBIn17[21] , \wAMid18[26] , \wBMid29[6] , \wBIn34[10] , \wBIn65[1] , 
        \wAMid92[0] , \ScanLink156[1] , \wBIn120[9] , \wRegInA35[8] , 
        \ScanLink199[8] , \wBIn41[20] , \wBIn122[11] , \wBIn62[11] , 
        \wRegInB121[2] , \wAIn16[19] , \wBIn101[20] , \wBMid117[3] , 
        \wRegInB59[29] , \wBIn21[24] , \wAMid27[1] , \wAIn35[31] , 
        \wBIn77[25] , \wBIn114[14] , \wAIn63[29] , \wAMid78[22] , 
        \wRegInB59[30] , \wBMid24[29] , \wAIn35[28] , \wAIn40[18] , 
        \wAIn67[5] , \wRegInA80[9] , \wBMid51[19] , \wBIn54[14] , \wAIn63[30] , 
        \wBMid72[31] , \wBMid81[8] , \wRegInA112[22] , \ScanLink253[30] , 
        \ScanLink253[29] , \ScanLink251[3] , \ScanLink205[28] , 
        \ScanLink226[19] , \ScanLink205[31] , \ScanLink38[30] , \wBMid72[28] , 
        \wRegInA107[16] , \ScanLink131[6] , \ScanLink38[29] , \wBIn4[6] , 
        \wBMid6[6] , \wBMid24[30] , \wAIn79[9] , \wBMid89[29] , \wRegInB31[9] , 
        \wRegInA124[27] , \ScanLink252[0] , \ScanLink132[5] , \ScanLink95[30] , 
        \wBMid89[30] , \ScanLink95[29] , \wAMid96[17] , \ScanLink9[16] , 
        \wBIn99[10] , \wBIn17[1] , \wAMid24[2] , \wAIn64[6] , \wAIn98[31] , 
        \wAMid107[20] , \wAMid124[11] , \wRegInB122[1] , \ScanLink11[8] , 
        \wRegInB81[19] , \wAMid83[23] , \wAMid112[14] , \wBMid114[0] , 
        \wAIn98[28] , \wAMid32[6] , \wBMid46[9] , \wAIn72[2] , \wBMid96[28] , 
        \wRegInA7[27] , \wRegInB115[26] , \wRegInB1[22] , \wRegInB123[23] , 
        \wBMid102[4] , \wBMid89[0] , \wBMid96[31] , \wRegInB100[12] , 
        \wBIn86[11] , \wAMid89[16] , \ScanLink244[4] , \wBMid101[10] , 
        \wAMid118[21] , \wBMid122[21] , \wAIn126[6] , \wBIn7[5] , 
        \wAMid12[13] , \wAMid24[16] , \wAMid51[26] , \wAIn87[30] , 
        \ScanLink124[1] , \wAIn87[29] , \wRegInA47[8] , \wRegInA88[1] , 
        \wBIn93[25] , \ScanLink3[23] , \wBMid114[24] , \ScanLink19[0] , 
        \wBMid58[5] , \wAMid67[23] , \wBIn68[24] , \wAMid72[17] , 
        \ScanLink247[7] , \wRegInB10[30] , \wRegInB33[18] , \wAMid44[12] , 
        \wRegInB46[28] , \wBIn14[2] , \wAIn125[5] , \ScanLink127[2] , 
        \wRegInB10[29] , \wBMid18[19] , \wAMid31[22] , \wAMid31[5] , 
        \wBMid101[7] , \wRegInB39[1] , \wRegInB46[31] , \wRegInB65[19] , 
        \ScanLink239[18] , \wRegInA118[17] , \ScanLink71[29] , 
        \ScanLink27[31] , \wAIn71[1] , \ScanLink71[30] , \ScanLink52[18] , 
        \ScanLink27[28] , \wBIn73[5] , \wAMid84[4] , \wBIn86[22] , 
        \wAMid89[25] , \wBIn93[16] , \wRegInA59[4] , \wRegInA101[3] , 
        \ScanLink3[10] , \wBMid114[17] , \wRegInB43[9] , \ScanLink220[0] , 
        \wRegInA78[19] , \wBMid101[23] , \wBMid122[12] , \wRegInB3[9] , 
        \ScanLink140[5] , \wAMid109[3] , \wAMid118[12] , \wRegInB1[11] , 
        \ScanLink151[28] , \ScanLink63[8] , \wRegInB100[21] , \wRegInB123[10] , 
        \ScanLink124[18] , \ScanLink107[30] , \ScanLink172[19] , 
        \ScanLink151[31] , \ScanLink107[29] , \wAMid0[24] , \wBIn2[8] , 
        \wBIn9[11] , \wAMid12[20] , \wAIn15[5] , \wAIn16[6] , \wAMid56[2] , 
        \wRegInA7[14] , \wRegInB115[15] , \ScanLink192[3] , \wAIn114[18] , 
        \wRegInA118[24] , \ScanLink191[0] , \ScanLink189[18] , \wAMid55[1] , 
        \ScanLink223[3] , \wAMid24[25] , \wAMid31[11] , \wAMid67[10] , 
        \wBIn68[17] , \wAMid44[21] , \wBIn70[6] , \wRegInA102[0] , 
        \ScanLink143[6] , \wAMid34[8] , \wBMid40[7] , \wAMid51[15] , 
        \wAMid72[24] , \wRegInA83[18] , \wAMid87[7] , \wRegInA13[11] , 
        \wRegInA30[20] , \wRegInA45[10] , \wRegInB95[27] , \wRegInA66[21] , 
        \wAMid82[29] , \wAIn99[22] , \wRegInA73[15] , \wAMid82[30] , 
        \wRegInA50[24] , \wBMid119[5] , \wRegInB21[3] , \wRegInA25[14] , 
        \wRegInB80[13] , \wRegInA93[0] , \ScanLink179[15] , \ScanLink81[17] , 
        \wAMid29[7] , \wBMid92[1] , \ScanLink94[23] , \wAIn120[8] , 
        \ScanLink119[11] , \wAIn4[20] , \wBMid45[27] , \wAIn69[3] , 
        \wRegInA41[6] , \wBMid88[23] , \ScanLink252[23] , \ScanLink241[9] , 
        \wBMid8[0] , \wBMid30[17] , \wRegInB22[0] , \wRegInA113[28] , 
        \wBMid66[16] , \ScanLink227[13] , \ScanLink182[14] , \wAMid0[17] , 
        \wAIn4[13] , \wBIn9[22] , \wBMid13[26] , \wRegInA113[31] , 
        \ScanLink59[27] , \wAIn17[13] , \wAIn21[16] , \wBMid25[23] , 
        \wBMid50[13] , \wBMid73[22] , \ScanLink204[22] , \wBMid91[2] , 
        \wRegInA42[5] , \ScanLink211[16] , \ScanLink39[23] , \ScanLink247[17] , 
        \ScanLink232[27] , \ScanLink197[20] , \wAIn77[17] , \wRegInB38[27] , 
        \wAIn34[22] , \wAIn54[26] , \wAIn41[12] , \wRegInA90[3] , 
        \wAMid79[31] , \wRegInB58[23] , \wBMid43[4] , \wAIn62[23] , 
        \wBMid107[9] , \wRegInA88[14] , \wAMid79[28] , \wRegInB45[7] , 
        \ScanLink119[22] , \ScanLink94[10] , \wAMid9[7] , \wAIn10[8] , 
        \wBIn68[4] , \wBMid88[10] , \ScanLink78[9] , \wAIn99[11] , 
        \wRegInB5[7] , \wRegInA25[2] , \ScanLink189[2] , \wRegInB58[8] , 
        \wRegInA73[26] , \ScanLink179[26] , \ScanLink81[24] , \wAMid106[19] , 
        \wRegInA25[27] , \wRegInB97[1] , \wRegInA50[17] , \wRegInB80[20] , 
        \ScanLink65[6] , \wAMid125[31] , \wBIn98[30] , \wAMid112[2] , 
        \wRegInA30[13] , \wRegInB95[14] , \wBMid24[3] , \wAMid125[28] , 
        \wRegInA45[23] , \wRegInA13[22] , \wAIn34[11] , \wAIn41[21] , 
        \wBIn98[29] , \wRegInA66[12] , \wRegInA119[1] , \ScanLink66[5] , 
        \wRegInA88[27] , \ScanLink238[2] , \wBIn16[18] , \wAIn17[20] , 
        \wAIn62[10] , \wRegInB58[10] , \wRegInB94[2] , \wBMid27[0] , 
        \wBIn63[28] , \wAIn77[24] , \wBIn100[19] , \wBIn123[31] , 
        \wRegInB38[14] , \wAIn21[25] , \wBIn35[30] , \wBIn40[19] , 
        \wAIn54[15] , \wBIn63[31] , \wBIn123[28] , \ScanLink158[7] , 
        \wBMid25[10] , \wBIn35[29] , \wBMid73[11] , \wAMid111[1] , 
        \ScanLink211[25] , \ScanLink232[14] , \ScanLink39[10] , 
        \ScanLink197[13] , \wBMid30[24] , \wBMid50[20] , \wRegInB46[4] , 
        \ScanLink247[24] , \wBMid45[14] , \ScanLink227[20] , \ScanLink182[27] , 
        \wAMid81[9] , \wRegInB6[4] , \ScanLink252[10] , \wBMid13[15] , 
        \ScanLink59[14] , \wBIn76[8] , \ScanLink204[11] , \ScanLink145[8] , 
        \wBIn12[30] , \wBIn12[29] , \wAIn13[11] , \wAIn30[20] , \wBMid66[25] , 
        \wBIn80[8] , \wRegInA26[1] , \wAIn45[10] , \wAIn66[21] , 
        \wRegInB29[11] , \wAMid77[9] , \wAIn25[14] , \wBIn31[18] , 
        \wBIn44[31] , \wBIn67[19] , \wRegInB49[15] , \wAIn73[15] , 
        \wBIn104[28] , \wRegInA99[22] , \ScanLink42[3] , \wBIn44[28] , 
        \wAIn50[24] , \wBMid77[20] , \wBIn104[31] , \wBIn127[19] , 
        \wBIn117[6] , \ScanLink215[14] , \ScanLink48[11] , \ScanLink243[15] , 
        \wAIn0[22] , \wBMid21[21] , \wBMid54[11] , \ScanLink236[25] , 
        \ScanLink193[22] , \wBMid41[25] , \wAIn0[11] , \wAMid4[26] , 
        \wBMid34[15] , \wRegInB62[2] , \ScanLink256[21] , \wBMid62[14] , 
        \ScanLink223[11] , \ScanLink186[16] , \ScanLink28[15] , \wBMid17[24] , 
        \ScanLink90[5] , \wAIn29[1] , \wAMid69[5] , \wRegInA120[8] , 
        \ScanLink200[20] , \ScanLink168[23] , \ScanLink90[21] , \wBIn114[5] , 
        \wBMid34[26] , \wAIn88[14] , \wBMid99[15] , \ScanLink93[6] , 
        \wAMid102[28] , \wRegInA21[16] , \wRegInA54[26] , \wRegInB61[1] , 
        \ScanLink202[8] , \ScanLink85[15] , \ScanLink108[27] , \wRegInA77[17] , 
        \wRegInA41[12] , \wRegInB84[11] , \ScanLink41[0] , \wRegInA34[22] , 
        \wRegInB91[25] , \wAMid102[31] , \wAMid121[19] , \wRegInA62[23] , 
        \wRegInA17[13] , \wRegInA117[19] , \wBMid41[16] , \ScanLink223[22] , 
        \ScanLink186[25] , \wBIn4[4] , \wAMid4[15] , \wBMid17[17] , 
        \ScanLink256[12] , \ScanLink200[13] , \wBIn7[7] , \wAIn8[9] , 
        \wAIn13[22] , \wBMid21[12] , \wBMid62[27] , \wRegInA66[3] , 
        \ScanLink28[26] , \wBMid77[13] , \ScanLink215[27] , \ScanLink48[22] , 
        \ScanLink236[16] , \ScanLink193[11] , \wAIn25[27] , \wAIn50[17] , 
        \wBMid54[22] , \ScanLink243[26] , \wBMid67[2] , \wAIn73[26] , 
        \wRegInB108[1] , \wRegInB49[26] , \wRegInA99[11] , \ScanLink118[5] , 
        \wAIn30[13] , \wAIn45[23] , \wAIn53[9] , \ScanLink26[7] , \wAIn66[12] , 
        \wRegInB29[22] , \wAMid16[11] , \wBIn19[16] , \wBMid18[7] , 
        \wBIn28[6] , \wAIn31[3] , \wBIn35[9] , \wBMid64[1] , \wAIn119[1] , 
        \wRegInA34[11] , \wRegInB91[16] , \wRegInA41[21] , \wAMid86[18] , 
        \wAIn88[27] , \wRegInA17[20] , \wRegInA62[10] , \wRegInA77[24] , 
        \wBMid99[26] , \wRegInA21[25] , \wRegInA54[15] , \wRegInB84[22] , 
        \ScanLink25[4] , \ScanLink106[9] , \wAMid71[7] , \wRegInA8[30] , 
        \wRegInA8[29] , \wRegInA65[0] , \ScanLink108[14] , \ScanLink85[26] , 
        \ScanLink168[10] , \ScanLink90[12] , \wRegInA9[3] , \wBIn86[6] , 
        \wAMid63[21] , \wAIn110[30] , \wAIn110[29] , \wRegInA19[6] , 
        \wRegInA109[21] , \ScanLink5[1] , \wRegInB79[3] , \wAMid20[14] , 
        \wAMid35[20] , \wAMid40[10] , \wBIn54[0] , \ScanLink167[0] , 
        \wAMid55[24] , \wBIn111[8] , \wRegInA87[30] , \ScanLink59[2] , 
        \wRegInA126[6] , \wBIn57[3] , \wAMid76[15] , \wRegInA87[29] , 
        \wBIn79[12] , \wAMid109[17] , \ScanLink207[5] , \ScanLink164[3] , 
        \wAMid12[11] , \wAMid15[3] , \wAMid16[22] , \wBIn19[25] , 
        \wAMid20[27] , \wBIn30[4] , \wAIn32[0] , \wBIn82[13] , \wBIn97[27] , 
        \wBMid110[26] , \wAMid98[20] , \ScanLink7[21] , \ScanLink204[6] , 
        \wBIn85[5] , \wBMid105[12] , \wBMid126[23] , \wRegInA125[5] , 
        \ScanLink95[8] , \wRegInB127[21] , \wRegInB5[20] , \ScanLink120[29] , 
        \ScanLink176[31] , \wAMid72[4] , \wRegInB104[10] , \ScanLink155[19] , 
        \ScanLink120[30] , \ScanLink103[18] , \wRegInA3[25] , \wRegInB111[24] , 
        \ScanLink219[9] , \ScanLink176[28] , \ScanLink88[7] , \ScanLink6[2] , 
        \wAIn101[3] , \ScanLink103[4] , \wAIn48[8] , \wAMid55[17] , 
        \wAIn87[1] , \wAMid76[26] , \wBIn79[21] , \wAMid35[13] , \wAMid63[12] , 
        \wRegInB42[19] , \wRegInB61[31] , \wAIn78[19] , \wRegInB37[29] , 
        \wAMid40[23] , \wRegInB61[28] , \wAIn55[7] , \wRegInB14[18] , 
        \wRegInB37[30] , \wBMid125[1] , \ScanLink248[19] , \wAMid16[0] , 
        \wBMid69[18] , \wRegInA109[12] , \wRegInB113[0] , \ScanLink75[18] , 
        \ScanLink56[30] , \wBMid126[2] , \ScanLink56[29] , \ScanLink23[19] , 
        \ScanLink20[9] , \wRegInA3[16] , \wRegInB111[17] , \wAMid31[7] , 
        \wBIn33[7] , \wAIn56[4] , \wBIn82[20] , \wBMid92[19] , \wRegInB5[13] , 
        \wRegInB127[12] , \wRegInB104[23] , \wRegInB110[3] , \wBMid105[21] , 
        \ScanLink100[7] , \wAIn83[18] , \wAIn84[2] , \wAIn102[0] , 
        \wBMid126[10] , \wBIn97[14] , \wAMid109[24] , \wBMid110[15] , 
        \wAMid98[13] , \ScanLink7[12] , \wBMid45[8] , \wRegInA118[15] , 
        \ScanLink189[29] , \wAIn71[3] , \wBMid101[5] , \wAIn114[30] , 
        \wAIn114[29] , \wRegInA59[6] , \ScanLink189[30] , \wRegInB39[3] , 
        \wAMid31[20] , \wBMid58[7] , \wAMid67[21] , \wBIn68[26] , 
        \wRegInA44[9] , \ScanLink127[0] , \wBIn14[0] , \wAMid44[10] , 
        \wBIn17[3] , \wAMid24[14] , \wAIn125[7] , \wAMid51[24] , 
        \wRegInA83[30] , \ScanLink19[2] , \wAMid72[15] , \wRegInA83[29] , 
        \ScanLink247[5] , \wRegInA88[3] , \wAIn126[4] , \ScanLink124[3] , 
        \wAMid12[22] , \wAMid24[27] , \wAMid32[4] , \wAIn72[0] , \wBIn86[13] , 
        \wBIn93[27] , \wBMid114[26] , \wRegInA78[28] , \ScanLink3[21] , 
        \wAMid89[14] , \wBMid101[12] , \wAMid118[23] , \wBMid122[23] , 
        \wRegInA78[31] , \ScanLink244[6] , \wRegInB1[20] , \ScanLink172[31] , 
        \ScanLink151[19] , \wRegInB123[21] , \ScanLink124[29] , \wAMid51[17] , 
        \wBMid89[2] , \wBMid102[6] , \ScanLink172[28] , \ScanLink107[18] , 
        \wRegInA7[25] , \wRegInB100[10] , \wRegInB115[24] , \ScanLink124[30] , 
        \wBIn70[4] , \wAMid67[12] , \wAMid72[26] , \wAMid87[5] , 
        \ScanLink143[4] , \wRegInB0[8] , \wBIn68[15] , \wRegInB33[29] , 
        \wRegInB40[8] , \wAIn15[7] , \wAMid31[13] , \wAMid44[23] , 
        \wRegInB46[19] , \ScanLink223[1] , \wRegInB65[31] , \wRegInB10[18] , 
        \wRegInB33[30] , \wRegInA102[2] , \wRegInB65[28] , \ScanLink239[30] , 
        \wBMid18[31] , \wAMid55[3] , \ScanLink191[2] , \ScanLink239[29] , 
        \ScanLink52[30] , \wBMid18[28] , \wRegInA118[26] , \ScanLink71[18] , 
        \ScanLink52[29] , \wAMid56[0] , \wAMid99[9] , \wRegInB115[17] , 
        \ScanLink60[9] , \ScanLink27[19] , \wRegInA7[16] , \wAIn0[20] , 
        \wAMid0[26] , \wBIn1[9] , \wAIn16[4] , \wBIn16[30] , \wBIn16[29] , 
        \wAIn17[11] , \wAIn34[20] , \wAIn41[10] , \wBIn73[7] , \wAMid84[6] , 
        \wBMid96[19] , \wRegInB1[13] , \ScanLink192[1] , \wRegInB100[23] , 
        \wRegInB123[12] , \wBIn86[20] , \wAMid89[27] , \wBMid101[21] , 
        \wAMid109[1] , \wAMid118[10] , \ScanLink140[7] , \wAIn87[18] , 
        \wBMid122[10] , \wRegInA101[1] , \wBIn93[14] , \wBMid114[15] , 
        \wRegInA90[1] , \ScanLink220[2] , \ScanLink3[12] , \wAMid37[9] , 
        \wRegInA88[16] , \wBMid43[6] , \wAIn62[21] , \wRegInB58[21] , 
        \wBIn40[31] , \wAIn77[15] , \wBIn63[19] , \wBIn100[28] , 
        \wRegInB38[25] , \wAIn21[14] , \wBIn40[28] , \wAIn54[24] , 
        \wBIn100[31] , \wBIn123[19] , \wBIn35[18] , \wRegInA42[7] , 
        \ScanLink211[14] , \wAIn4[22] , \wBMid8[2] , \wBMid25[21] , 
        \wBMid73[20] , \wAIn123[9] , \ScanLink39[21] , \ScanLink232[25] , 
        \ScanLink197[22] , \wBMid30[15] , \wBMid50[11] , \wBMid91[0] , 
        \ScanLink247[15] , \wRegInB22[2] , \ScanLink227[11] , 
        \ScanLink182[16] , \wBMid45[25] , \wBMid13[24] , \ScanLink252[21] , 
        \ScanLink204[20] , \ScanLink59[25] , \wAMid0[15] , \wAIn4[11] , 
        \wBIn9[13] , \wAMid29[5] , \wBMid66[14] , \ScanLink119[13] , 
        \wBMid92[3] , \wBMid119[7] , \ScanLink94[21] , \wBMid40[5] , 
        \wAIn69[1] , \wBMid88[21] , \wRegInA41[4] , \wBMid104[8] , 
        \wRegInB21[1] , \wRegInA73[17] , \ScanLink242[8] , \ScanLink179[17] , 
        \ScanLink81[15] , \wBMid45[16] , \wBIn98[18] , \wAIn99[20] , 
        \wAMid106[31] , \wAMid106[28] , \wRegInA25[16] , \wRegInB80[11] , 
        \wRegInA50[26] , \wRegInA93[2] , \wRegInA30[22] , \wRegInA45[12] , 
        \wRegInB95[25] , \wAMid125[19] , \wRegInA13[13] , \wRegInA66[23] , 
        \wBMid30[26] , \wRegInB6[6] , \ScanLink252[12] , \wBMid66[27] , 
        \wRegInA26[3] , \wRegInA113[19] , \ScanLink227[22] , \ScanLink182[25] , 
        \wBIn9[20] , \wAMid9[5] , \wAIn13[9] , \wBMid13[17] , \wAIn21[27] , 
        \wBMid25[12] , \wBMid50[22] , \wBMid73[13] , \ScanLink204[13] , 
        \ScanLink59[16] , \ScanLink39[12] , \ScanLink247[26] , 
        \ScanLink211[27] , \wRegInB46[6] , \ScanLink232[16] , 
        \ScanLink197[11] , \wBMid27[2] , \wAIn77[26] , \wRegInB38[16] , 
        \wAIn17[22] , \wAIn34[13] , \wAIn54[17] , \wAMid111[3] , 
        \ScanLink158[5] , \wAIn41[23] , \wRegInA119[3] , \ScanLink66[7] , 
        \wRegInB58[12] , \wRegInB94[0] , \wAIn62[12] , \wRegInA88[25] , 
        \ScanLink238[0] , \wBMid24[1] , \wBIn68[6] , \wAMid79[19] , 
        \wAMid112[0] , \wRegInA30[11] , \wRegInA45[21] , \wRegInB95[16] , 
        \wRegInA66[10] , \wBIn75[9] , \wAMid82[18] , \wAIn99[13] , 
        \wRegInA13[20] , \wRegInA73[24] , \wRegInB97[3] , \wRegInA25[25] , 
        \wRegInA50[15] , \wRegInB80[22] , \ScanLink65[4] , \wRegInA25[0] , 
        \ScanLink146[9] , \wAMid82[8] , \ScanLink189[0] , \ScanLink81[26] , 
        \wRegInB5[5] , \wRegInB45[5] , \ScanLink179[24] , \wAIn29[3] , 
        \wAMid69[7] , \wAMid74[8] , \wAIn88[16] , \wBMid88[12] , 
        \ScanLink119[20] , \ScanLink94[12] , \wRegInA17[11] , \wRegInA34[20] , 
        \wRegInA41[10] , \wRegInB91[27] , \ScanLink41[2] , \wRegInA62[21] , 
        \wBIn83[9] , \wAMid86[30] , \wAMid86[29] , \wRegInA77[15] , 
        \wBIn109[8] , \wRegInA21[14] , \wRegInB84[13] , \wRegInA54[24] , 
        \wBMid99[17] , \wRegInB61[3] , \wRegInA123[9] , \ScanLink93[4] , 
        \ScanLink108[25] , \ScanLink85[17] , \wBIn114[7] , \wRegInA8[18] , 
        \ScanLink168[21] , \ScanLink90[23] , \wBMid34[17] , \wRegInA117[28] , 
        \wBMid41[27] , \wRegInB62[0] , \ScanLink223[13] , \ScanLink186[14] , 
        \ScanLink256[23] , \wAIn0[13] , \wAMid4[24] , \wBMid17[26] , 
        \wRegInA117[31] , \ScanLink201[9] , \ScanLink200[22] , \wBIn12[18] , 
        \wAIn13[20] , \wAIn13[13] , \wBMid21[23] , \wBMid62[16] , 
        \wBMid77[22] , \wBIn117[4] , \ScanLink215[16] , \ScanLink90[7] , 
        \ScanLink28[17] , \ScanLink48[13] , \ScanLink236[27] , 
        \ScanLink193[20] , \wAIn25[16] , \wAIn50[26] , \wBMid54[13] , 
        \ScanLink243[17] , \wAIn73[17] , \wRegInB49[17] , \wRegInA99[20] , 
        \wAIn30[22] , \wAIn45[12] , \ScanLink42[1] , \wAIn66[23] , 
        \wRegInB29[13] , \wBIn28[4] , \wAIn50[8] , \wBMid99[24] , 
        \wRegInA65[2] , \ScanLink168[12] , \ScanLink90[10] , \ScanLink38[9] , 
        \wRegInB18[8] , \wRegInA77[26] , \ScanLink108[16] , \ScanLink85[24] , 
        \wRegInA21[27] , \wRegInA54[17] , \wRegInB84[20] , \ScanLink25[6] , 
        \wAMid102[19] , \wAMid121[31] , \wRegInA41[23] , \wAIn119[3] , 
        \wRegInA34[13] , \wRegInB91[14] , \wAIn30[11] , \wBMid64[3] , 
        \wAIn88[25] , \wAMid121[28] , \wRegInA62[12] , \wRegInA17[22] , 
        \wAIn45[21] , \ScanLink26[5] , \wBIn31[30] , \wAIn66[10] , 
        \wRegInB29[20] , \wBMid21[10] , \wAIn25[25] , \wBIn31[29] , 
        \wBIn67[28] , \wRegInB49[24] , \wBMid67[0] , \wAIn73[24] , 
        \wBIn104[19] , \wBIn127[31] , \wRegInA99[13] , \wBIn44[19] , 
        \wAIn50[15] , \wBIn67[31] , \wBMid54[20] , \wBMid77[11] , 
        \wBIn127[28] , \ScanLink118[7] , \wRegInB108[3] , \ScanLink243[24] , 
        \ScanLink215[25] , \ScanLink48[20] , \ScanLink236[14] , 
        \ScanLink193[13] , \wBMid41[14] , \ScanLink256[10] , \wAIn0[3] , 
        \wAIn1[19] , \wAMid4[17] , \wBMid34[24] , \wBMid62[25] , 
        \ScanLink223[20] , \ScanLink186[27] , \wRegInA66[1] , \ScanLink28[24] , 
        \wBMid4[25] , \wAMid15[1] , \wAMid16[13] , \wBMid17[15] , \wBIn36[8] , 
        \wAMid20[16] , \wAIn32[2] , \wRegInA3[27] , \wRegInB111[26] , 
        \ScanLink200[11] , \ScanLink105[8] , \ScanLink6[0] , \ScanLink88[5] , 
        \wBIn57[1] , \wAMid72[6] , \wBIn85[7] , \wBMid92[28] , \wRegInB5[22] , 
        \wRegInB127[23] , \wBIn82[11] , \wBMid92[31] , \wBMid105[10] , 
        \wRegInB104[12] , \wAIn83[30] , \wBIn112[9] , \wBMid126[21] , 
        \ScanLink204[4] , \wRegInA125[7] , \wAIn83[29] , \wBIn97[25] , 
        \wBIn98[8] , \wAMid109[15] , \ScanLink164[1] , \wAMid98[22] , 
        \ScanLink7[23] , \wBMid110[24] , \wRegInA126[4] , \wAMid55[26] , 
        \ScanLink59[0] , \wAMid76[17] , \wBIn79[10] , \ScanLink207[7] , 
        \ScanLink96[9] , \wAMid16[2] , \wBIn19[14] , \wBMid18[5] , 
        \wAMid63[23] , \wRegInB42[28] , \wAIn78[28] , \wAIn31[1] , 
        \wAMid35[22] , \wRegInB14[30] , \wRegInB37[18] , \wAMid40[12] , 
        \wRegInB42[31] , \wRegInB61[19] , \ScanLink167[2] , \wBIn54[2] , 
        \wAIn78[31] , \wBMid69[30] , \wRegInB14[29] , \wRegInB79[1] , 
        \ScanLink248[31] , \wRegInA109[23] , \ScanLink248[28] , \ScanLink5[3] , 
        \ScanLink23[31] , \wAMid71[5] , \wRegInA9[1] , \ScanLink75[29] , 
        \wBIn33[5] , \wBMid69[29] , \ScanLink23[28] , \wBIn82[22] , 
        \wBIn86[4] , \wRegInA19[4] , \ScanLink75[30] , \wBIn97[16] , 
        \wAMid98[11] , \wAMid109[26] , \ScanLink56[18] , \ScanLink7[10] , 
        \wBMid105[23] , \wBMid110[17] , \wAIn84[0] , \wAIn102[2] , 
        \ScanLink100[5] , \wBMid126[12] , \wRegInB127[10] , \wRegInB5[11] , 
        \ScanLink120[18] , \wRegInB104[21] , \wRegInB110[1] , 
        \ScanLink155[28] , \ScanLink103[30] , \ScanLink23[8] , 
        \wRegInB111[15] , \ScanLink176[19] , \ScanLink103[29] , 
        \ScanLink155[31] , \wAIn55[5] , \wAIn56[6] , \wBMid126[0] , 
        \wRegInA3[14] , \wRegInB113[2] , \wAIn110[18] , \wAMid16[20] , 
        \wAMid63[10] , \wBMid125[3] , \wRegInA109[10] , \wBIn19[27] , 
        \wAMid20[25] , \wBIn30[6] , \wAMid35[11] , \wAMid40[21] , 
        \wAMid55[15] , \wAIn87[3] , \wAIn101[1] , \wAMid76[24] , \wBIn79[23] , 
        \wRegInA87[18] , \ScanLink103[6] , \wRegInA103[25] , \wRegInB118[9] , 
        \ScanLink192[19] , \wBIn26[2] , \wAIn91[7] , \wRegInA120[14] , 
        \wAIn117[5] , \ScanLink115[2] , \wBIn13[21] , \wBIn13[12] , 
        \wBIn25[17] , \wBIn73[16] , \wBIn110[27] , \wRegInB105[6] , 
        \wRegInA116[11] , \wBIn30[23] , \wBIn50[27] , \wAIn43[1] , 
        \wBIn45[13] , \wBIn126[22] , \wBIn25[1] , \wAIn40[2] , \wBIn66[22] , 
        \wAMid69[25] , \wBMid74[9] , \wAMid87[10] , \wBIn105[13] , 
        \wAMid116[27] , \wRegInA98[19] , \wRegInB106[5] , \wBIn88[17] , 
        \wAMid92[24] , \wAMid120[22] , \wRegInA40[30] , \wRegInA63[18] , 
        \wRegInA16[28] , \wBMid69[6] , \wAMid103[13] , \wRegInA40[29] , 
        \wRegInA68[7] , \wAIn109[9] , \wRegInA16[31] , \wRegInA9[21] , 
        \wRegInA35[19] , \ScanLink169[18] , \ScanLink28[3] , \wAIn92[4] , 
        \wAIn114[6] , \wRegInA75[8] , \ScanLink116[1] , \wBIn30[10] , 
        \wBIn45[20] , \wBIn126[11] , \wBIn66[11] , \wAMid69[16] , 
        \wBIn105[20] , \wAIn67[29] , \wBIn110[14] , \wRegInB28[19] , 
        \wAMid67[1] , \wBIn73[25] , \wAIn3[0] , \wBMid4[16] , \wAIn12[19] , 
        \wAIn31[31] , \wBMid20[30] , \wBMid20[29] , \wBIn25[24] , \wAIn27[5] , 
        \wAIn31[28] , \wAIn44[18] , \wBIn50[14] , \wAIn67[30] , \wBIn90[0] , 
        \wRegInA103[16] , \wRegInA116[22] , \ScanLink201[28] , 
        \ScanLink222[19] , \ScanLink201[31] , \ScanLink211[3] , \wBMid55[19] , 
        \wBMid76[31] , \ScanLink49[19] , \wBIn42[6] , \wRegInA120[27] , 
        \ScanLink171[6] , \wAIn24[6] , \wAIn39[9] , \wBMid76[28] , 
        \wRegInB71[9] , \ScanLink212[0] , \wBIn41[5] , \wAMid92[17] , 
        \wAMid120[11] , \wRegInA1[9] , \wRegInA9[12] , \ScanLink172[5] , 
        \ScanLink91[30] , \ScanLink91[29] , \wAMid103[20] , \wAMid116[14] , 
        \wBIn119[2] , \ScanLink51[8] , \wRegInB85[19] , \wAMid64[2] , 
        \wBIn93[3] , \wAMid87[23] , \wAMid18[4] , \wAIn79[11] , \wBIn88[24] , 
        \wRegInB15[10] , \wRegInB60[20] , \wRegInB10[0] , \wRegInB36[21] , 
        \wRegInB43[11] , \wRegInA93[26] , \wAIn19[15] , \wBIn78[29] , 
        \wRegInB23[15] , \wRegInA86[12] , \wRegInB56[25] , \wAIn58[0] , 
        \wAIn97[9] , \wRegInA70[5] , \wBIn78[30] , \wRegInB75[14] , 
        \wBMid0[27] , \wBIn3[26] , \wBIn3[15] , \wBIn7[24] , \wBIn7[17] , 
        \wBMid68[10] , \ScanLink57[21] , \wBMid71[4] , \wAIn104[26] , 
        \ScanLink22[11] , \wAIn127[17] , \wRegInB103[8] , \ScanLink74[10] , 
        \ScanLink30[1] , \ScanLink229[15] , \ScanLink249[11] , 
        \ScanLink199[26] , \ScanLink61[24] , \wBMid86[25] , \wAIn89[5] , 
        \wBMid93[11] , \wAIn111[12] , \ScanLink42[15] , \ScanLink14[14] , 
        \ScanLink177[13] , \ScanLink102[23] , \ScanLink37[25] , 
        \ScanLink154[22] , \ScanLink121[12] , \ScanLink33[2] , 
        \ScanLink134[26] , \ScanLink162[27] , \ScanLink141[16] , 
        \ScanLink117[17] , \wBMid15[0] , \wBIn59[7] , \wBMid68[23] , 
        \wBMid72[7] , \wAIn82[10] , \wRegInB13[3] , \wBIn83[31] , 
        \wRegInA68[27] , \wRegInA73[6] , \wBIn83[28] , \wAIn97[24] , 
        \wBMid104[30] , \wAIn112[8] , \wBMid104[29] , \wAIn111[21] , 
        \wRegInA108[29] , \ScanLink249[22] , \ScanLink199[15] , 
        \ScanLink14[27] , \ScanLink61[17] , \wAMid123[1] , \wRegInA108[30] , 
        \ScanLink54[5] , \ScanLink37[16] , \ScanLink42[26] , \wAIn104[15] , 
        \ScanLink22[22] , \ScanLink57[12] , \wAIn127[24] , \ScanLink74[23] , 
        \wAMid17[19] , \wAIn19[26] , \wRegInB56[16] , \wRegInB74[4] , 
        \ScanLink229[26] , \ScanLink8[6] , \wAMid34[28] , \wRegInB23[26] , 
        \wRegInA86[21] , \wRegInB75[27] , \ScanLink86[3] , \wAMid41[18] , 
        \wBIn101[0] , \wRegInA14[1] , \wRegInB60[13] , \wBIn44[8] , 
        \wAMid62[30] , \wRegInB15[23] , \ScanLink177[8] , \wRegInA4[4] , 
        \wAMid34[31] , \wAMid62[29] , \wAIn79[22] , \wRegInB43[22] , 
        \wAIn82[23] , \wAIn97[17] , \wRegInB36[12] , \wRegInB77[7] , 
        \wRegInA93[15] , \ScanLink85[0] , \wBMid86[16] , \wBIn88[2] , 
        \wAMid99[31] , \wAMid99[28] , \ScanLink6[29] , \wBIn102[3] , 
        \wRegInA7[7] , \wRegInA68[14] , \wRegInA17[2] , \ScanLink6[30] , 
        \ScanLink141[25] , \ScanLink134[15] , \ScanLink162[14] , 
        \ScanLink57[6] , \wBMid16[3] , \ScanLink209[1] , \ScanLink177[20] , 
        \ScanLink117[24] , \wAIn22[8] , \wAMid120[2] , \wRegInB4[31] , 
        \wRegInB105[18] , \wRegInB126[30] , \ScanLink102[10] , \wBMid82[27] , 
        \wAIn86[12] , \wAIn93[26] , \wBMid93[22] , \wRegInB4[28] , 
        \ScanLink154[11] , \wBIn126[5] , \wRegInA33[4] , \wRegInB126[29] , 
        \ScanLink169[4] , \ScanLink121[21] , \wRegInA79[11] , \wRegInA19[15] , 
        \wRegInB53[1] , \ScanLink2[18] , \wAMid104[4] , \ScanLink230[8] , 
        \ScanLink130[24] , \wAMid89[3] , \ScanLink145[14] , \ScanLink166[25] , 
        \ScanLink113[15] , \wBIn9[1] , \wAMid13[31] , \wAIn18[2] , 
        \wBMid19[22] , \wBMid31[6] , \wBMid32[5] , \wAMid45[9] , \wBMid97[13] , 
        \wRegInB81[7] , \wRegInB101[29] , \ScanLink106[21] , \ScanLink173[11] , 
        \wRegInB0[19] , \wRegInB101[30] , \wRegInB122[18] , \ScanLink125[10] , 
        \ScanLink238[23] , \ScanLink150[20] , \ScanLink73[0] , 
        \ScanLink65[26] , \wBMid79[26] , \wAMid107[7] , \ScanLink46[17] , 
        \ScanLink10[16] , \wAIn115[10] , \ScanLink181[8] , \ScanLink33[27] , 
        \wAMid58[6] , \wAIn100[24] , \ScanLink70[3] , \ScanLink53[23] , 
        \ScanLink26[13] , \wAIn123[15] , \wRegInB82[4] , \ScanLink188[10] , 
        \ScanLink70[12] , \wAIn68[27] , \wRegInB27[17] , \wRegInA82[10] , 
        \wBIn125[6] , \wRegInA30[7] , \wRegInB52[27] , \wAMid30[19] , 
        \wAMid45[29] , \wRegInB71[16] , \wRegInB11[12] , \wRegInA112[8] , 
        \wAMid13[28] , \wAMid45[30] , \wAMid66[18] , \wRegInB64[22] , 
        \wRegInB32[23] , \wRegInB50[2] , \wRegInA97[24] , \wBMid56[1] , 
        \wRegInB47[13] , \ScanLink173[22] , \wBMid97[20] , \wBMid99[8] , 
        \wRegInA85[6] , \ScanLink150[13] , \ScanLink106[12] , \ScanLink129[6] , 
        \ScanLink125[23] , \wBMid82[14] , \ScanLink145[27] , \ScanLink130[17] , 
        \ScanLink166[16] , \ScanLink17[4] , \wBMid3[9] , \wBIn19[5] , 
        \wBMid19[11] , \wAIn61[9] , \wAIn68[14] , \wBMid84[7] , \wAIn86[21] , 
        \ScanLink249[3] , \ScanLink113[26] , \wBIn87[19] , \wBMid100[18] , 
        \wAMid119[29] , \wBMid123[29] , \wRegInA19[26] , \wRegInA57[0] , 
        \wRegInA98[9] , \ScanLink134[9] , \wRegInA79[22] , \wBMid87[4] , 
        \wAIn93[15] , \wBMid123[30] , \wAMid119[30] , \wRegInB37[5] , 
        \wRegInB11[21] , \wRegInA54[3] , \wRegInB64[11] , \wRegInB47[20] , 
        \wRegInB27[24] , \wRegInB32[10] , \wRegInB34[6] , \wRegInB52[14] , 
        \wRegInA97[17] , \wRegInA82[23] , \wRegInB71[25] , \wAIn100[17] , 
        \wRegInA86[5] , \ScanLink26[20] , \ScanLink53[10] , \wBMid55[2] , 
        \wAIn123[26] , \ScanLink70[21] , \wRegInB29[9] , \ScanLink188[23] , 
        \wAMid4[0] , \wAMid7[3] , \wBMid29[4] , \wBMid79[15] , \wAIn115[23] , 
        \ScanLink238[10] , \ScanLink10[25] , \ScanLink65[15] , 
        \ScanLink33[14] , \wAMid92[2] , \ScanLink46[24] , \ScanLink14[7] , 
        \wBIn65[3] , \ScanLink156[3] , \wBMid89[18] , \wRegInA117[5] , 
        \ScanLink68[1] , \ScanLink95[18] , \wAIn16[31] , \wAIn16[28] , 
        \wBIn17[10] , \wBIn34[21] , \wAMid40[4] , \wAMid96[26] , \wBIn99[21] , 
        \ScanLink236[6] , \wRegInB8[0] , \ScanLink9[27] , \wAMid83[12] , 
        \wAMid107[11] , \wAMid124[20] , \wRegInA28[5] , \wAMid112[25] , 
        \wRegInB81[28] , \ScanLink184[5] , \wRegInB48[0] , \wAIn98[19] , 
        \wRegInB81[31] , \wRegInB87[9] , \wBIn41[11] , \wAMid101[9] , 
        \wBIn122[20] , \ScanLink187[6] , \wAMid18[17] , \wBMid37[8] , 
        \wAMid43[7] , \wBIn62[20] , \wBIn101[11] , \wRegInB59[18] , 
        \wAIn40[30] , \wAMid78[13] , \wBIn114[25] , \wAIn63[18] , \wBIn77[14] , 
        \wBIn21[15] , \wBMid24[18] , \wAIn35[19] , \wRegInA109[9] , 
        \wAIn40[29] , \wBMid51[28] , \wBIn54[25] , \wBIn66[0] , \wBIn123[8] , 
        \wRegInA36[9] , \wAMid91[1] , \ScanLink226[31] , \ScanLink205[19] , 
        \ScanLink155[0] , \wRegInB99[5] , \wRegInA112[13] , \ScanLink253[18] , 
        \ScanLink226[28] , \ScanLink235[5] , \wBMid72[19] , \wRegInA107[27] , 
        \wBMid0[14] , \wBMid6[4] , \wAMid24[0] , \wBMid51[31] , 
        \wRegInA114[6] , \ScanLink38[18] , \wAIn64[4] , \wAMid112[16] , 
        \wRegInA124[16] , \wRegInA83[8] , \wAMid83[21] , \wBMid114[2] , 
        \wAMid124[13] , \wBIn8[19] , \wAMid96[15] , \wBIn99[12] , 
        \wRegInA12[19] , \wRegInA31[31] , \wRegInB122[3] , \wAMid107[22] , 
        \wRegInA67[29] , \ScanLink9[14] , \wRegInA31[28] , \wRegInA44[18] , 
        \wRegInA67[30] , \ScanLink132[7] , \ScanLink118[19] , \wBMid82[9] , 
        \wRegInA107[14] , \ScanLink252[2] , \ScanLink196[28] , 
        \wRegInA124[25] , \ScanLink196[31] , \ScanLink131[4] , \wAIn5[31] , 
        \wAIn5[28] , \wRegInB32[8] , \wRegInA112[20] , \wAIn5[7] , \wAIn6[4] , 
        \wBMid5[7] , \wBIn21[26] , \wAMid27[3] , \wAMid78[20] , \wBIn114[16] , 
        \ScanLink251[1] , \wBIn54[16] , \wAIn67[7] , \wBIn77[27] , 
        \wBMid117[1] , \wBIn34[12] , \wBIn41[22] , \wBIn122[13] , 
        \ScanLink12[9] , \wBIn62[13] , \wBIn101[22] , \wRegInB121[0] , 
        \wBIn17[23] , \wAMid18[24] , \wAIn21[2] , \wAMid61[6] , \wBIn96[7] , 
        \wAMid123[8] , \wBMid15[9] , \wAMid17[10] , \wAMid34[21] , 
        \wAIn111[31] , \wRegInB69[2] , \wAIn111[28] , \wRegInA108[20] , 
        \wAMid41[11] , \wBIn101[9] , \wRegInA14[8] , \ScanLink177[1] , 
        \wBIn44[1] , \wBIn18[17] , \wAMid21[15] , \wAMid62[20] , \wAMid77[14] , 
        \wBIn78[13] , \wRegInA86[28] , \ScanLink217[4] , \wBIn47[2] , 
        \wAMid54[25] , \wRegInA86[31] , \ScanLink49[3] , \wBIn96[26] , 
        \wAMid99[21] , \ScanLink6[20] , \wBMid111[27] , \wAMid62[5] , 
        \wBIn83[12] , \wBMid104[13] , \wAMid108[16] , \ScanLink174[2] , 
        \ScanLink85[9] , \ScanLink214[7] , \wRegInB105[11] , \ScanLink177[29] , 
        \ScanLink102[19] , \wAMid17[23] , \wBIn20[5] , \wAIn22[1] , 
        \ScanLink154[18] , \ScanLink121[31] , \wAMid54[16] , \wAIn58[9] , 
        \wAMid77[27] , \wBIn78[20] , \wBIn95[4] , \wRegInB4[21] , 
        \ScanLink177[30] , \wRegInA2[24] , \wRegInB110[25] , \wRegInB126[20] , 
        \ScanLink121[28] , \ScanLink98[6] , \ScanLink209[8] , \wAIn97[0] , 
        \wAIn111[2] , \wAMid21[26] , \wAMid34[12] , \wAMid41[22] , 
        \ScanLink113[5] , \wRegInB15[19] , \wRegInB36[31] , \wAMid62[13] , 
        \wAIn79[18] , \wRegInB60[29] , \wRegInB10[9] , \wRegInB36[28] , 
        \wBIn18[24] , \wAIn45[6] , \wRegInB43[18] , \wRegInB60[30] , 
        \wRegInA108[13] , \ScanLink249[18] , \ScanLink57[28] , \wAIn1[23] , 
        \wAMid5[27] , \wAIn12[10] , \wBIn23[6] , \wAIn46[5] , \wBMid68[19] , 
        \ScanLink22[18] , \wRegInB103[1] , \ScanLink74[19] , \ScanLink57[31] , 
        \ScanLink30[8] , \wAIn94[3] , \wBMid93[18] , \wRegInA2[17] , 
        \wRegInB110[16] , \wRegInB100[2] , \wRegInB105[22] , \wRegInB4[12] , 
        \wRegInB126[13] , \wAIn112[1] , \ScanLink110[6] , \wAIn67[20] , 
        \wAMid67[8] , \wAIn82[19] , \wBIn83[21] , \wBMid104[20] , \wBIn96[15] , 
        \wAMid99[12] , \ScanLink6[13] , \wAMid108[25] , \wBMid111[14] , 
        \wRegInB28[10] , \wBIn13[31] , \wBMid13[7] , \wAIn31[21] , 
        \wAIn44[11] , \wAMid125[6] , \wBIn90[9] , \wBIn45[29] , \wAIn51[25] , 
        \wBIn105[30] , \wBIn126[18] , \wBIn13[28] , \wAIn24[15] , \wBIn30[19] , 
        \ScanLink52[2] , \wBIn45[30] , \wBIn66[18] , \wAIn72[14] , 
        \wBIn105[29] , \wRegInA98[23] , \wBMid16[25] , \wBMid20[20] , 
        \wRegInA2[3] , \wRegInB48[14] , \ScanLink237[24] , \ScanLink192[23] , 
        \wBMid55[10] , \ScanLink242[14] , \wBMid76[21] , \wBIn107[7] , 
        \ScanLink214[15] , \wRegInA12[6] , \ScanLink49[10] , \ScanLink201[21] , 
        \wBMid35[14] , \wBMid63[15] , \ScanLink80[4] , \ScanLink29[14] , 
        \wBMid40[24] , \wRegInB72[3] , \ScanLink222[10] , \ScanLink187[17] , 
        \wAIn1[10] , \wAIn3[9] , \wBMid10[4] , \wAIn39[0] , \wBIn104[4] , 
        \wRegInA11[5] , \wAMid79[4] , \wBMid98[14] , \wRegInA1[0] , 
        \wRegInB71[0] , \ScanLink169[22] , \ScanLink91[20] , \ScanLink212[9] , 
        \ScanLink109[26] , \ScanLink84[14] , \wAMid126[5] , \wRegInA20[17] , 
        \ScanLink83[7] , \wRegInB85[10] , \wRegInA55[27] , \wRegInA76[16] , 
        \wAMid5[14] , \wBMid63[26] , \wAIn89[15] , \wAMid103[30] , 
        \wAMid120[18] , \wRegInA16[12] , \wAMid103[29] , \wRegInA63[22] , 
        \wRegInA35[23] , \wRegInB90[24] , \wRegInA40[13] , \ScanLink51[1] , 
        \wRegInA76[2] , \ScanLink29[27] , \wBMid16[16] , \wBMid40[17] , 
        \ScanLink201[12] , \wBMid35[27] , \wRegInA116[18] , \ScanLink242[27] , 
        \ScanLink222[23] , \ScanLink187[24] , \wBIn1[0] , \wBMid0[3] , 
        \wAMid1[25] , \wBIn8[10] , \wAIn12[23] , \wBMid20[13] , \wBMid55[23] , 
        \wRegInB16[7] , \wRegInB118[0] , \ScanLink237[17] , \ScanLink192[10] , 
        \wAIn24[26] , \wBMid76[12] , \ScanLink214[26] , \ScanLink49[23] , 
        \wAIn43[8] , \wAIn51[16] , \wAIn72[27] , \wBMid77[3] , \wRegInB48[27] , 
        \ScanLink108[4] , \wRegInA98[10] , \wAMid24[9] , \wBIn25[8] , 
        \wAIn31[12] , \wAIn67[13] , \wRegInB28[23] , \wBIn38[7] , \wAIn44[22] , 
        \ScanLink36[6] , \wBMid74[0] , \wAIn89[26] , \wRegInA16[21] , 
        \wRegInA63[11] , \wAIn109[0] , \wRegInA40[20] , \wRegInA35[10] , 
        \wRegInB90[17] , \wAMid87[19] , \wRegInA20[24] , \wRegInA55[14] , 
        \ScanLink35[5] , \wRegInA76[25] , \wRegInB85[23] , \wBMid98[27] , 
        \wRegInA75[1] , \ScanLink109[15] , \ScanLink84[27] , \ScanLink116[8] , 
        \wAMid83[31] , \wRegInA9[31] , \wRegInA9[28] , \wRegInB15[4] , 
        \ScanLink169[11] , \ScanLink91[13] , \wRegInA12[10] , \wRegInA24[15] , 
        \wRegInA31[21] , \wRegInA67[20] , \wRegInB94[26] , \wRegInA44[11] , 
        \ScanLink11[3] , \wRegInA51[25] , \wRegInB81[12] , \wRegInA83[1] , 
        \wAMid39[6] , \wBMid50[6] , \wRegInA72[14] , \wAIn79[2] , 
        \wAMid83[28] , \wBMid89[22] , \wAIn98[23] , \wRegInB31[2] , 
        \wRegInA51[7] , \ScanLink178[14] , \ScanLink80[16] , \ScanLink118[10] , 
        \wBMid82[0] , \wBMid109[4] , \ScanLink95[22] , \wBMid12[27] , 
        \wRegInA112[30] , \ScanLink205[23] , \ScanLink58[26] , \wAMid1[16] , 
        \wAMid4[9] , \wAIn5[21] , \wBMid31[16] , \wBMid67[17] , \wRegInB32[1] , 
        \wRegInA112[29] , \wBMid44[26] , \ScanLink226[12] , \ScanLink183[15] , 
        \ScanLink251[8] , \wBIn8[23] , \wAIn16[12] , \wAIn20[17] , 
        \wBMid24[22] , \ScanLink253[22] , \ScanLink233[26] , \ScanLink196[21] , 
        \wBMid51[12] , \wBMid81[3] , \ScanLink246[16] , \wAIn55[27] , 
        \wBMid72[23] , \wRegInA52[4] , \ScanLink210[17] , \ScanLink38[22] , 
        \wBMid53[5] , \wAIn63[22] , \wAIn76[16] , \wRegInB121[9] , 
        \ScanLink12[0] , \wAMid78[29] , \wRegInB39[26] , \wRegInA89[15] , 
        \wBMid117[8] , \wRegInB59[22] , \wAIn35[23] , \wAIn40[13] , 
        \wRegInA80[2] , \wAMid78[30] , \wBMid89[11] , \ScanLink68[8] , 
        \wRegInB55[6] , \wAIn16[21] , \wBMid34[2] , \wAIn98[10] , \wBIn120[2] , 
        \wRegInA35[3] , \ScanLink178[27] , \ScanLink118[23] , \ScanLink95[11] , 
        \ScanLink80[25] , \wRegInA24[26] , \wRegInA51[16] , \ScanLink199[3] , 
        \ScanLink75[7] , \wRegInB48[9] , \wRegInB81[21] , \wRegInA72[27] , 
        \wRegInB87[0] , \wBIn99[28] , \wRegInB8[9] , \wAMid124[29] , 
        \wRegInA67[13] , \wBIn78[5] , \wBIn99[31] , \wRegInA12[23] , 
        \wAMid102[3] , \wAMid107[18] , \wAMid124[30] , \wRegInA44[22] , 
        \wRegInA31[12] , \wRegInB94[15] , \wRegInB59[11] , \wRegInB84[3] , 
        \wBIn17[19] , \wAIn20[24] , \wBIn34[28] , \wAIn35[10] , \wAIn63[11] , 
        \wRegInA89[26] , \ScanLink228[3] , \wRegInA109[0] , \wAIn40[20] , 
        \ScanLink76[4] , \wBIn34[31] , \wBIn41[18] , \wAIn55[14] , 
        \wBIn62[30] , \wAMid101[0] , \wBIn122[29] , \ScanLink148[6] , 
        \wBMid37[1] , \wBIn62[29] , \wAIn76[25] , \wBMid51[21] , \wBIn101[18] , 
        \wRegInB39[15] , \wBIn122[30] , \ScanLink246[25] , \wRegInB56[5] , 
        \ScanLink233[15] , \ScanLink196[12] , \wBMid24[11] , \wBMid67[24] , 
        \wBMid72[10] , \ScanLink38[11] , \wRegInA36[0] , \ScanLink210[24] , 
        \wBIn123[1] , \wAIn5[12] , \wBMid12[14] , \wBIn66[9] , \wBMid44[15] , 
        \ScanLink205[10] , \ScanLink155[9] , \ScanLink58[15] , \wBMid31[25] , 
        \wAMid91[8] , \ScanLink253[11] , \ScanLink226[21] , \ScanLink183[26] , 
        \wAMid1[4] , \wBMid3[0] , \wBIn9[8] , \wAMid22[7] , \wRegInA6[26] , 
        \wRegInB114[27] , \wRegInB124[4] , \wBMid56[8] , \wBMid97[30] , 
        \wAIn62[3] , \wBMid99[1] , \wBMid112[5] , \wRegInB101[13] , 
        \wBMid97[29] , \wRegInB0[23] , \wAMid13[12] , \wAMid25[17] , 
        \wAMid73[16] , \wAIn86[31] , \wAIn86[28] , \wBIn87[10] , 
        \wAMid119[20] , \wBMid123[20] , \wRegInB122[22] , \wAMid88[17] , 
        \wBMid100[11] , \wBIn92[24] , \wBMid115[25] , \ScanLink254[5] , 
        \ScanLink2[22] , \wRegInA57[9] , \wRegInA98[0] , \ScanLink134[0] , 
        \wAMid30[23] , \wAMid50[27] , \wAMid45[13] , \wRegInB47[30] , 
        \wRegInB64[18] , \ScanLink137[3] , \wRegInB11[28] , \wBMid48[4] , 
        \wAMid66[22] , \wRegInB47[29] , \wBIn69[25] , \wRegInB32[19] , 
        \wRegInB127[7] , \wRegInB11[31] , \wRegInB29[0] , \wBMid19[18] , 
        \wAIn61[0] , \ScanLink238[19] , \ScanLink26[29] , \wRegInA49[5] , 
        \ScanLink70[31] , \ScanLink53[19] , \wAMid21[4] , \ScanLink26[30] , 
        \wBMid111[6] , \wRegInA119[16] , \ScanLink70[28] , \wRegInB53[8] , 
        \wBMid1[24] , \wAMid2[7] , \wAMid13[21] , \wAMid30[10] , \wAMid45[20] , 
        \wAMid45[0] , \wAMid46[3] , \wBIn63[4] , \wBIn92[17] , \wBMid115[16] , 
        \wAMid119[13] , \wAMid119[2] , \wRegInA111[2] , \ScanLink230[1] , 
        \ScanLink2[11] , \ScanLink150[4] , \wBIn87[23] , \wAMid94[5] , 
        \wBMid123[13] , \wRegInA79[18] , \wAMid88[24] , \wBMid100[22] , 
        \wRegInB0[10] , \wRegInB101[20] , \ScanLink106[28] , \ScanLink173[18] , 
        \ScanLink150[30] , \wRegInB114[14] , \wRegInB122[11] , 
        \ScanLink182[2] , \ScanLink150[29] , \ScanLink125[19] , 
        \ScanLink106[31] , \ScanLink73[9] , \wRegInA6[15] , \wRegInA119[25] , 
        \ScanLink188[19] , \wAIn115[19] , \ScanLink181[1] , \wRegInA112[1] , 
        \wAMid66[11] , \wBIn69[16] , \ScanLink233[2] , \wAMid25[24] , 
        \wAMid50[14] , \wAMid73[25] , \wAMid97[6] , \wRegInA82[19] , 
        \wBIn60[7] , \ScanLink153[7] , \wAIn4[18] , \wAMid81[2] , 
        \wRegInB89[6] , \wRegInA104[5] , \wRegInA125[15] , \wRegInA106[24] , 
        \ScanLink225[6] , \ScanLink197[18] , \wBIn9[30] , \wBIn9[29] , 
        \wAIn10[3] , \wAIn13[0] , \wBIn16[13] , \wBIn20[16] , \wBIn76[3] , 
        \wRegInA113[10] , \ScanLink145[3] , \wBIn55[26] , \wBIn76[17] , 
        \wAMid79[10] , \wBIn115[26] , \wRegInB94[9] , \ScanLink238[9] , 
        \wAMid19[14] , \wAMid53[4] , \wBIn35[22] , \wBIn63[23] , \wBIn100[12] , 
        \wBIn40[12] , \wAMid82[11] , \wBIn123[23] , \ScanLink197[5] , 
        \wRegInB58[3] , \wAMid112[9] , \wAMid113[26] , \wBMid24[8] , 
        \wAMid50[7] , \wAMid97[25] , \wBIn98[22] , \wAMid106[12] , 
        \wRegInA38[6] , \wRegInA45[28] , \wRegInA13[30] , \wRegInA30[18] , 
        \ScanLink194[6] , \ScanLink8[24] , \wAMid125[23] , \wRegInA45[31] , 
        \wRegInA66[19] , \wRegInA13[29] , \wRegInA107[6] , \ScanLink226[5] , 
        \ScanLink119[29] , \wBIn16[20] , \wBMid39[7] , \wBIn75[0] , 
        \wRegInA25[9] , \ScanLink119[30] , \ScanLink78[2] , \ScanLink189[9] , 
        \ScanLink146[0] , \wAMid82[1] , \wBIn63[10] , \wBIn100[21] , 
        \wAIn17[18] , \wAMid19[27] , \wBIn20[25] , \wAIn34[29] , \wBIn35[11] , 
        \wBIn40[21] , \wBIn123[10] , \wAIn41[19] , \wBIn55[15] , \wAIn77[4] , 
        \wRegInA90[8] , \wAIn62[31] , \wRegInB58[31] , \wAIn34[30] , 
        \wAMid37[0] , \wAIn62[28] , \wBIn115[15] , \wAMid79[23] , \wBIn76[24] , 
        \wRegInB58[28] , \wBMid25[31] , \wBMid107[2] , \wRegInA113[23] , 
        \wRegInA125[26] , \ScanLink252[31] , \ScanLink252[28] , 
        \ScanLink227[18] , \ScanLink204[30] , \ScanLink241[2] , 
        \ScanLink204[29] , \ScanLink121[7] , \wBIn2[3] , \wBMid1[17] , 
        \wBIn12[7] , \wBMid73[29] , \wBIn11[4] , \wBMid25[28] , \wAIn123[0] , 
        \ScanLink39[28] , \wRegInA106[17] , \wBMid50[18] , \wBMid91[9] , 
        \wAIn69[8] , \wBMid73[30] , \wBMid88[31] , \wRegInB21[8] , 
        \ScanLink39[31] , \ScanLink242[1] , \ScanLink94[28] , \wBMid88[28] , 
        \wAIn120[3] , \ScanLink122[4] , \wAMid34[3] , \wAMid97[16] , 
        \wBIn98[11] , \wAMid106[21] , \ScanLink94[31] , \wAMid125[10] , 
        \ScanLink8[17] , \wAIn74[7] , \wAMid82[22] , \wAIn99[29] , 
        \wBMid104[1] , \wRegInB80[18] , \wAIn99[30] , \wAMid113[15] , 
        \wRegInB10[11] , \wRegInB33[20] , \wRegInA96[27] , \wRegInB40[1] , 
        \wRegInB46[10] , \ScanLink223[8] , \wRegInA20[4] , \wRegInB65[21] , 
        \wBIn2[16] , \wBMid18[21] , \wAMid48[5] , \wRegInB70[15] , 
        \wAIn69[24] , \wRegInB26[14] , \wRegInA83[13] , \wAIn122[16] , 
        \wRegInB0[1] , \wRegInB53[24] , \wRegInB92[7] , \ScanLink189[13] , 
        \ScanLink71[11] , \wBMid21[5] , \wBMid78[25] , \wAIn101[27] , 
        \ScanLink60[0] , \ScanLink52[20] , \ScanLink27[10] , \wAIn114[13] , 
        \wAMid117[4] , \ScanLink47[14] , \ScanLink32[24] , \ScanLink239[20] , 
        \ScanLink64[25] , \wAMid56[9] , \wBMid96[10] , \ScanLink11[15] , 
        \wAMid99[0] , \wRegInB91[4] , \ScanLink151[23] , \ScanLink124[13] , 
        \ScanLink63[3] , \ScanLink107[22] , \ScanLink172[12] , 
        \ScanLink112[16] , \ScanLink167[26] , \wBMid18[12] , \wBMid22[6] , 
        \wBMid45[1] , \wBMid78[16] , \wBMid83[24] , \wAMid114[7] , 
        \ScanLink131[27] , \wBIn86[30] , \wBIn86[29] , \wAIn87[11] , 
        \wRegInA18[16] , \wRegInB43[2] , \wRegInA101[8] , \ScanLink192[8] , 
        \ScanLink144[17] , \wAIn92[25] , \wRegInB3[2] , \wRegInA78[12] , 
        \wBMid101[28] , \wBMid101[31] , \wAMid109[8] , \wAMid118[19] , 
        \wBMid122[19] , \wRegInA23[7] , \wAIn114[20] , \ScanLink32[17] , 
        \wAIn122[25] , \ScanLink239[13] , \ScanLink47[27] , \ScanLink11[26] , 
        \ScanLink64[16] , \ScanLink189[20] , \ScanLink71[22] , \wAIn101[14] , 
        \wRegInA96[6] , \ScanLink27[23] , \wRegInB70[26] , \ScanLink52[13] , 
        \wAIn0[30] , \wAIn0[29] , \wBIn2[25] , \wAMid12[18] , \wAIn69[17] , 
        \wRegInB24[5] , \wRegInB53[17] , \wRegInB26[27] , \wRegInA83[20] , 
        \wBIn14[9] , \wAMid31[30] , \wAMid31[29] , \wAMid67[28] , \wBMid97[7] , 
        \wRegInB46[23] , \wRegInB33[13] , \wRegInA96[14] , \wAMid44[19] , 
        \wRegInA44[0] , \wRegInB65[12] , \wAMid67[31] , \ScanLink127[9] , 
        \wRegInB10[22] , \wAIn87[22] , \wAIn92[16] , \wRegInA78[21] , 
        \wRegInB27[6] , \wRegInA47[3] , \ScanLink3[31] , \wBMid94[4] , 
        \ScanLink3[28] , \wRegInA18[25] , \ScanLink167[15] , \wBIn6[27] , 
        \wBIn6[14] , \wBMid46[2] , \wAIn72[9] , \wBMid83[17] , 
        \ScanLink144[24] , \ScanLink112[25] , \ScanLink131[14] , 
        \wRegInA95[5] , \ScanLink151[10] , \wBMid96[23] , \wRegInB1[29] , 
        \wRegInB123[28] , \ScanLink139[5] , \ScanLink124[20] , 
        \ScanLink172[21] , \wAIn83[13] , \wAIn84[9] , \wAIn96[27] , 
        \wRegInB1[30] , \wRegInB100[19] , \wRegInB123[31] , \ScanLink107[11] , 
        \wRegInA63[5] , \wAMid98[18] , \ScanLink7[19] , \wRegInA69[24] , 
        \ScanLink163[24] , \ScanLink116[14] , \wAMid15[8] , \wBMid62[4] , 
        \wBMid126[9] , \wBMid87[26] , \wAIn99[6] , \ScanLink135[25] , 
        \wBMid92[12] , \wRegInB5[18] , \ScanLink140[15] , \wAIn110[11] , 
        \wRegInB127[19] , \wRegInB104[31] , \wRegInB104[28] , \wRegInB110[8] , 
        \ScanLink155[21] , \ScanLink120[11] , \ScanLink23[1] , 
        \ScanLink103[20] , \ScanLink176[10] , \ScanLink43[16] , 
        \ScanLink198[25] , \ScanLink36[26] , \wAMid16[30] , \wAMid16[29] , 
        \wAIn18[16] , \wAIn48[3] , \wBMid61[7] , \wRegInA109[19] , 
        \ScanLink248[12] , \ScanLink60[27] , \wBMid69[13] , \wAIn126[14] , 
        \ScanLink228[16] , \ScanLink75[13] , \ScanLink15[17] , 
        \ScanLink56[22] , \wAIn105[25] , \ScanLink23[12] , \wRegInA60[6] , 
        \ScanLink20[2] , \wAIn101[8] , \wRegInB22[16] , \wRegInB74[17] , 
        \wRegInB57[26] , \wRegInA87[11] , \wAMid40[31] , \wAMid63[19] , 
        \wAIn78[12] , \wRegInB37[22] , \wRegInA92[25] , \wAMid35[18] , 
        \wAMid40[28] , \wRegInB42[12] , \wRegInB14[13] , \wBMid92[21] , 
        \wRegInB61[23] , \ScanLink155[12] , \ScanLink179[7] , 
        \ScanLink120[22] , \ScanLink176[23] , \ScanLink163[17] , 
        \ScanLink103[13] , \ScanLink6[9] , \wBMid5[26] , \wAIn8[2] , 
        \wBIn57[8] , \wBMid87[15] , \ScanLink219[2] , \ScanLink140[26] , 
        \ScanLink116[27] , \ScanLink135[16] , \wBIn112[0] , \ScanLink47[5] , 
        \wAIn83[20] , \wBIn98[1] , \ScanLink164[8] , \wRegInA69[17] , 
        \wAMid10[5] , \wAIn18[25] , \wAIn78[21] , \wBIn82[18] , \wAIn96[14] , 
        \wBMid105[19] , \wRegInB67[4] , \wBMid126[31] , \wBMid126[28] , 
        \wRegInB42[21] , \ScanLink95[3] , \wBIn111[3] , \wRegInB37[11] , 
        \wRegInA92[16] , \wRegInB14[20] , \wRegInB61[10] , \wRegInB57[15] , 
        \wRegInB64[7] , \wRegInB74[24] , \ScanLink96[0] , \ScanLink59[9] , 
        \wAIn31[8] , \wBMid69[20] , \wBIn79[19] , \wRegInB22[25] , 
        \wRegInA87[22] , \wAIn126[27] , \wRegInA9[8] , \ScanLink228[25] , 
        \ScanLink75[20] , \ScanLink23[21] , \wBIn35[2] , \wBIn49[4] , 
        \wAIn105[16] , \ScanLink56[11] , \wAIn82[7] , \wAIn110[22] , 
        \wRegInB79[8] , \ScanLink248[21] , \ScanLink44[6] , \ScanLink36[15] , 
        \ScanLink43[25] , \ScanLink198[16] , \ScanLink15[24] , 
        \ScanLink60[14] , \wAIn104[5] , \ScanLink106[2] , \wAIn50[1] , 
        \wBMid79[5] , \wRegInA8[22] , \ScanLink90[19] , \ScanLink38[0] , 
        \wAMid93[27] , \wAMid102[10] , \wRegInA78[4] , \wBIn12[11] , 
        \wAMid13[6] , \wAMid86[13] , \wBMid120[7] , \wAMid121[21] , 
        \wRegInB18[1] , \wRegInB116[6] , \wBIn89[14] , \wAMid117[24] , 
        \wRegInB84[30] , \wRegInB84[29] , \wAIn13[30] , \wBIn24[14] , 
        \wBIn31[20] , \wBIn67[21] , \wBMid67[9] , \wBMid123[4] , \wAMid68[26] , 
        \wBIn104[10] , \wBIn44[10] , \wAIn53[2] , \wBIn127[21] , \wAIn13[29] , 
        \wAIn30[18] , \wAIn45[28] , \wRegInB29[30] , \wBIn51[24] , 
        \wRegInB115[5] , \wBIn36[1] , \wAIn45[31] , \wBIn72[15] , 
        \wBIn111[24] , \wRegInB29[29] , \wAIn66[19] , \wAIn81[4] , 
        \wRegInA66[8] , \wRegInA117[12] , \ScanLink256[19] , \ScanLink223[29] , 
        \wAIn107[6] , \ScanLink223[30] , \ScanLink200[18] , \ScanLink105[1] , 
        \wBMid5[15] , \wBMid21[19] , \wBMid54[30] , \wBMid77[18] , 
        \wBMid54[29] , \wRegInA121[17] , \ScanLink48[29] , \wAIn34[5] , 
        \wAMid74[1] , \wRegInA102[26] , \ScanLink48[30] , \wAMid86[20] , 
        \wBIn89[27] , \wBIn109[1] , \wBIn51[6] , \wBIn83[0] , \wAMid117[17] , 
        \wAMid93[14] , \wAMid102[23] , \wAMid121[12] , \wRegInA34[29] , 
        \wRegInA41[19] , \wRegInA62[31] , \wRegInA17[18] , \wRegInA34[30] , 
        \ScanLink0[7] , \wRegInA8[11] , \wRegInA62[28] , \ScanLink168[28] , 
        \wBIn52[5] , \wRegInA121[24] , \wRegInA123[0] , \ScanLink168[31] , 
        \ScanLink162[6] , \ScanLink202[3] , \ScanLink193[30] , 
        \ScanLink161[5] , \wRegInB62[9] , \wRegInA102[15] , \ScanLink193[29] , 
        \wRegInA117[21] , \ScanLink201[0] , \wRegInA120[3] , \wAIn0[24] , 
        \wAIn0[7] , \wBMid0[23] , \wBIn12[22] , \wBIn24[27] , \wAIn37[6] , 
        \wBIn51[17] , \wBIn80[3] , \wBIn67[12] , \wBIn72[26] , \wBIn111[17] , 
        \wAMid77[2] , \wAMid68[15] , \wBIn104[23] , \wRegInA99[29] , 
        \ScanLink3[4] , \wBIn31[13] , \wBIn44[23] , \wBIn127[12] , 
        \wRegInA99[30] , \wRegInA114[2] , \ScanLink246[31] , \ScanLink42[8] , 
        \wBMid0[10] , \wAMid1[31] , \wAMid4[4] , \wRegInB56[8] , 
        \wRegInB99[1] , \wRegInA124[12] , \ScanLink210[29] , \ScanLink246[28] , 
        \ScanLink235[1] , \ScanLink233[18] , \ScanLink210[30] , \wBMid5[3] , 
        \wAMid7[7] , \wBMid12[19] , \wBMid31[28] , \wBMid44[18] , 
        \wRegInA107[23] , \wBMid67[30] , \wAMid91[5] , \wRegInA112[17] , 
        \wBMid67[29] , \wBIn17[14] , \wAMid18[13] , \wBIn21[11] , 
        \wBMid31[31] , \wBIn66[4] , \ScanLink58[18] , \ScanLink155[4] , 
        \wAMid43[3] , \wBIn54[21] , \ScanLink76[9] , \wBIn77[10] , 
        \wBIn114[21] , \wAMid78[17] , \wAIn20[30] , \wAIn20[29] , \wBIn62[24] , 
        \wAIn76[28] , \wBIn101[15] , \wRegInB39[18] , \wBIn34[25] , 
        \wAMid40[0] , \wBIn41[15] , \wAIn76[31] , \wAIn55[19] , \wBIn78[8] , 
        \wAMid83[16] , \wBIn122[24] , \ScanLink187[2] , \wRegInB48[4] , 
        \wAMid107[15] , \wAMid112[21] , \wRegInA28[1] , \wAMid96[22] , 
        \wRegInB94[18] , \ScanLink184[1] , \wBIn99[25] , \ScanLink9[23] , 
        \wRegInB8[4] , \wAMid124[24] , \wBMid29[0] , \wBIn65[7] , 
        \wRegInA117[1] , \ScanLink236[2] , \ScanLink156[7] , \ScanLink80[31] , 
        \ScanLink68[5] , \wAMid92[6] , \ScanLink80[28] , \wBIn62[17] , 
        \wBIn101[26] , \wRegInB121[4] , \wBIn17[27] , \wAMid18[20] , 
        \wBIn21[22] , \wBIn34[16] , \wBIn41[26] , \wBIn122[17] , \wBIn54[12] , 
        \wAIn67[3] , \wAMid27[7] , \wBIn77[23] , \wBIn114[12] , 
        \wRegInA89[18] , \wAMid78[24] , \wBMid53[8] , \wBMid117[5] , 
        \wRegInA112[24] , \ScanLink183[18] , \wAMid1[28] , \ScanLink251[5] , 
        \wRegInA52[9] , \wRegInA124[21] , \ScanLink131[0] , \wAMid1[9] , 
        \wBIn3[11] , \wBMid6[0] , \wAMid107[26] , \wBMid109[9] , 
        \wRegInA107[10] , \ScanLink252[6] , \ScanLink178[19] , 
        \ScanLink132[3] , \wAMid124[17] , \wAIn18[6] , \wAMid24[4] , 
        \wAMid96[11] , \wRegInB122[7] , \wBIn99[16] , \ScanLink9[10] , 
        \wAMid50[19] , \wAIn64[0] , \wAMid83[25] , \wBMid114[6] , 
        \wRegInA51[31] , \wRegInA72[19] , \wRegInA24[18] , \wAMid112[12] , 
        \wBIn125[2] , \wRegInB11[16] , \wRegInB32[27] , \wRegInA51[28] , 
        \wRegInB47[17] , \wRegInB50[6] , \wRegInA97[20] , \wRegInA30[3] , 
        \wRegInB64[26] , \wAMid73[31] , \wBMid19[26] , \wAMid25[30] , 
        \wAMid25[29] , \wRegInB71[12] , \wAMid58[2] , \wAIn68[23] , 
        \wRegInB27[13] , \wRegInA82[14] , \wAMid73[28] , \wRegInB52[23] , 
        \wAIn123[11] , \wRegInB82[0] , \wRegInA119[28] , \ScanLink70[16] , 
        \ScanLink188[14] , \wRegInA119[31] , \ScanLink53[27] , \wBMid31[2] , 
        \wBMid79[22] , \wAIn100[20] , \ScanLink26[17] , \wAMid107[3] , 
        \ScanLink70[7] , \ScanLink46[13] , \wAIn115[14] , \ScanLink238[27] , 
        \ScanLink33[23] , \ScanLink65[22] , \wAMid89[7] , \wBMid97[17] , 
        \ScanLink10[12] , \wRegInB81[3] , \ScanLink150[24] , \ScanLink125[14] , 
        \ScanLink73[4] , \ScanLink173[15] , \ScanLink106[25] , \wRegInA6[18] , 
        \wRegInB114[19] , \ScanLink113[11] , \ScanLink166[21] , \wBMid32[1] , 
        \wBMid82[23] , \wAMid104[0] , \ScanLink130[20] , \wRegInA19[11] , 
        \wRegInB53[5] , \ScanLink145[10] , \wAIn3[4] , \wBIn3[22] , 
        \wBIn19[1] , \wBMid19[15] , \wAMid21[9] , \wBIn63[9] , \wAIn86[16] , 
        \wAMid88[29] , \wAIn93[22] , \wAMid94[8] , \wRegInA79[15] , 
        \wBIn126[1] , \wRegInA33[0] , \ScanLink150[9] , \wBMid79[11] , 
        \wAMid88[30] , \wAIn115[27] , \ScanLink238[14] , \ScanLink46[20] , 
        \ScanLink33[10] , \ScanLink14[3] , \ScanLink10[21] , \ScanLink65[11] , 
        \wBMid55[6] , \wAIn123[22] , \ScanLink188[27] , \ScanLink70[25] , 
        \wAIn100[13] , \wRegInA49[8] , \wRegInA86[1] , \ScanLink26[24] , 
        \ScanLink53[14] , \wBMid48[9] , \wAIn68[10] , \wRegInB27[20] , 
        \wRegInB34[2] , \wRegInB52[10] , \wRegInB71[21] , \wRegInA82[27] , 
        \wBIn69[28] , \wBMid87[0] , \wRegInB47[24] , \wRegInB32[14] , 
        \wRegInA97[13] , \wBIn69[31] , \wRegInA54[7] , \wRegInB64[15] , 
        \wBMid84[3] , \wAIn86[25] , \wBIn92[30] , \wAIn93[11] , 
        \wRegInB11[25] , \wRegInA79[26] , \wRegInB37[1] , \ScanLink254[8] , 
        \wBMid115[31] , \wRegInA57[4] , \wBIn92[29] , \wBMid115[28] , 
        \wRegInA19[22] , \wRegInB124[9] , \ScanLink166[12] , \wBMid4[21] , 
        \wAMid5[19] , \wAIn6[9] , \wBIn7[20] , \wBIn7[13] , \wBIn9[5] , 
        \wBMid82[10] , \ScanLink249[7] , \ScanLink145[23] , \ScanLink113[22] , 
        \ScanLink130[13] , \wBMid97[24] , \wRegInA85[2] , \ScanLink17[0] , 
        \ScanLink150[17] , \ScanLink129[2] , \ScanLink125[27] , \wBMid56[5] , 
        \wBMid112[8] , \ScanLink173[26] , \wAIn82[14] , \wBIn96[18] , 
        \wAIn97[20] , \ScanLink106[16] , \wAMid108[31] , \wAMid108[28] , 
        \wRegInA73[2] , \wRegInB13[7] , \wBMid111[19] , \wRegInA68[23] , 
        \ScanLink162[23] , \ScanLink117[13] , \wBMid16[7] , \wBIn18[30] , 
        \wBIn18[29] , \wAMid18[0] , \wBIn20[8] , \wAIn46[8] , \wBMid72[3] , 
        \wAIn58[4] , \wBMid68[14] , \wBMid71[0] , \wBMid86[21] , 
        \ScanLink134[22] , \wAIn89[1] , \wBMid93[15] , \ScanLink141[12] , 
        \wAIn111[16] , \ScanLink177[17] , \ScanLink154[26] , \ScanLink121[16] , 
        \ScanLink33[6] , \ScanLink102[27] , \ScanLink42[11] , 
        \ScanLink249[15] , \ScanLink199[22] , \ScanLink37[21] , 
        \ScanLink61[20] , \wAIn127[13] , \ScanLink229[11] , \ScanLink74[14] , 
        \ScanLink14[10] , \ScanLink57[25] , \ScanLink22[15] , \wAIn104[22] , 
        \ScanLink30[5] , \wRegInA70[1] , \wRegInB75[10] , \ScanLink113[8] , 
        \wAIn19[11] , \wRegInB23[11] , \wRegInA86[16] , \wRegInB56[21] , 
        \wAIn79[15] , \wRegInB10[4] , \wRegInB36[25] , \wRegInA93[22] , 
        \wRegInB15[14] , \wRegInB43[15] , \wAMid62[8] , \wBMid93[26] , 
        \wAMid120[6] , \wRegInB60[24] , \ScanLink154[15] , \wBIn95[9] , 
        \ScanLink169[0] , \ScanLink121[25] , \ScanLink177[24] , 
        \ScanLink162[10] , \ScanLink102[14] , \wAIn19[22] , \wAMid21[18] , 
        \wAIn79[26] , \wAIn82[27] , \wBMid86[12] , \wRegInA2[29] , 
        \wRegInB110[28] , \ScanLink209[5] , \ScanLink117[20] , 
        \wRegInB110[31] , \ScanLink141[21] , \ScanLink134[11] , \wBIn88[6] , 
        \wBIn102[7] , \wRegInA2[30] , \ScanLink57[2] , \wRegInA17[6] , 
        \wAIn97[13] , \wRegInA7[3] , \wRegInA68[10] , \wRegInB77[3] , 
        \wRegInA4[0] , \ScanLink85[4] , \wRegInB43[26] , \wBIn101[4] , 
        \wRegInB36[16] , \wRegInA93[11] , \wRegInA14[5] , \wRegInB15[27] , 
        \wRegInB60[17] , \wRegInB75[23] , \wAMid54[28] , \wRegInB56[12] , 
        \wRegInB74[0] , \ScanLink86[7] , \ScanLink8[2] , \wAMid54[31] , 
        \wAMid77[19] , \wRegInB23[22] , \wRegInA86[25] , \wAIn127[20] , 
        \ScanLink217[9] , \wBIn13[16] , \wBMid15[4] , \ScanLink229[22] , 
        \ScanLink74[27] , \wBIn25[5] , \wBIn59[3] , \wBMid68[27] , 
        \wAMid123[5] , \ScanLink22[26] , \wAIn104[11] , \ScanLink57[16] , 
        \wAIn92[0] , \wAIn111[25] , \ScanLink249[26] , \ScanLink54[1] , 
        \ScanLink37[12] , \ScanLink42[22] , \ScanLink199[11] , 
        \ScanLink14[23] , \ScanLink61[13] , \wAIn114[2] , \ScanLink116[5] , 
        \wAIn40[6] , \wBMid69[2] , \ScanLink109[18] , \wRegInA9[25] , 
        \wRegInB15[9] , \ScanLink28[7] , \wAMid87[14] , \wBIn88[13] , 
        \wAMid92[20] , \wAMid103[17] , \wRegInA68[3] , \wAMid120[26] , 
        \wRegInA76[28] , \wRegInB106[1] , \wAMid116[23] , \wRegInA20[30] , 
        \wRegInA20[29] , \wRegInA55[19] , \wRegInA76[31] , \ScanLink35[8] , 
        \wBIn25[13] , \wBIn30[27] , \wBIn66[26] , \wAMid69[21] , \wBIn105[17] , 
        \wAIn43[5] , \wBIn45[17] , \wBIn126[26] , \ScanLink108[9] , 
        \wBIn50[23] , \wBIn73[12] , \wBIn110[23] , \wRegInB105[2] , 
        \wRegInA116[15] , \ScanLink187[29] , \wBIn26[6] , \wAIn91[3] , 
        \wAIn117[1] , \ScanLink187[30] , \ScanLink115[6] , \wBMid10[9] , 
        \wAMid64[6] , \wRegInA103[21] , \wRegInA120[10] , \wBIn88[20] , 
        \wBMid4[12] , \wAIn24[2] , \wAMid87[27] , \wBIn119[6] , \wBIn41[1] , 
        \wAMid79[9] , \wAIn89[18] , \wAMid92[13] , \wBIn93[7] , \wAMid116[10] , 
        \wAMid126[8] , \wAMid103[24] , \wAMid120[15] , \wRegInB90[29] , 
        \wRegInB90[30] , \wBIn104[9] , \wRegInA9[16] , \wRegInA11[8] , 
        \wBIn42[2] , \wBMid98[19] , \ScanLink172[1] , \wRegInA120[23] , 
        \ScanLink237[30] , \ScanLink212[4] , \ScanLink84[19] , 
        \ScanLink214[18] , \ScanLink171[2] , \wBMid16[31] , \wBMid35[19] , 
        \wRegInA103[12] , \ScanLink237[29] , \ScanLink242[19] , \wBMid16[28] , 
        \wBMid40[29] , \wRegInA116[26] , \ScanLink211[7] , \wBIn25[20] , 
        \wAIn27[1] , \wBMid40[30] , \wBMid63[18] , \ScanLink29[19] , 
        \ScanLink80[9] , \wBIn50[10] , \wBIn90[4] , \wAMid67[5] , 
        \wBIn110[10] , \wBIn73[21] , \wAMid4[20] , \wBIn6[19] , \wBIn13[25] , 
        \wAIn51[31] , \wBIn66[15] , \wAMid69[12] , \wAIn72[19] , \wBIn105[24] , 
        \wAMid15[5] , \wAMid16[24] , \wAMid16[17] , \wBIn19[10] , \wAIn24[18] , 
        \wBIn30[14] , \wBIn45[24] , \wAIn51[28] , \wRegInB48[19] , 
        \wBIn126[15] , \wAIn31[5] , \wAMid35[26] , \wBIn49[9] , \wBIn86[0] , 
        \wRegInA19[0] , \wAMid71[1] , \wRegInA9[5] , \ScanLink228[31] , 
        \wRegInB79[5] , \ScanLink228[28] , \ScanLink5[7] , \wRegInA109[27] , 
        \ScanLink43[31] , \ScanLink15[29] , \ScanLink60[19] , \ScanLink43[28] , 
        \ScanLink36[18] , \ScanLink15[30] , \wAMid40[16] , \ScanLink167[6] , 
        \wBIn54[6] , \wAIn18[31] , \wAIn18[28] , \wBMid18[1] , \wAMid63[27] , 
        \wRegInB57[18] , \wRegInB74[30] , \wAMid20[12] , \wAMid76[13] , 
        \wRegInB22[28] , \ScanLink207[3] , \wBIn79[14] , \wRegInB74[29] , 
        \wRegInA126[0] , \wBIn19[23] , \wAMid20[21] , \wBIn30[2] , \wAIn32[6] , 
        \wAMid55[22] , \wRegInB22[31] , \ScanLink59[4] , \wBIn57[5] , 
        \wBIn97[21] , \wAMid98[26] , \wBMid110[20] , \ScanLink7[27] , 
        \wAMid72[2] , \wBIn82[15] , \wAIn96[19] , \wAMid109[11] , 
        \wBMid126[25] , \ScanLink164[5] , \wRegInA125[3] , \wBMid105[14] , 
        \wRegInB67[9] , \ScanLink204[0] , \wRegInB104[16] , \wAMid55[11] , 
        \wAMid76[20] , \wBIn85[3] , \wRegInB5[26] , \wBMid87[18] , 
        \wRegInB127[27] , \ScanLink88[1] , \ScanLink47[8] , \wRegInA3[23] , 
        \wRegInB111[22] , \ScanLink6[4] , \wBIn79[27] , \wAIn87[7] , 
        \wAIn101[5] , \wAMid35[15] , \wAMid40[25] , \ScanLink103[2] , 
        \wRegInA92[31] , \wAMid63[14] , \wRegInA92[28] , \wAMid16[6] , 
        \wAIn55[1] , \wBMid125[7] , \wRegInA109[14] , \ScanLink198[28] , 
        \ScanLink198[31] , \wAIn56[2] , \wAIn105[31] , \wAIn105[28] , 
        \wAIn126[19] , \wRegInB113[6] , \ScanLink135[28] , \wRegInB111[11] , 
        \ScanLink163[30] , \ScanLink140[18] , \ScanLink116[19] , 
        \ScanLink135[31] , \wBMid62[9] , \wRegInA3[10] , \ScanLink163[29] , 
        \wBMid126[4] , \wBMid5[18] , \wAIn13[17] , \wBIn33[1] , \wAIn84[4] , 
        \wRegInB127[14] , \wRegInB5[15] , \wRegInB104[25] , \wRegInB110[5] , 
        \wAIn102[6] , \wRegInA63[8] , \ScanLink100[1] , \wAIn66[27] , 
        \wBIn82[26] , \wBMid105[27] , \wBMid126[16] , \wBIn97[12] , 
        \wAMid98[15] , \wBMid110[13] , \wAMid109[22] , \wRegInA69[29] , 
        \ScanLink7[14] , \wRegInB29[17] , \wRegInA69[30] , \wBMid21[27] , 
        \wAIn25[12] , \wAIn30[26] , \wAIn45[16] , \wAIn50[22] , \wAMid68[18] , 
        \wAIn73[13] , \ScanLink42[5] , \ScanLink3[9] , \wRegInB49[13] , 
        \wRegInA99[24] , \wRegInA121[30] , \ScanLink236[23] , 
        \ScanLink193[24] , \wBMid54[17] , \wRegInA102[18] , \ScanLink243[13] , 
        \wBIn117[0] , \ScanLink215[12] , \wRegInA121[29] , \ScanLink161[8] , 
        \ScanLink48[17] , \wBMid17[22] , \wBIn52[8] , \wBMid77[26] , 
        \ScanLink200[26] , \wBMid34[13] , \wBMid62[12] , \ScanLink28[13] , 
        \wRegInB62[4] , \ScanLink90[3] , \wBMid41[23] , \ScanLink223[17] , 
        \ScanLink186[10] , \wAIn0[17] , \wAMid4[13] , \wAIn29[7] , 
        \wBIn114[3] , \ScanLink256[27] , \wAIn34[8] , \wAMid69[3] , 
        \wBMid99[13] , \wRegInB61[7] , \ScanLink168[25] , \ScanLink108[21] , 
        \ScanLink90[27] , \ScanLink85[13] , \wRegInA21[10] , \wRegInB84[17] , 
        \ScanLink93[0] , \wBMid62[21] , \wAIn81[9] , \wAIn88[12] , 
        \wRegInA17[15] , \wRegInA54[20] , \wRegInA77[11] , \wAMid93[19] , 
        \wRegInA34[24] , \wRegInA62[25] , \wRegInA41[14] , \wRegInB91[23] , 
        \ScanLink41[6] , \wRegInA66[5] , \ScanLink28[20] , \wBMid17[11] , 
        \wBMid41[10] , \ScanLink200[15] , \wAMid0[22] , \wBIn9[17] , 
        \wAMid10[8] , \wAIn13[24] , \wBMid21[14] , \wBMid34[20] , 
        \ScanLink256[14] , \wBMid54[24] , \ScanLink243[20] , \ScanLink223[24] , 
        \ScanLink186[23] , \wRegInB108[7] , \ScanLink236[10] , 
        \ScanLink193[17] , \wAIn25[21] , \wBMid77[15] , \ScanLink215[21] , 
        \ScanLink48[24] , \wAIn50[11] , \wBMid67[4] , \wAIn73[20] , 
        \wRegInB49[20] , \ScanLink118[3] , \wBMid123[9] , \wRegInA99[17] , 
        \wBIn24[19] , \wAIn30[15] , \wBIn51[30] , \wAIn66[14] , \wBIn111[29] , 
        \wRegInB29[24] , \wRegInB115[8] , \wBIn72[18] , \wAIn45[25] , 
        \wBIn51[29] , \wBIn111[30] , \ScanLink26[1] , \wAIn88[21] , 
        \wRegInA62[16] , \wBIn11[9] , \wBIn28[0] , \wBMid64[7] , \wAIn119[7] , 
        \wRegInA17[26] , \wRegInA41[27] , \wRegInA78[9] , \wRegInA34[17] , 
        \wRegInB91[10] , \wBMid40[1] , \wBMid79[8] , \wBIn89[19] , 
        \wAMid117[29] , \wRegInA21[23] , \wRegInA54[13] , \wRegInB84[24] , 
        \ScanLink25[2] , \wRegInA77[22] , \wAMid117[30] , \ScanLink85[20] , 
        \wBMid99[20] , \wRegInA65[6] , \ScanLink108[12] , \wAIn104[8] , 
        \wAMid113[18] , \wRegInA13[17] , \ScanLink168[16] , \ScanLink90[14] , 
        \wRegInA25[12] , \wRegInA30[26] , \wRegInA66[27] , \wRegInA45[16] , 
        \wRegInB95[21] , \wRegInB80[15] , \wRegInA50[22] , \wRegInA93[6] , 
        \wAIn69[5] , \wAIn99[24] , \wRegInA73[13] , \wRegInB21[5] , 
        \wRegInA41[0] , \ScanLink179[13] , \ScanLink81[11] , \wBMid88[25] , 
        \wAMid29[1] , \ScanLink122[9] , \ScanLink119[17] , \wBMid92[7] , 
        \wBMid119[3] , \ScanLink94[25] , \wBMid13[20] , \ScanLink59[21] , 
        \ScanLink204[24] , \wAMid0[11] , \wBMid1[30] , \wAIn4[26] , 
        \wBMid8[6] , \wBMid30[11] , \wBMid66[10] , \wRegInB22[6] , 
        \ScanLink227[15] , \ScanLink182[12] , \wBMid45[21] , \ScanLink252[25] , 
        \wBIn9[24] , \wAIn17[15] , \wAIn21[10] , \wBMid25[25] , 
        \ScanLink232[21] , \ScanLink197[26] , \wBMid50[15] , \wBMid91[4] , 
        \ScanLink247[11] , \wAIn54[20] , \wBMid73[24] , \wRegInA42[3] , 
        \ScanLink211[10] , \ScanLink39[25] , \wAIn62[25] , \wBIn76[29] , 
        \wAIn77[11] , \wBIn115[18] , \wRegInB38[21] , \wRegInA88[12] , 
        \wRegInB58[25] , \wBIn20[31] , \wBMid43[2] , \wBIn20[28] , 
        \wAIn41[14] , \wAIn77[9] , \wRegInA90[5] , \wBIn55[18] , \wBIn76[30] , 
        \wAIn34[24] , \wBMid88[16] , \wRegInB45[1] , \wAMid9[1] , \wAIn17[26] , 
        \wBMid24[5] , \wAMid97[28] , \wAIn99[17] , \wRegInB5[1] , 
        \ScanLink226[8] , \ScanLink119[24] , \ScanLink94[16] , 
        \ScanLink81[22] , \wRegInA25[21] , \wRegInA25[4] , \ScanLink179[20] , 
        \wRegInA50[11] , \ScanLink189[4] , \wRegInB80[26] , \ScanLink65[0] , 
        \wRegInA73[20] , \wRegInB97[7] , \ScanLink8[29] , \wRegInA13[24] , 
        \wRegInA66[14] , \wBIn68[2] , \wAMid97[31] , \ScanLink8[30] , 
        \wAMid112[4] , \wRegInA30[15] , \wRegInA45[25] , \wRegInB95[12] , 
        \wRegInB58[16] , \wRegInB94[4] , \wAIn62[16] , \wRegInA88[21] , 
        \ScanLink238[4] , \wAMid19[19] , \wAIn21[23] , \wAIn34[17] , 
        \wRegInA119[7] , \wAIn41[27] , \ScanLink66[3] , \wAIn54[13] , 
        \wAMid111[7] , \ScanLink197[8] , \ScanLink158[1] , \wBMid27[6] , 
        \wAMid53[9] , \wBMid50[26] , \wAIn77[22] , \wRegInB38[12] , 
        \wRegInB46[2] , \ScanLink247[22] , \wBMid1[29] , \wBMid25[16] , 
        \wRegInA106[29] , \ScanLink232[12] , \ScanLink197[15] , \wBMid73[17] , 
        \wBMid66[23] , \wRegInA104[8] , \ScanLink39[16] , \wRegInA106[30] , 
        \ScanLink211[23] , \wRegInA125[18] , \wRegInA26[7] , \wBIn2[31] , 
        \wAIn4[15] , \wBMid13[13] , \ScanLink59[12] , \wBMid45[12] , 
        \ScanLink204[17] , \ScanLink252[16] , \wBMid30[22] , \wRegInB6[2] , 
        \ScanLink227[26] , \ScanLink182[21] , \ScanLink144[29] , \wBIn2[28] , 
        \ScanLink167[18] , \ScanLink131[19] , \ScanLink112[31] , 
        \ScanLink144[30] , \wBIn4[0] , \wBIn17[7] , \wAMid32[0] , 
        \wRegInA7[21] , \wRegInB115[20] , \ScanLink112[28] , \wAIn72[4] , 
        \wBMid89[6] , \wBMid102[2] , \wRegInB100[14] , \wBIn86[17] , 
        \wAMid89[10] , \wAMid118[27] , \wBMid122[27] , \wRegInB1[24] , 
        \wRegInA95[8] , \wRegInB123[25] , \ScanLink139[8] , \wBIn93[23] , 
        \wBMid101[16] , \wBMid114[22] , \ScanLink244[2] , \ScanLink3[25] , 
        \wBMid94[9] , \wRegInA18[28] , \wRegInA88[7] , \wAIn126[0] , 
        \ScanLink124[7] , \wBIn7[3] , \wAMid24[10] , \wAMid72[11] , 
        \wRegInA18[31] , \wRegInB24[8] , \ScanLink247[1] , \wAMid31[24] , 
        \wAMid51[20] , \ScanLink19[6] , \ScanLink127[4] , \wAMid12[15] , 
        \wBIn14[4] , \wAMid44[14] , \wAIn125[3] , \wAIn16[0] , \wAMid31[3] , 
        \wBMid58[3] , \wAMid67[25] , \wBIn68[22] , \wAIn71[7] , \wRegInB39[7] , 
        \wRegInA96[19] , \wAIn101[19] , \wAIn122[31] , \wAIn122[28] , 
        \wRegInA59[2] , \wBIn73[3] , \wBIn93[10] , \wBMid101[1] , 
        \wRegInA118[11] , \wBMid114[11] , \ScanLink3[16] , \wAMid109[5] , 
        \wRegInA101[5] , \ScanLink220[6] , \wAMid118[14] , \wBMid122[14] , 
        \ScanLink140[3] , \wAMid84[2] , \wAIn92[31] , \wBIn86[24] , 
        \wAMid89[23] , \wAIn92[28] , \wBMid101[25] , \wRegInB1[17] , 
        \wRegInB91[9] , \wRegInB100[27] , \wRegInB123[16] , \wAMid56[4] , 
        \wBMid83[30] , \wBMid83[29] , \wRegInB115[13] , \ScanLink192[5] , 
        \wRegInA7[12] , \wAMid12[26] , \wAIn15[3] , \wBMid21[8] , \wAMid55[7] , 
        \wRegInA118[22] , \ScanLink64[28] , \wBMid78[31] , \ScanLink32[30] , 
        \wAMid117[9] , \ScanLink11[18] , \ScanLink64[31] , \ScanLink47[19] , 
        \wAMid31[17] , \wAMid44[27] , \wBMid78[28] , \ScanLink191[6] , 
        \ScanLink32[29] , \wRegInA102[6] , \wAMid67[16] , \wBIn68[11] , 
        \wAMid48[8] , \wRegInB26[19] , \ScanLink223[5] , \wAIn69[29] , 
        \wAMid72[22] , \wAMid87[1] , \wAMid51[13] , \wAIn69[30] , 
        \wRegInA20[9] , \wRegInB53[29] , \wAMid4[30] , \wAMid4[29] , 
        \wBMid5[22] , \wAMid24[23] , \wBIn70[0] , \wRegInB70[18] , 
        \wRegInB53[30] , \wRegInA102[22] , \ScanLink243[29] , \ScanLink143[0] , 
        \ScanLink236[19] , \ScanLink215[31] , \ScanLink243[30] , \wAMid10[1] , 
        \wBIn12[15] , \wBMid17[18] , \wBMid62[28] , \wRegInA121[13] , 
        \ScanLink215[28] , \wAIn81[0] , \ScanLink28[29] , \wAIn107[2] , 
        \wBIn24[10] , \wBMid34[30] , \wBMid34[29] , \wBIn36[5] , \wBMid41[19] , 
        \ScanLink105[5] , \wBMid62[31] , \wRegInA117[16] , \ScanLink28[30] , 
        \wBIn72[11] , \wBIn111[20] , \wRegInB115[1] , \wAIn25[28] , 
        \wBIn51[20] , \ScanLink26[8] , \wBIn31[24] , \wBIn44[14] , \wAIn53[6] , 
        \wRegInB49[30] , \wAIn50[18] , \wAIn73[30] , \wBIn127[25] , 
        \wAMid13[2] , \wAIn25[31] , \wBIn67[25] , \wAMid68[22] , \wAIn73[29] , 
        \wBMid123[0] , \wRegInB49[29] , \wAMid86[17] , \wBIn89[10] , 
        \wBIn104[14] , \wAMid117[20] , \wRegInB18[5] , \wRegInB116[2] , 
        \wAIn88[28] , \wAMid93[23] , \wBIn12[26] , \wBIn28[9] , \wAIn50[5] , 
        \wAIn88[31] , \wBMid120[3] , \wAMid121[25] , \wAMid102[14] , 
        \wRegInA78[0] , \wBIn31[17] , \wBIn35[6] , \wBMid79[1] , \wBMid99[30] , 
        \wRegInA8[26] , \wRegInB91[19] , \ScanLink38[4] , \ScanLink85[29] , 
        \wAIn82[3] , \ScanLink85[30] , \wBMid99[29] , \ScanLink106[6] , 
        \wAIn104[1] , \wBIn44[27] , \wBIn127[16] , \wBIn67[16] , \wAMid68[11] , 
        \wBIn104[27] , \ScanLink3[0] , \wBIn24[23] , \wAIn37[2] , \wBIn72[22] , 
        \wAMid77[6] , \wBIn111[13] , \wBIn51[13] , \wBIn80[7] , 
        \wRegInA120[7] , \wRegInA117[25] , \ScanLink186[19] , \wBIn6[23] , 
        \wBIn6[10] , \wBMid5[11] , \wBIn52[1] , \wBIn117[9] , \wRegInA102[11] , 
        \ScanLink201[4] , \wRegInA121[20] , \ScanLink161[1] , \wAIn18[12] , 
        \wAIn34[1] , \wBIn51[2] , \wRegInA123[4] , \ScanLink202[7] , 
        \ScanLink108[28] , \ScanLink108[31] , \ScanLink93[9] , \wAMid93[10] , 
        \wAMid121[16] , \wRegInA8[15] , \ScanLink162[2] , \ScanLink0[3] , 
        \wAMid102[27] , \wBIn109[5] , \wAMid117[13] , \wRegInA21[19] , 
        \wAMid74[5] , \wBIn83[4] , \wRegInA54[29] , \wAMid76[29] , 
        \wAIn78[16] , \wAMid86[24] , \wBIn89[23] , \wRegInA54[30] , 
        \wRegInA77[18] , \wRegInB14[17] , \wRegInB61[27] , \wRegInB22[12] , 
        \wRegInB37[26] , \wRegInA92[21] , \wRegInB42[16] , \wRegInA87[15] , 
        \wRegInB57[22] , \wAMid20[31] , \wAMid20[28] , \wAIn48[7] , 
        \wAMid55[18] , \wRegInA60[2] , \wAMid76[30] , \wRegInB74[13] , 
        \wAIn55[8] , \wBMid61[3] , \wBMid69[17] , \ScanLink56[26] , 
        \ScanLink23[16] , \wAIn105[21] , \ScanLink20[6] , \wAIn126[10] , 
        \ScanLink228[12] , \ScanLink75[17] , \ScanLink248[16] , 
        \ScanLink198[21] , \ScanLink60[23] , \ScanLink43[12] , 
        \ScanLink15[13] , \wBMid87[22] , \wBMid92[16] , \wAIn110[15] , 
        \ScanLink176[14] , \ScanLink103[24] , \ScanLink36[22] , 
        \ScanLink155[25] , \ScanLink120[15] , \ScanLink23[5] , 
        \ScanLink135[21] , \wAIn99[2] , \wRegInA3[19] , \wRegInB111[18] , 
        \ScanLink140[11] , \ScanLink116[10] , \ScanLink163[20] , \wAIn8[6] , 
        \wAIn18[21] , \wBIn33[8] , \wBMid62[0] , \wAIn83[17] , \wRegInA63[1] , 
        \wRegInA69[20] , \ScanLink100[8] , \wBIn49[0] , \wBMid69[24] , 
        \wAIn96[23] , \wAIn110[26] , \ScanLink248[25] , \ScanLink198[12] , 
        \ScanLink15[20] , \ScanLink60[10] , \ScanLink44[2] , \ScanLink36[11] , 
        \ScanLink43[21] , \ScanLink23[25] , \wBIn86[9] , \wAIn105[12] , 
        \wRegInA19[9] , \ScanLink56[15] , \wAMid71[8] , \wAIn126[23] , 
        \wRegInB57[11] , \wRegInB64[3] , \ScanLink228[21] , \ScanLink75[24] , 
        \wBIn19[19] , \wBIn111[7] , \wRegInB22[21] , \wRegInB74[20] , 
        \wRegInA87[26] , \wRegInA126[9] , \ScanLink96[4] , \wRegInB14[24] , 
        \wRegInB61[14] , \wBMid18[8] , \wAIn78[25] , \wRegInB42[25] , 
        \wAIn83[24] , \wAIn96[10] , \wRegInB37[15] , \wRegInA92[12] , 
        \wRegInB67[0] , \ScanLink95[7] , \ScanLink204[9] , \wBIn97[28] , 
        \wBMid110[29] , \wRegInA69[13] , \wBMid87[11] , \wBIn97[31] , 
        \wBMid110[30] , \wBIn112[4] , \wBIn98[5] , \wAMid109[18] , 
        \ScanLink140[22] , \ScanLink135[12] , \ScanLink88[8] , 
        \ScanLink163[13] , \ScanLink47[1] , \wAIn16[9] , \wAIn87[15] , 
        \wAIn92[21] , \wBMid92[25] , \ScanLink219[6] , \ScanLink116[23] , 
        \ScanLink176[27] , \ScanLink155[16] , \ScanLink103[17] , \wRegInB3[6] , 
        \wRegInA23[3] , \ScanLink179[3] , \ScanLink120[26] , \wRegInA78[16] , 
        \wBIn93[19] , \wRegInA18[12] , \wRegInB43[6] , \wBMid114[18] , 
        \ScanLink131[23] , \wBMid83[20] , \wAMid114[3] , \wAMid99[4] , 
        \ScanLink144[13] , \ScanLink112[12] , \wBIn2[12] , \ScanLink167[22] , 
        \wBMid18[25] , \wBMid21[1] , \wBMid22[2] , \wBMid96[14] , 
        \wRegInB91[0] , \ScanLink172[16] , \ScanLink107[26] , 
        \ScanLink239[24] , \ScanLink151[27] , \ScanLink124[17] , 
        \ScanLink63[7] , \ScanLink64[21] , \wBMid78[21] , \wAIn114[17] , 
        \wAMid117[0] , \ScanLink47[10] , \ScanLink11[11] , \ScanLink52[24] , 
        \ScanLink32[20] , \wAMid48[1] , \wAIn101[23] , \ScanLink27[14] , 
        \wAIn122[12] , \wRegInB92[3] , \ScanLink60[4] , \ScanLink189[17] , 
        \ScanLink71[15] , \wAIn69[20] , \wRegInB26[10] , \wRegInA83[17] , 
        \wAMid87[8] , \wRegInB0[5] , \wRegInA20[0] , \wRegInB53[20] , 
        \wBIn2[21] , \wAMid32[9] , \wBIn68[18] , \wBIn70[9] , \wRegInB10[15] , 
        \wRegInB70[11] , \ScanLink143[9] , \wRegInB65[25] , \wRegInB33[24] , 
        \wRegInB40[5] , \wRegInA96[23] , \wRegInB46[14] , \wBMid46[6] , 
        \ScanLink172[25] , \wBMid83[13] , \wBMid96[27] , \wRegInA95[1] , 
        \ScanLink107[15] , \ScanLink151[14] , \wRegInB115[30] , 
        \ScanLink144[20] , \ScanLink139[1] , \ScanLink124[24] , 
        \ScanLink131[10] , \wRegInA7[31] , \ScanLink167[11] , \wBIn4[9] , 
        \wAIn87[26] , \wRegInA7[28] , \wRegInB115[29] , \ScanLink112[21] , 
        \wBMid94[0] , \wRegInA18[21] , \wAIn126[9] , \wRegInA47[7] , 
        \wAMid24[19] , \wAMid51[30] , \wAMid72[18] , \wAMid89[19] , 
        \wRegInA78[25] , \wAIn92[12] , \wBMid97[3] , \wRegInB10[26] , 
        \wRegInB27[2] , \wRegInA44[4] , \wRegInB65[16] , \wRegInB46[27] , 
        \wRegInB24[1] , \wRegInB33[17] , \wRegInA96[10] , \wRegInB53[13] , 
        \wRegInB26[23] , \wRegInA83[24] , \ScanLink247[8] , \wAIn69[13] , 
        \wRegInB70[22] , \wAMid0[18] , \wAMid9[8] , \wAIn10[7] , \wBMid18[16] , 
        \wAMid51[29] , \wAIn101[10] , \wRegInA96[2] , \ScanLink27[27] , 
        \ScanLink52[17] , \wBMid39[3] , \wBMid45[5] , \wBMid101[8] , 
        \wAIn122[21] , \wRegInA118[18] , \ScanLink71[26] , \wBMid78[12] , 
        \wAIn114[24] , \ScanLink239[17] , \ScanLink189[24] , \ScanLink11[22] , 
        \ScanLink64[12] , \wAMid82[5] , \ScanLink47[23] , \ScanLink32[13] , 
        \wRegInB5[8] , \ScanLink179[29] , \wAMid50[3] , \wBIn75[4] , 
        \ScanLink179[30] , \ScanLink146[4] , \wAMid97[21] , \wRegInB45[8] , 
        \wRegInA107[2] , \ScanLink78[6] , \ScanLink226[1] , \wBIn98[26] , 
        \ScanLink8[20] , \wAMid125[27] , \wAIn13[4] , \wBIn35[26] , 
        \wAMid82[15] , \wAMid106[16] , \wRegInA38[2] , \wAMid113[22] , 
        \wRegInA25[28] , \wRegInA50[18] , \wRegInA73[30] , \ScanLink194[2] , 
        \ScanLink65[9] , \wRegInB58[7] , \wRegInA73[29] , \wRegInA25[31] , 
        \wBIn16[17] , \wAMid19[10] , \wBIn40[16] , \wBIn123[27] , 
        \ScanLink197[1] , \ScanLink158[8] , \wAMid53[0] , \wBIn63[27] , 
        \wBIn76[13] , \wBIn100[16] , \wBIn115[22] , \wRegInA88[28] , 
        \wAMid79[14] , \wBIn20[12] , \wBIn55[22] , \wRegInA88[31] , 
        \wAIn1[27] , \wBIn1[4] , \wBIn2[7] , \wBMid1[20] , \wBIn76[7] , 
        \wAMid81[6] , \ScanLink182[31] , \ScanLink145[7] , \wRegInB89[2] , 
        \wRegInA113[14] , \ScanLink182[28] , \wRegInA104[1] , \wRegInA106[20] , 
        \ScanLink225[2] , \wBIn11[0] , \wAMid34[7] , \wAIn74[3] , 
        \wAMid113[11] , \wRegInA125[11] , \wBMid40[8] , \wAMid82[26] , 
        \wBMid104[5] , \wAMid97[12] , \wAMid125[14] , \wRegInB95[31] , 
        \wBIn98[15] , \ScanLink8[13] , \wAMid106[25] , \wRegInA41[9] , 
        \wRegInB95[28] , \wAIn120[7] , \ScanLink122[0] , \wAMid29[8] , 
        \wRegInA106[13] , \ScanLink242[5] , \ScanLink81[18] , 
        \ScanLink232[28] , \wRegInA125[22] , \ScanLink247[18] , 
        \ScanLink232[31] , \ScanLink211[19] , \ScanLink121[3] , \wBMid0[19] , 
        \wBMid0[7] , \wBMid1[13] , \wBIn12[3] , \wAIn123[4] , \wBMid3[4] , 
        \wBMid13[30] , \wBMid13[29] , \wBMid30[18] , \wBMid45[31] , 
        \wBMid66[19] , \ScanLink59[28] , \wRegInA113[27] , \wBIn16[24] , 
        \wAMid19[23] , \wBIn20[21] , \wAMid37[4] , \wBMid45[28] , 
        \ScanLink59[31] , \wBIn76[20] , \wBIn115[11] , \ScanLink241[6] , 
        \wAMid79[27] , \wBIn55[11] , \wAIn77[0] , \wBMid107[6] , \wAIn21[19] , 
        \wBIn35[15] , \wBIn40[25] , \wAIn54[29] , \wBIn123[14] , 
        \wRegInB38[31] , \wAIn54[30] , \wBIn63[14] , \wAIn77[18] , 
        \wBIn100[25] , \wRegInB38[28] , \wBIn19[8] , \wAMid21[0] , \wAIn61[4] , 
        \wBMid111[2] , \wRegInA119[12] , \wRegInA86[8] , \wRegInA49[1] , 
        \wBMid79[18] , \ScanLink33[19] , \ScanLink10[31] , \wRegInB127[3] , 
        \ScanLink46[29] , \wRegInB29[4] , \ScanLink10[28] , \wAMid13[16] , 
        \ScanLink65[18] , \ScanLink46[30] , \wAMid22[3] , \wAMid25[13] , 
        \wAMid30[27] , \wBMid48[0] , \wAMid66[26] , \wBIn69[21] , \wBMid87[9] , 
        \wAMid45[17] , \ScanLink137[7] , \wRegInB71[28] , \wAMid50[23] , 
        \wRegInB27[30] , \wAIn62[7] , \wAIn68[19] , \wRegInB27[29] , 
        \wRegInB52[19] , \wRegInB71[31] , \wAMid73[12] , \wBIn87[14] , 
        \wAMid88[13] , \wBIn92[20] , \wBMid115[21] , \wRegInA98[4] , 
        \ScanLink134[4] , \ScanLink2[26] , \wAIn93[18] , \wRegInB37[8] , 
        \wBMid100[15] , \wAMid119[24] , \wBMid123[24] , \ScanLink254[1] , 
        \wRegInB0[27] , \wRegInB122[26] , \wBMid99[5] , \wBMid112[1] , 
        \wRegInB101[17] , \wAMid1[0] , \wAMid2[3] , \wAMid13[25] , 
        \wAMid25[20] , \wAMid50[10] , \wBMid82[19] , \wRegInA6[22] , 
        \wRegInB114[23] , \wRegInB124[0] , \ScanLink17[9] , \wBIn60[3] , 
        \wAMid66[15] , \wBIn69[12] , \wAMid73[21] , \wAMid97[2] , 
        \ScanLink153[3] , \wRegInA97[29] , \ScanLink233[6] , \wBIn3[18] , 
        \wAMid30[14] , \wAMid45[24] , \wRegInA97[30] , \wRegInA112[5] , 
        \wBMid32[8] , \wAMid45[4] , \ScanLink181[5] , \wAMid46[7] , 
        \wAIn100[30] , \wAIn123[18] , \wRegInB82[9] , \wRegInA119[21] , 
        \wAIn100[29] , \wRegInB114[10] , \ScanLink130[30] , \ScanLink113[18] , 
        \wRegInA6[11] , \ScanLink166[28] , \wBIn63[0] , \wBIn87[27] , 
        \wAMid88[20] , \wAMid94[1] , \wAMid104[9] , \wRegInB0[14] , 
        \ScanLink182[6] , \ScanLink166[31] , \ScanLink145[19] , 
        \ScanLink130[29] , \wRegInB101[24] , \wRegInB122[15] , \wBMid100[26] , 
        \wAMid119[17] , \wAMid119[6] , \wBIn126[8] , \wBMid123[17] , 
        \wRegInA33[9] , \ScanLink150[0] , \wRegInA19[18] , \wRegInA111[6] , 
        \wAIn16[16] , \wAIn35[27] , \wAIn40[17] , \wBIn92[13] , \wBMid115[12] , 
        \ScanLink2[15] , \wRegInA80[6] , \ScanLink230[5] , \wAIn63[26] , 
        \wRegInA89[11] , \wRegInB59[26] , \wAMid18[30] , \wAMid18[29] , 
        \wBMid53[1] , \wAIn76[12] , \wRegInB39[22] , \wAIn20[13] , 
        \wAIn55[23] , \wBMid72[27] , \wRegInA52[0] , \wRegInA124[28] , 
        \ScanLink210[13] , \ScanLink12[4] , \ScanLink131[9] , \wAMid1[21] , 
        \wAIn5[25] , \wBMid24[26] , \ScanLink233[22] , \ScanLink38[26] , 
        \ScanLink196[25] , \wBMid31[12] , \wBMid51[16] , \wBMid81[7] , 
        \wRegInA107[19] , \wRegInA124[31] , \ScanLink246[12] , \wBMid44[22] , 
        \wRegInB32[5] , \ScanLink226[16] , \ScanLink183[11] , 
        \ScanLink253[26] , \wBMid12[23] , \ScanLink58[22] , \ScanLink205[27] , 
        \wAMid1[12] , \wAIn5[16] , \wBMid6[9] , \wBIn8[14] , \wAMid39[2] , 
        \wBMid67[13] , \ScanLink118[14] , \wBMid82[4] , \wBMid109[0] , 
        \ScanLink95[26] , \wBMid50[2] , \wAIn79[6] , \wRegInA51[3] , 
        \wBMid89[26] , \wRegInB31[6] , \ScanLink178[10] , \ScanLink80[12] , 
        \wAIn64[9] , \wAIn98[27] , \wRegInA72[10] , \wRegInA24[11] , 
        \wRegInB81[16] , \wRegInA83[5] , \wRegInA31[25] , \wRegInA51[21] , 
        \wRegInB94[22] , \wRegInA44[15] , \ScanLink11[7] , \wBMid44[11] , 
        \wAMid96[18] , \wRegInA12[14] , \ScanLink9[19] , \wRegInA67[24] , 
        \ScanLink253[15] , \wBMid31[21] , \wBMid67[20] , \ScanLink226[25] , 
        \ScanLink183[22] , \wRegInA36[4] , \wBIn8[27] , \wBMid12[10] , 
        \wBIn123[5] , \ScanLink58[11] , \wAIn16[25] , \wAIn20[20] , 
        \wBMid24[15] , \wBMid51[25] , \wBMid72[14] , \ScanLink205[14] , 
        \wRegInB56[1] , \wRegInB99[8] , \ScanLink246[21] , \ScanLink210[20] , 
        \ScanLink38[15] , \ScanLink235[8] , \ScanLink233[11] , 
        \ScanLink196[16] , \wBMid37[5] , \wAIn76[21] , \wRegInB39[11] , 
        \wBIn21[18] , \wAIn35[14] , \wAIn55[10] , \wAMid101[4] , 
        \ScanLink148[2] , \wRegInA109[4] , \wAIn40[24] , \wBIn54[28] , 
        \wBIn114[31] , \ScanLink76[0] , \wRegInB59[15] , \wRegInB84[7] , 
        \wBMid29[9] , \wBMid34[6] , \wAMid40[9] , \wBIn54[31] , \wBIn114[28] , 
        \wRegInA89[22] , \ScanLink228[7] , \wAIn63[15] , \wBIn77[19] , 
        \wBIn78[1] , \wAMid102[7] , \wRegInA28[8] , \wRegInA31[16] , 
        \wRegInA44[26] , \wRegInB94[11] , \ScanLink184[8] , \wRegInA67[17] , 
        \wRegInA12[27] , \wAIn98[14] , \wRegInA72[23] , \wRegInB87[4] , 
        \wAMid112[31] , \wAMid112[28] , \wRegInA24[22] , \wRegInA51[12] , 
        \ScanLink75[3] , \wRegInB81[25] , \wBIn120[6] , \wRegInA35[7] , 
        \ScanLink199[7] , \ScanLink178[23] , \ScanLink80[21] , \wRegInB55[2] , 
        \wBMid10[0] , \wAIn89[11] , \wBMid89[15] , \wRegInA117[8] , 
        \ScanLink118[27] , \ScanLink95[15] , \wRegInA16[16] , \wRegInA35[27] , 
        \wRegInB90[20] , \wRegInA40[17] , \ScanLink51[5] , \wRegInA63[26] , 
        \wRegInA76[12] , \wBMid35[10] , \wAIn39[4] , \wAMid79[0] , 
        \wBIn88[30] , \wBIn88[29] , \wAMid116[19] , \wAMid126[1] , 
        \wRegInA20[13] , \wRegInB85[14] , \wRegInA55[23] , \wBMid98[10] , 
        \wRegInB71[4] , \ScanLink109[22] , \ScanLink83[3] , \ScanLink84[10] , 
        \wBIn104[0] , \wRegInA1[4] , \ScanLink169[26] , \ScanLink91[24] , 
        \wRegInA11[1] , \wBIn41[8] , \wRegInB72[7] , \ScanLink172[8] , 
        \wBMid40[20] , \ScanLink222[14] , \ScanLink187[13] , \wAIn1[14] , 
        \wBMid4[31] , \wBMid4[28] , \wAMid5[23] , \wBMid16[21] , 
        \ScanLink201[25] , \wAIn12[27] , \wAIn12[14] , \wBMid13[3] , 
        \wBMid20[24] , \wBMid63[11] , \ScanLink29[10] , \wBMid76[25] , 
        \wBIn107[3] , \ScanLink214[11] , \ScanLink80[0] , \wRegInA12[2] , 
        \ScanLink49[14] , \wRegInA2[7] , \ScanLink237[20] , \ScanLink192[27] , 
        \wAIn24[11] , \wAIn51[21] , \wBMid55[14] , \ScanLink242[10] , 
        \wAIn72[10] , \wRegInB48[10] , \wRegInA98[27] , \wBIn25[30] , 
        \wBIn25[29] , \wAIn27[8] , \wAMid125[2] , \ScanLink52[6] , 
        \wAIn44[15] , \wBIn73[31] , \wBIn50[19] , \wAIn31[25] , \wAIn67[24] , 
        \wBIn73[28] , \wBIn110[19] , \wRegInB28[14] , \wAIn31[16] , 
        \wBIn38[3] , \wAIn92[9] , \wRegInB15[0] , \wRegInA75[5] , 
        \ScanLink169[15] , \ScanLink91[17] , \wAMid92[30] , \wBMid98[23] , 
        \wRegInA20[20] , \wRegInA55[10] , \wRegInA76[21] , \ScanLink109[11] , 
        \ScanLink84[23] , \wRegInB106[8] , \ScanLink35[1] , \wRegInB85[27] , 
        \wAIn109[4] , \wRegInA35[14] , \wRegInA40[24] , \wRegInB90[13] , 
        \wBMid74[4] , \wAIn89[22] , \wAMid92[29] , \wRegInA63[15] , 
        \wRegInA16[25] , \wAIn44[26] , \ScanLink36[2] , \wAIn24[22] , 
        \wAIn67[17] , \wRegInB28[27] , \wAMid69[28] , \wRegInB48[23] , 
        \wAIn72[23] , \wBMid77[7] , \wRegInA98[14] , \wAIn51[12] , 
        \wAMid69[31] , \ScanLink108[0] , \wBMid55[27] , \wBMid76[16] , 
        \wRegInA103[31] , \ScanLink214[22] , \wRegInA120[19] , 
        \ScanLink49[27] , \ScanLink242[23] , \wRegInB16[3] , \wRegInB118[4] , 
        \wBMid20[17] , \wRegInA103[28] , \ScanLink237[13] , \ScanLink192[14] , 
        \wBMid40[13] , \wAIn5[3] , \wAMid5[10] , \wBMid35[23] , \wBMid63[22] , 
        \wRegInA76[6] , \ScanLink222[27] , \ScanLink187[20] , \ScanLink29[23] , 
        \wBIn7[30] , \wBIn7[29] , \wBMid16[12] , \wAIn117[8] , 
        \ScanLink201[16] , \ScanLink162[19] , \ScanLink141[31] , 
        \wRegInA2[20] , \wRegInB110[21] , \ScanLink117[29] , \ScanLink141[28] , 
        \wAIn22[5] , \ScanLink134[18] , \ScanLink117[30] , \ScanLink98[2] , 
        \wAMid62[1] , \wBIn95[0] , \wRegInB4[25] , \wRegInB126[24] , 
        \ScanLink169[9] , \wRegInB105[15] , \wAIn6[0] , \wAMid17[14] , 
        \wBIn18[13] , \wAMid21[11] , \wBIn47[6] , \wBIn83[16] , \wBMid104[17] , 
        \ScanLink214[3] , \wBIn96[22] , \wAMid108[12] , \ScanLink174[6] , 
        \wAMid99[25] , \wBMid111[23] , \wRegInA68[19] , \ScanLink6[24] , 
        \wAMid54[21] , \ScanLink49[7] , \wAMid77[10] , \wRegInB74[9] , 
        \ScanLink217[0] , \wBIn78[17] , \wRegInA4[9] , \wAMid34[25] , 
        \wAMid62[24] , \wRegInA93[18] , \wAMid41[15] , \ScanLink177[5] , 
        \wBIn44[5] , \wAMid61[2] , \wRegInB69[6] , \ScanLink54[8] , 
        \wRegInA108[24] , \ScanLink199[18] , \wAIn127[29] , \wAIn21[6] , 
        \wBIn23[2] , \wBIn83[25] , \wBIn96[11] , \wBIn96[3] , \wAIn104[18] , 
        \wAIn127[30] , \wAMid108[21] , \wAMid99[16] , \wBMid111[10] , 
        \wBMid104[24] , \ScanLink6[17] , \wAIn94[7] , \wAIn97[29] , 
        \wAIn97[30] , \wAIn112[5] , \ScanLink110[2] , \wAIn46[1] , 
        \wBMid86[31] , \wRegInB4[16] , \wRegInB100[6] , \wRegInB126[17] , 
        \wRegInB105[26] , \wRegInB110[12] , \wRegInA2[13] , \wBMid86[28] , 
        \wAIn89[8] , \wRegInB103[5] , \ScanLink229[18] , \wAIn0[25] , 
        \wAIn0[6] , \wBMid0[22] , \wAMid1[8] , \wBIn3[10] , \wAMid17[27] , 
        \wBIn18[20] , \wAIn45[2] , \ScanLink61[30] , \wAMid62[17] , 
        \wBMid71[9] , \wRegInA108[17] , \ScanLink61[29] , \ScanLink42[18] , 
        \ScanLink37[28] , \ScanLink37[31] , \ScanLink14[19] , \wAMid18[9] , 
        \wBIn20[1] , \wAMid34[16] , \wAMid41[26] , \wAMid54[12] , \wAIn97[4] , 
        \wRegInA70[8] , \wAIn111[6] , \wRegInB56[31] , \wRegInB75[19] , 
        \wAMid21[22] , \wRegInB23[18] , \ScanLink113[1] , \wAIn19[18] , 
        \wAMid77[23] , \wBIn78[24] , \wRegInB56[28] , \wBMid82[22] , 
        \wAMid89[6] , \wAMid104[1] , \ScanLink130[21] , \wRegInA6[19] , 
        \ScanLink145[11] , \wRegInB114[18] , \ScanLink113[10] , \wBMid32[0] , 
        \wBIn63[8] , \wBMid97[16] , \wRegInB81[2] , \ScanLink166[20] , 
        \ScanLink106[24] , \ScanLink173[14] , \ScanLink125[15] , \wBIn126[0] , 
        \wRegInA33[1] , \ScanLink150[25] , \ScanLink73[5] , \wAIn86[17] , 
        \wAMid88[31] , \wAMid88[28] , \wAIn93[23] , \wAMid94[9] , 
        \ScanLink150[8] , \wRegInA19[10] , \wRegInA79[14] , \wRegInB53[4] , 
        \wBIn3[23] , \wBIn9[4] , \wAIn18[7] , \wAMid25[31] , \wAMid58[3] , 
        \wAIn68[22] , \wAMid73[29] , \wRegInB27[12] , \wRegInA82[15] , 
        \wAMid50[18] , \wRegInB52[22] , \wBMid19[27] , \wAMid25[28] , 
        \wAMid73[30] , \wBIn125[3] , \wRegInA30[2] , \wBMid31[3] , 
        \wRegInB11[17] , \wRegInB71[13] , \wRegInB32[26] , \wRegInB50[7] , 
        \wRegInB64[27] , \wRegInA97[21] , \wRegInB47[16] , \ScanLink238[26] , 
        \ScanLink65[23] , \ScanLink10[13] , \wBMid79[23] , \wAMid107[2] , 
        \ScanLink46[12] , \ScanLink33[22] , \wAIn115[15] , \wBMid56[4] , 
        \wBMid84[2] , \wAIn86[24] , \wAIn100[21] , \wRegInA119[30] , 
        \ScanLink70[6] , \ScanLink53[26] , \wAIn123[10] , \wRegInB82[1] , 
        \ScanLink188[15] , \ScanLink26[16] , \ScanLink70[17] , 
        \wRegInA119[29] , \wBIn92[28] , \wBMid115[29] , \wBIn92[31] , 
        \wBMid115[30] , \wRegInA19[23] , \wRegInA57[5] , \wAIn93[10] , 
        \wRegInB37[0] , \wRegInA79[27] , \ScanLink254[9] , \ScanLink173[27] , 
        \ScanLink106[17] , \wBMid112[9] , \wRegInA85[3] , \ScanLink150[16] , 
        \ScanLink129[3] , \ScanLink125[26] , \wBMid82[11] , \wBMid97[25] , 
        \ScanLink145[22] , \wRegInB124[8] , \ScanLink130[12] , \ScanLink17[1] , 
        \wAMid4[5] , \wAMid7[6] , \wBIn19[0] , \wAIn100[12] , \wRegInA49[9] , 
        \ScanLink249[6] , \ScanLink166[13] , \ScanLink113[23] , \wRegInA86[0] , 
        \ScanLink26[25] , \wBMid19[14] , \wAMid21[8] , \wAIn123[23] , 
        \ScanLink53[15] , \wBMid29[1] , \wAMid40[1] , \wBMid48[8] , 
        \wBMid55[7] , \wBIn69[30] , \wBMid79[10] , \ScanLink238[15] , 
        \ScanLink188[26] , \ScanLink70[24] , \ScanLink65[10] , 
        \ScanLink10[20] , \ScanLink33[11] , \wAIn115[26] , \wRegInB11[24] , 
        \wRegInA54[6] , \ScanLink46[21] , \ScanLink14[2] , \wRegInB64[14] , 
        \wRegInB47[25] , \wAIn68[11] , \wBIn69[29] , \wBMid87[1] , 
        \wRegInB32[15] , \wRegInA97[12] , \wRegInB34[3] , \wRegInB52[11] , 
        \wRegInB27[21] , \wRegInB71[20] , \wRegInA82[26] , \wBIn78[9] , 
        \wAMid96[23] , \wBIn99[24] , \wRegInB8[5] , \ScanLink9[22] , 
        \wAMid124[25] , \wRegInA28[0] , \wAMid83[17] , \wAMid107[14] , 
        \wRegInB94[19] , \ScanLink184[0] , \wAMid112[20] , \wAMid92[7] , 
        \wRegInB48[5] , \ScanLink80[29] , \wBIn65[6] , \ScanLink80[30] , 
        \wRegInA117[0] , \ScanLink156[6] , \ScanLink236[3] , \ScanLink68[4] , 
        \wBMid12[18] , \wBMid67[28] , \ScanLink155[5] , \ScanLink58[19] , 
        \wBMid31[30] , \wBMid31[29] , \wBMid44[19] , \wBIn66[5] , \wAMid91[4] , 
        \wBMid67[31] , \wRegInA112[16] , \wRegInB56[9] , \wRegInB99[0] , 
        \ScanLink246[29] , \wRegInA107[22] , \ScanLink235[0] , 
        \ScanLink210[31] , \ScanLink233[19] , \wBMid0[11] , \wBMid5[2] , 
        \wBMid6[1] , \wBIn17[15] , \wAIn20[28] , \wRegInA114[3] , 
        \wRegInA124[13] , \ScanLink246[30] , \ScanLink210[28] , \wBIn34[24] , 
        \wBIn41[14] , \wBIn122[25] , \wAIn55[18] , \wAIn76[30] , 
        \ScanLink187[3] , \wAMid18[12] , \wAIn20[31] , \wBIn21[10] , 
        \wAMid43[2] , \wBIn62[25] , \wAIn76[29] , \wBIn101[14] , 
        \wRegInB39[19] , \wBIn77[11] , \wAMid78[16] , \wBIn114[20] , 
        \wAMid24[5] , \wBIn54[20] , \wAIn64[1] , \wBMid109[8] , 
        \ScanLink132[2] , \ScanLink76[8] , \wAMid112[13] , \ScanLink252[7] , 
        \ScanLink178[18] , \wRegInA24[19] , \wRegInA51[29] , \wAMid83[24] , 
        \wBMid114[7] , \wRegInA51[30] , \wAMid124[16] , \wRegInA72[18] , 
        \wRegInB122[6] , \wBIn21[23] , \wAMid27[6] , \wAMid96[10] , 
        \wBIn99[17] , \ScanLink9[11] , \wAMid107[27] , \wBIn54[13] , 
        \wBMid53[9] , \wBIn77[22] , \wAMid78[25] , \wBIn114[13] , 
        \wBMid117[4] , \wRegInA89[19] , \wAIn67[2] , \wBIn34[17] , 
        \wBIn41[27] , \wBIn122[16] , \wBIn101[27] , \wBIn17[26] , \wBIn62[16] , 
        \wRegInB121[5] , \wAMid18[21] , \wRegInA52[8] , \wRegInA107[11] , 
        \wRegInA124[20] , \wAMid1[30] , \wAMid1[29] , \ScanLink131[1] , 
        \wRegInA112[25] , \ScanLink183[19] , \ScanLink251[4] , \wBMid4[20] , 
        \wBIn13[17] , \wBIn25[12] , \wBIn73[13] , \wRegInB105[3] , 
        \wBIn110[22] , \wBIn30[26] , \wAIn43[4] , \wBIn50[22] , \wBIn45[16] , 
        \wBIn126[27] , \ScanLink108[8] , \wBIn66[27] , \wBIn105[16] , 
        \wAMid69[20] , \wRegInA103[20] , \wBMid4[13] , \wAMid5[18] , 
        \wRegInA120[11] , \wBMid16[30] , \wBMid16[29] , \wBIn25[4] , 
        \wBIn26[7] , \wAIn91[2] , \wAIn117[0] , \ScanLink187[31] , 
        \ScanLink115[7] , \wBMid69[3] , \wRegInA9[24] , \wRegInB15[8] , 
        \wRegInA116[14] , \ScanLink187[28] , \ScanLink28[6] , \wAIn92[1] , 
        \ScanLink109[19] , \wAIn114[3] , \wAIn40[7] , \wAMid87[15] , 
        \wAMid116[22] , \wRegInA55[18] , \wRegInA76[30] , \ScanLink116[4] , 
        \wRegInA20[28] , \ScanLink35[9] , \wBIn88[12] , \wAMid92[21] , 
        \wRegInA20[31] , \wRegInA76[29] , \wRegInB106[0] , \wAMid120[27] , 
        \wRegInA68[2] , \wAMid103[16] , \wBMid35[18] , \wBMid40[31] , 
        \wBMid63[19] , \ScanLink80[8] , \ScanLink29[18] , \wRegInA116[27] , 
        \wBMid40[28] , \ScanLink211[6] , \wBIn42[3] , \wRegInA103[13] , 
        \wRegInA120[22] , \ScanLink242[18] , \ScanLink237[28] , 
        \ScanLink237[31] , \ScanLink214[19] , \wBIn13[24] , \wAIn24[19] , 
        \wBIn30[15] , \wBIn45[25] , \wAIn51[29] , \wBIn126[14] , 
        \ScanLink171[3] , \wAIn51[30] , \wBIn66[14] , \wBIn105[25] , 
        \wAMid69[13] , \wAIn72[18] , \wRegInB48[18] , \wAMid67[4] , 
        \wBIn73[20] , \wBIn110[11] , \wAIn3[5] , \wAIn24[3] , \wBIn25[21] , 
        \wAIn27[0] , \wBIn50[11] , \wAIn89[19] , \wBIn90[5] , \wAMid92[12] , 
        \wAMid120[14] , \wRegInB90[31] , \wAMid103[25] , \wRegInB90[28] , 
        \wAMid116[11] , \wAMid64[7] , \wBIn93[6] , \wBIn119[7] , \wAMid126[9] , 
        \wAMid87[26] , \wAIn6[8] , \wBIn7[12] , \wBMid10[8] , \wBIn88[21] , 
        \wBIn18[31] , \wBIn41[0] , \wBMid98[18] , \ScanLink212[5] , 
        \ScanLink84[18] , \wBIn104[8] , \wRegInA11[9] , \ScanLink172[0] , 
        \wBMid68[15] , \wAMid79[8] , \wRegInA9[17] , \wAIn104[23] , 
        \ScanLink57[24] , \ScanLink30[4] , \wBMid71[1] , \wAIn127[12] , 
        \ScanLink229[10] , \ScanLink22[14] , \ScanLink74[15] , 
        \ScanLink199[23] , \ScanLink61[21] , \ScanLink14[11] , \wAIn111[17] , 
        \ScanLink249[14] , \ScanLink42[10] , \ScanLink37[20] , \wRegInB15[15] , 
        \wRegInB60[25] , \wBIn18[28] , \wAIn79[14] , \wRegInB10[5] , 
        \wRegInB36[24] , \wRegInA93[23] , \wRegInB43[14] , \wAMid18[1] , 
        \wAIn19[10] , \wRegInB23[10] , \wRegInA86[17] , \wBIn20[9] , 
        \wAIn58[5] , \wRegInB56[20] , \wRegInA70[0] , \ScanLink113[9] , 
        \wAIn46[9] , \wAIn82[15] , \wBIn96[19] , \wAMid108[30] , 
        \wRegInB13[6] , \wRegInB75[11] , \wRegInA68[22] , \wBMid111[18] , 
        \wBMid86[20] , \wAIn89[0] , \wBMid93[14] , \wAIn97[21] , 
        \wAMid108[29] , \wRegInA73[3] , \ScanLink177[16] , \ScanLink102[26] , 
        \ScanLink121[17] , \ScanLink154[27] , \ScanLink33[7] , 
        \ScanLink134[23] , \ScanLink141[13] , \ScanLink117[12] , \wBMid15[5] , 
        \wAIn19[23] , \wBMid72[2] , \ScanLink162[22] , \wAMid21[19] , 
        \wAMid54[30] , \wAMid77[18] , \wRegInB56[13] , \ScanLink8[3] , 
        \wRegInB74[1] , \ScanLink217[8] , \wRegInB23[23] , \wRegInA86[24] , 
        \wAMid54[29] , \wRegInB75[22] , \wBIn59[2] , \wBMid68[26] , 
        \wAIn79[27] , \wBIn101[5] , \ScanLink86[6] , \wRegInA4[1] , 
        \wRegInA14[4] , \wRegInB60[16] , \wRegInB15[26] , \wRegInB43[27] , 
        \wRegInB36[17] , \wRegInA93[10] , \wAIn104[10] , \wAIn111[24] , 
        \ScanLink249[27] , \ScanLink14[22] , \ScanLink199[10] , 
        \ScanLink61[12] , \ScanLink37[13] , \ScanLink54[0] , \ScanLink42[23] , 
        \wAMid123[4] , \ScanLink22[27] , \wAIn127[21] , \ScanLink57[17] , 
        \ScanLink229[23] , \wBIn7[21] , \wBMid86[13] , \ScanLink141[20] , 
        \ScanLink74[26] , \wRegInA2[31] , \ScanLink57[3] , \wRegInB110[30] , 
        \ScanLink134[10] , \wAIn13[16] , \wBMid16[6] , \wAMid62[9] , 
        \wRegInA2[28] , \ScanLink162[11] , \wRegInB110[29] , \ScanLink209[4] , 
        \ScanLink117[21] , \ScanLink177[25] , \ScanLink102[15] , \wAIn25[13] , 
        \wAIn29[6] , \wAMid69[2] , \wAIn82[26] , \wBMid93[27] , \wBIn95[8] , 
        \wAMid120[7] , \ScanLink169[1] , \ScanLink154[14] , \ScanLink121[24] , 
        \wAIn97[12] , \ScanLink85[5] , \wRegInA7[2] , \wRegInB77[2] , 
        \wRegInA68[11] , \wBIn88[7] , \wBIn102[6] , \wRegInA17[7] , 
        \wBMid99[12] , \wRegInB61[6] , \ScanLink93[1] , \ScanLink108[20] , 
        \ScanLink85[12] , \ScanLink168[24] , \ScanLink90[26] , \wAIn34[9] , 
        \wAIn88[13] , \wBIn114[2] , \wRegInA17[14] , \wRegInA34[25] , 
        \wRegInB91[22] , \wRegInA41[15] , \ScanLink41[7] , \wRegInA62[24] , 
        \wAMid93[18] , \wRegInA77[10] , \wAIn50[23] , \wAMid68[19] , 
        \wAIn73[12] , \wRegInA21[11] , \wRegInA54[21] , \wRegInB84[16] , 
        \wRegInA99[25] , \ScanLink3[8] , \wRegInB49[12] , \wAIn30[27] , 
        \wAIn45[17] , \ScanLink42[4] , \wAIn66[26] , \wRegInB29[16] , 
        \wBMid34[12] , \ScanLink223[16] , \ScanLink186[11] , \wRegInB62[5] , 
        \ScanLink256[26] , \wAIn0[16] , \wAMid4[21] , \wBMid17[23] , 
        \wBMid41[22] , \ScanLink200[27] , \ScanLink90[2] , \wBMid5[19] , 
        \wBMid62[13] , \wBMid77[27] , \wBIn117[1] , \wRegInA121[28] , 
        \ScanLink28[12] , \ScanLink215[13] , \ScanLink48[16] , \wAMid10[9] , 
        \wBMid21[26] , \wBIn52[9] , \ScanLink161[9] , \wBIn28[1] , 
        \wBMid54[16] , \wRegInA102[19] , \wRegInA121[31] , \ScanLink236[22] , 
        \ScanLink193[25] , \wBIn89[18] , \ScanLink243[12] , \wAMid117[31] , 
        \wRegInA77[23] , \wAMid117[28] , \wRegInA54[12] , \wAIn119[6] , 
        \wRegInA21[22] , \ScanLink25[3] , \wRegInA34[16] , \wRegInA41[26] , 
        \wRegInB84[25] , \wRegInA78[8] , \wRegInB91[11] , \wRegInA62[17] , 
        \wBMid21[15] , \wBMid54[25] , \wBMid64[6] , \wAIn88[20] , 
        \wRegInA17[27] , \wBMid77[14] , \wBMid79[9] , \wBMid99[21] , 
        \wAIn104[9] , \wRegInA65[7] , \ScanLink168[17] , \ScanLink90[15] , 
        \ScanLink108[13] , \ScanLink85[21] , \wRegInB108[6] , 
        \ScanLink215[20] , \ScanLink48[25] , \ScanLink243[21] , 
        \ScanLink256[15] , \ScanLink236[11] , \ScanLink193[16] , \wBIn2[30] , 
        \wBIn2[29] , \wAMid4[12] , \wBMid34[21] , \wBMid41[11] , 
        \ScanLink223[25] , \ScanLink186[22] , \wBMid62[20] , \wAIn81[8] , 
        \wRegInA66[4] , \ScanLink28[21] , \wBIn6[18] , \wAIn13[25] , 
        \wBMid17[10] , \ScanLink200[14] , \wBIn24[18] , \wAIn30[14] , 
        \wAIn45[24] , \wBIn51[28] , \ScanLink26[0] , \wBIn111[31] , 
        \wRegInB115[9] , \wAMid16[16] , \wAIn18[30] , \wAIn25[20] , 
        \wBIn51[31] , \wAIn66[15] , \wBMid67[5] , \wBIn72[19] , \wBIn111[28] , 
        \wRegInB29[25] , \wRegInB49[21] , \wRegInA99[16] , \wAIn73[21] , 
        \wBMid123[8] , \wAIn31[4] , \wAIn32[7] , \wAIn50[10] , 
        \ScanLink118[2] , \wBIn57[4] , \wBIn82[14] , \wAIn96[18] , 
        \wRegInB67[8] , \wBMid105[15] , \wBMid126[24] , \ScanLink204[1] , 
        \wRegInA125[2] , \ScanLink164[4] , \wBMid87[19] , \wBIn97[20] , 
        \wAMid98[27] , \wAMid109[10] , \ScanLink7[26] , \wBMid110[21] , 
        \wRegInA3[22] , \ScanLink6[5] , \wRegInB111[23] , \ScanLink47[9] , 
        \ScanLink88[0] , \wAMid71[0] , \wAMid72[3] , \wBIn85[2] , 
        \wRegInB127[26] , \wRegInB5[27] , \wRegInB79[4] , \wRegInB104[17] , 
        \ScanLink43[29] , \ScanLink36[19] , \ScanLink15[31] , \ScanLink15[28] , 
        \wRegInA109[26] , \ScanLink5[6] , \ScanLink60[18] , \ScanLink43[30] , 
        \wRegInA9[4] , \wRegInA19[1] , \ScanLink228[29] , \wBIn49[8] , 
        \ScanLink228[30] , \wBIn86[1] , \wAIn18[29] , \wAMid20[13] , 
        \wAMid55[23] , \wRegInB74[28] , \wRegInA126[1] , \wRegInB22[30] , 
        \ScanLink59[5] , \wAMid76[12] , \wBIn79[15] , \wRegInB57[19] , 
        \wRegInB74[31] , \ScanLink207[2] , \wRegInB22[29] , \wAMid16[7] , 
        \wBIn19[11] , \wBMid18[0] , \wAMid35[27] , \wAMid63[26] , 
        \wAMid40[17] , \wBIn54[7] , \ScanLink167[7] , \wRegInB127[15] , 
        \wRegInB5[14] , \wRegInB104[24] , \wRegInB110[4] , \wBMid62[8] , 
        \wBMid126[5] , \wRegInA3[11] , \wRegInB111[10] , \ScanLink135[30] , 
        \ScanLink116[18] , \wBIn7[2] , \wAMid12[14] , \wAMid15[4] , 
        \wAMid16[25] , \wBIn33[0] , \wAIn56[3] , \ScanLink163[28] , 
        \wBIn82[27] , \wBIn97[13] , \wAMid98[14] , \wAMid109[23] , 
        \ScanLink163[31] , \ScanLink140[19] , \ScanLink135[29] , 
        \wRegInA69[31] , \wRegInA69[28] , \ScanLink7[15] , \wBMid110[12] , 
        \wAIn84[5] , \wBMid105[26] , \wRegInA63[9] , \wAIn102[7] , 
        \wBMid126[17] , \wAMid63[15] , \wRegInA92[29] , \ScanLink100[0] , 
        \wBIn19[22] , \wAMid20[20] , \wAMid35[14] , \wAMid40[24] , 
        \wRegInA92[30] , \wAMid55[10] , \wAIn87[6] , \wBIn30[3] , \wAIn101[4] , 
        \ScanLink103[3] , \wAIn55[0] , \wAMid76[21] , \wBIn79[26] , 
        \wAIn105[30] , \wAIn126[18] , \wRegInB113[7] , \wAIn105[29] , 
        \wRegInA109[15] , \ScanLink198[30] , \wBMid125[6] , \ScanLink198[29] , 
        \wBIn14[5] , \wAMid31[25] , \wBMid58[2] , \wRegInA96[18] , 
        \wAMid67[24] , \wBIn68[23] , \wAMid44[15] , \wAIn125[2] , 
        \ScanLink127[5] , \wAMid24[11] , \wAMid31[2] , \wAMid51[21] , 
        \wAMid72[10] , \wRegInB24[9] , \ScanLink19[7] , \ScanLink247[0] , 
        \wAMid32[1] , \wAIn71[6] , \wAIn101[18] , \wBMid101[0] , \wAIn122[29] , 
        \wRegInA118[10] , \wAIn122[30] , \wRegInA59[3] , \wAIn72[5] , 
        \wRegInB39[6] , \wRegInA95[9] , \wRegInB1[25] , \wRegInB123[24] , 
        \ScanLink139[9] , \wBMid89[7] , \wRegInB100[15] , \wBMid102[3] , 
        \wRegInA7[20] , \ScanLink167[19] , \ScanLink144[31] , \wRegInB115[21] , 
        \ScanLink112[29] , \wBIn4[1] , \wRegInA18[30] , \wRegInA88[6] , 
        \ScanLink144[28] , \ScanLink131[18] , \ScanLink112[30] , 
        \ScanLink124[6] , \wAIn15[2] , \wBIn17[6] , \wBIn86[16] , \wBIn93[22] , 
        \wAIn126[1] , \wBMid94[8] , \wBMid114[23] , \wRegInA18[29] , 
        \ScanLink3[24] , \wBMid101[17] , \wAMid89[11] , \wAMid117[8] , 
        \wAMid118[26] , \wBMid122[26] , \ScanLink244[3] , \ScanLink64[30] , 
        \wBMid21[9] , \wAMid55[6] , \wBMid78[29] , \ScanLink47[18] , 
        \ScanLink191[7] , \ScanLink32[28] , \ScanLink64[29] , \wBMid78[30] , 
        \ScanLink32[31] , \ScanLink11[19] , \wRegInA118[23] , \wAMid24[22] , 
        \wAMid51[12] , \wAIn69[31] , \wRegInA20[8] , \wBIn70[1] , 
        \wRegInB70[19] , \ScanLink143[1] , \wAMid72[23] , \wRegInB53[31] , 
        \wAMid87[0] , \wAMid12[27] , \wAMid48[9] , \wAIn69[28] , 
        \wRegInB26[18] , \wAMid67[17] , \wRegInB53[28] , \wBIn68[10] , 
        \wAMid31[16] , \wAMid44[26] , \wRegInA102[7] , \ScanLink223[4] , 
        \wAMid56[5] , \wBIn73[2] , \wAMid84[3] , \wBIn86[25] , \wBMid101[24] , 
        \wAMid89[22] , \wAIn92[30] , \wAIn92[29] , \wAMid109[4] , 
        \wAMid118[15] , \wBIn93[11] , \wBMid122[15] , \wRegInA101[4] , 
        \ScanLink140[2] , \ScanLink220[7] , \wBMid114[10] , \ScanLink3[17] , 
        \wBMid83[31] , \wRegInA7[13] , \wRegInB115[12] , \wAMid0[23] , 
        \wAIn4[27] , \wBMid8[7] , \wAIn16[1] , \wBMid83[28] , \wBMid25[24] , 
        \wBMid73[25] , \wRegInB1[16] , \wRegInB123[17] , \ScanLink192[4] , 
        \wRegInA42[2] , \wRegInB91[8] , \wRegInB100[26] , \ScanLink211[11] , 
        \ScanLink39[24] , \wBMid50[14] , \ScanLink232[20] , \ScanLink197[27] , 
        \wBMid91[5] , \ScanLink247[10] , \ScanLink227[14] , \ScanLink182[13] , 
        \wBMid30[10] , \wRegInB22[7] , \wBMid13[21] , \wBMid45[20] , 
        \ScanLink252[24] , \ScanLink204[25] , \ScanLink59[20] , \wAMid0[19] , 
        \wAMid0[10] , \wAIn4[14] , \wBIn9[16] , \wAIn17[14] , \wBIn20[30] , 
        \wBIn20[29] , \wAIn41[15] , \wBMid66[11] , \wBIn76[31] , \wBIn55[19] , 
        \wAIn77[8] , \wRegInA90[4] , \wAIn34[25] , \wAIn62[24] , \wBIn76[28] , 
        \wBIn115[19] , \wRegInA88[13] , \wBMid43[3] , \wAIn21[11] , 
        \wAIn54[21] , \wAIn77[10] , \wRegInB38[20] , \wRegInB58[24] , 
        \wAMid29[0] , \wBMid40[0] , \wAIn99[25] , \wRegInA73[12] , 
        \wAMid113[19] , \wRegInA93[7] , \wRegInA13[16] , \wRegInA25[13] , 
        \wRegInA30[27] , \wRegInA50[23] , \wRegInB80[14] , \wRegInB95[20] , 
        \wRegInA45[17] , \wRegInA66[26] , \ScanLink119[16] , \wBMid92[6] , 
        \ScanLink94[24] , \wAMid9[0] , \wBIn11[8] , \wAIn69[4] , \wBMid88[24] , 
        \wBMid119[2] , \wRegInA41[1] , \ScanLink122[8] , \wAIn17[27] , 
        \wAMid19[18] , \wAMid53[8] , \wRegInB21[4] , \ScanLink179[12] , 
        \ScanLink81[10] , \wAIn21[22] , \wBMid27[7] , \wAIn77[23] , 
        \wRegInB38[13] , \wAMid111[6] , \wAIn34[16] , \wAIn54[12] , 
        \ScanLink158[0] , \ScanLink197[9] , \wAIn41[26] , \wRegInA119[6] , 
        \ScanLink66[2] , \wRegInB58[17] , \wRegInB94[5] , \wAIn62[17] , 
        \wRegInA88[20] , \ScanLink238[5] , \wBMid30[23] , \wBMid45[13] , 
        \wRegInB6[3] , \ScanLink252[17] , \ScanLink227[27] , \ScanLink182[20] , 
        \wBMid66[22] , \wRegInA26[6] , \wBMid1[31] , \wBMid1[28] , 
        \wBMid13[12] , \ScanLink204[16] , \wRegInA104[9] , \ScanLink59[13] , 
        \ScanLink39[17] , \wBMid50[27] , \wBMid73[16] , \wRegInA106[31] , 
        \wRegInA125[19] , \ScanLink211[22] , \wRegInB46[3] , \wBMid1[21] , 
        \wAMid4[31] , \wBIn6[22] , \wBIn6[11] , \wBIn9[25] , \wBMid25[17] , 
        \wRegInA106[28] , \ScanLink247[23] , \wRegInB5[0] , \wRegInA25[5] , 
        \ScanLink232[13] , \ScanLink197[14] , \ScanLink189[5] , 
        \ScanLink179[21] , \ScanLink81[23] , \wBMid24[4] , \wBIn68[3] , 
        \wBMid88[17] , \wRegInB45[0] , \ScanLink94[17] , \ScanLink226[9] , 
        \ScanLink119[25] , \wAMid97[30] , \wRegInA45[24] , \wAMid112[5] , 
        \ScanLink8[31] , \wRegInA30[14] , \wRegInB95[13] , \wAMid97[29] , 
        \wRegInA66[15] , \ScanLink8[28] , \wAIn99[16] , \wRegInA13[25] , 
        \wRegInA3[18] , \wRegInA25[20] , \wRegInA50[10] , \wRegInA73[21] , 
        \wRegInB97[6] , \ScanLink65[1] , \wRegInB80[27] , \wRegInB111[19] , 
        \ScanLink116[11] , \wAIn8[7] , \wAIn18[13] , \wAMid20[30] , 
        \wAMid20[29] , \wBIn33[9] , \wBMid62[1] , \wBMid87[23] , \wAIn99[3] , 
        \ScanLink163[21] , \wBMid92[17] , \ScanLink140[10] , \ScanLink135[20] , 
        \ScanLink120[14] , \wAIn96[22] , \ScanLink176[15] , \ScanLink155[24] , 
        \ScanLink103[25] , \ScanLink23[4] , \wRegInA63[0] , \wAIn48[6] , 
        \wAMid55[19] , \wAIn83[16] , \wRegInA69[21] , \ScanLink100[9] , 
        \wAMid76[31] , \wRegInA60[3] , \wAMid76[28] , \wRegInB74[12] , 
        \wRegInB22[13] , \wRegInA87[14] , \wAIn55[9] , \wAIn78[17] , 
        \wRegInB37[27] , \wRegInB57[23] , \wRegInA92[20] , \wRegInB14[16] , 
        \wRegInB42[17] , \wRegInB61[26] , \wBMid61[2] , \wAIn110[14] , 
        \ScanLink43[13] , \ScanLink36[23] , \ScanLink198[20] , 
        \ScanLink60[22] , \ScanLink15[12] , \wBMid69[16] , \wAIn105[20] , 
        \wAIn126[11] , \ScanLink248[17] , \ScanLink228[13] , \ScanLink75[16] , 
        \ScanLink56[27] , \ScanLink20[7] , \wAIn83[25] , \wBIn97[30] , 
        \wBIn112[5] , \ScanLink23[17] , \wBIn98[4] , \wBMid110[31] , 
        \wAMid109[19] , \wRegInA69[12] , \wBIn97[29] , \wBMid110[28] , 
        \wBMid92[24] , \wAIn96[11] , \wRegInB67[1] , \ScanLink204[8] , 
        \ScanLink179[2] , \ScanLink155[17] , \ScanLink95[6] , 
        \ScanLink120[27] , \ScanLink176[26] , \ScanLink103[16] , \wBMid5[23] , 
        \wAMid10[0] , \wAIn18[20] , \wBIn19[18] , \wBIn49[1] , \wBMid69[25] , 
        \wAMid71[9] , \wBMid87[10] , \ScanLink219[7] , \ScanLink163[12] , 
        \ScanLink140[23] , \ScanLink116[22] , \ScanLink135[13] , 
        \ScanLink88[9] , \ScanLink47[0] , \wAIn105[13] , \wAIn126[22] , 
        \wRegInA19[8] , \ScanLink228[20] , \ScanLink75[25] , \ScanLink23[24] , 
        \wBIn86[8] , \ScanLink56[14] , \wAIn110[27] , \ScanLink36[10] , 
        \wRegInB42[24] , \ScanLink248[24] , \ScanLink44[3] , \ScanLink43[20] , 
        \ScanLink15[21] , \ScanLink198[13] , \ScanLink60[11] , \wBMid18[9] , 
        \wRegInB37[14] , \wRegInA92[13] , \wAIn78[24] , \wBIn111[6] , 
        \wRegInB14[25] , \wRegInB61[15] , \wRegInB74[21] , \wRegInA126[8] , 
        \ScanLink96[5] , \wBIn28[8] , \wAIn50[4] , \wAIn88[30] , 
        \wRegInB22[20] , \wRegInB57[10] , \wRegInB64[2] , \wRegInA87[27] , 
        \wRegInA78[1] , \wAMid102[15] , \wRegInB91[18] , \wBMid17[19] , 
        \wBIn35[7] , \wAIn82[2] , \wAMid86[16] , \wAIn88[29] , \wAMid93[22] , 
        \wBMid120[2] , \wAMid121[24] , \wBIn89[11] , \wAMid117[21] , 
        \wRegInB18[4] , \wRegInB116[3] , \wAIn104[0] , \ScanLink85[31] , 
        \wBMid34[28] , \wBMid41[18] , \wBMid79[0] , \wBMid99[28] , 
        \ScanLink106[7] , \ScanLink85[28] , \wBMid99[31] , \wRegInA8[27] , 
        \ScanLink38[5] , \wBMid62[30] , \ScanLink28[31] , \wRegInA117[17] , 
        \wBMid62[29] , \wAIn81[1] , \ScanLink28[28] , \ScanLink105[4] , 
        \wBMid34[31] , \wBIn36[4] , \wAIn107[3] , \wBMid5[10] , \wBIn12[27] , 
        \wBIn12[14] , \wAMid13[3] , \wRegInB49[28] , \wRegInA102[23] , 
        \wRegInA121[12] , \ScanLink243[31] , \ScanLink243[28] , 
        \ScanLink215[29] , \ScanLink236[18] , \ScanLink215[30] , \wAIn25[30] , 
        \wBIn24[22] , \wBIn24[11] , \wAIn25[29] , \wAIn53[7] , \wBIn67[24] , 
        \wAIn73[28] , \wBIn104[15] , \wBMid123[1] , \wAMid68[23] , 
        \wRegInB49[31] , \wBIn31[25] , \wBIn44[15] , \wAIn73[31] , 
        \wBIn127[24] , \wAIn50[19] , \wAIn34[0] , \wBIn51[21] , 
        \ScanLink26[9] , \wBIn51[3] , \wBIn72[10] , \wRegInB115[0] , 
        \wBIn111[21] , \wRegInA8[14] , \ScanLink162[3] , \wAMid74[4] , 
        \wRegInA123[5] , \ScanLink108[30] , \ScanLink202[6] , 
        \ScanLink108[29] , \ScanLink93[8] , \wAMid86[25] , \wBIn89[22] , 
        \wRegInA54[31] , \wRegInA77[19] , \wAIn37[3] , \wBIn51[12] , 
        \wBIn83[5] , \wBIn109[4] , \wAMid117[12] , \wRegInA21[18] , 
        \wAMid93[11] , \wAMid102[26] , \wRegInA54[28] , \wAMid121[17] , 
        \ScanLink0[2] , \wBIn67[17] , \wBIn72[23] , \wBIn80[6] , \wAMid77[7] , 
        \wBIn104[26] , \wBIn111[12] , \wAMid68[10] , \ScanLink3[1] , 
        \wBIn31[16] , \wBIn44[26] , \wBIn127[17] , \wBIn52[0] , \wBIn117[8] , 
        \wRegInA121[21] , \wRegInA102[10] , \ScanLink161[0] , \wRegInA117[24] , 
        \ScanLink186[18] , \ScanLink201[5] , \wAMid4[28] , \wRegInA120[6] , 
        \wAMid9[9] , \wBIn20[13] , \wBIn55[23] , \wBIn76[12] , \wAMid79[15] , 
        \wRegInA88[30] , \wAIn13[5] , \wBIn16[16] , \wBIn115[23] , 
        \wRegInA88[29] , \wAMid19[11] , \wAMid53[1] , \wBIn63[26] , 
        \wBIn100[17] , \wBIn35[27] , \wBIn40[17] , \wBIn123[26] , 
        \ScanLink158[9] , \ScanLink197[0] , \wAMid81[7] , \wRegInB89[3] , 
        \wRegInA104[0] , \wRegInA125[10] , \wRegInA106[21] , \ScanLink225[3] , 
        \wRegInA113[15] , \ScanLink182[29] , \wBIn1[5] , \wBMid1[12] , 
        \wAIn10[6] , \wBMid39[2] , \wBIn75[5] , \wBIn76[6] , \ScanLink182[30] , 
        \ScanLink145[6] , \wRegInB45[9] , \wRegInA107[3] , \ScanLink226[0] , 
        \ScanLink179[31] , \ScanLink78[7] , \wAMid82[4] , \wRegInB5[9] , 
        \ScanLink179[28] , \ScanLink146[5] , \wAMid82[14] , \wAMid113[23] , 
        \wRegInA25[30] , \wRegInB58[6] , \wRegInA73[28] , \wRegInA50[19] , 
        \wRegInA73[31] , \wRegInA25[29] , \wRegInA38[3] , \ScanLink65[8] , 
        \wBIn12[2] , \wBMid13[31] , \wBMid30[19] , \wAMid50[2] , 
        \wAMid106[17] , \ScanLink194[3] , \wAMid97[20] , \wBIn98[27] , 
        \ScanLink8[21] , \wAMid125[26] , \ScanLink59[30] , \wBMid13[28] , 
        \wBMid45[29] , \wRegInA113[26] , \ScanLink241[7] , \ScanLink59[29] , 
        \wBMid45[30] , \wBMid66[18] , \wRegInA125[23] , \ScanLink232[30] , 
        \ScanLink211[18] , \wAIn123[5] , \ScanLink121[2] , \wBIn2[6] , 
        \wBIn16[25] , \wAIn54[31] , \wBIn100[24] , \wRegInB38[29] , 
        \wRegInA106[12] , \ScanLink247[19] , \ScanLink232[29] , \wBIn63[15] , 
        \wAIn77[19] , \wAMid19[22] , \wBIn20[20] , \wAIn21[18] , \wBIn35[14] , 
        \wBIn40[24] , \wAIn54[28] , \wBIn123[15] , \wRegInB38[30] , 
        \wBIn55[10] , \wAIn77[1] , \wAMid29[9] , \wAMid34[6] , \wAMid37[5] , 
        \wBIn76[21] , \wAMid79[26] , \wAMid97[13] , \wBIn98[14] , 
        \wAMid106[24] , \wBMid107[7] , \wBIn115[10] , \wRegInB95[29] , 
        \wAMid125[15] , \wRegInB95[30] , \ScanLink8[12] , \wBMid40[9] , 
        \wAMid82[27] , \wBMid104[4] , \wAIn74[2] , \wAMid113[10] , 
        \ScanLink242[4] , \ScanLink81[19] , \wRegInA41[8] , \ScanLink122[1] , 
        \wBIn11[1] , \wBMid18[24] , \wAIn120[6] , \wAIn122[13] , 
        \wRegInB92[2] , \ScanLink189[16] , \ScanLink71[14] , \wBMid21[0] , 
        \wBMid78[20] , \wAIn101[22] , \ScanLink60[5] , \ScanLink52[25] , 
        \wAMid117[1] , \ScanLink47[11] , \ScanLink27[15] , \ScanLink32[21] , 
        \wAIn114[16] , \ScanLink239[25] , \ScanLink64[20] , \ScanLink11[10] , 
        \wBIn68[19] , \wRegInB33[25] , \wRegInB40[4] , \wRegInA96[22] , 
        \wRegInB10[14] , \wRegInB46[15] , \wRegInB65[24] , \wBIn2[13] , 
        \wAMid48[0] , \wAIn69[21] , \wBIn70[8] , \wRegInA20[1] , 
        \ScanLink143[8] , \wRegInB70[10] , \wAMid87[9] , \wRegInB0[4] , 
        \wAIn87[14] , \wBIn93[18] , \wBMid114[19] , \wRegInA18[13] , 
        \wRegInB26[11] , \wRegInA83[16] , \wRegInB53[21] , \wRegInB43[7] , 
        \wAIn92[20] , \wRegInB3[7] , \wBMid96[15] , \wRegInA23[2] , 
        \wRegInA78[17] , \ScanLink124[16] , \wAMid99[5] , \wRegInB91[1] , 
        \ScanLink151[26] , \ScanLink107[27] , \ScanLink63[6] , 
        \ScanLink172[17] , \ScanLink112[13] , \wBMid22[3] , \ScanLink167[23] , 
        \wAIn16[8] , \wBMid83[21] , \wAMid24[18] , \wAMid114[2] , 
        \ScanLink131[22] , \ScanLink144[12] , \wAMid51[28] , \wRegInB70[23] , 
        \wBMid0[18] , \wAMid1[20] , \wBIn2[20] , \wBMid18[17] , \wBMid45[4] , 
        \wAMid51[31] , \wAIn69[12] , \wAMid72[19] , \wRegInB24[0] , 
        \wRegInB53[12] , \wBMid78[13] , \wBMid97[2] , \wRegInB26[22] , 
        \wRegInA83[25] , \ScanLink247[9] , \wRegInB33[16] , \wRegInB46[26] , 
        \wRegInA96[11] , \wRegInB10[27] , \wRegInA44[5] , \wRegInB65[17] , 
        \ScanLink32[12] , \wAIn114[25] , \wAIn122[20] , \ScanLink239[16] , 
        \ScanLink64[13] , \ScanLink47[22] , \ScanLink11[23] , 
        \ScanLink189[25] , \wAIn101[11] , \wBMid101[9] , \wRegInA118[19] , 
        \ScanLink71[27] , \wRegInA96[3] , \ScanLink27[26] , \ScanLink52[16] , 
        \wBIn4[8] , \wAMid32[8] , \wBMid83[12] , \wRegInA7[29] , 
        \ScanLink167[10] , \wRegInB115[28] , \ScanLink144[21] , 
        \ScanLink112[20] , \wBMid96[26] , \wRegInA7[30] , \wRegInA95[0] , 
        \wRegInB115[31] , \ScanLink151[15] , \ScanLink131[11] , 
        \ScanLink139[0] , \ScanLink124[25] , \ScanLink172[24] , \wBMid46[7] , 
        \ScanLink107[14] , \wAMid89[18] , \wAIn92[13] , \wRegInB27[3] , 
        \wRegInA47[6] , \wRegInA78[24] , \wBMid6[8] , \wBIn8[15] , 
        \wAMid39[3] , \wAIn79[7] , \wAIn87[27] , \wAIn126[8] , \wBMid89[27] , 
        \wBMid94[1] , \wRegInA18[20] , \wRegInB31[7] , \ScanLink178[11] , 
        \ScanLink80[13] , \wRegInA51[2] , \ScanLink118[15] , \wBMid82[5] , 
        \ScanLink95[27] , \wBMid109[1] , \wRegInA12[15] , \wBMid12[22] , 
        \wAIn16[17] , \wAMid18[31] , \wBMid50[3] , \wAIn64[8] , \wAMid96[19] , 
        \wRegInA67[25] , \wRegInA31[24] , \ScanLink9[18] , \wRegInA44[14] , 
        \wRegInB94[23] , \ScanLink11[6] , \wAIn98[26] , \wRegInA24[10] , 
        \wRegInB81[17] , \wRegInA83[4] , \wRegInA51[20] , \wRegInA72[11] , 
        \wAIn55[22] , \wAMid18[28] , \wAIn20[12] , \wAIn76[13] , 
        \wRegInB39[23] , \ScanLink12[5] , \wBMid53[0] , \wAIn63[27] , 
        \wRegInA89[10] , \wAIn35[26] , \wAIn40[16] , \wRegInB59[27] , 
        \wRegInA80[7] , \ScanLink205[26] , \ScanLink58[23] , \wAIn5[24] , 
        \wBMid31[13] , \wBMid67[12] , \wRegInB32[4] , \ScanLink226[17] , 
        \ScanLink183[10] , \wBMid24[27] , \wBMid44[23] , \ScanLink253[27] , 
        \wRegInA124[30] , \wBMid51[17] , \wRegInA107[18] , \ScanLink233[23] , 
        \ScanLink196[24] , \wBMid81[6] , \wRegInA52[1] , \wRegInA124[29] , 
        \ScanLink246[13] , \ScanLink210[12] , \ScanLink38[27] , \wBMid0[6] , 
        \wAMid1[13] , \wBIn8[26] , \wBMid34[7] , \wAMid40[8] , \wBMid72[26] , 
        \wAIn98[15] , \wAMid112[29] , \wRegInA51[13] , \ScanLink131[8] , 
        \wRegInA24[23] , \wRegInB81[24] , \ScanLink75[2] , \wAMid112[30] , 
        \wRegInA72[22] , \wRegInB87[5] , \wRegInA67[16] , \wBIn78[0] , 
        \wAMid102[6] , \wRegInA12[26] , \wRegInA28[9] , \wRegInA44[27] , 
        \wRegInA31[17] , \wRegInB94[10] , \ScanLink184[9] , \wBMid89[14] , 
        \wRegInA117[9] , \wBMid24[14] , \wBMid29[8] , \wRegInB55[3] , 
        \ScanLink95[14] , \ScanLink178[22] , \ScanLink118[26] , 
        \ScanLink80[20] , \wBMid51[24] , \wBIn120[7] , \wRegInA35[6] , 
        \ScanLink199[6] , \wRegInB56[0] , \wRegInB99[9] , \ScanLink246[20] , 
        \wBMid67[21] , \wBMid72[15] , \ScanLink235[9] , \ScanLink233[10] , 
        \ScanLink196[17] , \ScanLink38[14] , \wRegInA36[5] , \ScanLink210[21] , 
        \wBIn123[4] , \wAIn5[17] , \wBMid12[11] , \ScanLink205[15] , 
        \ScanLink58[10] , \wAIn16[24] , \wBMid31[20] , \wBMid44[10] , 
        \ScanLink253[14] , \ScanLink226[24] , \ScanLink183[23] , \wAIn20[21] , 
        \wBIn21[19] , \wAIn35[15] , \wBIn54[30] , \wAIn63[14] , 
        \wRegInB59[14] , \wRegInB84[6] , \wBIn77[18] , \wBIn114[29] , 
        \wRegInA89[23] , \ScanLink228[6] , \wRegInA109[5] , \wAIn40[25] , 
        \wBIn54[29] , \ScanLink76[1] , \wAMid101[5] , \wBIn114[30] , 
        \wBMid37[4] , \wAIn55[11] , \ScanLink148[3] , \wAIn76[20] , 
        \wRegInB39[10] , \wBMid82[18] , \wBIn87[15] , \wAIn93[19] , 
        \wAMid119[25] , \wBMid123[25] , \wBMid100[14] , \wRegInB37[9] , 
        \wAMid88[12] , \wBIn92[21] , \ScanLink254[0] , \wBMid115[20] , 
        \wRegInA98[5] , \ScanLink2[27] , \ScanLink134[5] , \ScanLink17[8] , 
        \wRegInB124[1] , \wAMid1[1] , \wBIn3[19] , \wBMid3[5] , \wAMid22[2] , 
        \wRegInA6[23] , \wRegInB114[22] , \wAIn62[6] , \wBMid99[4] , 
        \wRegInB101[16] , \wBMid112[0] , \wRegInB0[26] , \wRegInB122[27] , 
        \ScanLink10[29] , \wAMid13[17] , \wBIn19[9] , \wAIn61[5] , 
        \wBMid79[19] , \wRegInB127[2] , \wRegInB29[5] , \ScanLink65[19] , 
        \ScanLink46[31] , \ScanLink10[30] , \wRegInA49[0] , \ScanLink46[28] , 
        \ScanLink33[18] , \wRegInA86[9] , \wAMid21[1] , \wAMid25[12] , 
        \wAIn68[18] , \wBMid111[3] , \wRegInB52[18] , \wRegInA119[13] , 
        \wRegInB71[30] , \wAMid73[13] , \wRegInB27[28] , \wAMid30[26] , 
        \wAMid50[22] , \wRegInB71[29] , \wRegInB27[31] , \wAMid45[16] , 
        \ScanLink137[6] , \wBMid32[9] , \wAMid46[6] , \wBMid48[1] , 
        \wAMid66[27] , \wBIn69[20] , \wBMid87[8] , \wAMid104[8] , 
        \wRegInB0[15] , \wRegInB101[25] , \wRegInB122[14] , \ScanLink182[7] , 
        \ScanLink130[28] , \ScanLink166[30] , \ScanLink145[18] , 
        \wRegInA6[10] , \wRegInB114[11] , \ScanLink113[19] , \ScanLink130[31] , 
        \wRegInA19[19] , \ScanLink166[29] , \ScanLink230[4] , \wAMid2[2] , 
        \wAMid30[15] , \wAMid45[25] , \wBIn63[1] , \wBIn92[12] , 
        \wBMid115[13] , \wAMid119[16] , \wBIn126[9] , \wRegInA111[7] , 
        \ScanLink2[14] , \wRegInA33[8] , \wAMid119[7] , \wBIn87[26] , 
        \wAMid94[0] , \wBMid123[16] , \ScanLink150[1] , \wBMid100[27] , 
        \wAMid88[21] , \wRegInA97[31] , \wRegInA112[4] , \wAMid66[14] , 
        \wRegInA97[28] , \wBIn69[13] , \wAIn5[2] , \wAIn6[1] , \wAMid13[24] , 
        \wAMid17[15] , \wAMid25[21] , \wAMid50[11] , \wAMid73[20] , 
        \ScanLink233[7] , \wAMid97[3] , \wAMid34[24] , \wAMid45[5] , 
        \wBIn60[2] , \ScanLink153[2] , \wAIn100[31] , \wAIn100[28] , 
        \wAIn123[19] , \wRegInB82[8] , \wRegInA119[20] , \ScanLink181[4] , 
        \wAMid41[14] , \wBIn44[4] , \ScanLink177[4] , \wBIn18[12] , 
        \wRegInA4[8] , \wAIn21[7] , \wAMid21[10] , \wAMid62[25] , 
        \wRegInA93[19] , \wAMid77[11] , \wBIn78[16] , \wRegInB74[8] , 
        \ScanLink217[1] , \wAMid54[20] , \wAIn104[19] , \ScanLink49[6] , 
        \wAIn127[31] , \wAMid61[3] , \wBIn96[2] , \wAIn127[28] , \wAMid62[0] , 
        \wRegInB69[7] , \wRegInA108[25] , \ScanLink199[19] , \ScanLink54[9] , 
        \wRegInB105[14] , \wBIn7[31] , \wAIn22[4] , \wBIn95[1] , 
        \wRegInB4[24] , \wRegInB126[25] , \ScanLink169[8] , \wBIn7[28] , 
        \ScanLink141[29] , \ScanLink134[19] , \ScanLink117[31] , 
        \ScanLink98[3] , \wAIn45[3] , \wBIn47[7] , \wBIn96[23] , \wAMid99[24] , 
        \wRegInA2[21] , \ScanLink162[18] , \ScanLink141[30] , \wRegInA68[18] , 
        \wRegInB110[20] , \ScanLink117[28] , \ScanLink6[25] , \wBMid111[22] , 
        \ScanLink174[7] , \wBMid71[8] , \wBIn83[17] , \wAMid108[13] , 
        \wBMid104[16] , \wRegInA108[16] , \ScanLink214[2] , \ScanLink61[28] , 
        \ScanLink37[30] , \ScanLink14[18] , \ScanLink61[31] , \ScanLink42[19] , 
        \ScanLink37[29] , \wAMid0[27] , \wAIn1[26] , \wAMid5[22] , 
        \wBMid16[20] , \wAMid17[26] , \wAMid18[8] , \wAMid77[22] , 
        \wBIn78[25] , \wRegInB103[4] , \ScanLink229[19] , \wRegInB23[19] , 
        \wAIn19[19] , \wBIn20[0] , \wAMid21[23] , \wAMid54[13] , 
        \wRegInB56[29] , \wAIn97[5] , \wRegInA70[9] , \wAIn111[7] , 
        \ScanLink113[0] , \wRegInB56[30] , \wRegInB75[18] , \wAMid34[17] , 
        \wAMid41[27] , \wAMid62[16] , \wBIn18[21] , \wBMid20[25] , \wBIn23[3] , 
        \wAIn94[6] , \wAIn112[4] , \wAIn46[0] , \wBIn83[24] , \wAIn97[31] , 
        \ScanLink110[3] , \wBMid86[29] , \wBIn96[10] , \wAIn97[28] , 
        \wBMid104[25] , \wAMid99[17] , \ScanLink6[16] , \wBMid111[11] , 
        \wAMid108[20] , \wAIn89[9] , \wBMid86[30] , \wRegInA2[12] , 
        \wRegInB4[17] , \wRegInB100[7] , \wRegInB105[27] , \wRegInB110[13] , 
        \wRegInB126[16] , \wBMid55[15] , \wRegInA2[6] , \ScanLink237[21] , 
        \ScanLink192[26] , \wBMid76[24] , \wBIn107[2] , \ScanLink242[11] , 
        \wRegInA12[3] , \ScanLink49[15] , \ScanLink214[10] , \ScanLink201[24] , 
        \ScanLink80[1] , \wBMid35[11] , \wBMid63[10] , \ScanLink222[15] , 
        \ScanLink29[11] , \ScanLink187[12] , \wRegInB72[6] , \wAIn1[15] , 
        \wAMid5[11] , \wBMid10[1] , \wAIn12[15] , \wBMid40[21] , \wAIn67[25] , 
        \wBIn73[29] , \wBIn110[18] , \wRegInB28[15] , \wBMid13[2] , 
        \wAIn24[10] , \wBIn25[31] , \wBIn25[28] , \wAIn27[9] , \wAIn44[14] , 
        \wBIn50[18] , \wBIn73[30] , \wAMid125[3] , \wAIn31[24] , \wAIn51[20] , 
        \wAIn72[11] , \wRegInA98[26] , \ScanLink52[7] , \wBIn88[31] , 
        \wAMid116[18] , \wAMid126[0] , \wRegInB48[11] , \wRegInA20[12] , 
        \wRegInB85[15] , \wBIn88[28] , \wRegInA55[22] , \wAIn12[26] , 
        \wAIn24[23] , \wAIn39[5] , \wAIn89[10] , \wRegInA16[17] , 
        \wRegInA76[13] , \wRegInA63[27] , \wRegInA35[26] , \wRegInA40[16] , 
        \wRegInB90[21] , \ScanLink51[4] , \wBIn41[9] , \wBIn104[1] , 
        \wRegInA11[0] , \ScanLink172[9] , \wAMid79[1] , \wRegInA1[5] , 
        \wBMid98[11] , \wRegInB71[5] , \ScanLink169[27] , \ScanLink91[25] , 
        \ScanLink109[23] , \ScanLink84[11] , \ScanLink83[2] , \wAIn51[13] , 
        \ScanLink108[1] , \wAMid69[30] , \wAMid69[29] , \wRegInB48[22] , 
        \wRegInA98[15] , \wAIn72[22] , \wBMid77[6] , \wAIn31[17] , 
        \wAIn67[16] , \wRegInB28[26] , \wAIn44[27] , \ScanLink36[3] , 
        \wBMid63[23] , \wRegInA76[7] , \ScanLink29[22] , \wBMid16[13] , 
        \wAIn117[9] , \ScanLink201[17] , \wBMid4[30] , \wBMid35[22] , 
        \wBMid40[12] , \ScanLink222[26] , \ScanLink187[21] , \wBMid55[26] , 
        \wRegInB16[2] , \wRegInB118[5] , \wBMid4[29] , \wBMid20[16] , 
        \wRegInA103[29] , \ScanLink242[22] , \wBMid76[17] , \ScanLink237[12] , 
        \ScanLink192[15] , \wBIn9[12] , \wAMid29[4] , \wBIn38[2] , 
        \wBMid74[5] , \wAIn89[23] , \wAIn92[8] , \wRegInA103[30] , 
        \ScanLink49[26] , \wRegInA120[18] , \ScanLink214[23] , 
        \ScanLink109[10] , \ScanLink84[22] , \wAMid92[28] , \wBMid98[22] , 
        \wRegInA75[4] , \wRegInB15[1] , \ScanLink169[14] , \ScanLink91[16] , 
        \wRegInA63[14] , \wRegInA16[24] , \wAMid92[31] , \wRegInA40[25] , 
        \wAIn109[5] , \wRegInA35[15] , \wRegInB90[12] , \wAIn69[0] , 
        \wRegInA20[21] , \wRegInA55[11] , \wRegInB85[26] , \ScanLink35[0] , 
        \wRegInB21[0] , \wRegInA76[20] , \wRegInB106[9] , \ScanLink242[9] , 
        \ScanLink179[16] , \ScanLink81[14] , \wBMid88[20] , \wRegInA41[5] , 
        \ScanLink119[12] , \wBMid92[2] , \ScanLink94[20] , \wBMid13[25] , 
        \wBIn16[31] , \wBIn40[29] , \wBMid40[4] , \wBIn98[19] , \wAMid106[30] , 
        \wBMid119[6] , \wRegInA13[12] , \wAMid125[18] , \wRegInA66[22] , 
        \wAIn99[21] , \wAMid106[29] , \wRegInA30[23] , \wRegInB95[24] , 
        \wRegInA25[17] , \wRegInA45[13] , \wRegInA93[3] , \wRegInA50[27] , 
        \wRegInB80[10] , \wBIn100[30] , \wBMid104[9] , \wBIn123[18] , 
        \wRegInA73[16] , \wAIn54[25] , \wBIn16[28] , \wAIn21[15] , 
        \wBIn35[19] , \wBIn40[30] , \wBIn100[29] , \wRegInB38[24] , 
        \wBIn63[18] , \wAIn77[14] , \wAIn17[10] , \wAMid37[8] , \wAIn62[20] , 
        \wRegInA88[17] , \wAIn34[21] , \wAIn41[11] , \wBMid43[7] , 
        \wRegInB58[20] , \wRegInA90[0] , \ScanLink204[21] , \ScanLink59[24] , 
        \wAMid0[14] , \wBIn1[8] , \wAIn4[23] , \wBMid8[3] , \wBMid66[15] , 
        \ScanLink227[10] , \ScanLink182[17] , \wBMid30[14] , \wRegInB22[3] , 
        \ScanLink252[20] , \wBMid25[20] , \wBMid45[24] , \wBMid50[10] , 
        \ScanLink232[24] , \ScanLink197[23] , \wBMid73[21] , \wBMid91[1] , 
        \wRegInA42[6] , \ScanLink247[14] , \ScanLink211[15] , \wAIn123[8] , 
        \ScanLink39[20] , \wBIn9[21] , \wBMid24[0] , \wAMid82[19] , 
        \wAIn99[12] , \wRegInA25[24] , \wRegInA50[14] , \ScanLink65[5] , 
        \wRegInB80[23] , \wRegInB97[2] , \wRegInA13[21] , \wRegInA66[11] , 
        \wRegInA73[25] , \wBIn68[7] , \wAMid112[1] , \wRegInA45[20] , 
        \wRegInA30[10] , \wRegInB95[17] , \wBMid88[13] , \wBMid25[13] , 
        \wBMid50[23] , \wBIn75[8] , \wAMid82[9] , \wRegInB5[4] , 
        \wRegInB45[4] , \ScanLink94[13] , \ScanLink179[25] , \ScanLink119[21] , 
        \ScanLink81[27] , \wRegInA25[1] , \wRegInB46[7] , \ScanLink189[1] , 
        \ScanLink146[8] , \ScanLink247[27] , \wBMid66[26] , \wBMid73[12] , 
        \ScanLink232[17] , \ScanLink197[10] , \ScanLink211[26] , 
        \ScanLink39[13] , \wRegInA26[2] , \wAIn4[10] , \wBMid13[16] , 
        \ScanLink204[12] , \ScanLink59[17] , \ScanLink252[13] , \wBIn4[5] , 
        \wAMid9[4] , \wAIn17[23] , \wBMid30[27] , \wBMid45[17] , \wRegInB6[7] , 
        \ScanLink227[23] , \ScanLink182[24] , \wRegInA113[18] , 
        \wRegInB58[13] , \wRegInB94[1] , \wAIn13[8] , \wAIn34[12] , 
        \wAIn62[13] , \wAMid79[18] , \wRegInA88[24] , \ScanLink238[1] , 
        \wRegInA119[2] , \wAIn41[22] , \ScanLink66[6] , \wAIn21[26] , 
        \wAMid111[2] , \wBMid27[3] , \wAIn54[16] , \ScanLink158[4] , 
        \wRegInB38[17] , \wAIn77[27] , \wBIn86[12] , \wAMid89[15] , 
        \wAMid118[22] , \wBMid122[22] , \wRegInA78[30] , \wBMid101[13] , 
        \wBIn93[26] , \wRegInA78[29] , \ScanLink244[7] , \ScanLink3[20] , 
        \wBMid114[27] , \wRegInA88[2] , \ScanLink124[2] , \wBIn7[6] , 
        \wBIn14[1] , \wBIn17[2] , \wAMid24[15] , \wAMid31[6] , \wAMid32[5] , 
        \wAIn126[5] , \wRegInA7[24] , \wRegInB115[25] , \ScanLink172[29] , 
        \wAIn71[2] , \wAIn72[1] , \wBMid89[3] , \wRegInB100[11] , 
        \wBMid102[7] , \ScanLink124[31] , \ScanLink107[19] , \ScanLink151[18] , 
        \wAIn114[31] , \wRegInB1[21] , \wRegInB123[20] , \ScanLink172[30] , 
        \ScanLink124[28] , \wRegInB39[2] , \wAIn114[28] , \wRegInA59[7] , 
        \ScanLink189[31] , \wBMid45[9] , \wBMid101[4] , \wAMid72[14] , 
        \wRegInA118[14] , \ScanLink189[28] , \ScanLink247[4] , \wRegInA83[28] , 
        \wAMid31[21] , \wAMid51[25] , \wRegInA44[8] , \wRegInA83[31] , 
        \ScanLink19[3] , \wAMid44[11] , \wAIn125[6] , \ScanLink127[1] , 
        \wAMid12[10] , \wAIn16[5] , \wBMid58[6] , \wAMid67[20] , \wBIn68[27] , 
        \wBMid96[18] , \wRegInB100[22] , \wRegInB123[13] , \wRegInB1[12] , 
        \wAMid56[1] , \ScanLink192[0] , \wAMid99[8] , \wRegInA7[17] , 
        \wRegInB115[16] , \wAIn0[21] , \wAMid4[25] , \wAMid12[23] , 
        \wAMid31[12] , \wAMid44[22] , \wBIn73[6] , \wAIn87[19] , 
        \ScanLink220[3] , \wBIn93[15] , \ScanLink3[13] , \wAMid109[0] , 
        \wBMid114[14] , \wAMid118[11] , \wRegInA101[0] , \wBMid122[11] , 
        \wAMid84[7] , \ScanLink140[6] , \wBIn86[21] , \wAMid89[26] , 
        \wBMid101[20] , \wRegInB10[19] , \wRegInA102[3] , \wRegInB33[31] , 
        \wRegInB65[29] , \wAMid67[13] , \wBIn68[14] , \wRegInB33[28] , 
        \wRegInB40[9] , \wRegInB46[18] , \wRegInB65[30] , \wAIn15[6] , 
        \wBMid18[30] , \wBMid18[29] , \wAMid24[26] , \wAMid51[16] , 
        \wAMid72[27] , \wRegInB0[9] , \ScanLink223[0] , \wAMid87[4] , 
        \wBIn70[5] , \ScanLink143[5] , \wRegInA118[27] , \ScanLink60[8] , 
        \ScanLink52[28] , \ScanLink27[18] , \wAMid55[2] , \ScanLink71[19] , 
        \ScanLink52[31] , \ScanLink239[28] , \wAMid15[0] , \wAMid16[12] , 
        \wBIn19[15] , \wAMid35[23] , \wRegInB42[30] , \wRegInB61[18] , 
        \ScanLink239[31] , \ScanLink191[3] , \wAMid40[13] , \wBIn54[3] , 
        \wAIn78[30] , \wRegInB14[28] , \ScanLink167[3] , \wRegInB42[29] , 
        \wBMid18[4] , \wRegInB37[19] , \wAMid20[17] , \wAMid63[22] , 
        \wRegInB14[31] , \wAMid76[16] , \wAIn78[29] , \ScanLink207[6] , 
        \wBIn79[11] , \wAIn31[0] , \wAMid55[27] , \wRegInA126[5] , 
        \wBMid69[28] , \wRegInA19[5] , \ScanLink96[8] , \ScanLink59[1] , 
        \ScanLink23[29] , \wAIn32[3] , \wBMid69[31] , \wAMid71[4] , 
        \wBIn86[5] , \ScanLink75[31] , \ScanLink56[19] , \wRegInA9[0] , 
        \wAMid72[7] , \wRegInB79[0] , \ScanLink248[29] , \ScanLink75[28] , 
        \ScanLink23[30] , \ScanLink5[2] , \wRegInA109[22] , \ScanLink248[30] , 
        \wBMid92[30] , \wRegInB104[13] , \wBIn57[0] , \wAIn83[31] , 
        \wAIn83[28] , \wBIn85[6] , \wBMid92[29] , \wRegInB127[22] , 
        \wRegInB5[23] , \wBIn97[24] , \wBMid110[25] , \wRegInA3[26] , 
        \ScanLink88[4] , \ScanLink6[1] , \wRegInB111[27] , \wAMid98[23] , 
        \ScanLink7[22] , \wBIn98[9] , \wBIn112[8] , \ScanLink164[0] , 
        \wBIn82[10] , \wAMid109[14] , \wBMid126[20] , \wRegInA125[6] , 
        \wBMid105[11] , \wRegInA109[11] , \ScanLink204[5] , \wAMid16[21] , 
        \wBIn19[26] , \wAMid20[24] , \wAIn55[4] , \wBMid125[2] , \wAMid55[14] , 
        \wAMid76[25] , \wAIn110[19] , \wRegInB113[3] , \wBIn79[22] , 
        \wRegInA87[19] , \wAIn87[2] , \wBIn30[7] , \wAIn101[0] , 
        \ScanLink103[7] , \wAMid35[10] , \wAMid40[20] , \wAMid63[11] , 
        \wAMid16[3] , \wBIn33[4] , \wAIn84[1] , \wAIn102[3] , \wAIn56[7] , 
        \wBIn82[23] , \wBMid126[13] , \ScanLink100[4] , \wBIn97[17] , 
        \wBMid105[22] , \wBMid110[16] , \wAMid98[10] , \ScanLink7[11] , 
        \wAMid109[27] , \wBMid17[27] , \wBMid21[22] , \wBMid126[1] , 
        \wRegInA3[15] , \wRegInB111[14] , \wRegInB127[11] , \wRegInB104[20] , 
        \ScanLink103[28] , \wRegInB110[0] , \ScanLink176[18] , 
        \ScanLink155[30] , \wRegInB5[10] , \ScanLink120[19] , 
        \ScanLink103[31] , \ScanLink155[29] , \ScanLink23[9] , \wBMid54[12] , 
        \ScanLink236[26] , \ScanLink193[21] , \wBMid77[23] , \wBIn117[5] , 
        \ScanLink243[16] , \ScanLink215[17] , \ScanLink48[12] , 
        \ScanLink200[23] , \wRegInA117[30] , \ScanLink90[6] , \wBMid34[16] , 
        \wBMid62[17] , \ScanLink28[16] , \wRegInB62[1] , \wRegInA117[29] , 
        \ScanLink223[12] , \ScanLink186[15] , \ScanLink201[8] , \wAIn0[12] , 
        \wAMid4[16] , \wBIn12[19] , \wAIn13[12] , \wBMid41[26] , 
        \ScanLink256[22] , \wAIn66[22] , \wRegInB29[12] , \wAIn25[24] , 
        \wAIn25[17] , \wAIn30[23] , \wAIn45[13] , \wAIn50[27] , \wAIn29[2] , 
        \wAIn73[16] , \wRegInA99[21] , \ScanLink42[0] , \wAMid74[9] , 
        \wBIn83[8] , \wAMid86[31] , \wBIn109[9] , \wRegInA21[15] , 
        \wRegInB49[16] , \wRegInB84[12] , \wRegInA54[25] , \wAMid86[28] , 
        \wAIn88[17] , \wRegInA17[10] , \wRegInA77[14] , \wRegInA62[20] , 
        \wRegInA34[21] , \wRegInB91[26] , \wRegInA41[11] , \ScanLink41[3] , 
        \wBIn31[28] , \wAMid69[6] , \wBIn114[6] , \wRegInA8[19] , 
        \wBMid99[16] , \wRegInB61[2] , \ScanLink168[20] , \ScanLink90[22] , 
        \ScanLink108[24] , \wRegInA123[8] , \ScanLink85[16] , \ScanLink93[5] , 
        \wBIn31[31] , \wBIn44[18] , \wAIn50[14] , \wBIn67[30] , \wBIn127[29] , 
        \ScanLink118[6] , \wRegInB49[25] , \wAIn13[21] , \wBIn67[29] , 
        \wBIn104[18] , \wRegInA99[12] , \wBIn127[30] , \wBMid67[1] , 
        \wAIn73[25] , \wAIn30[10] , \wAIn66[11] , \wRegInB29[21] , 
        \wAIn45[20] , \ScanLink26[4] , \wBMid62[24] , \wRegInA66[0] , 
        \ScanLink28[25] , \wBMid17[14] , \wBIn36[9] , \ScanLink200[10] , 
        \ScanLink105[9] , \wBIn7[16] , \wBMid21[11] , \wBMid34[25] , 
        \wBMid41[15] , \ScanLink256[11] , \ScanLink223[21] , \ScanLink186[26] , 
        \wBMid54[21] , \wRegInB108[2] , \ScanLink243[25] , \wBIn28[5] , 
        \wAIn50[9] , \wBMid64[2] , \wBMid77[10] , \ScanLink236[15] , 
        \ScanLink193[12] , \wAIn88[24] , \wBMid99[25] , \wRegInA65[3] , 
        \ScanLink215[24] , \ScanLink48[21] , \ScanLink108[17] , 
        \ScanLink85[25] , \wRegInA62[13] , \ScanLink168[13] , \ScanLink90[11] , 
        \ScanLink38[8] , \wAMid121[29] , \wRegInA17[23] , \wRegInA41[22] , 
        \wAIn119[2] , \wRegInA34[12] , \wRegInB91[15] , \wAMid102[18] , 
        \wAMid121[30] , \wRegInB18[9] , \wRegInA21[26] , \wRegInA54[16] , 
        \ScanLink25[7] , \wRegInA77[27] , \wRegInB84[21] , \ScanLink117[16] , 
        \wAMid18[5] , \wAIn58[1] , \wBMid72[6] , \wBIn78[31] , \wAIn82[11] , 
        \wBIn83[30] , \wBIn83[29] , \wBMid86[24] , \ScanLink162[26] , 
        \wAIn89[4] , \wBMid93[10] , \ScanLink141[17] , \ScanLink134[27] , 
        \ScanLink121[13] , \wAIn97[25] , \ScanLink177[12] , \ScanLink154[23] , 
        \ScanLink102[22] , \ScanLink33[3] , \wBMid104[28] , \wBMid104[31] , 
        \wAIn112[9] , \wRegInA73[7] , \wRegInB13[2] , \wRegInA68[26] , 
        \wBIn78[28] , \wAIn97[8] , \wRegInA70[4] , \wRegInB75[15] , 
        \wAIn19[14] , \wRegInB23[14] , \wRegInA86[13] , \wBMid71[5] , 
        \wAIn79[10] , \wRegInB10[1] , \wRegInB36[20] , \wRegInB56[24] , 
        \wRegInA93[27] , \wAIn111[13] , \wRegInB15[11] , \wRegInB43[10] , 
        \wRegInB60[21] , \ScanLink42[14] , \ScanLink37[24] , \ScanLink199[27] , 
        \ScanLink61[25] , \ScanLink14[15] , \wAIn127[16] , \wRegInB103[9] , 
        \ScanLink249[10] , \ScanLink229[14] , \ScanLink74[11] , \wAIn0[2] , 
        \wAIn1[18] , \wBIn7[25] , \wBMid16[2] , \wAIn22[9] , \wBMid68[11] , 
        \wAIn104[27] , \ScanLink57[20] , \ScanLink30[0] , \ScanLink22[10] , 
        \wAIn82[22] , \wBIn88[3] , \wAMid99[30] , \wBIn102[2] , \wRegInA17[3] , 
        \ScanLink6[31] , \wRegInA7[6] , \wRegInA68[15] , \wAIn97[16] , 
        \wAMid99[29] , \ScanLink6[28] , \wAMid120[3] , \wRegInB77[6] , 
        \ScanLink85[1] , \ScanLink154[10] , \wBMid93[23] , \wRegInB126[28] , 
        \ScanLink169[5] , \ScanLink121[20] , \wRegInB4[29] , \wRegInB105[19] , 
        \wRegInB126[31] , \ScanLink177[21] , \ScanLink102[11] , \wRegInB4[30] , 
        \wBMid15[1] , \wBMid86[17] , \ScanLink209[0] , \ScanLink162[15] , 
        \ScanLink117[25] , \ScanLink141[24] , \wAIn127[25] , \ScanLink134[14] , 
        \ScanLink57[7] , \ScanLink229[27] , \wAMid17[18] , \wBIn59[6] , 
        \wBMid68[22] , \wAIn104[14] , \ScanLink74[22] , \wAMid123[0] , 
        \ScanLink22[23] , \wAIn111[20] , \ScanLink57[13] , \ScanLink37[17] , 
        \wRegInB43[23] , \wRegInA108[31] , \wRegInA108[28] , \ScanLink249[23] , 
        \ScanLink54[4] , \ScanLink42[27] , \ScanLink14[26] , \ScanLink61[16] , 
        \ScanLink199[14] , \wAIn19[27] , \wAMid34[30] , \wRegInA4[5] , 
        \wAMid34[29] , \wAMid62[28] , \wAIn79[23] , \wRegInB36[13] , 
        \wRegInA93[14] , \wBIn101[1] , \wRegInA14[0] , \wRegInB60[12] , 
        \wAMid41[19] , \wBIn44[9] , \wRegInB15[22] , \wAMid62[31] , 
        \ScanLink177[9] , \wRegInB75[26] , \ScanLink86[2] , \wBIn25[0] , 
        \wAIn40[3] , \wRegInB23[27] , \wRegInB56[17] , \wRegInB74[5] , 
        \ScanLink8[7] , \wRegInA40[28] , \wRegInA68[6] , \wRegInA86[20] , 
        \wBMid74[8] , \wAMid92[25] , \wAMid103[12] , \wAIn109[8] , 
        \wRegInA16[30] , \wRegInA35[18] , \wRegInA40[31] , \wRegInA63[19] , 
        \wRegInA16[29] , \wAMid87[11] , \wBIn88[16] , \wAMid120[23] , 
        \wAIn92[5] , \wAMid116[26] , \wRegInB106[4] , \wRegInA75[9] , 
        \wAIn114[7] , \wBMid69[7] , \ScanLink116[0] , \wRegInA9[20] , 
        \ScanLink169[19] , \ScanLink28[2] , \wAIn3[1] , \wBMid4[24] , 
        \wBIn26[3] , \wAIn91[6] , \wRegInA116[10] , \wAIn117[4] , 
        \ScanLink115[3] , \wBIn13[13] , \wRegInA103[24] , \wRegInB118[8] , 
        \wRegInA120[15] , \ScanLink192[18] , \wBIn25[16] , \wBIn30[22] , 
        \wAIn43[0] , \wBIn66[23] , \wAMid69[24] , \wBIn105[12] , 
        \wRegInA98[18] , \wBIn45[12] , \wBIn126[23] , \wAIn39[8] , 
        \wBIn50[26] , \wBIn73[17] , \wRegInB105[7] , \wBIn110[26] , 
        \wRegInA1[8] , \wRegInA9[13] , \ScanLink91[28] , \wBIn41[4] , 
        \ScanLink172[4] , \ScanLink91[31] , \wAMid64[3] , \wRegInB71[8] , 
        \ScanLink212[1] , \wBIn88[25] , \wAIn12[18] , \wAIn24[7] , 
        \wAMid87[22] , \wBIn25[25] , \wAIn27[4] , \wAIn44[19] , \wBIn50[15] , 
        \wAMid92[16] , \wBIn93[2] , \wAMid116[15] , \wBIn119[3] , 
        \wRegInB85[18] , \wAMid103[21] , \wAMid120[10] , \ScanLink51[9] , 
        \wAIn67[31] , \wAIn31[29] , \wAIn31[30] , \wAIn67[28] , \wBIn90[1] , 
        \wAMid67[0] , \wBIn73[24] , \wBIn110[15] , \wRegInB28[18] , 
        \wAIn1[22] , \wBMid0[26] , \wBMid4[17] , \wBIn13[20] , \wBIn66[10] , 
        \wAMid69[17] , \wBIn105[21] , \wBMid20[31] , \wBIn30[11] , 
        \wBIn45[21] , \wBIn126[10] , \wRegInA120[26] , \ScanLink49[18] , 
        \wBIn42[7] , \wBMid76[29] , \wAIn16[30] , \wBIn21[14] , \wBMid20[28] , 
        \wRegInA103[17] , \ScanLink171[7] , \wBMid55[18] , \wBMid76[30] , 
        \wRegInA116[23] , \ScanLink222[18] , \ScanLink201[30] , 
        \ScanLink211[2] , \ScanLink201[29] , \wAIn16[29] , \wAIn35[18] , 
        \wAIn40[28] , \wRegInA109[8] , \wBIn54[24] , \wBIn17[11] , 
        \wAMid18[16] , \wAIn40[31] , \wBIn77[15] , \wRegInB59[19] , 
        \wAMid43[6] , \wAIn63[19] , \wAMid78[12] , \wBIn114[24] , \wBIn34[20] , 
        \wBMid37[9] , \wBIn101[10] , \wBIn62[21] , \wAMid101[8] , \wBIn41[10] , 
        \wBIn122[21] , \wRegInA114[7] , \ScanLink187[7] , \ScanLink38[19] , 
        \wBMid0[15] , \wAMid4[1] , \wBMid51[30] , \wBMid72[18] , \wBMid51[29] , 
        \wRegInA124[17] , \wRegInB99[4] , \wAIn5[30] , \wAIn5[29] , 
        \wAMid7[2] , \wBMid24[19] , \wBIn66[1] , \wAMid91[0] , 
        \wRegInA107[26] , \ScanLink235[4] , \wBIn123[9] , \wRegInA112[12] , 
        \ScanLink253[19] , \ScanLink226[29] , \wRegInA36[8] , 
        \ScanLink226[30] , \ScanLink205[18] , \ScanLink155[1] , 
        \ScanLink236[7] , \ScanLink95[19] , \wBMid29[5] , \wBIn65[2] , 
        \wBMid89[19] , \wRegInA117[4] , \ScanLink68[0] , \wAMid92[3] , 
        \ScanLink156[2] , \wAMid40[5] , \wAMid83[13] , \wAIn98[18] , 
        \wRegInB87[8] , \wAMid107[10] , \wAMid112[24] , \wRegInB48[1] , 
        \wRegInB81[30] , \wRegInA28[4] , \wRegInB81[29] , \ScanLink184[4] , 
        \wAMid96[27] , \ScanLink9[26] , \wBIn99[20] , \wRegInB8[1] , 
        \wAMid124[21] , \wRegInB32[9] , \wRegInA112[21] , \ScanLink251[0] , 
        \wRegInA124[24] , \ScanLink196[30] , \wAIn3[8] , \wBIn3[27] , 
        \wBIn3[14] , \wBMid5[6] , \wBIn101[23] , \wRegInA107[15] , 
        \ScanLink131[5] , \ScanLink196[29] , \wBMid6[5] , \wBIn17[22] , 
        \wAMid18[25] , \wBIn62[12] , \wRegInB121[1] , \wBIn21[27] , 
        \wBIn34[13] , \wBIn41[23] , \wBIn122[12] , \wBIn54[17] , 
        \ScanLink12[8] , \wAIn67[6] , \wAMid27[2] , \wBIn77[26] , 
        \wAMid78[21] , \wAMid107[23] , \wBIn114[17] , \wBMid117[0] , 
        \wRegInA31[29] , \wAMid124[12] , \wRegInA12[18] , \wRegInA31[30] , 
        \wRegInA44[19] , \wRegInA67[31] , \wRegInB122[2] , \wBIn8[18] , 
        \wAMid24[1] , \wAMid96[14] , \wRegInA67[28] , \ScanLink9[15] , 
        \wBIn99[13] , \wAIn64[5] , \wAMid83[20] , \wBMid114[3] , 
        \wRegInA83[9] , \wAMid112[17] , \ScanLink252[3] , \ScanLink118[18] , 
        \wAMid13[30] , \wAMid13[29] , \wBMid19[23] , \wBMid82[8] , 
        \wAIn123[14] , \wRegInB82[5] , \ScanLink188[11] , \ScanLink132[6] , 
        \ScanLink70[13] , \ScanLink53[22] , \wBMid31[7] , \wAMid45[8] , 
        \wBMid79[27] , \wAIn100[25] , \wAMid107[6] , \ScanLink70[2] , 
        \ScanLink46[16] , \ScanLink26[12] , \wAIn115[11] , \ScanLink181[9] , 
        \ScanLink33[26] , \ScanLink238[22] , \ScanLink65[27] , 
        \ScanLink10[17] , \wAMid45[31] , \wAMid66[19] , \wRegInB32[22] , 
        \wRegInA97[25] , \wRegInB50[3] , \wRegInB47[12] , \wAMid30[18] , 
        \wAMid45[28] , \wRegInB11[13] , \wRegInA112[9] , \wRegInB64[23] , 
        \wAIn18[3] , \wAMid58[7] , \wAIn68[26] , \wBIn125[7] , \wRegInA30[6] , 
        \wRegInB71[17] , \wAIn86[13] , \wRegInA19[14] , \wRegInB27[16] , 
        \wRegInB52[26] , \wRegInA82[11] , \wRegInB53[0] , \ScanLink230[9] , 
        \ScanLink2[19] , \wAMid89[2] , \wAIn93[27] , \wBMid97[12] , 
        \wBIn126[4] , \wRegInA33[5] , \wRegInA79[10] , \wRegInB0[18] , 
        \wRegInB101[31] , \wRegInB122[19] , \ScanLink125[11] , \wRegInB81[6] , 
        \ScanLink150[21] , \ScanLink73[1] , \wRegInB101[28] , 
        \ScanLink106[20] , \ScanLink173[10] , \ScanLink113[14] , \wBMid3[8] , 
        \wBMid32[4] , \wAIn68[15] , \wBMid82[26] , \ScanLink166[24] , 
        \wAMid104[5] , \ScanLink130[25] , \wRegInB34[7] , \wRegInB71[24] , 
        \ScanLink145[15] , \wRegInB52[15] , \wBMid79[14] , \wBMid87[5] , 
        \wRegInB27[25] , \wRegInB32[11] , \wRegInB47[21] , \wRegInA82[22] , 
        \wRegInA97[16] , \wRegInB11[20] , \wRegInA54[2] , \wRegInB64[10] , 
        \wAIn115[22] , \ScanLink33[15] , \ScanLink46[25] , \ScanLink14[6] , 
        \wBIn19[4] , \wBMid55[3] , \wAIn123[27] , \wRegInB29[8] , 
        \ScanLink10[24] , \ScanLink238[11] , \ScanLink65[14] , 
        \ScanLink188[22] , \wAIn61[8] , \wAIn100[16] , \ScanLink70[20] , 
        \wRegInA86[4] , \ScanLink26[21] , \wBMid19[10] , \ScanLink53[11] , 
        \wBIn9[0] , \wBMid82[15] , \ScanLink249[2] , \ScanLink166[17] , 
        \ScanLink145[26] , \ScanLink113[27] , \wRegInA85[7] , 
        \ScanLink130[16] , \ScanLink17[5] , \ScanLink150[12] , 
        \ScanLink129[7] , \ScanLink125[22] , \wAIn39[1] , \wBMid56[0] , 
        \wBMid97[21] , \wBMid99[9] , \ScanLink173[23] , \ScanLink106[13] , 
        \wAMid79[5] , \wBMid84[6] , \wAIn86[20] , \wBIn87[18] , \wAIn93[14] , 
        \wBMid100[19] , \wRegInB37[4] , \wAMid119[31] , \wBMid123[31] , 
        \wRegInA79[23] , \wAMid119[28] , \wBMid123[28] , \wRegInA57[1] , 
        \wRegInA98[8] , \ScanLink134[8] , \wRegInA19[27] , \wBMid98[15] , 
        \wRegInA1[1] , \wRegInB71[1] , \ScanLink109[27] , \ScanLink83[6] , 
        \ScanLink212[8] , \ScanLink84[15] , \ScanLink169[23] , 
        \ScanLink91[21] , \wAIn89[14] , \wAMid103[31] , \wAMid103[28] , 
        \wBIn104[5] , \wRegInA11[4] , \wRegInA35[22] , \wRegInB90[25] , 
        \wRegInA16[13] , \wRegInA40[12] , \ScanLink51[0] , \wAMid120[19] , 
        \wRegInA63[23] , \wBMid10[5] , \wRegInA76[17] , \wAIn12[11] , 
        \wBIn13[30] , \wBIn13[29] , \wBIn45[31] , \wAIn72[15] , \wBIn105[28] , 
        \wAMid126[4] , \wRegInA20[16] , \wRegInB85[11] , \wRegInA55[26] , 
        \wRegInA98[22] , \wBIn66[19] , \wRegInB48[15] , \wAIn24[14] , 
        \wBIn45[28] , \wBIn105[31] , \wBIn126[19] , \wAIn51[24] , \wBMid13[6] , 
        \wBIn30[18] , \wAIn31[20] , \wAIn44[10] , \ScanLink52[3] , 
        \wAMid125[7] , \wAIn67[21] , \wAMid67[9] , \wBIn90[8] , 
        \wRegInB28[11] , \wBMid35[15] , \wRegInB72[2] , \ScanLink222[11] , 
        \ScanLink187[16] , \wAIn1[11] , \wAMid5[26] , \wBMid16[24] , 
        \wBMid40[25] , \ScanLink201[20] , \ScanLink80[5] , \wBMid20[21] , 
        \wBMid63[14] , \ScanLink29[15] , \wBMid76[20] , \wBIn107[6] , 
        \wRegInA12[7] , \ScanLink49[11] , \ScanLink214[14] , \wBMid20[12] , 
        \wBIn25[9] , \wBIn38[6] , \wBMid55[11] , \wRegInA2[2] , 
        \ScanLink237[25] , \ScanLink192[22] , \wAMid87[18] , \ScanLink242[15] , 
        \wAIn109[1] , \wRegInA20[25] , \wRegInA55[15] , \wRegInA76[24] , 
        \wRegInB85[22] , \ScanLink35[4] , \wRegInA35[11] , \wRegInA40[21] , 
        \wRegInB90[16] , \wBMid74[1] , \wAIn89[27] , \wRegInA63[10] , 
        \wRegInA9[30] , \wRegInA9[29] , \wRegInB15[5] , \wRegInA16[20] , 
        \ScanLink91[12] , \ScanLink169[10] , \wRegInA75[0] , \wBMid55[22] , 
        \wBMid76[13] , \wBMid98[26] , \ScanLink116[9] , \ScanLink109[14] , 
        \ScanLink84[26] , \ScanLink214[27] , \ScanLink49[22] , \wRegInB16[6] , 
        \wRegInB118[1] , \ScanLink242[26] , \ScanLink237[16] , 
        \ScanLink192[11] , \wAIn5[6] , \wAMid5[15] , \wBMid35[26] , 
        \wBMid40[16] , \ScanLink222[22] , \ScanLink187[25] , \wBMid63[27] , 
        \wRegInA76[3] , \wRegInA116[19] , \ScanLink29[26] , \wAIn12[22] , 
        \wBMid16[17] , \ScanLink201[13] , \wAIn31[13] , \wAIn44[23] , 
        \ScanLink36[7] , \wAIn22[0] , \wAIn24[27] , \wAIn43[9] , \wAIn67[12] , 
        \wAIn72[26] , \wRegInB28[22] , \wRegInB48[26] , \wRegInA98[11] , 
        \wBMid77[2] , \wBIn47[3] , \wAIn51[17] , \ScanLink108[5] , 
        \wBIn83[13] , \wBMid104[12] , \ScanLink214[6] , \ScanLink174[3] , 
        \ScanLink85[8] , \wBIn96[27] , \wAMid108[17] , \wBMid111[26] , 
        \wAMid99[20] , \ScanLink6[21] , \wRegInA2[25] , \wRegInB110[24] , 
        \ScanLink209[9] , \ScanLink98[7] , \wAMid62[4] , \wBIn95[5] , 
        \ScanLink177[31] , \ScanLink154[19] , \wRegInB4[20] , \wRegInB126[21] , 
        \ScanLink121[29] , \ScanLink177[28] , \wRegInB105[10] , 
        \ScanLink102[18] , \ScanLink121[30] , \wAIn6[5] , \wBMid15[8] , 
        \wAMid61[7] , \wAIn111[30] , \wAIn111[29] , \wRegInB69[3] , 
        \wRegInA108[21] , \wAMid17[22] , \wAMid17[11] , \wBIn18[16] , 
        \wAIn21[3] , \wAMid21[14] , \wBIn96[6] , \wAMid123[9] , \wAMid54[24] , 
        \wAMid77[15] , \wRegInA86[30] , \ScanLink217[5] , \ScanLink49[2] , 
        \wBIn78[12] , \wRegInA86[29] , \wBIn18[25] , \wBIn23[7] , 
        \wAMid34[20] , \wAMid62[21] , \wBIn101[8] , \wRegInA14[9] , 
        \wAMid41[10] , \wBIn44[0] , \ScanLink177[0] , \wAIn46[4] , 
        \wBMid93[19] , \wRegInB4[13] , \wRegInB126[12] , \wRegInA2[16] , 
        \wRegInB100[3] , \wRegInB105[23] , \wRegInB110[17] , \wAIn82[18] , 
        \wAMid108[24] , \wBIn83[20] , \wBIn96[14] , \wBMid111[15] , 
        \wAMid99[13] , \ScanLink6[12] , \wAIn94[2] , \wBMid104[21] , 
        \wAIn112[0] , \wAMid62[12] , \wAIn79[19] , \wRegInB10[8] , 
        \wRegInB36[29] , \ScanLink110[7] , \wRegInB43[19] , \wRegInB60[31] , 
        \wBIn20[4] , \wAMid21[27] , \wAMid34[13] , \wAMid41[23] , 
        \wRegInB15[18] , \wRegInB36[30] , \wRegInB60[28] , \wAMid54[17] , 
        \wAIn58[8] , \wAIn97[1] , \wAIn111[3] , \ScanLink113[4] , 
        \wAMid77[26] , \wBIn78[21] , \wRegInB103[0] , \ScanLink74[18] , 
        \ScanLink57[30] , \ScanLink57[29] , \wBMid0[2] , \wBMid3[1] , 
        \wAMid13[13] , \wAIn45[7] , \wBMid68[18] , \ScanLink30[9] , 
        \ScanLink22[19] , \wRegInB47[28] , \wRegInA108[12] , \ScanLink249[19] , 
        \wBMid19[19] , \wAMid21[5] , \wAMid25[16] , \wAMid30[22] , 
        \wBMid48[5] , \wAMid66[23] , \wBIn69[24] , \wRegInB11[30] , 
        \wRegInB32[18] , \wRegInB47[31] , \wRegInB64[19] , \wAMid45[12] , 
        \wRegInB11[29] , \ScanLink137[2] , \wAMid50[26] , \wAMid73[17] , 
        \wAIn61[1] , \wBMid111[7] , \ScanLink26[31] , \wRegInA49[4] , 
        \wRegInA119[17] , \ScanLink70[29] , \ScanLink70[30] , \ScanLink26[28] , 
        \ScanLink53[18] , \wBIn9[9] , \wAIn62[2] , \wRegInB127[6] , 
        \wRegInB29[1] , \ScanLink238[18] , \wAMid22[6] , \wBMid97[28] , 
        \wRegInB122[23] , \wRegInB0[22] , \wBMid56[9] , \wBMid97[31] , 
        \wBMid99[0] , \wRegInB101[12] , \wBMid112[4] , \wRegInB124[5] , 
        \wAMid1[24] , \wAMid1[5] , \wAMid2[6] , \wAMid25[25] , \wAMid45[1] , 
        \wAIn86[30] , \wRegInA6[27] , \wRegInA57[8] , \wRegInA98[1] , 
        \wRegInB114[26] , \wAIn86[29] , \wBIn92[25] , \ScanLink134[1] , 
        \ScanLink2[23] , \wBMid115[24] , \wBIn87[11] , \wAMid88[16] , 
        \wBMid100[10] , \wAIn115[18] , \wAMid119[21] , \wBMid123[21] , 
        \ScanLink254[4] , \ScanLink181[0] , \wAMid50[15] , \wRegInA119[24] , 
        \ScanLink188[18] , \wBIn60[6] , \ScanLink153[6] , \wAMid66[10] , 
        \wBIn69[17] , \wAMid73[24] , \wAMid97[7] , \wRegInA82[18] , 
        \wAMid13[20] , \wAMid30[11] , \wAMid45[21] , \wRegInA112[0] , 
        \ScanLink233[3] , \wBIn63[5] , \wBIn87[22] , \wAMid88[25] , 
        \wAMid94[4] , \wBMid100[23] , \wAMid119[12] , \wRegInA79[19] , 
        \wAMid119[3] , \wBMid123[12] , \wRegInB53[9] , \wRegInA111[3] , 
        \ScanLink150[5] , \ScanLink230[0] , \wAIn5[20] , \wBMid24[23] , 
        \wAMid46[2] , \wBIn92[16] , \ScanLink2[10] , \wBMid115[17] , 
        \wBMid72[22] , \wRegInB0[11] , \wRegInA6[14] , \wRegInB114[15] , 
        \wRegInB122[10] , \ScanLink182[3] , \ScanLink125[18] , 
        \ScanLink106[30] , \wRegInA52[5] , \wRegInB101[21] , \ScanLink150[28] , 
        \ScanLink73[8] , \ScanLink173[19] , \ScanLink106[29] , 
        \ScanLink150[31] , \ScanLink210[16] , \ScanLink38[23] , \wBMid31[17] , 
        \wBMid51[13] , \ScanLink233[27] , \ScanLink196[20] , \wBMid81[2] , 
        \wRegInA112[28] , \ScanLink246[17] , \ScanLink226[13] , 
        \ScanLink183[14] , \wRegInB32[0] , \ScanLink253[23] , \wBMid12[26] , 
        \wBMid44[27] , \ScanLink251[9] , \wRegInA112[31] , \ScanLink205[22] , 
        \ScanLink58[27] , \wAMid1[17] , \wAIn5[13] , \wBIn8[11] , \wAIn16[13] , 
        \wAIn35[22] , \wAIn40[12] , \wBMid67[16] , \wAMid78[31] , 
        \wRegInA80[3] , \wAIn63[23] , \wAMid78[28] , \wRegInA89[14] , 
        \wAIn20[16] , \wBMid53[4] , \wAIn55[26] , \wAIn76[17] , \wBMid117[9] , 
        \wRegInB39[27] , \wRegInB59[23] , \wRegInB121[8] , \wAMid24[8] , 
        \ScanLink12[1] , \wAMid39[7] , \wBMid50[7] , \wAMid83[29] , 
        \wAIn98[22] , \wAMid83[30] , \wRegInA24[14] , \wRegInA72[15] , 
        \wRegInB81[13] , \wRegInA83[0] , \wRegInA12[11] , \wRegInA31[20] , 
        \wRegInA51[24] , \wRegInA44[10] , \wRegInB94[27] , \ScanLink11[2] , 
        \wRegInA67[21] , \ScanLink118[11] , \wBMid82[1] , \ScanLink95[23] , 
        \wAIn16[20] , \wBIn17[18] , \wBIn34[30] , \wAIn79[3] , \wBMid109[5] , 
        \wBMid89[23] , \wRegInB31[3] , \wRegInA51[6] , \ScanLink178[15] , 
        \ScanLink80[17] , \wAIn20[25] , \wBIn34[29] , \wBMid37[0] , 
        \wBIn62[28] , \wBIn101[19] , \wRegInB39[14] , \wBIn122[31] , 
        \wAIn76[24] , \wAMid101[1] , \wAIn35[11] , \wBIn41[19] , \wAIn55[15] , 
        \wBIn122[28] , \ScanLink148[7] , \wBIn62[31] , \wAIn40[21] , 
        \wRegInA109[1] , \ScanLink76[5] , \wAIn63[10] , \wRegInB59[10] , 
        \wRegInB84[2] , \wRegInA89[27] , \ScanLink228[2] , \ScanLink253[10] , 
        \wBMid31[24] , \wBMid44[14] , \wAMid91[9] , \ScanLink226[20] , 
        \ScanLink183[27] , \wBMid67[25] , \wRegInA36[1] , \wBIn2[17] , 
        \wAMid4[8] , \wBMid12[15] , \wBIn66[8] , \wBIn123[0] , 
        \ScanLink205[11] , \ScanLink155[8] , \ScanLink58[14] , \wBMid24[10] , 
        \wBMid51[20] , \wBMid72[11] , \wRegInB56[4] , \ScanLink210[25] , 
        \ScanLink38[10] , \ScanLink246[24] , \wBIn8[22] , \wBIn120[3] , 
        \wRegInA35[2] , \ScanLink233[14] , \ScanLink196[13] , \ScanLink199[2] , 
        \ScanLink178[26] , \ScanLink80[24] , \wBMid34[3] , \wBIn78[4] , 
        \wBMid89[10] , \wRegInB55[7] , \ScanLink95[10] , \ScanLink118[22] , 
        \wBIn99[30] , \wRegInA44[23] , \ScanLink68[9] , \wAMid102[2] , 
        \wRegInA31[13] , \wRegInB94[14] , \wBIn99[29] , \wAMid107[19] , 
        \wAMid124[31] , \wRegInA67[12] , \wRegInB8[8] , \wRegInA12[22] , 
        \wAMid56[8] , \wBMid83[25] , \wAIn98[11] , \wAMid124[28] , 
        \wRegInA24[27] , \wRegInB48[8] , \wRegInB87[1] , \wRegInA51[17] , 
        \wRegInA72[26] , \wRegInB81[20] , \ScanLink75[6] , \wAMid114[6] , 
        \ScanLink131[26] , \ScanLink192[9] , \ScanLink144[16] , \wAMid99[1] , 
        \ScanLink112[17] , \wBMid22[7] , \wAMid48[4] , \wAIn69[25] , 
        \wBIn86[31] , \wBMid96[11] , \wRegInB91[5] , \ScanLink167[27] , 
        \ScanLink172[13] , \ScanLink107[23] , \ScanLink124[12] , \wAMid109[9] , 
        \wAMid118[18] , \wRegInA23[6] , \ScanLink151[22] , \ScanLink63[2] , 
        \wBMid122[18] , \wBIn86[28] , \wAIn92[24] , \wBMid101[30] , 
        \wRegInB3[3] , \wAIn87[10] , \wBMid101[29] , \wRegInA18[17] , 
        \wRegInA78[13] , \wRegInB43[3] , \wRegInA101[9] , \wRegInB0[0] , 
        \wRegInB26[15] , \wRegInA83[12] , \wRegInB53[25] , \wBIn2[24] , 
        \wBMid18[20] , \wBMid21[4] , \wRegInB10[10] , \wRegInA20[5] , 
        \wRegInB70[14] , \wRegInB33[21] , \wRegInB40[0] , \wRegInB65[20] , 
        \wRegInB46[11] , \wRegInA96[26] , \ScanLink239[21] , \ScanLink223[9] , 
        \ScanLink64[24] , \ScanLink11[14] , \wBMid78[24] , \wAMid117[5] , 
        \ScanLink47[15] , \wAIn114[12] , \ScanLink32[25] , \ScanLink52[21] , 
        \wBMid46[3] , \wAIn87[23] , \wAIn101[26] , \wAIn122[17] , 
        \wRegInB92[6] , \ScanLink189[12] , \ScanLink60[1] , \ScanLink27[11] , 
        \ScanLink71[10] , \wAIn92[17] , \wBMid94[5] , \wRegInA18[24] , 
        \ScanLink3[29] , \wRegInB27[7] , \wRegInA47[2] , \ScanLink3[30] , 
        \wRegInA78[20] , \wRegInB100[18] , \wRegInB123[30] , \ScanLink172[20] , 
        \ScanLink107[10] , \wAIn72[8] , \wRegInB1[31] , \wBMid83[16] , 
        \wBMid96[22] , \wRegInB1[28] , \wRegInA95[4] , \wRegInB123[29] , 
        \ScanLink151[11] , \ScanLink139[4] , \ScanLink124[21] , 
        \ScanLink144[25] , \ScanLink131[15] , \wAMid12[19] , \wBIn14[8] , 
        \wBMid18[13] , \wAIn101[15] , \ScanLink167[14] , \ScanLink112[24] , 
        \wRegInA96[7] , \ScanLink52[12] , \ScanLink27[22] , \wAMid31[28] , 
        \wBMid45[0] , \wAIn122[24] , \wBMid78[17] , \ScanLink239[12] , 
        \ScanLink189[21] , \ScanLink71[23] , \ScanLink64[17] , 
        \ScanLink11[27] , \wAIn114[21] , \ScanLink32[16] , \wRegInA44[1] , 
        \ScanLink47[26] , \wRegInB65[13] , \wRegInB10[23] , \wAMid44[18] , 
        \wAMid67[30] , \wRegInB46[22] , \ScanLink127[8] , \wAMid31[31] , 
        \wAMid67[29] , \wBMid97[6] , \wRegInB33[12] , \wRegInA96[15] , 
        \wAIn69[16] , \wRegInB24[4] , \wRegInB53[16] , \wRegInB26[26] , 
        \wRegInA83[21] , \wRegInB70[27] , \wAIn0[31] , \wBIn1[1] , \wBIn2[2] , 
        \wBMid1[25] , \wAIn4[19] , \wBIn9[31] , \wAIn10[2] , \wBMid24[9] , 
        \wAMid50[6] , \wRegInA45[30] , \wAMid97[24] , \wRegInA66[18] , 
        \ScanLink8[25] , \wBIn98[23] , \wAMid112[8] , \wAMid125[22] , 
        \wRegInA13[28] , \wRegInA38[7] , \wRegInA45[29] , \wBMid39[6] , 
        \wAMid82[10] , \wAMid106[13] , \wRegInA13[31] , \wRegInA30[19] , 
        \ScanLink194[7] , \wAMid113[27] , \wAMid82[0] , \wRegInB58[2] , 
        \wBIn75[1] , \wRegInA25[8] , \ScanLink189[8] , \ScanLink146[1] , 
        \wBIn9[28] , \wRegInA107[7] , \ScanLink119[31] , \ScanLink78[3] , 
        \wBIn76[2] , \ScanLink226[4] , \ScanLink145[2] , \ScanLink119[28] , 
        \wAMid81[3] , \wRegInB89[7] , \wRegInA113[11] , \wRegInA104[4] , 
        \wRegInA106[25] , \ScanLink225[7] , \ScanLink197[19] , \wAIn13[1] , 
        \wRegInA125[14] , \wBIn16[12] , \wAMid19[15] , \wBIn35[23] , 
        \wBIn40[13] , \wBIn123[22] , \ScanLink197[4] , \wAMid53[5] , 
        \wBIn20[17] , \wBIn63[22] , \wBIn100[13] , \wBIn76[16] , 
        \wRegInB94[8] , \wAMid79[11] , \wBIn115[27] , \ScanLink238[8] , 
        \wBIn55[27] , \wAIn69[9] , \wBMid88[29] , \ScanLink122[5] , 
        \ScanLink94[30] , \wBMid1[16] , \wBIn11[5] , \wBIn12[6] , \wBIn16[21] , 
        \wAIn17[19] , \wAIn34[31] , \wAMid34[2] , \wAIn74[6] , \wBMid88[30] , 
        \wAIn120[2] , \wAMid113[14] , \wRegInB21[9] , \ScanLink94[29] , 
        \ScanLink242[0] , \wAIn99[31] , \wRegInB80[19] , \wAMid37[1] , 
        \wAIn62[29] , \wAMid82[23] , \wAIn99[28] , \wAMid97[17] , 
        \wBMid104[0] , \wAMid125[11] , \ScanLink8[16] , \wBIn98[10] , 
        \wAMid106[20] , \wBIn76[25] , \wAMid79[22] , \wBIn115[14] , 
        \wBMid107[3] , \wAMid19[26] , \wBIn20[24] , \wAIn34[28] , \wAIn41[18] , 
        \wBIn55[14] , \wAIn62[30] , \wRegInB58[29] , \wAIn77[5] , 
        \wRegInA90[9] , \wBIn35[10] , \wBIn40[20] , \wBIn123[11] , 
        \wRegInB58[30] , \wBIn63[11] , \wBIn100[20] , \wBMid25[30] , 
        \wBMid25[29] , \wRegInA106[16] , \wBMid50[19] , \wBMid73[31] , 
        \ScanLink39[30] , \wBMid91[8] , \wRegInA125[27] , \wAIn123[1] , 
        \ScanLink39[29] , \wBMid73[28] , \ScanLink121[6] , \wBMid5[27] , 
        \wBIn12[10] , \wAIn13[31] , \wAIn13[28] , \wRegInA113[22] , 
        \ScanLink252[30] , \ScanLink204[28] , \ScanLink227[19] , 
        \ScanLink204[31] , \ScanLink252[29] , \ScanLink241[3] , \wAIn45[30] , 
        \wRegInB115[4] , \wAIn66[18] , \wBIn72[14] , \wBIn111[25] , 
        \wRegInB29[28] , \wBIn24[15] , \wAIn30[19] , \wBIn31[21] , 
        \wAIn45[29] , \wBIn51[25] , \wAIn53[3] , \wRegInB29[31] , \wBIn44[11] , 
        \wBIn127[20] , \wAMid13[7] , \wBMid21[18] , \wBMid54[28] , 
        \wBIn67[20] , \wBMid67[8] , \wBIn104[11] , \wBMid123[5] , 
        \wAMid68[27] , \wBMid77[19] , \wRegInA102[27] , \ScanLink48[31] , 
        \wAMid10[4] , \wBIn35[3] , \wBIn36[0] , \wBMid54[31] , \wAIn81[5] , 
        \wRegInA121[16] , \ScanLink48[28] , \wAIn107[7] , \wRegInA66[9] , 
        \ScanLink223[31] , \ScanLink200[19] , \ScanLink105[0] , \wBMid79[4] , 
        \wRegInA8[23] , \wRegInA117[13] , \ScanLink256[18] , \ScanLink223[28] , 
        \ScanLink90[18] , \ScanLink38[1] , \wAIn82[6] , \wAIn104[4] , 
        \wAMid86[12] , \wBIn89[15] , \wAMid117[25] , \ScanLink106[3] , 
        \wRegInB84[28] , \wRegInB18[0] , \wRegInB84[31] , \wRegInB116[7] , 
        \wAIn50[0] , \wAMid93[26] , \wBMid120[6] , \wAMid121[20] , 
        \wRegInA78[5] , \wAMid102[11] , \wRegInA120[2] , \wAIn0[28] , 
        \wRegInB62[8] , \wRegInA117[20] , \wBIn6[26] , \wBIn6[15] , 
        \wBMid5[14] , \wBIn52[4] , \wRegInA102[14] , \ScanLink201[1] , 
        \wRegInA121[25] , \ScanLink193[28] , \ScanLink193[31] , \wBIn12[23] , 
        \wBIn31[12] , \wBIn44[22] , \wBIn127[13] , \wRegInA99[31] , 
        \ScanLink161[4] , \ScanLink42[9] , \wBIn67[13] , \wAMid68[14] , 
        \wBIn104[22] , \wRegInA99[28] , \ScanLink3[5] , \wAMid15[9] , 
        \wBIn24[26] , \wAIn37[7] , \wBIn51[16] , \wBIn72[27] , \wAMid77[3] , 
        \wBIn111[16] , \wAIn34[4] , \wBIn80[2] , \wAMid93[15] , \wAMid121[13] , 
        \wRegInA17[19] , \wRegInA34[31] , \ScanLink0[6] , \wRegInA62[29] , 
        \wAMid102[22] , \wRegInA34[28] , \wAMid117[16] , \wRegInA41[18] , 
        \wRegInA62[30] , \wBIn51[7] , \wAMid74[0] , \wBIn83[1] , \wBIn109[0] , 
        \wAMid86[21] , \wBIn89[26] , \wRegInA123[1] , \ScanLink202[2] , 
        \ScanLink168[30] , \ScanLink162[7] , \wBMid69[12] , \wAIn105[24] , 
        \wRegInA8[10] , \ScanLink168[29] , \ScanLink56[23] , \ScanLink20[3] , 
        \ScanLink23[13] , \wAIn126[15] , \ScanLink228[17] , \ScanLink75[12] , 
        \wRegInA109[18] , \ScanLink198[24] , \ScanLink60[26] , \wAMid16[31] , 
        \wAMid35[19] , \wAMid40[29] , \wBMid61[6] , \ScanLink15[16] , 
        \wAIn110[10] , \ScanLink248[13] , \ScanLink43[17] , \ScanLink36[27] , 
        \wRegInB14[12] , \wRegInB61[22] , \wAMid16[28] , \wAMid40[30] , 
        \wAMid63[18] , \wRegInB37[23] , \wRegInA92[24] , \wAIn78[13] , 
        \wRegInB42[13] , \wAIn18[17] , \wRegInB22[17] , \wRegInA87[10] , 
        \wAIn48[2] , \wRegInB57[27] , \wAIn83[12] , \wAMid98[19] , 
        \wAIn101[9] , \wRegInA60[7] , \wRegInA69[25] , \wRegInB74[16] , 
        \ScanLink7[18] , \wAIn84[8] , \wBMid87[27] , \wBMid92[13] , 
        \wAIn96[26] , \wRegInA63[4] , \wRegInB127[18] , \wRegInB104[30] , 
        \wRegInB104[29] , \wRegInB110[9] , \ScanLink103[21] , 
        \ScanLink176[11] , \ScanLink120[10] , \wRegInB5[19] , 
        \ScanLink155[20] , \ScanLink23[0] , \wAIn99[7] , \ScanLink140[14] , 
        \ScanLink135[24] , \ScanLink116[15] , \wAIn18[24] , \wBMid62[5] , 
        \wBMid126[8] , \ScanLink163[25] , \wAIn31[9] , \wAIn78[20] , 
        \wBIn79[18] , \wRegInB57[14] , \wRegInB64[6] , \wBIn111[2] , 
        \wRegInB22[24] , \wRegInA87[23] , \wRegInB74[25] , \ScanLink96[1] , 
        \ScanLink59[8] , \wRegInB14[21] , \wRegInB61[11] , \wRegInB37[10] , 
        \wRegInB42[20] , \wRegInA92[17] , \wAIn105[17] , \wAIn110[23] , 
        \wRegInB79[9] , \ScanLink15[25] , \ScanLink248[20] , \ScanLink198[17] , 
        \ScanLink60[15] , \ScanLink36[14] , \ScanLink44[7] , \ScanLink43[24] , 
        \wBIn49[5] , \wBMid69[21] , \ScanLink23[20] , \wBMid87[14] , 
        \wAIn126[26] , \ScanLink56[10] , \wRegInA9[9] , \ScanLink228[24] , 
        \ScanLink140[27] , \ScanLink75[21] , \ScanLink135[17] , 
        \ScanLink47[4] , \ScanLink6[8] , \wAIn8[3] , \wBIn82[19] , 
        \wBMid92[20] , \ScanLink219[3] , \ScanLink163[16] , \ScanLink116[26] , 
        \ScanLink179[6] , \ScanLink176[22] , \ScanLink155[13] , 
        \ScanLink103[12] , \ScanLink120[23] , \wBMid105[18] , \wBMid126[29] , 
        \ScanLink95[2] , \wAIn83[21] , \wAIn96[15] , \wBMid126[30] , 
        \wRegInB67[5] , \wRegInA69[16] , \wAMid12[31] , \wBMid18[22] , 
        \wBIn57[9] , \wBIn98[0] , \wBIn112[1] , \ScanLink164[9] , 
        \wAIn101[24] , \ScanLink60[3] , \ScanLink27[13] , \wBMid21[6] , 
        \wAIn122[15] , \ScanLink52[23] , \wRegInB92[4] , \ScanLink189[10] , 
        \ScanLink71[12] , \ScanLink11[16] , \wAMid55[9] , \ScanLink64[26] , 
        \wBMid78[26] , \ScanLink239[23] , \ScanLink32[27] , \wAIn114[10] , 
        \wAMid117[7] , \ScanLink191[8] , \wRegInB65[22] , \ScanLink47[17] , 
        \wAMid12[28] , \wAMid31[19] , \wAMid44[29] , \wRegInB10[12] , 
        \wRegInA102[8] , \wRegInB46[13] , \wAMid44[30] , \wRegInB33[23] , 
        \wRegInA96[24] , \wRegInB40[2] , \wAMid48[6] , \wAMid67[18] , 
        \wAIn69[27] , \wRegInB0[2] , \wRegInB53[27] , \wRegInB26[17] , 
        \wRegInA83[10] , \wRegInB70[16] , \wBIn2[15] , \wBMid22[5] , 
        \wBMid83[27] , \wAIn87[12] , \wRegInA20[7] , \ScanLink220[8] , 
        \wAIn92[26] , \wRegInA18[15] , \ScanLink3[18] , \wRegInA23[4] , 
        \wRegInB43[1] , \wBMid96[13] , \wRegInB3[1] , \wRegInA78[11] , 
        \wRegInB91[7] , \wRegInB100[29] , \ScanLink172[11] , \ScanLink107[21] , 
        \wRegInB100[30] , \wRegInB123[18] , \ScanLink151[20] , 
        \ScanLink124[10] , \ScanLink63[0] , \wRegInB1[19] , \ScanLink144[14] , 
        \wAMid114[4] , \ScanLink131[24] , \wAIn69[14] , \wAMid99[3] , 
        \ScanLink167[25] , \ScanLink112[15] , \wRegInB24[6] , \wRegInB26[24] , 
        \wRegInB53[14] , \wRegInA83[23] , \wAIn0[19] , \wBIn1[3] , \wBIn2[26] , 
        \wBMid18[11] , \wBMid78[15] , \wBMid97[4] , \wRegInB10[21] , 
        \wRegInB70[25] , \ScanLink19[8] , \wRegInB33[10] , \wRegInA44[3] , 
        \wRegInB65[11] , \wRegInA96[17] , \wRegInB39[9] , \wRegInB46[20] , 
        \ScanLink239[10] , \ScanLink64[15] , \ScanLink11[25] , 
        \ScanLink47[24] , \ScanLink32[14] , \wAIn114[23] , \wBMid45[2] , 
        \wAIn71[9] , \wAIn101[17] , \ScanLink52[10] , \wRegInA96[5] , 
        \ScanLink27[20] , \ScanLink189[23] , \wBMid83[14] , \wAIn122[26] , 
        \ScanLink71[21] , \ScanLink144[27] , \ScanLink131[17] , 
        \ScanLink112[26] , \wBMid1[27] , \wAIn13[3] , \wAIn17[31] , 
        \wAIn17[28] , \wBIn17[9] , \wBMid46[1] , \wBMid89[8] , 
        \ScanLink167[16] , \ScanLink107[12] , \wBIn86[19] , \wAIn92[15] , 
        \wBMid96[20] , \ScanLink172[22] , \ScanLink139[6] , \ScanLink124[23] , 
        \wAMid118[30] , \wAMid118[29] , \wRegInA95[6] , \ScanLink151[13] , 
        \wBMid122[29] , \wBMid122[30] , \wBMid101[18] , \wRegInB27[5] , 
        \wAIn87[21] , \wBMid94[7] , \wRegInA78[22] , \wRegInA18[26] , 
        \ScanLink124[9] , \wAIn41[30] , \wAIn62[18] , \wRegInA47[0] , 
        \wRegInA88[9] , \wBIn76[14] , \wAMid79[13] , \wBIn115[25] , 
        \wAIn34[19] , \wAIn41[29] , \wBIn55[25] , \wRegInB58[18] , 
        \wRegInA119[9] , \wBIn20[15] , \wBIn40[11] , \wBIn123[20] , 
        \ScanLink197[6] , \wBIn16[10] , \wBMid27[8] , \wBIn35[21] , 
        \wAMid111[9] , \wBIn63[20] , \wBIn100[11] , \wAMid19[17] , 
        \wAMid53[7] , \wBMid25[18] , \wRegInA106[27] , \wBMid50[31] , 
        \wBMid50[28] , \ScanLink225[5] , \wRegInB89[5] , \wRegInA125[16] , 
        \wBMid1[14] , \wAIn4[31] , \wAIn10[0] , \wBMid39[4] , \wBMid73[19] , 
        \wBIn76[0] , \wRegInA104[6] , \ScanLink227[31] , \ScanLink204[19] , 
        \ScanLink39[18] , \ScanLink145[0] , \wAMid81[1] , \wRegInA26[9] , 
        \wRegInA113[13] , \ScanLink227[28] , \ScanLink252[18] , \wBMid88[18] , 
        \wRegInA107[5] , \ScanLink78[1] , \ScanLink226[6] , \ScanLink94[18] , 
        \wAMid50[4] , \wBIn75[3] , \wAMid82[2] , \wAMid82[12] , \wAIn99[19] , 
        \wAMid113[25] , \ScanLink146[3] , \wRegInB80[31] , \wRegInB80[28] , 
        \wRegInB97[9] , \wAMid125[20] , \wRegInB58[0] , \wAMid97[26] , 
        \wBIn98[21] , \wAMid106[11] , \ScanLink194[5] , \ScanLink8[27] , 
        \wRegInA38[5] , \wAIn4[28] , \ScanLink241[1] , \wBMid8[8] , 
        \wRegInB22[8] , \wRegInA113[20] , \wRegInA106[14] , \ScanLink197[28] , 
        \wBIn12[4] , \wAIn123[3] , \wBIn2[0] , \wBIn16[23] , \wBIn35[12] , 
        \wRegInA125[25] , \ScanLink121[4] , \ScanLink197[31] , \wBIn40[22] , 
        \wBIn123[13] , \wAMid19[24] , \wBIn20[26] , \wAMid37[3] , \wBIn63[13] , 
        \wBIn100[22] , \wAMid79[20] , \wBMid107[1] , \wBIn76[27] , 
        \wBIn115[16] , \wAMid34[0] , \wBIn55[16] , \wAIn74[4] , \wAIn77[7] , 
        \wAMid97[15] , \wBIn98[12] , \wRegInA66[29] , \wAMid106[22] , 
        \wAMid125[13] , \wRegInA13[19] , \ScanLink8[14] , \wRegInA30[31] , 
        \wRegInA30[28] , \wRegInA45[18] , \wRegInA66[30] , \wRegInA93[8] , 
        \wAMid82[21] , \wAMid113[16] , \wBMid104[2] , \ScanLink242[2] , 
        \wBIn9[19] , \wBIn11[7] , \wAIn120[0] , \ScanLink122[7] , \wBMid92[9] , 
        \wAMid10[6] , \wBMid64[9] , \ScanLink119[19] , \wBMid120[4] , 
        \wAMid121[22] , \wRegInA17[28] , \wRegInA41[30] , \wRegInA62[18] , 
        \wBIn35[1] , \wAIn50[2] , \wAMid93[24] , \wAMid102[13] , \wAIn119[9] , 
        \wRegInA34[19] , \wRegInA17[31] , \wRegInA41[29] , \wRegInA78[7] , 
        \wBMid79[6] , \wAMid86[10] , \wAMid117[27] , \wBIn89[17] , 
        \wRegInB18[2] , \wRegInB116[5] , \wBIn36[2] , \wAIn82[4] , 
        \wAIn104[6] , \wRegInA65[8] , \ScanLink106[1] , \wRegInA8[21] , 
        \ScanLink38[3] , \ScanLink168[18] , \ScanLink105[2] , \wAIn81[7] , 
        \wAIn107[5] , \wRegInA117[11] , \wAIn0[9] , \wAIn1[20] , \wBIn6[24] , 
        \wBIn6[17] , \wBMid5[25] , \wRegInA102[25] , \wRegInB108[9] , 
        \ScanLink193[19] , \wRegInA121[14] , \wBMid5[16] , \wBIn12[21] , 
        \wBIn12[12] , \wAMid13[5] , \wBIn31[23] , \wBIn44[13] , \wBIn127[22] , 
        \wAIn53[1] , \wBIn67[22] , \wBIn104[13] , \wRegInA99[19] , 
        \wAMid68[25] , \wBMid123[7] , \wAIn13[19] , \wBIn24[17] , \wBIn51[27] , 
        \wBIn72[16] , \wBIn111[27] , \wRegInB115[6] , \wAIn29[9] , \wBIn51[5] , 
        \ScanLink162[5] , \ScanLink90[30] , \wAIn34[6] , \wBIn83[3] , 
        \wRegInA8[12] , \ScanLink90[29] , \wRegInB61[9] , \ScanLink202[0] , 
        \wRegInA123[3] , \wAMid74[2] , \wAMid86[23] , \wBIn109[2] , 
        \wAMid117[14] , \wRegInB84[19] , \wBIn89[24] , \wAMid93[17] , 
        \wAMid102[20] , \wAMid121[11] , \ScanLink0[4] , \ScanLink41[8] , 
        \wBIn24[24] , \wAIn30[31] , \wAIn66[29] , \wBIn72[25] , \wAMid77[1] , 
        \wBIn111[14] , \wRegInB29[19] , \wAIn30[28] , \wBIn31[10] , 
        \wAIn37[5] , \wAIn45[18] , \wBIn80[0] , \wBIn51[14] , \wAIn66[30] , 
        \wBIn44[20] , \wBIn127[11] , \wBMid21[29] , \wBMid54[19] , 
        \wBIn67[11] , \wBIn104[20] , \ScanLink3[7] , \wAMid68[16] , 
        \wBMid77[31] , \wBMid77[28] , \wRegInA102[16] , \wBMid21[30] , 
        \wBIn52[6] , \ScanLink161[6] , \wBMid62[7] , \wBMid87[25] , 
        \wAIn99[5] , \wRegInA117[22] , \wRegInA120[0] , \wRegInA121[27] , 
        \ScanLink256[30] , \ScanLink48[19] , \ScanLink200[28] , 
        \ScanLink256[29] , \ScanLink201[3] , \ScanLink223[19] , 
        \ScanLink200[31] , \ScanLink140[16] , \ScanLink135[26] , \wAIn8[1] , 
        \wAMid16[8] , \ScanLink163[27] , \wAIn18[15] , \wBIn82[31] , 
        \wBMid92[11] , \ScanLink176[13] , \ScanLink116[17] , \ScanLink155[22] , 
        \ScanLink103[23] , \ScanLink120[12] , \ScanLink23[2] , \wBIn82[28] , 
        \wAIn102[8] , \wBMid105[30] , \wBMid126[18] , \wRegInA63[6] , 
        \wAIn83[10] , \wAIn96[24] , \wBMid105[29] , \wRegInA69[27] , 
        \wAIn48[0] , \wBIn79[29] , \wRegInB57[25] , \wRegInB22[15] , 
        \wRegInB74[14] , \wRegInA87[12] , \wBMid61[4] , \wAIn78[11] , 
        \wBIn79[30] , \wAIn87[9] , \wRegInA60[5] , \wRegInB14[10] , 
        \wRegInB61[20] , \wRegInB37[21] , \wRegInB42[11] , \wRegInA92[26] , 
        \wBMid125[9] , \ScanLink15[14] , \ScanLink248[11] , \wBMid69[10] , 
        \wAIn105[26] , \wAIn110[12] , \ScanLink198[26] , \ScanLink60[24] , 
        \ScanLink36[25] , \ScanLink43[15] , \ScanLink20[1] , \wAIn126[17] , 
        \ScanLink56[21] , \ScanLink23[11] , \wRegInB113[8] , \ScanLink228[15] , 
        \ScanLink75[10] , \wAIn32[8] , \wAIn83[23] , \wAMid98[28] , 
        \wRegInA69[14] , \ScanLink7[29] , \wBMid92[22] , \wAIn96[17] , 
        \wBIn98[2] , \wAMid98[31] , \ScanLink7[30] , \wBIn112[3] , 
        \wRegInB67[7] , \ScanLink95[0] , \wRegInB127[30] , \wRegInB104[18] , 
        \ScanLink103[10] , \wRegInB127[29] , \wRegInB5[31] , \ScanLink176[20] , 
        \wRegInB5[28] , \ScanLink179[4] , \ScanLink120[21] , \wBMid87[16] , 
        \ScanLink155[11] , \ScanLink47[6] , \ScanLink219[1] , 
        \ScanLink140[25] , \ScanLink135[15] , \ScanLink116[24] , \wAMid16[19] , 
        \wAMid35[31] , \wAMid35[28] , \wAMid40[18] , \wBIn49[7] , 
        \ScanLink163[14] , \wBIn54[8] , \wBMid69[23] , \wAIn105[15] , 
        \ScanLink56[12] , \wAIn110[21] , \wAIn126[24] , \ScanLink228[26] , 
        \ScanLink23[22] , \ScanLink75[23] , \wRegInA109[30] , \wRegInA109[29] , 
        \ScanLink248[22] , \ScanLink198[15] , \ScanLink60[17] , 
        \ScanLink15[27] , \ScanLink5[9] , \ScanLink43[26] , \ScanLink44[5] , 
        \ScanLink36[16] , \wAMid63[30] , \wRegInB14[23] , \ScanLink167[8] , 
        \wBIn111[0] , \wRegInB61[13] , \wAMid63[29] , \wRegInB37[12] , 
        \wRegInA92[15] , \wAIn78[22] , \wRegInB42[22] , \wAIn18[26] , 
        \wRegInB22[26] , \wRegInA87[21] , \wBMid20[23] , \wBMid55[13] , 
        \wBMid76[22] , \wRegInB57[16] , \wRegInB64[4] , \wRegInB74[27] , 
        \ScanLink96[3] , \wBIn107[4] , \wRegInA12[5] , \ScanLink49[13] , 
        \ScanLink214[16] , \ScanLink242[17] , \wRegInA2[0] , \ScanLink237[27] , 
        \ScanLink192[20] , \ScanLink211[9] , \wAMid5[24] , \wBMid35[17] , 
        \wBMid40[27] , \ScanLink222[13] , \ScanLink187[14] , \wBMid63[16] , 
        \wRegInB72[0] , \wRegInA116[28] , \ScanLink80[7] , \ScanLink29[17] , 
        \wAIn12[13] , \wBMid16[26] , \wRegInA116[31] , \ScanLink201[22] , 
        \wAIn31[22] , \wAIn44[12] , \wAMid125[5] , \wBMid13[4] , \wAIn1[13] , 
        \wBMid10[7] , \wAIn24[16] , \wAIn67[23] , \wAIn72[17] , 
        \wRegInB28[13] , \wRegInB48[17] , \wRegInA98[20] , \ScanLink52[1] , 
        \wAIn51[26] , \wAMid87[29] , \wAIn12[20] , \wBIn13[18] , \wAIn39[3] , 
        \wAMid64[8] , \wRegInA76[15] , \wAMid79[7] , \wAMid87[30] , 
        \wBIn93[9] , \wAIn89[16] , \wBIn119[8] , \wAMid126[6] , 
        \wRegInA55[24] , \wRegInA20[14] , \wRegInA35[20] , \wRegInA40[10] , 
        \wRegInB85[13] , \ScanLink51[2] , \wRegInB90[27] , \wRegInA63[21] , 
        \wRegInA1[3] , \wRegInA9[18] , \wRegInA16[11] , \ScanLink169[21] , 
        \ScanLink91[23] , \wBIn66[28] , \wAIn72[24] , \wBMid77[0] , 
        \wBMid98[17] , \wBIn104[7] , \wRegInA11[6] , \ScanLink83[4] , 
        \wBIn105[19] , \wBIn126[31] , \wRegInB71[3] , \ScanLink84[17] , 
        \ScanLink109[25] , \wRegInA98[13] , \wRegInB48[24] , \wAIn24[25] , 
        \wBIn30[30] , \wBIn45[19] , \wBIn126[28] , \ScanLink108[7] , 
        \wAIn51[15] , \wBIn66[31] , \wBIn30[29] , \wAIn31[11] , \wAIn44[21] , 
        \ScanLink36[5] , \wAIn67[10] , \wRegInB28[20] , \wBMid35[24] , 
        \ScanLink222[20] , \ScanLink187[27] , \wAIn5[4] , \wAMid5[17] , 
        \wBMid16[15] , \wBMid40[14] , \ScanLink201[11] , \ScanLink115[8] , 
        \wBIn26[8] , \wAIn6[7] , \wAMid17[13] , \wBMid20[10] , \wBMid63[25] , 
        \wBMid76[11] , \wRegInA76[1] , \ScanLink29[24] , \ScanLink214[25] , 
        \ScanLink49[20] , \wBIn38[4] , \wBMid55[20] , \wRegInB16[4] , 
        \wRegInB118[3] , \ScanLink237[14] , \ScanLink192[13] , \wBMid98[24] , 
        \ScanLink242[24] , \wRegInB15[7] , \wRegInA75[2] , \ScanLink169[12] , 
        \ScanLink109[16] , \ScanLink91[10] , \ScanLink84[24] , \ScanLink28[9] , 
        \wAIn40[8] , \wAMid103[19] , \wAIn109[3] , \wRegInA35[13] , 
        \wRegInB90[14] , \wAMid120[31] , \wRegInA40[23] , \wAMid62[23] , 
        \wBMid74[3] , \wRegInA16[22] , \wAIn79[28] , \wAIn89[25] , 
        \wAMid120[28] , \wRegInA63[12] , \wRegInB15[30] , \wRegInA20[27] , 
        \wRegInA76[26] , \wRegInA55[17] , \wRegInB85[20] , \ScanLink35[6] , 
        \wRegInB36[18] , \wRegInB43[28] , \wBIn18[14] , \wAMid21[16] , 
        \wAMid34[22] , \wAMid41[12] , \wBIn44[2] , \wRegInB15[29] , 
        \wAIn79[31] , \wRegInB43[31] , \ScanLink177[2] , \wRegInB60[19] , 
        \wAMid54[26] , \ScanLink86[9] , \ScanLink49[0] , \wAMid77[17] , 
        \wBIn78[10] , \ScanLink217[7] , \wAIn21[1] , \wAMid61[5] , 
        \ScanLink74[29] , \wBMid68[30] , \ScanLink22[31] , \wBIn96[4] , 
        \ScanLink57[18] , \ScanLink74[30] , \ScanLink22[28] , \wAIn22[2] , 
        \wBMid68[29] , \wBMid93[28] , \wBIn95[7] , \wRegInB69[1] , 
        \wRegInA108[23] , \ScanLink249[31] , \wRegInB126[23] , 
        \ScanLink249[28] , \wAMid120[8] , \wRegInB4[22] , \wBMid16[9] , 
        \wRegInB105[12] , \wAIn45[5] , \wBIn47[1] , \wAMid62[6] , 
        \wBMid93[31] , \wBIn88[8] , \wRegInA2[27] , \wRegInB110[26] , 
        \ScanLink98[5] , \wAMid108[15] , \ScanLink174[1] , \wAIn82[30] , 
        \wBIn102[9] , \wAIn82[29] , \wRegInA17[8] , \wBIn83[11] , \wBIn96[25] , 
        \wAMid99[22] , \ScanLink6[23] , \wBMid104[10] , \wBMid111[24] , 
        \ScanLink214[4] , \wAIn111[18] , \wRegInB103[2] , \wRegInA108[10] , 
        \wAIn0[0] , \wAIn1[30] , \wAIn1[29] , \wBMid0[0] , \wAMid17[20] , 
        \wBIn20[6] , \wAMid21[25] , \ScanLink113[6] , \wAMid54[15] , 
        \wAIn111[1] , \wAMid77[24] , \wBIn78[23] , \wAIn97[3] , 
        \wRegInA86[18] , \wBIn18[27] , \wBIn23[5] , \wAMid34[11] , 
        \wAMid62[10] , \wAMid41[21] , \wBIn83[22] , \wBMid104[23] , 
        \wAIn46[6] , \wAIn94[0] , \wAIn112[2] , \ScanLink110[5] , \wBIn96[16] , 
        \wAMid99[11] , \wAMid108[26] , \ScanLink6[10] , \wBMid111[17] , 
        \wRegInA2[14] , \wRegInB13[9] , \wRegInB110[15] , \wBIn87[13] , 
        \wRegInB4[11] , \wRegInB126[10] , \ScanLink154[28] , \ScanLink121[18] , 
        \ScanLink102[30] , \ScanLink33[8] , \wRegInB100[1] , \wRegInB105[21] , 
        \ScanLink177[19] , \ScanLink154[31] , \ScanLink102[29] , 
        \ScanLink254[6] , \wAMid88[14] , \wBMid100[12] , \wBIn92[27] , 
        \wBMid115[26] , \wAMid119[23] , \wRegInA79[28] , \wBMid123[23] , 
        \wRegInA79[31] , \wRegInA98[3] , \ScanLink134[3] , \wRegInA6[25] , 
        \ScanLink2[21] , \wRegInB114[24] , \ScanLink249[9] , \wRegInB124[7] , 
        \wAMid1[26] , \wAMid1[7] , \wBMid3[3] , \wAMid22[4] , \wAIn62[0] , 
        \wRegInB0[20] , \wRegInB122[21] , \ScanLink125[29] , \ScanLink173[31] , 
        \wBMid99[2] , \wRegInB101[10] , \ScanLink150[19] , \ScanLink125[30] , 
        \ScanLink106[18] , \wBMid112[6] , \ScanLink173[28] , \wAIn115[29] , 
        \wAMid13[11] , \wAMid21[7] , \wBMid55[8] , \wAIn115[30] , 
        \wRegInB127[4] , \wRegInB29[3] , \wBMid111[5] , \ScanLink188[29] , 
        \wRegInA119[15] , \wAMid25[14] , \wAMid50[24] , \wAIn61[3] , 
        \wRegInA49[6] , \ScanLink188[30] , \wRegInA82[30] , \wBMid48[7] , 
        \wAMid73[15] , \wRegInA82[29] , \wAMid66[21] , \wBIn69[26] , 
        \wAMid30[20] , \wAMid45[10] , \wRegInA54[9] , \ScanLink137[0] , 
        \wAMid46[0] , \wBMid97[19] , \wRegInB0[13] , \wRegInB122[12] , 
        \wRegInA6[16] , \wRegInB101[23] , \wAIn86[18] , \wAMid89[9] , 
        \wBIn92[14] , \wBMid115[15] , \wRegInA111[1] , \wRegInB114[17] , 
        \ScanLink182[1] , \ScanLink230[2] , \ScanLink2[12] , \wAMid2[4] , 
        \wBIn63[7] , \wBIn87[20] , \wAMid88[27] , \wBMid100[21] , \wAMid94[6] , 
        \wAMid119[10] , \wBMid123[10] , \ScanLink150[7] , \wAMid119[1] , 
        \wRegInB47[19] , \wRegInB64[31] , \wAIn5[22] , \wBIn8[13] , 
        \wAMid13[22] , \ScanLink233[1] , \wAIn18[8] , \wAMid25[27] , 
        \wAMid30[13] , \wAMid66[12] , \wRegInB32[29] , \wRegInB50[8] , 
        \wBIn69[15] , \wRegInB64[28] , \wAMid45[23] , \wRegInB11[18] , 
        \wRegInB32[30] , \wRegInA112[2] , \ScanLink153[4] , \wAMid50[17] , 
        \wBIn60[4] , \wBMid19[31] , \wAMid73[26] , \wAMid97[5] , 
        \ScanLink70[18] , \ScanLink53[30] , \wBMid19[28] , \wRegInA119[26] , 
        \ScanLink70[9] , \ScanLink53[29] , \ScanLink26[19] , \wAMid45[3] , 
        \ScanLink238[30] , \ScanLink181[2] , \ScanLink238[29] , \wRegInB31[1] , 
        \ScanLink252[8] , \ScanLink178[17] , \ScanLink80[15] , \wAIn16[11] , 
        \wBIn17[30] , \wBIn17[29] , \wAMid39[5] , \wBMid82[3] , \wBMid109[7] , 
        \ScanLink95[21] , \wBMid50[5] , \wAIn79[1] , \wBMid89[21] , 
        \ScanLink118[13] , \wAIn98[20] , \wBIn99[18] , \wAMid107[28] , 
        \wRegInA31[22] , \wRegInA44[12] , \wRegInA51[4] , \ScanLink11[0] , 
        \wRegInB94[25] , \wRegInA67[23] , \wAMid107[31] , \wAMid124[19] , 
        \wRegInA12[13] , \wRegInB122[9] , \wBMid114[8] , \wRegInA72[17] , 
        \wRegInA24[16] , \wRegInA51[26] , \wRegInA83[2] , \wRegInB81[11] , 
        \wAIn20[14] , \wBIn34[18] , \wBIn41[31] , \wBIn62[19] , \wBIn101[28] , 
        \wRegInB39[25] , \wAIn76[15] , \ScanLink12[3] , \wAIn35[20] , 
        \wBIn41[28] , \wAIn55[24] , \wBIn101[31] , \wBIn122[19] , \wAIn40[10] , 
        \wBMid53[6] , \wRegInA80[1] , \wAMid27[9] , \wAIn63[21] , 
        \wRegInB59[21] , \wRegInA89[16] , \wBMid31[15] , \wBMid44[25] , 
        \ScanLink253[21] , \wRegInB32[2] , \ScanLink226[11] , 
        \ScanLink183[16] , \wBMid67[14] , \wAMid1[15] , \wAIn5[11] , 
        \wAMid7[9] , \wBMid12[24] , \ScanLink205[20] , \wBMid24[21] , 
        \wBMid51[11] , \wBMid72[20] , \ScanLink58[25] , \ScanLink38[21] , 
        \wRegInA52[7] , \ScanLink210[14] , \wBMid81[0] , \ScanLink246[15] , 
        \wBMid34[1] , \wBIn78[6] , \wAMid83[18] , \ScanLink233[25] , 
        \ScanLink196[22] , \wAIn98[13] , \wRegInB87[3] , \wRegInA24[25] , 
        \wRegInA72[24] , \wRegInA51[15] , \wRegInB81[22] , \ScanLink75[4] , 
        \wAMid102[0] , \wRegInA31[11] , \wRegInB94[16] , \wRegInA44[21] , 
        \wRegInA12[20] , \wRegInA67[10] , \ScanLink118[20] , \wBIn8[20] , 
        \ScanLink95[12] , \wBMid24[12] , \wBIn65[9] , \wBMid89[12] , 
        \wRegInB55[5] , \ScanLink199[0] , \wBMid72[13] , \wAMid92[8] , 
        \wBIn120[1] , \ScanLink156[9] , \wRegInA35[0] , \ScanLink178[24] , 
        \ScanLink210[27] , \ScanLink80[26] , \ScanLink38[12] , \wBMid31[26] , 
        \wBMid51[22] , \ScanLink233[16] , \ScanLink196[11] , \wRegInB56[6] , 
        \wRegInA112[19] , \ScanLink246[26] , \ScanLink226[22] , 
        \ScanLink183[25] , \wBMid12[17] , \wBMid44[16] , \ScanLink253[12] , 
        \ScanLink205[13] , \wBIn123[2] , \ScanLink58[16] , \wBMid4[26] , 
        \wBIn7[27] , \wBIn7[14] , \wAIn16[22] , \wAIn35[13] , \wAIn40[23] , 
        \wBMid67[27] , \wRegInA36[3] , \wRegInA109[3] , \ScanLink76[7] , 
        \wAIn63[12] , \wAMid78[19] , \wRegInA89[25] , \ScanLink228[0] , 
        \wAMid17[30] , \wAMid17[29] , \wAIn20[27] , \wBMid37[2] , \wAIn76[26] , 
        \wRegInB39[16] , \wRegInB59[12] , \wRegInB84[0] , \wAIn55[17] , 
        \ScanLink148[5] , \wAMid101[3] , \wBMid68[13] , \wAIn104[25] , 
        \wAIn127[14] , \ScanLink229[16] , \ScanLink74[13] , \ScanLink30[2] , 
        \wBMid71[7] , \wAIn111[11] , \ScanLink57[22] , \ScanLink22[12] , 
        \ScanLink37[26] , \ScanLink249[12] , \ScanLink42[16] , 
        \ScanLink14[17] , \wRegInB43[12] , \wRegInA108[19] , \ScanLink61[27] , 
        \ScanLink199[25] , \wAMid41[31] , \wRegInB10[3] , \wRegInB36[22] , 
        \wRegInA93[25] , \wAMid62[19] , \wAIn79[12] , \wRegInB60[23] , 
        \wAMid18[7] , \wAIn19[16] , \wAMid34[18] , \wAMid41[28] , 
        \wRegInB15[13] , \wAIn58[3] , \wAIn111[8] , \wRegInB75[17] , 
        \wRegInA70[6] , \wRegInB23[16] , \wRegInB56[26] , \wRegInA86[11] , 
        \wBMid72[4] , \wAIn82[13] , \wRegInA68[24] , \wAIn94[9] , \wAIn97[27] , 
        \wAMid99[18] , \ScanLink6[19] , \wRegInB13[0] , \wBMid93[12] , 
        \wRegInB4[18] , \wRegInA73[5] , \wRegInB105[31] , \wRegInB126[19] , 
        \ScanLink154[21] , \ScanLink33[1] , \ScanLink121[11] , \wRegInB100[8] , 
        \wRegInB105[28] , \ScanLink177[10] , \ScanLink102[20] , \wBMid15[3] , 
        \wAIn19[25] , \wBIn78[19] , \wBMid86[26] , \wAIn89[6] , 
        \ScanLink162[24] , \ScanLink141[15] , \ScanLink117[14] , 
        \wRegInB75[24] , \ScanLink134[25] , \ScanLink86[0] , \ScanLink49[9] , 
        \wRegInB23[25] , \wRegInA86[22] , \wAIn79[21] , \wRegInB36[11] , 
        \wRegInB56[15] , \wRegInB74[7] , \ScanLink8[5] , \wRegInA93[16] , 
        \wBIn101[3] , \wRegInA4[7] , \wRegInB43[21] , \wRegInA14[2] , 
        \wRegInB15[20] , \wRegInB60[10] , \wAIn111[22] , \ScanLink54[6] , 
        \ScanLink42[25] , \ScanLink37[15] , \wRegInB69[8] , \ScanLink249[21] , 
        \ScanLink199[16] , \ScanLink61[14] , \ScanLink14[24] , \wAIn21[8] , 
        \wBIn59[4] , \wAIn127[27] , \ScanLink229[25] , \ScanLink74[20] , 
        \wBMid68[20] , \wAIn104[16] , \ScanLink57[11] , \wAMid123[2] , 
        \ScanLink22[21] , \ScanLink209[2] , \ScanLink117[27] , \wAIn12[30] , 
        \wBMid16[0] , \wBMid86[15] , \ScanLink162[17] , \ScanLink57[5] , 
        \wBMid93[21] , \ScanLink169[7] , \ScanLink141[26] , \ScanLink134[16] , 
        \ScanLink121[22] , \wAMid120[1] , \ScanLink154[12] , \ScanLink102[13] , 
        \wBIn25[14] , \wAIn31[18] , \wAIn44[28] , \wBIn47[8] , \wBIn83[18] , 
        \wAIn97[14] , \wRegInB77[4] , \ScanLink177[23] , \wBIn88[1] , 
        \wBMid104[19] , \ScanLink174[8] , \ScanLink85[3] , \wBIn50[24] , 
        \wAIn82[20] , \wBIn102[0] , \wRegInA17[1] , \wRegInA7[4] , 
        \wRegInA68[17] , \wRegInB28[30] , \wAIn12[29] , \wAIn44[31] , 
        \wAIn67[19] , \wBIn73[15] , \wBIn110[24] , \wRegInB28[29] , 
        \wRegInB105[5] , \wBIn13[11] , \wBIn66[21] , \wBIn105[10] , 
        \wAMid69[26] , \wBMid77[9] , \wBIn30[20] , \wAIn43[2] , \wBIn45[10] , 
        \wBIn126[21] , \wBMid55[30] , \wRegInA120[17] , \ScanLink49[29] , 
        \wBMid76[18] , \wBMid20[19] , \wRegInA103[26] , \ScanLink49[30] , 
        \wBIn25[2] , \wBIn26[1] , \wBMid55[29] , \wRegInA116[12] , 
        \ScanLink222[29] , \ScanLink222[30] , \ScanLink201[18] , 
        \ScanLink115[1] , \wAIn91[4] , \wAIn117[6] , \wRegInA9[22] , 
        \wRegInA76[8] , \ScanLink91[19] , \ScanLink28[0] , \wAIn40[1] , 
        \wBMid69[5] , \wAIn92[7] , \wAIn114[5] , \ScanLink116[2] , 
        \wAMid87[13] , \wRegInB85[30] , \wBIn88[14] , \wAMid103[10] , 
        \wAMid116[24] , \wRegInB106[6] , \wRegInB85[29] , \wRegInA68[4] , 
        \wAMid92[27] , \wAMid120[21] , \wRegInB72[9] , \wRegInA116[21] , 
        \ScanLink211[0] , \wBMid4[15] , \wBIn13[22] , \wBIn42[5] , 
        \wRegInA2[9] , \wRegInA103[15] , \wRegInA120[24] , \ScanLink171[5] , 
        \ScanLink192[30] , \ScanLink192[29] , \wBIn25[27] , \wBIn30[13] , 
        \wBIn66[12] , \wBIn105[23] , \wRegInA98[29] , \wAMid69[15] , 
        \wBIn45[23] , \wBIn126[12] , \ScanLink52[8] , \wRegInA98[30] , 
        \wAIn27[6] , \wBIn50[17] , \wBIn90[3] , \wAMid0[25] , \wBMid0[24] , 
        \wAIn3[3] , \wAMid67[2] , \wBIn73[26] , \wAMid87[20] , \wAMid92[14] , 
        \wAMid103[23] , \wBIn110[17] , \wRegInA35[29] , \wRegInA40[19] , 
        \wRegInA63[31] , \wRegInA63[28] , \wAMid120[12] , \wRegInA16[18] , 
        \wRegInA35[30] , \wAIn5[18] , \wAMid7[0] , \wAIn24[5] , \wAMid64[1] , 
        \wBIn88[27] , \wBIn93[0] , \wAMid116[17] , \wBMid29[7] , \wBMid34[8] , 
        \wBIn41[6] , \wBIn119[1] , \wRegInA9[11] , \ScanLink212[3] , 
        \ScanLink169[28] , \ScanLink172[6] , \wAMid102[9] , \wAMid107[12] , 
        \wRegInA12[30] , \wRegInA31[18] , \ScanLink169[31] , \ScanLink184[6] , 
        \wRegInA28[6] , \wRegInA44[28] , \wRegInA12[29] , \wAMid40[7] , 
        \wAMid124[23] , \wRegInA44[31] , \wRegInA67[19] , \wBIn65[0] , 
        \wAMid83[11] , \wAMid96[25] , \wBIn99[22] , \wRegInB8[3] , 
        \ScanLink9[24] , \wAMid112[26] , \wRegInB48[3] , \wBIn120[8] , 
        \wRegInA35[9] , \ScanLink199[9] , \ScanLink156[0] , \wAMid92[1] , 
        \ScanLink236[5] , \wBIn8[30] , \wBIn8[29] , \ScanLink118[29] , 
        \ScanLink118[30] , \ScanLink68[2] , \wRegInA112[10] , \wRegInA117[6] , 
        \wBIn66[3] , \wAMid91[2] , \ScanLink155[3] , \wRegInA124[15] , 
        \wBMid0[17] , \wAMid4[3] , \wRegInA107[24] , \wRegInA114[5] , 
        \wBMid5[4] , \wBMid6[7] , \wBIn17[13] , \wBIn62[23] , \wBIn101[12] , 
        \wRegInB99[6] , \ScanLink235[6] , \ScanLink196[18] , \wAMid18[14] , 
        \wBIn21[16] , \wBIn34[22] , \wBIn41[12] , \wAMid43[4] , \wBIn122[23] , 
        \ScanLink187[5] , \wBIn54[26] , \wAMid24[3] , \wBIn77[17] , 
        \wAMid78[10] , \wAIn79[8] , \wBMid89[31] , \wBIn114[26] , 
        \ScanLink228[9] , \wRegInB84[9] , \ScanLink95[28] , \ScanLink132[4] , 
        \ScanLink95[31] , \wAMid83[22] , \wBMid89[28] , \wRegInB31[8] , 
        \ScanLink252[1] , \wAIn98[29] , \wBMid114[1] , \wAIn64[7] , 
        \wAIn98[30] , \wAMid112[15] , \wAMid96[16] , \wBIn99[11] , 
        \wAMid107[21] , \wRegInB81[18] , \ScanLink11[9] , \wRegInB122[0] , 
        \ScanLink9[17] , \wAIn16[18] , \wBIn21[25] , \wAMid124[10] , 
        \wAIn35[29] , \wAIn40[19] , \wRegInB59[31] , \wBIn54[15] , 
        \wAIn63[31] , \wAIn67[4] , \wRegInA80[8] , \wBIn17[20] , \wAMid27[0] , 
        \wAIn35[30] , \wBMid117[2] , \wAMid78[23] , \wRegInB59[28] , 
        \wAIn63[28] , \wBIn77[24] , \wBIn114[15] , \wAMid18[27] , \wBIn34[11] , 
        \wBIn62[10] , \wBIn101[21] , \wRegInB121[3] , \wBIn41[21] , 
        \wBIn122[10] , \wBMid0[9] , \wBIn3[25] , \wBIn3[16] , \wBMid24[31] , 
        \wBMid72[29] , \wRegInA124[26] , \ScanLink131[7] , \ScanLink38[28] , 
        \wBMid24[28] , \wBMid51[18] , \wBMid72[30] , \ScanLink38[31] , 
        \wBMid81[9] , \wBMid32[6] , \wRegInA107[17] , \wRegInA112[23] , 
        \ScanLink253[28] , \ScanLink251[2] , \ScanLink226[18] , 
        \ScanLink205[30] , \ScanLink253[31] , \ScanLink205[29] , \wBIn9[2] , 
        \wAIn18[1] , \wAMid46[9] , \ScanLink166[26] , \wBMid82[24] , 
        \wAMid89[0] , \ScanLink113[16] , \ScanLink182[8] , \ScanLink145[17] , 
        \wAIn86[11] , \wBIn87[30] , \wBIn87[29] , \wBMid97[10] , \wAMid104[7] , 
        \ScanLink150[23] , \ScanLink130[27] , \ScanLink125[13] , 
        \ScanLink73[3] , \wBMid100[28] , \wRegInB81[4] , \ScanLink173[12] , 
        \ScanLink106[22] , \wAIn93[25] , \wBMid100[31] , \wRegInA79[12] , 
        \wAMid119[19] , \wBMid123[19] , \wBIn126[6] , \wRegInA33[7] , 
        \wAMid119[8] , \wRegInA111[8] , \wRegInA19[16] , \wRegInB53[2] , 
        \wRegInB71[15] , \wBMid19[21] , \wBMid31[5] , \wAMid58[5] , 
        \wAIn68[24] , \wBIn125[5] , \wRegInA30[4] , \wRegInB52[24] , 
        \wRegInB27[14] , \wRegInA82[13] , \wBMid79[25] , \wRegInB11[11] , 
        \wRegInB32[20] , \wRegInB47[10] , \wRegInB50[1] , \ScanLink233[8] , 
        \wRegInB64[21] , \wRegInA97[27] , \ScanLink33[24] , \wAMid107[4] , 
        \wAIn115[13] , \ScanLink46[14] , \ScanLink10[15] , \wAIn100[27] , 
        \wAIn123[16] , \ScanLink238[20] , \ScanLink65[25] , \wRegInB82[7] , 
        \ScanLink188[13] , \ScanLink70[11] , \ScanLink70[0] , \ScanLink26[10] , 
        \wBMid84[4] , \wRegInA57[3] , \ScanLink53[20] , \ScanLink2[31] , 
        \wAIn86[22] , \wRegInA19[25] , \ScanLink2[28] , \wAIn93[16] , 
        \wRegInB37[6] , \wRegInA79[21] , \wBMid56[2] , \wAIn62[9] , 
        \wBMid97[23] , \wRegInB122[28] , \ScanLink129[5] , \ScanLink125[20] , 
        \wRegInB0[29] , \ScanLink150[10] , \wRegInB0[30] , \wRegInA85[5] , 
        \wRegInB101[19] , \wRegInB122[31] , \ScanLink106[11] , 
        \ScanLink249[0] , \ScanLink173[21] , \ScanLink113[25] , 
        \ScanLink166[15] , \wAMid13[18] , \wBIn19[6] , \wBMid55[1] , 
        \wBMid82[17] , \ScanLink17[7] , \ScanLink145[24] , \ScanLink130[14] , 
        \wAIn123[25] , \ScanLink188[20] , \ScanLink70[22] , \wBMid19[12] , 
        \wAMid30[30] , \wAMid66[28] , \wBMid79[16] , \wAIn100[14] , 
        \ScanLink53[13] , \wRegInA86[6] , \ScanLink46[27] , \ScanLink26[23] , 
        \ScanLink33[17] , \ScanLink14[4] , \wAIn115[20] , \wRegInB32[13] , 
        \ScanLink238[13] , \ScanLink65[16] , \ScanLink10[26] , \wRegInA97[14] , 
        \wBMid87[7] , \wRegInB47[23] , \wBMid25[22] , \wAMid30[29] , 
        \wAMid45[19] , \wAMid66[31] , \wRegInB11[22] , \ScanLink137[9] , 
        \wRegInA54[0] , \wRegInB64[12] , \wBMid50[12] , \wAIn68[17] , 
        \wRegInB71[26] , \wRegInB27[27] , \wRegInA82[20] , \wRegInB34[5] , 
        \wRegInB52[17] , \wBMid91[3] , \ScanLink247[16] , \wBMid66[17] , 
        \wBMid73[23] , \ScanLink232[26] , \ScanLink197[21] , \ScanLink39[22] , 
        \wRegInA42[4] , \ScanLink211[17] , \wBIn2[9] , \wAIn4[21] , 
        \wBMid13[27] , \ScanLink204[23] , \wRegInA113[30] , \ScanLink59[26] , 
        \wBMid8[1] , \wBMid45[26] , \ScanLink252[22] , \ScanLink241[8] , 
        \wAIn17[12] , \wBMid30[16] , \wRegInB22[1] , \ScanLink227[12] , 
        \ScanLink182[15] , \wBMid43[5] , \wBMid107[8] , \wRegInA113[29] , 
        \wAIn21[17] , \wAIn34[23] , \wAIn62[22] , \wRegInB58[22] , 
        \wAMid79[29] , \wRegInA88[15] , \wAIn41[13] , \wAMid79[30] , 
        \wRegInA90[2] , \wAMid34[9] , \wBMid40[6] , \wAIn54[27] , \wAIn77[16] , 
        \wRegInB38[26] , \wAMid82[31] , \wAMid82[28] , \wAIn99[23] , 
        \wRegInA25[15] , \wRegInA50[25] , \wRegInB80[12] , \wRegInA93[1] , 
        \wRegInA73[14] , \wRegInA13[10] , \wRegInA66[20] , \wRegInA30[21] , 
        \wRegInA45[11] , \wRegInB95[26] , \wAIn69[2] , \wBMid88[22] , 
        \wAIn120[9] , \wRegInA41[7] , \wAMid0[16] , \wBIn9[10] , \wAMid9[6] , 
        \wBIn16[19] , \wAIn21[24] , \wAMid29[6] , \wBMid92[0] , \wBMid119[4] , 
        \ScanLink94[22] , \wBIn40[18] , \wBIn123[29] , \wRegInB21[2] , 
        \ScanLink179[14] , \ScanLink119[10] , \ScanLink81[16] , 
        \ScanLink158[6] , \wAIn54[14] , \wBIn63[30] , \wAMid111[0] , 
        \wBMid27[1] , \wBIn35[28] , \wAIn77[25] , \wBIn100[18] , \wBIn123[30] , 
        \wRegInB38[15] , \wBIn63[29] , \wBIn35[31] , \wAIn62[11] , 
        \wBMid13[14] , \wAIn17[21] , \wRegInA88[26] , \ScanLink238[3] , 
        \wAIn34[10] , \wAIn41[20] , \wRegInB58[11] , \wRegInB94[3] , 
        \ScanLink66[4] , \wRegInA119[0] , \ScanLink204[10] , \ScanLink145[9] , 
        \wBIn76[9] , \ScanLink59[15] , \wAIn4[12] , \wBMid30[25] , 
        \wBMid66[24] , \wRegInA26[0] , \ScanLink227[21] , \ScanLink182[26] , 
        \wAMid81[8] , \wRegInB6[5] , \wBIn4[7] , \wBIn7[4] , \wBIn9[23] , 
        \wBMid25[11] , \wBMid45[15] , \ScanLink252[11] , \wBMid50[21] , 
        \ScanLink232[15] , \ScanLink197[12] , \wBMid73[10] , \wRegInB46[5] , 
        \ScanLink247[25] , \ScanLink211[24] , \ScanLink39[11] , \wBMid88[11] , 
        \wRegInB5[6] , \ScanLink179[27] , \wRegInA25[3] , \ScanLink189[3] , 
        \ScanLink81[25] , \ScanLink119[23] , \ScanLink78[8] , \ScanLink94[11] , 
        \wAIn10[9] , \wBMid24[2] , \wRegInB45[6] , \wBIn68[5] , \wBIn98[28] , 
        \wAMid125[29] , \wRegInA13[23] , \wRegInA66[13] , \wAMid106[18] , 
        \wRegInA30[12] , \wRegInB95[15] , \wAMid112[3] , \wAMid125[30] , 
        \wRegInA45[22] , \wBIn14[3] , \wBIn98[31] , \wAIn99[10] , 
        \wRegInA25[26] , \wRegInB80[21] , \wRegInA50[16] , \ScanLink65[7] , 
        \wRegInB97[0] , \wAIn125[4] , \wRegInB10[28] , \wRegInB58[9] , 
        \wRegInA73[27] , \wAMid12[12] , \wAMid31[23] , \wAMid44[13] , 
        \wRegInB46[30] , \ScanLink127[3] , \wRegInB65[18] , \wBMid58[4] , 
        \wRegInB10[31] , \wRegInB33[19] , \wAMid67[22] , \wBIn68[25] , 
        \wRegInB46[29] , \wBMid18[18] , \wAMid24[17] , \wAMid51[27] , 
        \wAMid72[16] , \ScanLink247[6] , \ScanLink19[1] , \ScanLink52[19] , 
        \wAMid31[4] , \wAIn71[0] , \wRegInA59[5] , \ScanLink71[31] , 
        \wBMid101[6] , \ScanLink27[29] , \wRegInA118[16] , \ScanLink71[28] , 
        \wAMid32[7] , \wBMid46[8] , \wBMid89[1] , \wRegInB39[0] , 
        \ScanLink239[19] , \ScanLink27[30] , \wRegInB100[13] , \wBMid96[30] , 
        \wBMid102[5] , \wAIn72[3] , \wBMid96[29] , \wRegInB1[23] , 
        \wRegInB123[22] , \wAIn87[28] , \wRegInA7[26] , \wRegInB115[27] , 
        \wBIn93[24] , \wBMid114[25] , \ScanLink3[22] , \wAMid12[21] , 
        \wAIn15[4] , \wBIn17[0] , \wAIn126[7] , \ScanLink124[0] , \wAMid55[0] , 
        \wBIn86[10] , \wAIn87[31] , \wRegInA88[0] , \wAMid118[20] , 
        \wRegInA47[9] , \wBMid122[20] , \ScanLink244[5] , \wAMid89[17] , 
        \wBMid101[11] , \wAIn114[19] , \ScanLink191[1] , \wAMid24[24] , 
        \wAMid72[25] , \wAMid87[6] , \wRegInA118[25] , \ScanLink189[19] , 
        \wRegInA83[19] , \ScanLink143[7] , \wAMid31[10] , \wAMid51[14] , 
        \wBIn70[7] , \wAMid44[20] , \wRegInA102[1] , \ScanLink223[2] , 
        \wAIn16[7] , \wAMid67[11] , \wBIn68[16] , \wBIn73[4] , \wAMid84[5] , 
        \wBIn86[23] , \wAMid109[2] , \wAMid118[13] , \wBMid122[13] , 
        \ScanLink140[4] , \wAMid89[24] , \wBMid101[22] , \wRegInB3[8] , 
        \wRegInA78[18] , \wBIn93[17] , \wBMid114[16] , \ScanLink220[1] , 
        \wRegInB43[8] , \ScanLink3[11] , \wRegInA101[2] , \ScanLink192[2] , 
        \wAIn0[23] , \wAMid4[27] , \wAIn8[8] , \wAMid56[3] , \wRegInA7[15] , 
        \wBIn82[12] , \wBMid105[13] , \wBMid126[22] , \wRegInB1[10] , 
        \wRegInB100[20] , \wRegInB115[14] , \ScanLink172[18] , 
        \ScanLink151[30] , \ScanLink107[28] , \wRegInB123[11] , 
        \ScanLink151[29] , \ScanLink107[31] , \ScanLink63[9] , 
        \ScanLink124[19] , \wRegInA125[4] , \ScanLink95[9] , \ScanLink204[7] , 
        \wBIn12[31] , \wAMid15[2] , \wAMid16[23] , \wAMid16[10] , \wBMid18[6] , 
        \wAMid20[15] , \wAIn31[2] , \wAIn32[1] , \wBIn57[2] , \wBIn97[26] , 
        \wAMid98[21] , \ScanLink7[20] , \wAMid109[16] , \wBMid110[27] , 
        \ScanLink164[2] , \wAMid72[5] , \wRegInA3[24] , \ScanLink88[6] , 
        \wRegInB104[11] , \wRegInB111[25] , \ScanLink219[8] , 
        \ScanLink120[31] , \ScanLink6[3] , \ScanLink176[29] , 
        \ScanLink103[19] , \wBIn85[4] , \wRegInB127[20] , \ScanLink120[28] , 
        \wRegInB5[21] , \ScanLink176[30] , \ScanLink155[18] , \wBIn86[7] , 
        \wAIn110[31] , \wRegInB79[2] , \wRegInA109[20] , \wAIn110[28] , 
        \ScanLink5[0] , \wRegInA19[7] , \wAMid55[25] , \wAMid71[6] , 
        \wAMid76[14] , \wBIn79[13] , \wRegInA9[2] , \wRegInA87[28] , 
        \ScanLink207[4] , \wRegInA87[31] , \ScanLink59[3] , \wAMid35[21] , 
        \wAMid40[11] , \wBIn54[1] , \wRegInA126[7] , \wBIn111[9] , 
        \ScanLink167[1] , \wAMid63[20] , \wAMid16[1] , \wBIn19[17] , 
        \wAIn56[5] , \wBMid92[18] , \wRegInB127[13] , \wRegInB104[22] , 
        \wRegInB110[2] , \wRegInB5[12] , \wBMid126[3] , \wRegInA3[17] , 
        \wBIn33[6] , \wAIn83[19] , \wBIn97[15] , \wAMid98[12] , 
        \wRegInB111[16] , \ScanLink7[13] , \wBMid110[14] , \wAMid109[25] , 
        \wBMid126[11] , \wAMid35[12] , \wBIn82[21] , \wAIn84[3] , \wAIn102[1] , 
        \ScanLink100[6] , \wBMid105[20] , \wRegInB61[29] , \wAMid40[22] , 
        \wRegInB14[19] , \wRegInB37[31] , \wRegInB42[18] , \wRegInB61[30] , 
        \wBIn19[24] , \wAMid20[26] , \wAMid63[13] , \wRegInB37[28] , 
        \wAMid76[27] , \wAIn78[18] , \wBIn79[20] , \ScanLink103[5] , 
        \wBIn30[5] , \wAIn48[9] , \wAMid55[16] , \wAIn101[2] , \wBMid69[19] , 
        \wAIn87[0] , \ScanLink23[18] , \ScanLink20[8] , \wBMid125[0] , 
        \wRegInB113[1] , \ScanLink56[28] , \ScanLink248[18] , \ScanLink75[19] , 
        \ScanLink56[31] , \wRegInA109[13] , \wAIn29[0] , \wAIn55[6] , 
        \wBMid99[14] , \wRegInB61[0] , \ScanLink202[9] , \ScanLink85[14] , 
        \ScanLink108[26] , \ScanLink93[7] , \wBIn31[19] , \wAMid69[4] , 
        \wBIn114[4] , \ScanLink168[22] , \ScanLink90[20] , \wAIn88[15] , 
        \wRegInA62[22] , \wAMid102[30] , \wAMid121[18] , \wRegInA17[12] , 
        \wAMid102[29] , \wRegInA34[23] , \wRegInA41[13] , \ScanLink41[1] , 
        \wRegInB91[24] , \wRegInA21[17] , \wRegInA54[27] , \wRegInB84[10] , 
        \wRegInA77[16] , \ScanLink42[2] , \wBIn12[28] , \wAIn25[15] , 
        \wBIn44[29] , \wAIn50[25] , \wBIn104[30] , \wBIn127[18] , 
        \wRegInB49[14] , \wAIn13[10] , \wBIn44[30] , \wBIn67[18] , 
        \wBIn104[29] , \wRegInA99[23] , \wAIn73[14] , \wAIn30[21] , 
        \wAIn66[20] , \wAMid77[8] , \wRegInB29[10] , \wAIn45[11] , \wBIn80[9] , 
        \wBMid62[15] , \ScanLink90[4] , \ScanLink28[14] , \wBMid17[25] , 
        \wRegInA120[9] , \ScanLink200[21] , \ScanLink256[20] , \wAIn0[10] , 
        \wAMid4[14] , \wBMid17[16] , \wBMid21[20] , \wBMid34[14] , 
        \wBMid41[24] , \ScanLink223[10] , \ScanLink186[17] , \wBMid54[10] , 
        \wRegInB62[3] , \ScanLink243[14] , \wBMid21[13] , \wBIn28[7] , 
        \wBMid64[0] , \wBMid77[21] , \ScanLink236[24] , \ScanLink193[23] , 
        \wAMid86[19] , \wBIn117[7] , \ScanLink48[10] , \wRegInA21[24] , 
        \wRegInB84[23] , \ScanLink215[15] , \wRegInA54[14] , \ScanLink25[5] , 
        \wRegInA17[21] , \wRegInA77[25] , \wAIn88[26] , \wRegInA62[11] , 
        \wBIn35[8] , \wAIn119[0] , \wRegInA34[10] , \wRegInB91[17] , 
        \wRegInA8[31] , \wRegInA41[20] , \wRegInA8[28] , \ScanLink168[11] , 
        \ScanLink90[13] , \ScanLink108[15] , \ScanLink85[27] , \wBMid99[27] , 
        \ScanLink106[8] , \wRegInA65[1] , \wBMid54[23] , \wRegInB108[0] , 
        \ScanLink236[17] , \ScanLink193[10] , \wBMid77[12] , \ScanLink243[27] , 
        \ScanLink215[26] , \ScanLink48[23] , \ScanLink200[12] , \wBMid34[27] , 
        \wBMid62[26] , \wRegInA66[2] , \ScanLink28[27] , \wRegInA117[18] , 
        \ScanLink223[23] , \ScanLink186[24] , \ScanLink256[13] , \wBMid0[30] , 
        \wAMid1[22] , \wAIn13[23] , \wBMid41[17] , \wAIn66[13] , 
        \wRegInB29[23] , \wAIn25[26] , \wAIn30[12] , \wAIn45[22] , 
        \ScanLink26[6] , \wAIn50[16] , \ScanLink118[4] , \wAIn53[8] , 
        \wBMid24[25] , \wBMid51[15] , \wBMid67[3] , \wRegInA99[10] , 
        \wAIn73[27] , \wRegInB49[27] , \wBMid81[4] , \ScanLink246[11] , 
        \wBMid67[10] , \wBMid72[24] , \ScanLink233[21] , \ScanLink196[26] , 
        \wRegInA52[3] , \ScanLink38[25] , \ScanLink210[10] , \wAMid1[11] , 
        \wAIn5[26] , \wBMid12[20] , \ScanLink205[24] , \ScanLink58[21] , 
        \ScanLink253[25] , \wBMid5[9] , \wAIn16[15] , \wBMid31[11] , 
        \wBMid44[21] , \ScanLink226[15] , \ScanLink183[12] , \wRegInB32[6] , 
        \wAIn20[10] , \wBIn21[31] , \wBIn21[28] , \wAIn35[24] , \wBMid53[2] , 
        \wAIn63[25] , \wRegInB59[25] , \wBIn77[29] , \wBIn114[18] , 
        \wRegInA89[12] , \wAIn40[14] , \wBIn54[18] , \wAIn67[9] , \wBIn77[30] , 
        \wRegInA80[5] , \ScanLink12[7] , \wAIn55[20] , \wRegInB39[21] , 
        \wBIn8[17] , \wBMid50[1] , \wAIn76[11] , \wAIn98[24] , \wAMid112[18] , 
        \wRegInA51[22] , \wRegInA83[6] , \wRegInA24[12] , \wRegInB81[15] , 
        \wAIn79[5] , \wRegInA12[17] , \wRegInA67[27] , \wRegInA72[13] , 
        \wRegInA31[26] , \wRegInA44[16] , \ScanLink11[4] , \wRegInB94[21] , 
        \ScanLink132[9] , \wBMid89[25] , \wRegInA51[0] , \wBMid12[13] , 
        \wAIn16[26] , \wAMid18[19] , \wAIn20[23] , \wAMid39[1] , \wBMid82[7] , 
        \ScanLink95[25] , \wBMid109[3] , \wAIn55[13] , \wRegInB31[5] , 
        \ScanLink178[13] , \ScanLink118[17] , \ScanLink80[11] , 
        \ScanLink148[1] , \wAMid101[7] , \ScanLink187[8] , \wBMid37[6] , 
        \wRegInB39[12] , \wAMid43[9] , \wAIn76[22] , \wAIn63[16] , 
        \wRegInA89[21] , \ScanLink228[4] , \wAIn35[17] , \wAIn40[27] , 
        \wRegInB59[16] , \wRegInB84[4] , \ScanLink76[3] , \wRegInA109[7] , 
        \ScanLink205[17] , \ScanLink58[12] , \wAIn5[15] , \wBMid31[22] , 
        \wBMid67[23] , \wBIn123[6] , \wRegInA36[7] , \ScanLink226[26] , 
        \ScanLink183[21] , \ScanLink253[16] , \wBMid24[16] , \wBMid44[12] , 
        \wRegInA107[29] , \ScanLink233[12] , \ScanLink196[15] , \wBMid0[29] , 
        \wBMid51[26] , \wRegInB56[2] , \wRegInA107[30] , \wRegInA124[18] , 
        \ScanLink246[22] , \ScanLink210[23] , \wBMid0[4] , \wBIn3[31] , 
        \wBMid3[7] , \wBIn8[24] , \wBMid72[17] , \wBMid89[16] , \wBIn120[5] , 
        \wRegInA114[8] , \ScanLink199[4] , \ScanLink178[20] , \ScanLink38[16] , 
        \ScanLink80[22] , \wRegInA35[4] , \ScanLink236[8] , \ScanLink118[24] , 
        \ScanLink95[16] , \wAMid13[15] , \wAMid30[24] , \wBMid34[5] , 
        \wRegInA12[24] , \wRegInB55[1] , \wAMid45[14] , \wBIn78[2] , 
        \wAMid96[28] , \wRegInA67[14] , \ScanLink9[29] , \wAMid96[31] , 
        \wAMid102[4] , \wRegInA31[15] , \wRegInB94[12] , \wRegInA44[25] , 
        \ScanLink9[30] , \wAIn98[17] , \wRegInA24[21] , \wRegInA51[11] , 
        \wRegInB81[26] , \ScanLink75[0] , \wRegInB87[7] , \wRegInA72[20] , 
        \ScanLink137[4] , \wBMid48[3] , \wAMid66[25] , \wBIn69[22] , 
        \wRegInA97[19] , \wAMid21[3] , \wAMid25[10] , \wAMid50[20] , 
        \wAMid73[11] , \wRegInB34[8] , \wAIn61[7] , \wAIn100[19] , 
        \wAIn123[31] , \wRegInA49[2] , \wBMid111[1] , \wAIn123[28] , 
        \wRegInA119[11] , \wAMid22[0] , \wBMid99[6] , \wRegInB127[0] , 
        \wRegInB29[7] , \wRegInB101[14] , \ScanLink14[9] , \wBMid112[2] , 
        \wAIn62[4] , \wRegInB0[24] , \wRegInB122[25] , \ScanLink129[8] , 
        \wRegInA85[8] , \ScanLink130[19] , \ScanLink113[31] , \wBIn3[28] , 
        \wRegInA6[21] , \ScanLink145[29] , \wRegInB114[20] , \wRegInB124[3] , 
        \ScanLink113[28] , \ScanLink145[30] , \wAMid1[3] , \wAMid2[0] , 
        \wAMid25[23] , \wBMid31[8] , \wBMid79[31] , \wBMid84[9] , 
        \ScanLink166[18] , \wBIn87[17] , \wAMid88[10] , \wBIn92[23] , 
        \wBMid115[22] , \wRegInA19[28] , \ScanLink2[25] , \wAMid119[27] , 
        \wRegInA19[31] , \wRegInA98[7] , \ScanLink134[7] , \wBMid123[27] , 
        \ScanLink254[2] , \wBMid100[16] , \ScanLink33[30] , \ScanLink10[18] , 
        \wAMid45[7] , \ScanLink65[28] , \wAMid58[8] , \wAIn68[29] , 
        \wBMid79[28] , \ScanLink33[29] , \wAMid107[9] , \ScanLink181[6] , 
        \ScanLink65[31] , \ScanLink46[19] , \wRegInB52[29] , \wRegInA119[22] , 
        \wAMid73[22] , \wAMid97[1] , \wRegInB27[19] , \ScanLink153[0] , 
        \wAMid30[17] , \wAMid50[13] , \wBIn60[0] , \wRegInB52[30] , 
        \wRegInB71[18] , \wAIn68[30] , \wBIn125[8] , \wRegInA30[9] , 
        \wAMid45[27] , \wRegInA112[6] , \wAMid13[26] , \ScanLink233[5] , 
        \wBIn63[3] , \wAMid66[16] , \wBIn69[11] , \wAIn93[31] , \wBMid123[14] , 
        \wBIn87[24] , \wAMid88[23] , \wAIn93[28] , \wAMid119[14] , 
        \ScanLink150[3] , \wAMid119[5] , \wBIn92[10] , \wAMid94[2] , 
        \wBMid100[25] , \wBMid115[11] , \ScanLink230[6] , \ScanLink2[16] , 
        \wAIn5[0] , \wAMid46[4] , \wBMid82[30] , \wBMid82[29] , 
        \wRegInA111[5] , \ScanLink182[5] , \wRegInA6[12] , \wBIn47[5] , 
        \wBIn83[15] , \wBMid104[14] , \wRegInB0[17] , \wRegInB81[9] , 
        \wRegInB101[27] , \wRegInB114[13] , \wRegInB122[16] , \ScanLink214[0] , 
        \wBIn96[21] , \wAIn97[19] , \wRegInA7[9] , \wRegInB77[9] , 
        \wAMid99[26] , \wBMid111[20] , \wAMid108[11] , \ScanLink174[5] , 
        \ScanLink6[27] , \wBMid86[18] , \wRegInA2[23] , \ScanLink98[1] , 
        \ScanLink57[8] , \wRegInB110[22] , \wAIn6[3] , \wAIn21[5] , 
        \wAIn22[6] , \wAMid62[2] , \wRegInB105[16] , \wBIn95[3] , 
        \wRegInB126[27] , \wRegInB4[26] , \wBIn59[9] , \wRegInB69[5] , 
        \wRegInA108[27] , \ScanLink61[19] , \ScanLink42[31] , \ScanLink14[29] , 
        \ScanLink42[28] , \ScanLink37[18] , \ScanLink14[30] , \wBIn96[0] , 
        \ScanLink229[31] , \ScanLink229[28] , \wBIn7[19] , \wAMid17[17] , 
        \wBIn18[10] , \wAIn19[31] , \wAIn19[28] , \wAMid61[1] , \wAMid77[13] , 
        \wBIn78[14] , \wRegInB23[28] , \ScanLink217[3] , \wAMid54[22] , 
        \wRegInB56[18] , \wRegInB75[30] , \ScanLink8[8] , \wRegInB23[31] , 
        \ScanLink49[4] , \wAMid21[12] , \wAMid34[26] , \wAMid41[16] , 
        \wBIn44[6] , \wRegInB75[29] , \ScanLink177[6] , \wAMid62[27] , 
        \wAIn46[2] , \wRegInB4[15] , \wRegInB100[5] , \wRegInB105[25] , 
        \wRegInB126[14] , \ScanLink162[30] , \ScanLink141[18] , 
        \ScanLink134[28] , \wAMid17[24] , \wBIn18[23] , \wBIn23[1] , 
        \wBMid72[9] , \wBIn96[12] , \wRegInA2[10] , \ScanLink162[29] , 
        \wRegInA68[29] , \wRegInB110[11] , \ScanLink134[31] , 
        \ScanLink117[19] , \wAMid99[15] , \wBMid111[13] , \wAMid108[22] , 
        \wRegInA68[30] , \ScanLink6[14] , \wAMid34[15] , \wBIn83[26] , 
        \wAIn94[4] , \wAIn112[6] , \wRegInA73[8] , \ScanLink110[1] , 
        \wBMid104[27] , \wAMid41[25] , \wRegInA93[31] , \wBIn20[2] , 
        \wAMid21[21] , \wAMid62[14] , \wRegInA93[28] , \wAMid77[20] , 
        \wBIn78[27] , \ScanLink113[2] , \wAMid54[11] , \wAIn111[5] , 
        \wAIn97[7] , \wAIn104[28] , \wAMid0[31] , \wAIn1[24] , \wAMid5[20] , 
        \wBMid10[3] , \wAIn24[8] , \wAIn39[7] , \wAIn45[1] , \wAIn104[31] , 
        \wAIn127[19] , \wRegInB103[6] , \wRegInA108[14] , \ScanLink199[28] , 
        \wBMid98[13] , \wRegInB71[7] , \ScanLink199[31] , \ScanLink109[21] , 
        \ScanLink84[13] , \ScanLink83[0] , \wAMid79[3] , \wBIn104[3] , 
        \wRegInA11[2] , \wRegInA1[7] , \ScanLink169[25] , \ScanLink91[27] , 
        \wAIn89[12] , \wAMid92[19] , \wRegInA63[25] , \wRegInA16[15] , 
        \wRegInA35[24] , \wRegInA40[14] , \ScanLink51[6] , \wRegInB90[23] , 
        \wRegInA55[20] , \wAMid126[2] , \wRegInA20[10] , \wRegInA76[11] , 
        \wRegInB85[17] , \wAIn12[17] , \wBMid13[0] , \wAIn24[12] , 
        \ScanLink52[5] , \wAIn51[22] , \wAMid69[18] , \wRegInB48[13] , 
        \wRegInA98[24] , \wAIn72[13] , \wAIn31[26] , \wAIn67[27] , 
        \wRegInB28[17] , \wAIn44[16] , \wBMid63[12] , \wAMid125[1] , 
        \ScanLink80[3] , \ScanLink29[13] , \wBMid16[22] , \ScanLink201[26] , 
        \wAIn1[17] , \wBMid4[18] , \wBMid20[27] , \wBMid35[13] , \wBMid40[23] , 
        \wRegInB72[4] , \ScanLink222[17] , \ScanLink187[10] , \wBMid55[17] , 
        \wRegInA103[18] , \ScanLink242[13] , \wRegInA120[30] , \wBIn42[8] , 
        \wRegInA2[4] , \ScanLink237[23] , \ScanLink192[24] , \wBMid76[26] , 
        \wAMid5[13] , \wBMid16[11] , \wBMid20[14] , \wBIn38[0] , \wBMid74[7] , 
        \wBIn88[19] , \wBIn107[0] , \wRegInA12[1] , \ScanLink171[8] , 
        \wRegInA120[29] , \ScanLink49[17] , \wAMid116[30] , \wAMid116[29] , 
        \ScanLink214[12] , \wRegInA20[23] , \wRegInA55[13] , \wRegInB85[24] , 
        \ScanLink35[2] , \wRegInA76[22] , \wAIn89[21] , \wRegInA16[26] , 
        \wRegInA63[16] , \wBMid69[8] , \wAIn109[7] , \wRegInA35[17] , 
        \wRegInB90[10] , \wRegInB15[3] , \wRegInA40[27] , \wRegInA68[9] , 
        \ScanLink91[14] , \ScanLink169[16] , \wBMid98[20] , \wAIn114[8] , 
        \ScanLink109[12] , \ScanLink84[20] , \wRegInA75[6] , \wBMid55[24] , 
        \ScanLink237[10] , \ScanLink192[17] , \wBMid76[15] , \wRegInB16[0] , 
        \wRegInB118[7] , \ScanLink242[20] , \ScanLink214[21] , 
        \ScanLink49[24] , \ScanLink201[15] , \wBMid35[20] , \wBMid63[21] , 
        \wAIn91[9] , \wRegInA76[5] , \ScanLink29[20] , \ScanLink222[24] , 
        \ScanLink187[23] , \wBIn1[7] , \wBIn2[4] , \wBMid1[23] , \wAMid4[19] , 
        \wBIn6[20] , \wBIn6[13] , \wAIn12[24] , \wBMid40[10] , \wBIn50[30] , 
        \wAIn67[14] , \wBIn73[18] , \wBIn110[29] , \wRegInB28[24] , 
        \wAIn18[11] , \wBIn19[30] , \wBIn19[29] , \wAIn24[21] , \wBIn25[19] , 
        \wAIn44[25] , \wRegInB105[8] , \wBIn50[29] , \ScanLink36[1] , 
        \wBIn110[30] , \wAIn31[15] , \wAIn51[11] , \ScanLink108[3] , 
        \wBMid61[0] , \wBMid69[14] , \wAIn72[20] , \wRegInA98[17] , 
        \wBMid77[4] , \wAIn105[22] , \wAIn126[13] , \wRegInB48[20] , 
        \ScanLink228[11] , \ScanLink75[14] , \ScanLink20[5] , \ScanLink23[15] , 
        \wAIn110[16] , \ScanLink56[25] , \ScanLink36[21] , \ScanLink248[15] , 
        \ScanLink43[11] , \ScanLink15[10] , \wRegInB42[15] , \ScanLink198[22] , 
        \ScanLink60[20] , \wAIn78[15] , \wRegInB37[25] , \wRegInA92[22] , 
        \wRegInB61[24] , \wBIn30[8] , \wRegInB14[14] , \wRegInB74[10] , 
        \ScanLink103[8] , \wAIn48[4] , \wRegInA60[1] , \wBMid62[3] , 
        \wAIn83[14] , \wAMid109[28] , \wRegInB22[11] , \wRegInB57[21] , 
        \wRegInA87[16] , \wRegInA69[23] , \wBMid92[15] , \wAIn96[20] , 
        \wBIn97[18] , \wBMid110[19] , \wAMid109[31] , \wRegInA63[2] , 
        \ScanLink155[26] , \ScanLink120[16] , \ScanLink23[6] , 
        \ScanLink176[17] , \ScanLink103[27] , \wAIn18[22] , \wAMid20[18] , 
        \wAMid55[28] , \wAIn56[8] , \wBMid87[21] , \ScanLink163[23] , 
        \ScanLink140[12] , \ScanLink116[13] , \wAIn99[1] , \ScanLink135[22] , 
        \ScanLink96[7] , \wAMid55[31] , \wRegInB74[23] , \ScanLink207[9] , 
        \wAMid76[19] , \wRegInB22[22] , \wRegInA87[25] , \wBIn49[3] , 
        \wAIn78[26] , \wRegInB37[16] , \wRegInB57[12] , \wRegInB64[0] , 
        \wRegInA92[11] , \wAIn110[25] , \wBIn111[4] , \wRegInB14[27] , 
        \wRegInB42[26] , \wRegInB61[17] , \ScanLink44[1] , \ScanLink43[22] , 
        \ScanLink36[12] , \wAIn126[20] , \ScanLink248[26] , \ScanLink198[11] , 
        \ScanLink60[13] , \ScanLink15[23] , \ScanLink228[22] , 
        \ScanLink75[27] , \wBMid69[27] , \wAIn105[11] , \ScanLink56[16] , 
        \ScanLink23[26] , \wRegInA3[29] , \wRegInB111[28] , \ScanLink219[5] , 
        \ScanLink116[20] , \wBMid5[21] , \wAIn8[5] , \wAMid72[8] , \wBIn85[9] , 
        \wBMid87[12] , \wRegInA3[30] , \ScanLink163[10] , \ScanLink47[2] , 
        \wRegInB111[31] , \ScanLink135[11] , \ScanLink140[21] , \wBMid92[26] , 
        \ScanLink179[0] , \ScanLink120[25] , \ScanLink176[24] , 
        \ScanLink155[15] , \ScanLink103[14] , \wAIn96[13] , \wRegInB67[3] , 
        \wBIn98[6] , \wRegInA125[9] , \ScanLink95[4] , \wBIn112[7] , 
        \wBIn12[16] , \wBIn24[13] , \wBIn51[23] , \wAIn83[27] , 
        \wRegInA69[10] , \wBIn67[26] , \wAMid68[21] , \wBIn72[12] , 
        \wBIn104[17] , \wBIn111[23] , \wRegInB115[2] , \wBMid123[3] , 
        \wAMid13[1] , \wBIn31[27] , \wBIn44[17] , \wBIn127[26] , 
        \ScanLink118[9] , \wAIn53[5] , \wRegInA121[10] , \wBIn36[6] , 
        \wRegInA102[21] , \wRegInA117[15] , \ScanLink186[29] , 
        \ScanLink186[30] , \ScanLink105[6] , \wAIn81[3] , \wAIn107[1] , 
        \wBMid5[12] , \wAMid10[2] , \wBIn35[5] , \wRegInA8[25] , 
        \ScanLink38[7] , \wAIn50[6] , \wBMid79[2] , \wAIn82[0] , \wAIn104[2] , 
        \ScanLink106[5] , \ScanLink108[18] , \wAMid86[14] , \wBIn89[13] , 
        \wRegInA21[30] , \wAMid102[17] , \wAMid117[23] , \wRegInB18[6] , 
        \wRegInA77[28] , \wRegInB116[1] , \wRegInA21[29] , \ScanLink25[8] , 
        \wRegInA54[19] , \wRegInA77[31] , \wRegInA78[3] , \wBMid120[0] , 
        \wAMid121[26] , \wBMid17[31] , \wBMid41[29] , \wAMid93[20] , 
        \ScanLink201[7] , \wBMid17[28] , \wBMid34[19] , \wRegInA117[26] , 
        \wBMid41[30] , \ScanLink90[9] , \wBMid62[18] , \wRegInA120[4] , 
        \ScanLink28[19] , \wAIn10[4] , \wBIn12[25] , \wBIn52[2] , 
        \wRegInB49[19] , \wRegInA102[12] , \wRegInA121[23] , \ScanLink161[2] , 
        \ScanLink243[19] , \ScanLink236[30] , \ScanLink215[18] , 
        \ScanLink236[29] , \wBIn24[20] , \wAIn25[18] , \wAIn50[31] , 
        \wAMid68[12] , \wAIn73[19] , \wBIn104[24] , \ScanLink3[3] , 
        \wBIn67[15] , \wBIn31[14] , \wBIn44[24] , \wBIn127[15] , \wAIn50[28] , 
        \wAIn34[2] , \wAIn37[1] , \wBIn51[10] , \wBIn80[4] , \wBIn72[21] , 
        \wAMid77[5] , \wAMid74[6] , \wAMid86[27] , \wAIn88[18] , 
        \wAMid102[24] , \wBIn111[10] , \wRegInB91[29] , \wBIn89[20] , 
        \wAMid93[13] , \wAMid121[15] , \wRegInB91[30] , \ScanLink0[0] , 
        \wBIn83[7] , \wAMid117[10] , \wBIn51[1] , \wAMid69[9] , \wBMid99[19] , 
        \wBIn109[6] , \wRegInA123[7] , \wRegInA8[16] , \ScanLink202[4] , 
        \ScanLink85[19] , \ScanLink162[1] , \wBIn68[8] , \wBIn114[9] , 
        \wRegInB95[18] , \ScanLink194[1] , \wAMid106[15] , \wRegInA38[1] , 
        \wBMid13[19] , \wBMid30[31] , \wBMid30[28] , \wBMid39[0] , 
        \wAMid50[0] , \wAMid125[24] , \wBIn75[7] , \wAMid82[16] , 
        \wAMid97[22] , \wBIn98[25] , \ScanLink8[23] , \wAMid113[21] , 
        \wRegInB58[4] , \ScanLink146[7] , \ScanLink81[31] , \wAMid82[6] , 
        \ScanLink81[28] , \wRegInA107[1] , \ScanLink226[2] , \ScanLink78[5] , 
        \wBMid45[18] , \wBMid66[30] , \wAMid81[5] , \wRegInB6[8] , 
        \wRegInA113[17] , \wBIn76[4] , \ScanLink145[4] , \wBMid66[29] , 
        \ScanLink59[18] , \wRegInA104[2] , \wRegInA125[12] , \ScanLink211[29] , 
        \wAIn13[7] , \wBIn16[14] , \wAMid19[13] , \wAIn21[30] , \wBIn63[24] , 
        \wBIn100[15] , \wRegInB38[18] , \wRegInB46[8] , \wRegInA106[23] , 
        \ScanLink247[31] , \ScanLink232[18] , \ScanLink225[1] , 
        \ScanLink211[30] , \wRegInB89[1] , \ScanLink247[28] , \wAIn77[28] , 
        \wAMid53[3] , \wBIn40[15] , \wAIn54[19] , \wBIn123[24] , 
        \ScanLink197[2] , \wAIn77[31] , \wBIn20[11] , \wAIn21[29] , 
        \wBIn35[25] , \wBIn55[21] , \ScanLink66[9] , \wBIn76[10] , 
        \wAMid79[17] , \wBIn115[21] , \wBMid119[9] , \wBMid1[10] , \wBIn11[3] , 
        \wAIn120[4] , \ScanLink122[3] , \wBIn16[27] , \wAMid19[20] , 
        \wBIn20[22] , \wAMid34[4] , \wAMid82[25] , \ScanLink242[6] , 
        \ScanLink179[19] , \wBMid104[6] , \wRegInA73[19] , \wRegInA50[31] , 
        \wAIn74[0] , \wAMid113[12] , \wRegInA50[28] , \wAMid97[11] , 
        \wAMid106[26] , \wRegInA25[18] , \wBIn98[16] , \ScanLink8[10] , 
        \wAMid125[17] , \wAMid37[7] , \wBMid43[8] , \wBIn55[12] , \wAIn77[3] , 
        \wBIn76[23] , \wBMid107[5] , \wAMid79[24] , \wBIn115[12] , 
        \wRegInA88[18] , \wBIn35[16] , \wBIn63[17] , \wBIn100[26] , 
        \wBIn40[26] , \wBIn123[17] , \wAIn123[7] , \wBIn12[0] , \wRegInA42[9] , 
        \wRegInA125[21] , \ScanLink121[0] , \wRegInA106[10] , \ScanLink241[5] , 
        \wAMid0[28] , \wRegInA113[24] , \ScanLink182[18] , \wBIn2[11] , 
        \wBMid22[1] , \wAMid24[29] , \wBIn73[9] , \wBMid83[23] , \wAMid99[7] , 
        \wRegInA7[18] , \ScanLink167[21] , \wRegInB115[19] , \ScanLink112[11] , 
        \ScanLink144[10] , \wAMid84[8] , \wAMid89[29] , \wBMid96[17] , 
        \wAMid114[0] , \ScanLink151[24] , \ScanLink131[20] , \ScanLink124[14] , 
        \ScanLink63[4] , \wRegInB91[3] , \ScanLink172[15] , \ScanLink107[25] , 
        \wAIn92[22] , \wRegInB3[5] , \wRegInA78[15] , \wAMid89[30] , 
        \wAIn87[16] , \wRegInA23[0] , \ScanLink140[9] , \wRegInA18[11] , 
        \wRegInB43[5] , \wAMid51[19] , \wAMid72[31] , \wRegInB70[12] , 
        \wBIn2[22] , \wAIn15[9] , \wAMid24[30] , \wRegInA20[3] , \wAMid48[2] , 
        \wAIn69[23] , \wAMid72[28] , \wRegInB53[23] , \wRegInB0[6] , 
        \wRegInB26[13] , \wRegInA83[14] , \wBMid78[22] , \wRegInB10[16] , 
        \wRegInB33[27] , \wRegInB40[6] , \wRegInB46[17] , \wRegInA96[20] , 
        \wRegInB65[26] , \wAIn114[14] , \ScanLink32[23] , \wAMid117[3] , 
        \wBMid18[26] , \wBMid21[2] , \ScanLink47[13] , \ScanLink11[12] , 
        \wAIn101[20] , \wAIn122[11] , \ScanLink239[27] , \ScanLink64[22] , 
        \wRegInB92[0] , \wRegInA118[28] , \ScanLink189[14] , \ScanLink71[16] , 
        \wRegInA118[31] , \ScanLink60[7] , \ScanLink52[27] , \ScanLink27[17] , 
        \wBMid46[5] , \wAIn87[25] , \wBIn93[30] , \wBIn93[29] , \wBMid94[3] , 
        \wBMid114[31] , \wRegInA18[22] , \wRegInA47[4] , \wBMid114[28] , 
        \wAIn92[11] , \ScanLink244[8] , \wBMid96[24] , \wRegInB27[1] , 
        \wRegInA78[26] , \ScanLink139[2] , \ScanLink124[27] , \wBMid102[8] , 
        \wRegInA95[2] , \ScanLink151[17] , \ScanLink107[16] , 
        \ScanLink172[26] , \ScanLink112[22] , \wBIn7[9] , \wBMid18[15] , 
        \wAMid31[9] , \wBMid45[6] , \wBMid83[10] , \ScanLink167[12] , 
        \ScanLink144[23] , \ScanLink131[13] , \ScanLink189[27] , 
        \ScanLink71[25] , \wAIn122[22] , \ScanLink52[14] , \wBMid58[9] , 
        \wBMid78[11] , \wAIn101[13] , \wRegInA59[8] , \wRegInA96[1] , 
        \ScanLink47[20] , \ScanLink27[24] , \wAIn114[27] , \ScanLink32[10] , 
        \wRegInB33[14] , \wRegInA96[13] , \ScanLink239[14] , \ScanLink64[11] , 
        \ScanLink11[21] , \wBIn68[31] , \wBIn68[28] , \wBMid97[0] , 
        \wAIn125[9] , \wRegInB46[24] , \wRegInB10[25] , \wRegInA44[7] , 
        \wRegInB65[15] , \wAIn0[27] , \wBMid21[24] , \wBMid54[14] , 
        \wAIn69[10] , \wRegInB70[21] , \wBMid77[25] , \wRegInB24[2] , 
        \wRegInB26[20] , \wRegInB53[10] , \wRegInA83[27] , \wBIn117[3] , 
        \ScanLink48[14] , \ScanLink215[11] , \ScanLink243[10] , 
        \ScanLink236[20] , \ScanLink193[27] , \wAIn0[14] , \wAMid4[23] , 
        \wBMid34[10] , \wBMid41[20] , \ScanLink256[24] , \wRegInB62[7] , 
        \ScanLink223[14] , \ScanLink186[13] , \wBMid62[11] , \ScanLink90[0] , 
        \ScanLink28[10] , \wAIn13[27] , \wAIn13[14] , \wBMid17[21] , 
        \ScanLink200[25] , \wBIn24[30] , \wBIn24[29] , \wAIn30[25] , 
        \wAIn37[8] , \wAIn45[15] , \wBIn51[19] , \wBIn72[31] , \wAMid13[8] , 
        \wAIn25[11] , \wAIn66[24] , \wBIn72[28] , \wAIn73[10] , \wBIn111[19] , 
        \wRegInB29[14] , \wRegInB49[10] , \wRegInA99[27] , \ScanLink42[6] , 
        \wAIn29[4] , \wAIn50[21] , \wBIn51[8] , \wAMid69[0] , \wAIn88[11] , 
        \wBIn89[30] , \wBIn89[29] , \wRegInA77[12] , \wAMid117[19] , 
        \wRegInA54[23] , \wRegInA21[13] , \wRegInB84[14] , \wRegInA34[27] , 
        \wRegInA41[17] , \ScanLink41[5] , \wRegInA62[26] , \wRegInB91[20] , 
        \wRegInA17[16] , \ScanLink0[9] , \ScanLink168[26] , \ScanLink90[24] , 
        \ScanLink162[8] , \wBMid67[7] , \wAIn73[23] , \wBMid99[10] , 
        \wBIn114[0] , \ScanLink93[3] , \wRegInB61[4] , \ScanLink108[22] , 
        \ScanLink85[10] , \wRegInA99[14] , \wAMid68[28] , \wRegInB49[23] , 
        \wAIn25[22] , \wAIn50[12] , \ScanLink118[0] , \wAMid68[31] , 
        \wAIn30[16] , \wAIn45[26] , \ScanLink26[2] , \wAIn66[17] , 
        \wRegInB29[27] , \wBMid34[23] , \ScanLink223[27] , \ScanLink186[20] , 
        \wBIn4[3] , \wAMid4[10] , \wBMid17[12] , \wBMid41[13] , 
        \ScanLink256[17] , \ScanLink200[16] , \wAIn107[8] , \wBIn6[30] , 
        \wBIn6[29] , \wBMid5[31] , \wBMid5[28] , \wBMid62[22] , \wRegInA66[6] , 
        \ScanLink28[23] , \wBMid77[16] , \wRegInA102[31] , \wRegInA121[19] , 
        \ScanLink215[22] , \ScanLink48[27] , \wBMid21[17] , \wRegInA102[28] , 
        \ScanLink236[13] , \ScanLink193[14] , \wAMid16[14] , \wBIn19[13] , 
        \wBMid18[2] , \wBIn28[3] , \wBMid54[27] , \wAIn82[9] , \wBMid99[23] , 
        \wRegInB108[4] , \ScanLink243[23] , \wRegInA65[5] , \ScanLink168[15] , 
        \ScanLink108[11] , \ScanLink90[17] , \ScanLink85[23] , \wBMid64[4] , 
        \wAMid93[30] , \wAIn119[4] , \wRegInA34[14] , \wRegInA41[24] , 
        \wRegInB91[13] , \wBMid120[9] , \wAIn88[22] , \wRegInA17[25] , 
        \wRegInA62[15] , \wAMid93[29] , \wRegInA21[20] , \wRegInA77[21] , 
        \wRegInB84[27] , \wRegInB116[8] , \wRegInA54[10] , \ScanLink25[1] , 
        \wRegInA92[18] , \wAMid63[24] , \wAMid20[11] , \wAMid35[25] , 
        \wAMid40[15] , \wBIn54[5] , \ScanLink167[5] , \wAMid55[21] , 
        \ScanLink59[7] , \wAIn31[6] , \wAMid71[2] , \wAMid76[10] , 
        \wRegInA126[3] , \wBIn79[17] , \wRegInB64[9] , \ScanLink207[0] , 
        \wBIn86[3] , \wAIn126[29] , \wRegInA9[6] , \wAIn105[18] , 
        \wAIn126[30] , \wRegInA19[3] , \wAIn32[5] , \wBIn85[0] , 
        \wRegInB127[24] , \wRegInB79[6] , \wRegInA109[24] , \ScanLink44[8] , 
        \ScanLink198[18] , \ScanLink5[4] , \ScanLink179[9] , \wRegInB5[25] , 
        \wAMid72[1] , \wRegInB104[15] , \wRegInA3[20] , \wRegInB111[21] , 
        \ScanLink116[29] , \ScanLink6[7] , \ScanLink163[19] , 
        \ScanLink140[31] , \ScanLink135[18] , \ScanLink116[30] , 
        \ScanLink88[2] , \wAMid15[6] , \wAIn55[2] , \wBIn57[6] , 
        \wAMid109[12] , \ScanLink164[6] , \ScanLink140[28] , \wBIn82[16] , 
        \wBIn97[22] , \wRegInA69[19] , \wAMid98[25] , \wBMid110[23] , 
        \wBMid105[17] , \ScanLink204[3] , \ScanLink7[24] , \wBMid126[26] , 
        \wRegInA125[0] , \ScanLink36[28] , \wBMid61[9] , \ScanLink60[30] , 
        \ScanLink43[18] , \ScanLink36[31] , \ScanLink15[19] , \wBMid125[4] , 
        \wRegInA109[17] , \ScanLink60[29] , \wAMid16[27] , \wAIn18[18] , 
        \wAMid20[22] , \wRegInB113[5] , \ScanLink228[18] , \ScanLink103[1] , 
        \wBIn30[1] , \wRegInB57[31] , \wAMid55[12] , \wAIn101[6] , 
        \wRegInB74[19] , \wAIn87[4] , \wRegInA60[8] , \wBIn19[20] , 
        \wAMid76[23] , \wRegInB57[28] , \wBIn79[24] , \wRegInB22[18] , 
        \wAMid16[5] , \wBIn33[2] , \wAMid35[16] , \wAMid63[17] , \wAMid40[26] , 
        \wBIn82[25] , \wAIn96[29] , \wBMid105[24] , \wAIn84[7] , \wAIn96[30] , 
        \wAIn102[5] , \wBMid126[15] , \ScanLink100[2] , \wBIn97[11] , 
        \wAMid109[21] , \wAMid98[16] , \wBMid110[10] , \wBMid126[7] , 
        \ScanLink7[17] , \wRegInA3[13] , \wAIn56[1] , \wBMid87[31] , 
        \wBMid87[28] , \wAIn99[8] , \wRegInB111[12] , \wBIn86[14] , 
        \wAMid89[13] , \wRegInB127[17] , \wRegInB5[16] , \wRegInB104[26] , 
        \wRegInB110[6] , \ScanLink244[1] , \wAIn92[18] , \wBMid101[15] , 
        \wRegInB27[8] , \wAMid118[24] , \wBMid122[24] , \wBIn17[4] , 
        \wAIn126[3] , \ScanLink124[4] , \wAMid31[0] , \wAMid32[3] , 
        \wAIn72[7] , \wBMid83[19] , \wBIn93[20] , \wBMid114[21] , 
        \wRegInA88[4] , \ScanLink3[26] , \wRegInA7[22] , \wRegInB115[23] , 
        \wRegInB1[27] , \wRegInB123[26] , \wBMid89[5] , \wRegInB100[17] , 
        \wBMid102[1] , \wBMid78[18] , \ScanLink47[29] , \ScanLink32[19] , 
        \wBMid101[2] , \wRegInB39[4] , \ScanLink64[18] , \ScanLink11[31] , 
        \ScanLink47[30] , \ScanLink11[28] , \wRegInA118[12] , \wAIn71[4] , 
        \wRegInA59[1] , \wRegInA96[8] , \wBIn2[18] , \wBIn7[0] , \wAMid12[16] , 
        \wAMid24[13] , \wAMid51[23] , \wRegInB26[30] , \ScanLink19[5] , 
        \wBMid58[0] , \wAIn69[19] , \wAMid72[12] , \wRegInB70[28] , 
        \ScanLink247[2] , \wRegInB26[29] , \wRegInB53[19] , \wRegInB70[31] , 
        \wAMid67[26] , \wBIn68[21] , \wBMid97[9] , \wBIn14[7] , \wAIn125[0] , 
        \wAMid31[27] , \wAMid44[17] , \ScanLink127[7] , \wRegInB1[14] , 
        \wRegInB123[15] , \wRegInB100[24] , \wBMid22[8] , \ScanLink167[28] , 
        \wAIn0[4] , \wAMid0[21] , \wAIn4[25] , \wBIn9[14] , \wAMid12[25] , 
        \wAIn16[3] , \wAMid56[7] , \wRegInA7[11] , \wRegInB115[10] , 
        \ScanLink131[30] , \ScanLink192[6] , \ScanLink112[18] , 
        \ScanLink167[31] , \ScanLink144[19] , \wBIn73[0] , \wAMid84[1] , 
        \wBIn86[27] , \wAMid89[20] , \wBIn93[13] , \wAMid114[9] , 
        \ScanLink131[29] , \wBMid114[12] , \wRegInA101[6] , \ScanLink220[5] , 
        \ScanLink3[15] , \wRegInA18[18] , \wBMid101[26] , \wBMid122[17] , 
        \wAMid109[6] , \wAMid118[17] , \wRegInA23[9] , \ScanLink140[0] , 
        \ScanLink223[6] , \wAIn15[0] , \wAMid24[20] , \wAMid31[14] , 
        \wAMid67[15] , \wBIn68[12] , \wRegInA96[29] , \wAMid44[24] , 
        \wRegInA96[30] , \wRegInA102[5] , \ScanLink143[3] , \wAMid51[10] , 
        \wBIn70[3] , \wAMid72[21] , \wAMid87[2] , \wAIn101[30] , \wAIn101[29] , 
        \wAIn122[18] , \wRegInB92[9] , \wRegInA118[21] , \ScanLink191[5] , 
        \wAMid55[4] , \wRegInB21[6] , \ScanLink179[10] , \ScanLink81[12] , 
        \wAIn17[16] , \wAMid19[30] , \wAMid19[29] , \wAMid29[2] , \wBMid92[4] , 
        \ScanLink94[26] , \wBMid119[0] , \wBMid40[2] , \wAIn69[6] , 
        \ScanLink119[14] , \wBMid88[26] , \wAMid97[18] , \wRegInA30[25] , 
        \wRegInA41[3] , \wRegInA45[15] , \wRegInA66[24] , \wRegInB95[22] , 
        \ScanLink8[19] , \wAIn99[27] , \wRegInA13[14] , \wAIn74[9] , 
        \wRegInA50[21] , \wRegInA73[10] , \wRegInA25[11] , \wRegInB80[16] , 
        \wRegInA93[5] , \wAIn77[12] , \wRegInB38[22] , \wAIn21[13] , 
        \wAIn34[27] , \wAIn54[23] , \wAIn41[17] , \wRegInA90[6] , \wBMid43[1] , 
        \wAIn62[26] , \wRegInB58[26] , \wRegInA88[11] , \ScanLink252[26] , 
        \wBMid8[5] , \wBMid45[22] , \wBMid30[12] , \ScanLink227[16] , 
        \ScanLink182[11] , \wBMid66[13] , \wRegInB22[5] , \wAMid0[12] , 
        \wBMid1[19] , \wBIn12[9] , \wBMid13[23] , \ScanLink204[27] , 
        \ScanLink59[22] , \wAIn4[16] , \wBIn9[27] , \wBMid24[6] , 
        \wBMid25[26] , \wBMid50[16] , \wBMid73[27] , \wRegInA42[0] , 
        \ScanLink121[9] , \ScanLink39[26] , \wRegInA125[28] , 
        \ScanLink211[13] , \wBMid91[7] , \ScanLink247[12] , \wRegInA106[19] , 
        \wBIn68[1] , \wAIn99[14] , \wAMid113[31] , \wRegInA125[31] , 
        \ScanLink232[22] , \ScanLink197[25] , \wRegInB97[4] , \wAMid113[28] , 
        \wRegInA73[23] , \wRegInA25[22] , \wRegInB80[25] , \wRegInA50[12] , 
        \ScanLink65[3] , \wAMid112[7] , \wRegInA30[16] , \wRegInA38[8] , 
        \wRegInA45[26] , \wRegInB95[11] , \ScanLink194[8] , \wRegInA13[27] , 
        \wAMid50[9] , \wRegInA66[17] , \ScanLink119[27] , \ScanLink94[15] , 
        \wBMid25[15] , \wBMid39[9] , \wBMid88[15] , \wRegInB45[2] , 
        \wRegInA25[7] , \wRegInA107[8] , \ScanLink189[7] , \wBMid73[14] , 
        \wRegInB5[2] , \ScanLink179[23] , \ScanLink211[20] , \ScanLink81[21] , 
        \ScanLink39[15] , \wBMid30[21] , \wBMid50[25] , \wRegInB46[1] , 
        \ScanLink232[11] , \ScanLink225[8] , \ScanLink197[16] , \wRegInB89[8] , 
        \ScanLink247[21] , \ScanLink227[25] , \ScanLink182[22] , \wRegInB6[1] , 
        \ScanLink252[15] , \wBMid13[10] , \wBMid45[11] , \ScanLink204[14] , 
        \ScanLink59[11] , \wBMid0[20] , \wAMid2[9] , \wAMid9[2] , \wBIn20[18] , 
        \wAIn41[24] , \wBMid66[20] , \wRegInA26[4] , \wBIn55[28] , 
        \wBIn115[31] , \ScanLink66[0] , \wAIn34[14] , \wRegInA119[4] , 
        \wBIn55[31] , \wBIn76[19] , \wAIn62[15] , \wAIn17[25] , \wBIn115[28] , 
        \wRegInA88[22] , \ScanLink238[7] , \wBMid19[25] , \wAIn21[20] , 
        \wBMid27[5] , \wRegInB38[11] , \wRegInB58[15] , \wRegInB94[7] , 
        \wAIn54[10] , \wAIn77[21] , \ScanLink158[2] , \wAMid111[4] , 
        \wAIn100[23] , \ScanLink70[4] , \ScanLink53[24] , \ScanLink26[14] , 
        \wBMid31[1] , \wAIn123[12] , \wRegInB82[3] , \ScanLink188[17] , 
        \ScanLink70[15] , \ScanLink10[11] , \wBMid79[21] , \ScanLink238[24] , 
        \ScanLink65[21] , \wAMid107[0] , \wAIn115[17] , \ScanLink33[20] , 
        \wRegInB11[15] , \wRegInB64[25] , \ScanLink46[10] , \wBIn3[21] , 
        \wBIn3[12] , \wAIn18[5] , \wAMid58[1] , \wAIn68[20] , \wBIn69[18] , 
        \wRegInB32[24] , \wRegInB47[14] , \wRegInB50[5] , \wRegInA97[23] , 
        \wAMid97[8] , \wRegInB52[20] , \wRegInB27[10] , \wRegInA82[17] , 
        \wBIn60[9] , \wRegInB71[11] , \ScanLink153[9] , \wBMid32[2] , 
        \wBMid82[20] , \wAIn86[15] , \wBIn125[1] , \wRegInA30[0] , 
        \wBIn92[19] , \wAIn93[21] , \wBMid115[18] , \wBIn126[2] , 
        \wRegInA19[12] , \wRegInB53[6] , \wRegInA33[3] , \wBMid97[14] , 
        \wRegInA79[16] , \wRegInB81[0] , \ScanLink173[16] , \ScanLink150[27] , 
        \ScanLink106[26] , \ScanLink125[17] , \ScanLink73[7] , 
        \ScanLink145[13] , \wAMid104[3] , \ScanLink130[23] , \wBIn19[2] , 
        \wAMid25[19] , \wAMid50[30] , \wAIn68[13] , \wAMid89[4] , 
        \ScanLink166[22] , \ScanLink113[12] , \wAMid50[29] , \wAMid73[18] , 
        \wRegInB27[23] , \wRegInA82[24] , \wRegInB34[1] , \wRegInB52[13] , 
        \wBMid79[12] , \wBMid87[3] , \wRegInB11[26] , \wRegInB71[22] , 
        \wRegInB32[17] , \wRegInA54[4] , \wRegInB64[16] , \wRegInA97[10] , 
        \wRegInB127[9] , \wRegInB47[27] , \ScanLink238[17] , \ScanLink65[12] , 
        \ScanLink10[22] , \ScanLink46[23] , \ScanLink14[0] , \wAIn115[24] , 
        \ScanLink33[13] , \wBMid19[16] , \ScanLink53[17] , \wBMid55[5] , 
        \wAIn100[10] , \wBMid111[8] , \wRegInA86[2] , \ScanLink26[27] , 
        \ScanLink188[24] , \wBMid82[13] , \wAIn123[21] , \wRegInA119[18] , 
        \ScanLink70[26] , \wRegInA6[31] , \ScanLink17[3] , \wRegInA6[28] , 
        \wRegInB114[30] , \ScanLink130[10] , \ScanLink145[20] , 
        \wRegInB114[29] , \ScanLink249[4] , \ScanLink113[21] , \wAMid4[7] , 
        \wBIn9[6] , \wAMid22[9] , \wBMid56[6] , \ScanLink166[11] , 
        \ScanLink106[15] , \ScanLink173[25] , \wBIn17[17] , \wAMid18[10] , 
        \wBIn21[12] , \wBIn54[22] , \wBIn77[13] , \wBMid84[0] , \wAMid88[19] , 
        \wAIn93[12] , \wBMid97[27] , \ScanLink129[1] , \ScanLink125[24] , 
        \wRegInA85[1] , \ScanLink150[14] , \wRegInB37[2] , \wRegInA19[21] , 
        \wRegInA79[25] , \wAIn86[26] , \wRegInA57[7] , \wAMid78[14] , 
        \wBIn114[22] , \wRegInA89[28] , \wRegInA89[31] , \wBIn34[26] , 
        \wBIn41[16] , \wBIn122[27] , \ScanLink148[8] , \ScanLink187[1] , 
        \wAMid43[0] , \wBIn62[27] , \wBIn101[16] , \wRegInA107[20] , 
        \wRegInB99[2] , \ScanLink235[2] , \wRegInA114[1] , \wRegInA124[11] , 
        \wBMid0[13] , \wAMid1[18] , \wBIn66[7] , \ScanLink183[31] , 
        \ScanLink155[7] , \wAMid7[4] , \wAMid91[6] , \wRegInA112[14] , 
        \ScanLink183[28] , \wRegInA117[2] , \ScanLink68[6] , \ScanLink236[1] , 
        \wBMid12[30] , \wBMid12[29] , \wBMid29[3] , \wRegInB55[8] , 
        \wAMid40[3] , \wBIn65[4] , \wAMid92[5] , \ScanLink178[29] , 
        \wAMid83[15] , \wAMid112[22] , \ScanLink178[30] , \ScanLink156[4] , 
        \wRegInA24[31] , \wRegInA24[28] , \ScanLink75[9] , \wRegInA51[18] , 
        \wRegInA72[30] , \wAMid124[27] , \wRegInB48[7] , \wRegInA72[29] , 
        \wBMid44[31] , \wAMid96[21] , \wBIn99[26] , \ScanLink9[20] , 
        \wAMid107[16] , \wRegInB8[7] , \ScanLink184[2] , \wRegInA28[2] , 
        \wBMid67[19] , \wBMid44[28] , \ScanLink251[6] , \ScanLink58[28] , 
        \wRegInA112[27] , \wBMid31[18] , \ScanLink58[31] , \wRegInA107[13] , 
        \ScanLink246[18] , \ScanLink233[28] , \wAIn3[7] , \wBMid4[22] , 
        \wBMid5[0] , \wBIn17[24] , \wAMid18[23] , \wAIn20[19] , 
        \wRegInA124[22] , \ScanLink131[3] , \ScanLink233[31] , 
        \ScanLink210[19] , \wBIn34[15] , \wBIn41[25] , \wBIn122[14] , 
        \wRegInB39[31] , \wAIn55[29] , \wBMid6[3] , \wBIn21[21] , \wAMid27[4] , 
        \wAIn55[30] , \wBIn62[14] , \wAIn76[18] , \wBIn101[25] , 
        \wRegInB39[28] , \wRegInB121[7] , \wBIn77[20] , \wBMid117[6] , 
        \wAMid78[27] , \wBIn114[11] , \wBIn54[11] , \wAIn67[0] , \wAMid96[12] , 
        \wBIn99[15] , \ScanLink9[13] , \wRegInB94[31] , \wRegInB122[4] , 
        \wBMid16[18] , \wAMid24[7] , \wBMid50[8] , \wAIn64[3] , \wAMid107[25] , 
        \wAMid124[14] , \wRegInB94[28] , \wAMid83[26] , \wAMid112[11] , 
        \wBMid114[5] , \wBIn25[6] , \wBIn38[9] , \wAMid39[8] , \wRegInA51[9] , 
        \ScanLink252[5] , \ScanLink132[0] , \ScanLink80[18] , \wAIn89[28] , 
        \wAMid92[23] , \wAMid120[25] , \wRegInB90[19] , \wAIn40[5] , 
        \wAMid103[14] , \wRegInA68[0] , \wBMid69[1] , \wAMid87[17] , 
        \wBIn88[10] , \wAIn89[31] , \wAMid116[20] , \wRegInB106[2] , 
        \wBMid98[30] , \ScanLink84[29] , \wBIn26[5] , \wBMid35[30] , 
        \wAIn92[3] , \wBMid98[29] , \wAIn114[1] , \ScanLink116[6] , 
        \wRegInA9[26] , \ScanLink84[30] , \ScanLink28[4] , \ScanLink115[5] , 
        \wAIn117[2] , \wBMid35[29] , \wBMid63[28] , \wAIn91[0] , 
        \ScanLink29[29] , \wBMid40[19] , \wBMid63[31] , \wRegInA116[16] , 
        \ScanLink29[30] , \wRegInB16[9] , \wRegInA103[22] , \ScanLink237[19] , 
        \ScanLink214[31] , \wRegInA120[13] , \ScanLink242[29] , 
        \ScanLink214[28] , \wBIn13[15] , \wAIn24[28] , \wBIn30[24] , 
        \wAIn43[6] , \wBIn45[14] , \wAIn51[18] , \wBIn126[25] , 
        \ScanLink242[30] , \wAIn72[30] , \wRegInB48[30] , \wBIn66[25] , 
        \wAMid69[22] , \wBIn105[14] , \wAIn72[29] , \wRegInB48[29] , 
        \wAIn24[31] , \wAIn24[1] , \wBIn25[10] , \wBIn50[20] , \wBIn73[11] , 
        \wBIn110[20] , \wRegInB105[1] , \ScanLink36[8] , \wBIn41[2] , 
        \ScanLink172[2] , \wBIn93[4] , \wRegInA9[15] , \ScanLink212[7] , 
        \ScanLink109[31] , \ScanLink109[28] , \ScanLink83[9] , \wRegInA55[29] , 
        \wBIn88[23] , \wAMid116[13] , \wBIn119[5] , \wRegInA20[19] , 
        \wBMid13[9] , \wAMid64[5] , \wAMid87[24] , \wRegInA55[30] , 
        \wRegInA76[18] , \wAMid92[10] , \wAMid103[27] , \wAMid120[16] , 
        \wRegInA0[3] , \wBIn1[27] , \wAIn5[9] , \wBMid4[11] , \wBIn13[26] , 
        \wBIn25[23] , \wAMid67[6] , \wBIn73[22] , \wBIn110[13] , \wAIn27[2] , 
        \wBIn50[13] , \wBIn90[7] , \wAMid125[8] , \wBIn30[17] , \wBIn45[27] , 
        \wBIn126[16] , \wBIn66[16] , \wAMid69[11] , \wBIn105[27] , 
        \wRegInA103[11] , \wAMid5[30] , \wAMid5[29] , \wBIn42[1] , 
        \wBIn107[9] , \ScanLink171[1] , \wRegInA12[8] , \wRegInA120[20] , 
        \ScanLink211[4] , \wBIn7[10] , \wBMid72[0] , \wBMid86[22] , 
        \wRegInA116[25] , \ScanLink187[19] , \ScanLink141[11] , \wAIn89[2] , 
        \ScanLink134[21] , \wAMid18[3] , \wAIn19[12] , \wAMid21[31] , 
        \wBIn23[8] , \wBMid93[16] , \wRegInA2[19] , \ScanLink162[20] , 
        \wRegInB110[18] , \ScanLink177[14] , \ScanLink117[10] , 
        \ScanLink154[25] , \ScanLink102[24] , \ScanLink121[15] , 
        \ScanLink33[5] , \wAIn82[17] , \wAIn97[23] , \wRegInA73[1] , 
        \ScanLink110[8] , \wRegInA68[20] , \wRegInB13[4] , \wAMid77[29] , 
        \wRegInB56[22] , \wRegInB23[12] , \wRegInA86[15] , \wAMid21[28] , 
        \wAIn45[8] , \wAMid54[18] , \wAIn58[7] , \wRegInB75[13] , 
        \wAMid77[30] , \wBMid71[3] , \wAIn79[16] , \wRegInB10[7] , 
        \wRegInB15[17] , \wRegInB60[27] , \wRegInA70[2] , \wRegInB36[26] , 
        \wRegInB43[16] , \wRegInA93[21] , \ScanLink249[16] , \ScanLink14[13] , 
        \wAIn111[15] , \ScanLink199[21] , \ScanLink61[23] , \ScanLink37[22] , 
        \ScanLink42[12] , \wBMid68[17] , \wAIn104[21] , \ScanLink30[6] , 
        \ScanLink22[16] , \wAIn82[24] , \wBIn96[28] , \wBMid111[29] , 
        \wAIn127[10] , \ScanLink57[26] , \wRegInA7[0] , \wRegInA68[13] , 
        \ScanLink229[12] , \ScanLink74[17] , \wBIn88[5] , \wBIn96[31] , 
        \wAMid108[18] , \wBMid111[30] , \wRegInA17[5] , \wAIn97[10] , 
        \wBIn102[4] , \wRegInB77[0] , \ScanLink214[9] , \ScanLink85[7] , 
        \ScanLink102[17] , \wBIn7[23] , \wBMid16[4] , \wBMid86[11] , 
        \wBMid93[25] , \ScanLink177[27] , \ScanLink169[3] , \ScanLink121[26] , 
        \wAMid120[5] , \ScanLink154[16] , \ScanLink57[1] , \ScanLink209[6] , 
        \ScanLink141[22] , \ScanLink134[12] , \ScanLink98[8] , 
        \ScanLink117[23] , \wAMid8[12] , \wBMid15[7] , \wBIn59[0] , 
        \ScanLink162[13] , \wBMid68[24] , \wBIn96[9] , \wAIn104[12] , 
        \ScanLink57[15] , \ScanLink22[25] , \wAMid123[6] , \ScanLink229[21] , 
        \wBIn18[19] , \wAMid61[8] , \wAIn127[23] , \ScanLink74[24] , 
        \wAIn79[25] , \wBIn101[7] , \wAIn111[26] , \ScanLink249[25] , 
        \ScanLink199[12] , \ScanLink61[10] , \ScanLink14[20] , \ScanLink54[2] , 
        \ScanLink42[21] , \ScanLink37[11] , \wRegInA14[6] , \wRegInB15[24] , 
        \wRegInB60[14] , \wRegInB36[15] , \wRegInA93[12] , \wRegInA4[3] , 
        \wRegInB43[25] , \wAIn19[21] , \wRegInB23[21] , \wRegInA86[26] , 
        \wBIn28[18] , \wAIn29[20] , \wRegInB13[20] , \wRegInB56[11] , 
        \wRegInB74[3] , \wRegInB75[20] , \ScanLink86[4] , \ScanLink8[1] , 
        \wAIn49[24] , \wRegInB14[7] , \wRegInB25[25] , \wRegInB30[11] , 
        \wRegInB66[10] , \wRegInA74[2] , \wRegInB45[21] , \wRegInA95[16] , 
        \wRegInA80[22] , \wRegInB50[15] , \ScanLink29[9] , \wRegInB73[24] , 
        \wBIn39[4] , \ScanLink51[11] , \wAIn108[3] , \wBMid38[21] , 
        \wAIn41[8] , \wAIn102[16] , \ScanLink24[21] , \wBMid58[25] , 
        \wBMid75[3] , \ScanLink72[20] , \wAIn121[27] , \ScanLink67[14] , 
        \ScanLink12[24] , \wBMid76[0] , \wAIn117[22] , \ScanLink219[20] , 
        \ScanLink44[25] , \ScanLink34[6] , \ScanLink31[15] , \wBMid80[15] , 
        \wBMid95[21] , \ScanLink171[23] , \ScanLink104[13] , \ScanLink89[21] , 
        \ScanLink152[12] , \ScanLink127[22] , \ScanLink109[7] , 
        \ScanLink132[16] , \ScanLink164[17] , \ScanLink147[26] , 
        \ScanLink37[5] , \ScanLink111[27] , \wAMid8[21] , \wBMid9[19] , 
        \wBMid11[7] , \wBIn27[8] , \wAIn84[20] , \wBIn85[18] , \wBMid121[28] , 
        \wRegInA38[16] , \wRegInA58[12] , \wRegInA77[1] , \ScanLink114[8] , 
        \wRegInB88[25] , \wAIn91[14] , \wBMid102[19] , \wRegInB17[4] , 
        \wBMid121[31] , \wRegInB119[3] , \wBMid58[16] , \ScanLink12[17] , 
        \wAMid65[8] , \wBIn92[9] , \wAIn117[11] , \ScanLink67[27] , 
        \wBIn118[8] , \ScanLink31[26] , \ScanLink219[13] , \ScanLink44[16] , 
        \ScanLink24[12] , \wBMid38[12] , \wAIn102[25] , \wAIn121[14] , 
        \ScanLink51[22] , \ScanLink50[2] , \wAMid78[7] , \wRegInB50[26] , 
        \ScanLink72[13] , \wRegInB25[16] , \wRegInA80[11] , \wAMid0[7] , 
        \wAIn1[9] , \wAMid11[30] , \wAMid32[18] , \wAIn38[3] , \wBIn105[7] , 
        \wRegInA10[6] , \wRegInB73[17] , \wAIn49[17] , \ScanLink82[4] , 
        \wAMid11[29] , \wAIn29[13] , \wAMid47[28] , \wRegInB66[23] , 
        \wRegInB13[13] , \wAMid47[31] , \wAMid64[19] , \wRegInB45[12] , 
        \wBMid80[26] , \wAIn84[13] , \wAIn91[27] , \wBIn106[4] , 
        \wRegInA13[5] , \wRegInB30[22] , \wRegInB70[3] , \wRegInA58[21] , 
        \wRegInA95[25] , \wRegInB88[16] , \wRegInA3[0] , \ScanLink0[19] , 
        \wAMid124[5] , \wRegInA38[25] , \wRegInB73[0] , \ScanLink210[9] , 
        \ScanLink81[7] , \ScanLink147[15] , \ScanLink132[25] , 
        \ScanLink164[24] , \wBIn1[14] , \wBMid2[26] , \wBMid2[15] , 
        \wBMid12[4] , \wBIn22[5] , \wBMid95[12] , \wRegInB2[18] , 
        \wRegInB103[28] , \ScanLink171[10] , \ScanLink111[14] , 
        \ScanLink89[12] , \ScanLink104[20] , \ScanLink152[21] , 
        \ScanLink53[1] , \wRegInB103[31] , \wRegInA105[15] , \wRegInB120[19] , 
        \ScanLink194[29] , \ScanLink127[11] , \ScanLink111[5] , \wAIn113[2] , 
        \wAIn4[4] , \wAIn7[30] , \wAIn95[0] , \ScanLink194[30] , 
        \wRegInA126[24] , \wAIn7[29] , \wAIn109[29] , \wBIn15[22] , 
        \wBIn23[27] , \wBIn75[26] , \wAIn109[30] , \wBIn116[17] , 
        \wRegInB12[9] , \wRegInA110[21] , \wBIn36[13] , \wAIn47[6] , 
        \wBIn56[17] , \wAMid59[10] , \wAMid39[14] , \wBIn43[23] , 
        \ScanLink32[8] , \wBIn120[12] , \wBMid17[9] , \wBIn21[6] , \wAIn44[5] , 
        \wBIn60[12] , \wBIn103[23] , \wRegInB101[1] , \wAMid110[17] , 
        \wAMid81[20] , \wAMid94[14] , \wBMid109[26] , \wAMid105[23] , 
        \wAMid126[12] , \wRegInA65[28] , \wRegInA10[18] , \wRegInA33[30] , 
        \wRegInA46[19] , \wRegInA65[31] , \wRegInB102[2] , \wRegInA33[29] , 
        \wAIn23[2] , \wBIn36[20] , \wBIn43[10] , \wAIn96[3] , \wAIn110[1] , 
        \ScanLink112[6] , \wRegInB9[14] , \wRegInB108[24] , \ScanLink139[30] , 
        \ScanLink139[29] , \wBIn94[7] , \wBIn120[21] , \wAMid39[27] , 
        \wAMid121[8] , \wBIn60[21] , \wAIn14[30] , \wAIn14[29] , \wBIn15[11] , 
        \wAMid63[6] , \wBIn103[10] , \wAIn42[31] , \wBIn75[15] , \wBIn116[24] , 
        \wAIn61[19] , \wRegInB78[31] , \wBIn23[14] , \wAIn42[28] , 
        \ScanLink99[5] , \wBIn56[24] , \wAMid59[23] , \wRegInB78[28] , 
        \wBMid26[19] , \wAIn37[18] , \wBIn46[1] , \wBIn89[8] , 
        \ScanLink224[30] , \wBIn103[9] , \ScanLink207[18] , \ScanLink175[1] , 
        \wRegInA16[8] , \wRegInA110[12] , \ScanLink251[19] , \ScanLink224[29] , 
        \ScanLink215[4] , \wBMid53[29] , \wRegInA105[26] , \wBMid70[18] , 
        \wRegInA126[17] , \ScanLink19[28] , \wAMid3[4] , \wAIn7[7] , 
        \wBIn45[2] , \wBMid53[30] , \wRegInB9[27] , \wRegInB108[17] , 
        \ScanLink19[31] , \ScanLink176[2] , \ScanLink216[7] , \ScanLink87[9] , 
        \ScanLink48[0] , \ScanLink97[19] , \wAIn20[1] , \wAMid60[5] , 
        \wAMid94[27] , \wAMid126[21] , \wBIn97[4] , \wAMid105[10] , 
        \wAMid81[13] , \wAMid110[24] , \wRegInB83[29] , \wRegInB68[1] , 
        \wRegInB83[30] , \wBMid109[15] , \ScanLink232[1] , \wAIn10[18] , 
        \wBIn11[20] , \wAIn19[8] , \wBIn61[4] , \wRegInB51[8] , 
        \wRegInA113[2] , \ScanLink152[4] , \ScanLink93[31] , \wBIn32[11] , 
        \wAMid44[3] , \wAMid85[22] , \wAMid90[16] , \wAMid96[5] , 
        \wRegInB119[12] , \ScanLink93[28] , \wBMid118[10] , \wAMid101[21] , 
        \wAMid122[10] , \ScanLink71[9] , \wAMid114[15] , \wRegInB87[18] , 
        \ScanLink180[2] , \wBIn47[21] , \wAMid48[26] , \wBIn124[10] , 
        \wAIn33[30] , \wBIn64[10] , \wBIn107[21] , \wBIn27[25] , \wAMid28[22] , 
        \wAIn33[29] , \wAMid47[0] , \wAIn65[28] , \wAMid88[9] , \wBIn112[15] , 
        \wBIn71[24] , \ScanLink183[1] , \wAIn46[19] , \wBIn52[15] , 
        \wAIn65[31] , \wRegInA110[1] , \ScanLink255[31] , \ScanLink203[29] , 
        \wBMid1[0] , \wAIn3[18] , \wBMid2[3] , \wBMid6[17] , \wBMid22[28] , 
        \wBMid57[18] , \wRegInA114[23] , \ScanLink255[28] , \ScanLink231[2] , 
        \ScanLink220[18] , \ScanLink203[30] , \wBMid74[30] , \wAMid95[6] , 
        \wRegInA101[17] , \wBIn62[7] , \ScanLink151[7] , \ScanLink68[29] , 
        \wBMid22[31] , \wBMid74[29] , \wAMid118[1] , \wRegInA122[26] , 
        \wAMid114[26] , \ScanLink68[30] , \wRegInB28[3] , \wRegInB126[4] , 
        \wBMid6[24] , \wAMid20[7] , \wBMid54[8] , \wAMid85[11] , \wBMid110[5] , 
        \wAMid122[23] , \wRegInA14[29] , \wAMid90[25] , \wBMid118[23] , 
        \wBMid49[7] , \wAIn60[3] , \wAMid101[12] , \wRegInA42[31] , 
        \wRegInA61[19] , \wRegInA14[30] , \wRegInA37[18] , \wRegInA42[28] , 
        \wRegInA48[6] , \wRegInB119[21] , \ScanLink148[28] , \ScanLink256[5] , 
        \ScanLink148[31] , \wRegInA55[9] , \ScanLink136[0] , \wRegInA101[24] , 
        \ScanLink255[6] , \ScanLink190[18] , \wRegInA122[15] , \wRegInA99[3] , 
        \ScanLink135[3] , \wRegInA114[10] , \wBIn71[17] , \wBIn112[26] , 
        \ScanLink248[9] , \wBIn5[25] , \wBIn11[13] , \wBIn27[16] , 
        \wAMid28[11] , \wBIn52[26] , \wRegInB125[7] , \wBIn32[22] , 
        \wBIn47[12] , \wAMid48[15] , \wBIn124[23] , \wAIn63[0] , \wBIn64[23] , 
        \wBMid113[6] , \wBMid98[2] , \wBIn107[12] , \wAMid23[4] , \wAIn80[22] , 
        \wAIn95[16] , \wRegInA29[20] , \wRegInB57[6] , \wBMid84[17] , 
        \wBIn122[2] , \wRegInB99[13] , \ScanLink4[28] , \wRegInA37[3] , 
        \ScanLink4[31] , \wRegInA49[24] , \ScanLink136[14] , \wRegInB85[0] , 
        \wRegInA108[3] , \ScanLink143[24] , \ScanLink77[7] , \ScanLink229[0] , 
        \ScanLink115[25] , \ScanLink160[15] , \ScanLink98[17] , \wAMid6[9] , 
        \wAIn8[14] , \wBMid29[17] , \wBMid36[2] , \wBMid91[23] , 
        \wRegInB6[30] , \wRegInB107[19] , \wRegInB124[31] , \ScanLink175[21] , 
        \ScanLink100[11] , \wAMid100[3] , \wRegInB6[29] , \wRegInB124[28] , 
        \ScanLink149[5] , \ScanLink123[20] , \ScanLink156[10] , 
        \ScanLink63[16] , \wBMid35[1] , \wBIn79[6] , \wAIn113[20] , 
        \wRegInB86[3] , \ScanLink16[26] , \ScanLink74[4] , \ScanLink40[27] , 
        \ScanLink55[13] , \ScanLink35[17] , \wAMid103[0] , \ScanLink208[16] , 
        \wAIn106[14] , \ScanLink20[23] , \ScanLink76[22] , \wBMid49[13] , 
        \wAIn125[25] , \wRegInA84[20] , \wAMid15[18] , \wAMid36[29] , 
        \wAIn38[16] , \wRegInB21[27] , \wRegInB54[17] , \wRegInB54[5] , 
        \wRegInB77[26] , \wAMid43[19] , \wAIn58[12] , \wAMid60[31] , 
        \wBIn64[9] , \wRegInB17[22] , \ScanLink198[0] , \ScanLink157[9] , 
        \wAMid60[28] , \wBIn121[1] , \wRegInA34[0] , \wRegInB62[12] , 
        \wAMid93[8] , \wRegInB34[13] , \wRegInA91[14] , \wAMid36[30] , 
        \wRegInB41[23] , \ScanLink175[12] , \ScanLink100[22] , \ScanLink13[3] , 
        \wBIn0[3] , \wAIn2[21] , \wAIn2[12] , \wBIn5[16] , \wBMid84[24] , 
        \wBMid91[10] , \ScanLink156[23] , \wRegInA81[1] , \ScanLink143[17] , 
        \ScanLink123[13] , \ScanLink136[27] , \ScanLink160[26] , \wAIn8[27] , 
        \wAMid26[9] , \wBMid52[6] , \ScanLink115[16] , \ScanLink98[24] , 
        \wAIn38[25] , \wAMid38[5] , \wAIn58[21] , \wAIn80[11] , \wBIn81[30] , 
        \wBMid106[31] , \wBMid125[19] , \wRegInB33[2] , \wRegInA49[17] , 
        \wRegInB99[20] , \wBIn81[29] , \wBMid80[0] , \wRegInA29[13] , 
        \wRegInA53[7] , \wAIn95[25] , \wBMid106[28] , \wRegInB62[21] , 
        \wBMid83[3] , \wBMid108[7] , \wRegInB17[11] , \wRegInB30[1] , 
        \wRegInB41[10] , \ScanLink253[8] , \wRegInB34[20] , \wRegInB54[24] , 
        \wRegInA91[27] , \wBIn119[19] , \wRegInA84[13] , \wRegInB21[14] , 
        \wRegInB77[15] , \wBMid49[20] , \wBIn59[19] , \wRegInA50[4] , 
        \wAIn78[1] , \wAIn106[27] , \ScanLink20[10] , \ScanLink10[0] , 
        \ScanLink208[25] , \ScanLink55[20] , \wBIn10[19] , \wAIn11[21] , 
        \wBMid29[24] , \wBMid51[5] , \wAIn125[16] , \wRegInB123[9] , 
        \ScanLink76[11] , \wBMid115[8] , \ScanLink63[25] , \ScanLink16[15] , 
        \wAIn32[10] , \wAIn47[20] , \wAIn113[13] , \wRegInA82[2] , 
        \ScanLink35[24] , \ScanLink40[14] , \wAIn64[11] , \wBIn33[31] , 
        \wBMid47[1] , \wBIn65[29] , \wAIn71[25] , \wBMid88[8] , \wBIn106[18] , 
        \wBIn125[30] , \wBMid23[11] , \wAIn27[24] , \wBIn33[28] , \wBIn46[18] , 
        \wAIn52[14] , \wBIn65[30] , \wBIn125[29] , \ScanLink138[6] , 
        \wBMid75[10] , \wAIn119[26] , \wRegInB68[14] , \wRegInA94[6] , 
        \ScanLink217[24] , \ScanLink234[15] , \ScanLink191[12] , 
        \ScanLink69[10] , \wBMid36[25] , \wBMid56[21] , \ScanLink241[25] , 
        \wRegInB26[5] , \wBMid43[15] , \wBMid95[7] , \ScanLink221[21] , 
        \ScanLink184[26] , \wAMid6[16] , \wBIn16[9] , \ScanLink254[11] , 
        \wBMid15[14] , \wBMid60[24] , \wRegInA46[0] , \ScanLink202[10] , 
        \ScanLink125[9] , \wBMid43[26] , \wBMid44[2] , \wAIn70[9] , 
        \wBMid96[4] , \wRegInB25[6] , \wRegInA89[9] , \wRegInA45[3] , 
        \ScanLink149[22] , \ScanLink92[11] , \ScanLink18[8] , 
        \ScanLink129[26] , \wAMid100[18] , \wAMid123[30] , \wRegInA23[26] , 
        \wRegInB38[9] , \ScanLink87[25] , \wRegInA75[27] , \wRegInB86[21] , 
        \wRegInA56[16] , \wRegInA36[12] , \wRegInB93[15] , \wRegInA97[5] , 
        \wBMid119[30] , \wAMid123[29] , \wRegInA43[22] , \wBMid119[29] , 
        \wRegInA15[23] , \wRegInA60[13] , \wBIn3[0] , \wAMid6[25] , 
        \wBMid36[16] , \wRegInB42[1] , \wRegInA115[29] , \ScanLink254[22] , 
        \ScanLink221[8] , \ScanLink221[12] , \ScanLink184[15] , \wBIn10[7] , 
        \wAIn11[12] , \wBMid15[27] , \wBMid60[17] , \wBMid23[22] , 
        \wBMid56[12] , \wBMid75[23] , \wAIn119[15] , \wRegInA115[30] , 
        \ScanLink202[23] , \wRegInA22[4] , \ScanLink217[17] , 
        \ScanLink241[16] , \wRegInB2[1] , \ScanLink234[26] , \ScanLink191[21] , 
        \ScanLink69[23] , \wBMid23[5] , \wAIn27[17] , \wAIn71[16] , 
        \wRegInB90[7] , \wAMid29[28] , \wAIn52[27] , \wRegInB68[27] , 
        \ScanLink62[0] , \wAIn32[23] , \wAIn47[13] , \wAMid115[4] , 
        \wAMid29[31] , \wAMid14[21] , \wBMid20[6] , \wAIn64[22] , \wAMid98[3] , 
        \wRegInA15[10] , \wRegInA36[21] , \wRegInA43[11] , \ScanLink61[3] , 
        \wRegInA60[20] , \wRegInB93[26] , \wRegInB93[4] , \wRegInA75[14] , 
        \wAMid35[0] , \wAMid49[6] , \wAMid54[9] , \wAMid84[28] , \wAMid84[31] , 
        \wRegInA56[25] , \ScanLink190[8] , \wAMid116[7] , \wRegInA23[15] , 
        \wRegInB86[12] , \wRegInB41[2] , \wRegInA103[8] , \ScanLink129[15] , 
        \ScanLink87[16] , \wRegInB118[18] , \ScanLink92[22] , \wAIn75[4] , 
        \wAIn112[19] , \wRegInB1[2] , \wRegInA21[7] , \ScanLink149[11] , 
        \wRegInA92[8] , \wBMid105[2] , \wAMid37[10] , \wAMid61[11] , 
        \ScanLink243[2] , \wBIn38[17] , \wAMid42[20] , \wAIn121[0] , 
        \wAMid22[24] , \wBMid9[8] , \wAMid57[14] , \wBIn58[13] , 
        \ScanLink123[7] , \wAMid74[25] , \wBMid93[9] , \wBIn118[13] , 
        \wRegInA85[19] , \wBIn95[17] , \wBMid112[16] , \wRegInB23[8] , 
        \ScanLink240[1] , \ScanLink5[11] , \wBIn80[23] , \wBMid107[22] , 
        \wAIn2[31] , \wAIn2[28] , \wAMid2[27] , \wAMid2[14] , \wAIn6[10] , 
        \wAIn9[1] , \wBMid8[20] , \wBMid8[13] , \wAMid10[23] , \wAIn11[0] , 
        \wBIn13[4] , \wAIn122[3] , \ScanLink120[4] , \wAMid14[12] , 
        \wAMid22[17] , \wAMid36[3] , \wBMid106[1] , \wBMid124[13] , 
        \wRegInB7[10] , \wRegInA28[19] , \ScanLink157[29] , \wRegInB106[20] , 
        \wRegInB125[11] , \ScanLink174[18] , \ScanLink122[19] , 
        \ScanLink101[31] , \ScanLink157[30] , \ScanLink101[28] , 
        \wRegInB113[14] , \wAMid57[27] , \wBIn58[20] , \wAIn76[7] , 
        \wRegInA1[15] , \ScanLink79[1] , \wRegInA106[5] , \wBMid38[4] , 
        \wAMid61[22] , \wAMid74[16] , \wBIn118[20] , \ScanLink227[6] , 
        \wRegInB35[19] , \wRegInB16[31] , \wAMid37[23] , \wAMid42[13] , 
        \wAIn59[18] , \wAMid83[2] , \wRegInB40[29] , \ScanLink147[3] , 
        \wBIn74[3] , \wRegInB16[28] , \wBIn38[24] , \wBMid48[19] , 
        \wRegInB40[30] , \wRegInB63[18] , \wRegInB59[0] , \wRegInB96[9] , 
        \ScanLink77[28] , \ScanLink21[30] , \wAMid51[4] , \ScanLink195[5] , 
        \ScanLink77[31] , \ScanLink54[19] , \wAIn12[3] , \wBMid90[29] , 
        \wRegInA1[26] , \wRegInA39[5] , \ScanLink21[29] , \wRegInB113[27] , 
        \wRegInB7[23] , \wRegInA118[9] , \ScanLink196[6] , \wRegInB125[22] , 
        \wAMid26[26] , \wBMid26[8] , \wBMid90[30] , \wAMid110[9] , 
        \wBIn29[21] , \wAIn36[5] , \wAMid52[7] , \wRegInB106[13] , 
        \wAMid76[1] , \wBIn77[0] , \wBIn80[10] , \wRegInB88[5] , 
        \ScanLink224[5] , \wBMid107[11] , \wBMid124[20] , \wRegInA105[6] , 
        \wAMid80[1] , \wAIn81[31] , \wRegInA27[9] , \wRegInB98[19] , 
        \ScanLink144[0] , \wAIn81[28] , \wBIn95[24] , \wBMid112[25] , 
        \ScanLink5[22] , \wRegInB117[16] , \wBIn81[0] , \wRegInA5[17] , 
        \wBIn50[5] , \wBIn53[6] , \wBIn84[21] , \wBMid94[18] , \wBMid103[20] , 
        \wRegInB3[12] , \wRegInB102[22] , \wRegInB121[13] , \ScanLink88[18] , 
        \ScanLink2[7] , \wBMid120[11] , \ScanLink160[6] , \wAIn85[19] , 
        \wRegInA121[0] , \wBIn91[15] , \ScanLink1[13] , \wBMid116[14] , 
        \ScanLink200[3] , \wAIn28[9] , \ScanLink163[5] , \wAMid53[16] , 
        \wAMid70[27] , \wAIn28[19] , \wAMid65[13] , \wRegInB44[18] , 
        \ScanLink203[0] , \wRegInB67[30] , \wBIn109[25] , \wRegInB31[28] , 
        \wRegInB60[9] , \wAMid33[12] , \wAMid46[22] , \wRegInB67[29] , 
        \wBIn49[25] , \wRegInB12[19] , \wRegInB31[31] , \wRegInA122[3] , 
        \wAMid9[18] , \wAMid11[6] , \wAMid12[5] , \wAIn35[6] , \wBIn82[3] , 
        \wBIn108[2] , \ScanLink218[19] , \wBIn37[2] , \wBMid39[18] , 
        \wAMid75[2] , \ScanLink73[19] , \ScanLink50[31] , \ScanLink50[28] , 
        \ScanLink40[8] , \ScanLink25[18] , \ScanLink1[4] , \wAIn52[1] , 
        \wAIn80[7] , \wAIn106[5] , \ScanLink104[2] , \wBIn84[12] , 
        \wBIn91[26] , \ScanLink1[20] , \wBMid103[13] , \wBMid116[27] , 
        \wRegInB109[9] , \wBMid120[22] , \wRegInA59[18] , \wRegInB3[21] , 
        \wRegInB121[20] , \ScanLink126[28] , \ScanLink153[18] , \wBMid122[7] , 
        \ScanLink170[30] , \wRegInB102[11] , \ScanLink126[31] , 
        \ScanLink105[19] , \wBMid65[9] , \wBMid121[4] , \wRegInA5[24] , 
        \wRegInB117[25] , \ScanLink170[29] , \wRegInB114[6] , \wAIn51[2] , 
        \wAIn118[9] , \wAIn116[28] , \wRegInA79[7] , \wAMid10[10] , 
        \wAMid65[20] , \wAIn116[31] , \wRegInB19[2] , \wRegInB117[5] , 
        \wBMid78[6] , \wBIn109[16] , \wAMid26[15] , \wBIn29[12] , 
        \wAMid33[21] , \wBIn34[1] , \wAMid46[11] , \ScanLink107[1] , 
        \wBIn49[16] , \wAIn105[6] , \wAMid53[25] , \wAIn83[4] , \wRegInA64[8] , 
        \wRegInA81[31] , \ScanLink39[3] , \wBMid32[27] , \wBIn48[7] , 
        \wAMid70[14] , \wRegInA81[28] , \wRegInA32[10] , \wRegInB97[17] , 
        \wBIn55[8] , \wAMid80[19] , \wRegInA11[21] , \wRegInA47[20] , 
        \wRegInA64[11] , \wRegInA71[25] , \ScanLink4[9] , \wRegInA27[24] , 
        \wRegInB82[23] , \ScanLink45[5] , \wRegInA52[14] , \ScanLink166[8] , 
        \wBIn110[0] , \ScanLink158[14] , \wRegInB65[4] , \ScanLink83[27] , 
        \ScanLink138[10] , \ScanLink96[13] , \ScanLink97[3] , \wRegInA111[18] , 
        \ScanLink78[26] , \wBMid47[17] , \ScanLink225[23] , \ScanLink180[24] , 
        \ScanLink250[13] , \wBMid11[16] , \wBMid64[26] , \wBIn99[2] , 
        \ScanLink206[12] , \wAIn6[23] , \wBIn14[31] , \wBIn14[28] , 
        \wAIn15[23] , \wAIn23[26] , \wBMid27[13] , \wBMid71[12] , 
        \wAIn108[10] , \wBIn113[3] , \ScanLink213[26] , \ScanLink94[0] , 
        \ScanLink230[17] , \ScanLink195[10] , \wBMid52[23] , \wRegInB66[7] , 
        \ScanLink245[27] , \ScanLink18[22] , \wAIn56[16] , \wAIn75[27] , 
        \wRegInB19[26] , \ScanLink178[4] , \wAIn33[8] , \wAIn36[12] , 
        \wAIn43[22] , \wAMid58[29] , \ScanLink46[6] , \wRegInB79[22] , 
        \wAMid58[30] , \wAIn60[13] , \ScanLink218[1] , \wAIn15[10] , 
        \wAIn36[21] , \wAIn49[0] , \wAIn86[9] , \wRegInA61[5] , 
        \ScanLink138[23] , \ScanLink96[20] , \wBMid60[4] , \ScanLink158[27] , 
        \ScanLink83[14] , \wAMid104[30] , \wAMid104[29] , \wBMid124[9] , 
        \wRegInA27[17] , \wRegInA52[27] , \wRegInA71[16] , \wRegInB82[10] , 
        \wRegInA47[13] , \ScanLink21[1] , \wRegInA32[23] , \wRegInA64[22] , 
        \wRegInB97[24] , \wRegInA11[12] , \wRegInB112[8] , \wRegInB79[11] , 
        \wAIn43[11] , \wAIn98[5] , \wAMid17[8] , \wBMid63[7] , \wAIn60[20] , 
        \wBIn42[30] , \wBIn61[18] , \wAIn75[14] , \wBIn102[29] , \wAIn23[15] , 
        \wBMid27[20] , \wBIn37[19] , \ScanLink22[2] , \wBIn42[29] , 
        \wBMid52[10] , \wAIn56[25] , \wBMid71[21] , \wBIn102[30] , 
        \wBIn121[18] , \wRegInB19[15] , \wAIn103[8] , \wRegInA62[6] , 
        \ScanLink213[15] , \ScanLink245[14] , \ScanLink18[11] , 
        \ScanLink230[24] , \ScanLink195[23] , \wBMid47[24] , \ScanLink250[20] , 
        \wBMid32[14] , \ScanLink225[10] , \ScanLink78[15] , \ScanLink180[17] , 
        \wBIn3[9] , \wBIn4[26] , \wAMid8[6] , \wAIn9[17] , \wBMid11[25] , 
        \wBMid64[15] , \wAIn108[23] , \wBMid25[2] , \wAIn39[15] , \wBIn58[29] , 
        \wAIn59[11] , \wRegInB4[6] , \wRegInB35[10] , \wRegInA90[17] , 
        \ScanLink206[21] , \wRegInB40[20] , \wBIn118[30] , \wRegInB16[21] , 
        \ScanLink188[3] , \wRegInA24[3] , \wRegInB63[11] , \ScanLink79[8] , 
        \wRegInB76[25] , \wBIn58[30] , \wBIn118[29] , \wRegInB20[24] , 
        \wRegInA85[23] , \wRegInB44[6] , \wRegInB55[14] , \ScanLink77[21] , 
        \wBMid48[10] , \wAIn124[26] , \wAIn11[9] , \wBIn69[5] , 
        \ScanLink54[10] , \wAMid113[3] , \ScanLink209[15] , \ScanLink21[20] , 
        \wBMid26[1] , \wBMid28[14] , \wAIn107[17] , \wAIn112[23] , 
        \ScanLink64[7] , \ScanLink41[24] , \ScanLink62[15] , \ScanLink34[14] , 
        \wBMid90[20] , \wRegInB59[9] , \wRegInB96[0] , \ScanLink17[25] , 
        \wAMid110[0] , \ScanLink159[6] , \ScanLink122[23] , \ScanLink157[13] , 
        \ScanLink239[3] , \ScanLink174[22] , \ScanLink101[12] , 
        \ScanLink114[26] , \wRegInB95[3] , \ScanLink161[16] , \ScanLink99[14] , 
        \wAIn9[24] , \wBMid28[27] , \wAMid35[9] , \wBMid41[6] , \wBIn77[9] , 
        \wBMid85[14] , \ScanLink137[17] , \wRegInA118[0] , \ScanLink142[27] , 
        \ScanLink67[4] , \wBIn80[19] , \wAMid80[8] , \wAIn81[21] , 
        \wRegInA27[0] , \wRegInB98[10] , \ScanLink144[9] , \wRegInA48[27] , 
        \wRegInB7[5] , \wBMid107[18] , \wAIn94[15] , \wBMid124[30] , 
        \wAIn112[10] , \wBMid124[29] , \wRegInA28[23] , \wRegInB47[5] , 
        \wRegInA92[1] , \ScanLink34[27] , \ScanLink41[17] , \ScanLink17[16] , 
        \ScanLink62[26] , \wBMid48[23] , \wAIn39[26] , \wAIn107[24] , 
        \wAIn124[15] , \ScanLink77[12] , \ScanLink21[13] , \wAIn121[9] , 
        \ScanLink209[26] , \ScanLink54[23] , \wRegInB76[16] , \wBIn4[15] , 
        \wBMid9[1] , \wAMid14[31] , \wAMid14[28] , \wAMid28[6] , \wAIn68[2] , 
        \wRegInA40[7] , \wBMid93[0] , \wBMid118[4] , \wRegInB55[27] , 
        \wRegInB20[17] , \wRegInA85[10] , \wAMid37[19] , \wAMid42[30] , 
        \wAMid61[18] , \wRegInB40[13] , \wRegInB20[2] , \wRegInB35[23] , 
        \wRegInA90[24] , \wAMid42[29] , \wAIn59[22] , \wRegInB63[22] , 
        \wAIn81[12] , \wBMid90[3] , \wRegInB16[12] , \wAIn94[26] , 
        \wRegInA28[10] , \wRegInA43[4] , \wRegInA48[14] , \wRegInB98[23] , 
        \ScanLink5[18] , \wRegInB23[1] , \ScanLink240[8] , \ScanLink161[25] , 
        \wBMid7[14] , \wBMid42[5] , \wBIn72[4] , \wBMid85[27] , \wBMid106[8] , 
        \wRegInA91[2] , \ScanLink142[14] , \ScanLink114[15] , \ScanLink99[27] , 
        \ScanLink137[24] , \wBMid90[13] , \ScanLink157[20] , \wRegInB7[19] , 
        \wRegInB106[30] , \wRegInB106[29] , \wRegInB125[18] , 
        \ScanLink122[10] , \ScanLink174[11] , \ScanLink141[4] , 
        \ScanLink101[21] , \wAMid85[5] , \wAMid108[2] , \wRegInB2[8] , 
        \wRegInA123[25] , \ScanLink191[31] , \ScanLink191[28] , 
        \wRegInA100[14] , \ScanLink221[1] , \wRegInB42[8] , \wRegInA115[20] , 
        \wBMid3[16] , \wBIn5[7] , \wBIn10[23] , \wAIn17[7] , \wBIn26[26] , 
        \wAMid29[21] , \wRegInA100[2] , \ScanLink193[2] , \wBIn53[16] , 
        \wAMid57[3] , \wBIn113[16] , \wBIn70[27] , \wBIn10[10] , \wAIn14[4] , 
        \wBIn33[12] , \wBIn65[13] , \wBIn106[22] , \ScanLink62[9] , 
        \wBIn46[22] , \wAMid49[25] , \wAMid54[0] , \wAMid84[21] , 
        \wBIn125[13] , \ScanLink190[1] , \wBMid47[8] , \wBIn71[7] , 
        \wAMid86[6] , \wAMid91[15] , \wAMid100[22] , \wAMid115[16] , 
        \wRegInA43[18] , \wRegInA60[30] , \wBMid119[13] , \wRegInA36[28] , 
        \wAMid123[13] , \wRegInA60[29] , \wRegInA15[19] , \wRegInA36[31] , 
        \wRegInB118[11] , \wBMid103[5] , \wRegInA103[1] , \ScanLink149[18] , 
        \ScanLink142[7] , \ScanLink222[2] , \wBIn65[20] , \wBMid88[1] , 
        \wBIn106[11] , \wAIn11[31] , \wBIn33[21] , \wAMid33[7] , \wBIn46[11] , 
        \wAMid49[16] , \wBIn125[20] , \wAIn47[29] , \wAIn73[3] , \wBIn53[25] , 
        \wAIn11[28] , \wBIn26[15] , \wAMid29[12] , \wAIn32[19] , \wAIn47[30] , 
        \wBIn113[25] , \wAIn64[18] , \wBIn70[14] , \wBIn16[0] , \wAIn127[7] , 
        \wRegInA115[13] , \ScanLink254[18] , \ScanLink221[28] , \wBIn6[4] , 
        \wBMid7[27] , \wRegInA46[9] , \ScanLink221[31] , \ScanLink202[19] , 
        \ScanLink125[0] , \wRegInA89[0] , \wRegInA123[16] , \wBMid23[18] , 
        \wBMid56[31] , \wBMid75[19] , \ScanLink245[5] , \wBMid56[28] , 
        \wRegInA100[27] , \ScanLink69[19] , \wBIn14[21] , \wAMid14[2] , 
        \wBIn15[3] , \wAIn124[4] , \ScanLink126[3] , \wAMid30[4] , 
        \wBMid59[4] , \wAIn70[0] , \wAMid100[11] , \wRegInB118[22] , 
        \ScanLink246[6] , \ScanLink92[18] , \ScanLink18[1] , \wAMid91[26] , 
        \wBMid100[6] , \wAMid123[20] , \wRegInA58[5] , \wBMid119[20] , 
        \wBIn31[5] , \wAMid84[12] , \wRegInB38[0] , \wRegInB86[31] , 
        \wAMid115[25] , \wRegInB86[28] , \wRegInB8[17] , \wRegInB109[27] , 
        \ScanLink96[29] , \wAIn49[9] , \wAIn86[0] , \wAIn100[2] , 
        \ScanLink102[5] , \ScanLink96[30] , \wAMid80[23] , \wAMid95[17] , 
        \wAMid104[20] , \ScanLink21[8] , \wBMid124[0] , \wRegInB112[1] , 
        \wBMid108[25] , \wAIn54[6] , \wRegInB82[19] , \wAMid111[14] , 
        \wAIn15[19] , \wBIn22[24] , \wAIn36[28] , \wBIn37[10] , \wBIn61[11] , 
        \wBIn102[20] , \wRegInB111[2] , \wAMid38[17] , \wBIn42[20] , 
        \wBIn121[11] , \wRegInB79[18] , \wAIn36[31] , \wAIn43[18] , 
        \wAIn57[5] , \wBIn57[14] , \wAMid58[13] , \wAIn60[30] , \wAMid17[1] , 
        \wAIn60[29] , \wBIn117[14] , \wBIn74[25] , \wBIn32[6] , 
        \wRegInA111[22] , \ScanLink250[29] , \ScanLink250[30] , 
        \ScanLink225[19] , \ScanLink206[31] , \ScanLink206[28] , 
        \ScanLink101[6] , \wBMid71[28] , \wAIn103[1] , \wBMid27[30] , 
        \wAIn85[3] , \wBMid27[29] , \wBMid52[19] , \wRegInA127[27] , 
        \wBMid71[31] , \ScanLink18[18] , \wRegInA104[16] , \wAMid80[10] , 
        \wRegInB78[2] , \ScanLink4[0] , \wBIn0[24] , \wBMid3[25] , 
        \wBMid19[6] , \wAIn30[2] , \wBIn87[7] , \wAMid104[13] , \wBMid108[16] , 
        \wAMid111[27] , \wRegInA11[31] , \wRegInA32[19] , \wBIn55[1] , 
        \wAMid70[6] , \wAMid95[24] , \wRegInA11[28] , \wRegInA18[7] , 
        \wRegInA47[29] , \wRegInA8[2] , \wRegInB8[24] , \wRegInA47[30] , 
        \wRegInA64[18] , \wRegInA127[7] , \ScanLink206[4] , \ScanLink138[19] , 
        \ScanLink58[3] , \ScanLink166[1] , \wBIn110[9] , \wRegInB109[14] , 
        \wRegInA124[4] , \wRegInA127[14] , \ScanLink94[9] , \wAIn6[19] , 
        \wAIn9[8] , \wRegInA104[25] , \ScanLink205[7] , \ScanLink195[19] , 
        \wRegInA111[11] , \wBIn14[12] , \wBIn22[17] , \wBIn56[2] , 
        \wBIn57[27] , \wAMid58[20] , \wAIn108[19] , \ScanLink165[2] , 
        \ScanLink89[6] , \wBIn61[22] , \wBIn74[16] , \wBIn117[27] , 
        \ScanLink218[8] , \ScanLink7[3] , \wAMid73[5] , \wBIn102[13] , 
        \wAIn33[1] , \wBIn37[23] , \wBIn42[13] , \wBIn84[4] , \wBIn121[22] , 
        \wAMid38[24] , \wAIn85[23] , \wAIn90[17] , \wRegInB109[0] , 
        \wRegInA39[15] , \wRegInA59[11] , \wRegInB89[26] , \wRegInA67[2] , 
        \ScanLink1[30] , \ScanLink165[14] , \ScanLink110[24] , \ScanLink1[29] , 
        \wBIn0[17] , \wBMid8[30] , \wBMid8[29] , \wAIn52[8] , \wBMid81[16] , 
        \ScanLink133[15] , \wBMid94[22] , \wRegInB3[28] , \ScanLink146[25] , 
        \ScanLink27[6] , \wRegInB121[29] , \ScanLink126[21] , \ScanLink119[4] , 
        \wBMid66[3] , \ScanLink153[11] , \wAIn116[21] , \wRegInB3[31] , 
        \wRegInB102[18] , \wRegInB121[30] , \ScanLink105[10] , 
        \ScanLink218[23] , \ScanLink170[20] , \ScanLink88[22] , 
        \ScanLink45[26] , \ScanLink24[5] , \ScanLink66[17] , \ScanLink30[16] , 
        \wAMid9[11] , \wBIn29[7] , \wBMid39[22] , \wBMid59[26] , 
        \ScanLink13[27] , \wBMid65[0] , \ScanLink73[23] , \wAIn120[24] , 
        \ScanLink50[12] , \wAIn118[0] , \wAMid10[19] , \wAIn48[27] , 
        \wAIn103[15] , \ScanLink25[22] , \wAMid65[29] , \wRegInB24[26] , 
        \wRegInB72[27] , \wRegInB51[16] , \wRegInA81[21] , \wRegInB31[12] , 
        \wRegInA94[15] , \wAIn28[23] , \wAMid33[31] , \wBIn34[8] , 
        \wAMid46[18] , \wRegInB44[22] , \wAMid65[30] , \ScanLink107[8] , 
        \wRegInB12[23] , \wAMid33[28] , \wBMid94[11] , \wRegInA64[1] , 
        \wRegInB67[13] , \ScanLink153[22] , \ScanLink43[2] , \ScanLink170[13] , 
        \ScanLink126[12] , \ScanLink88[11] , \ScanLink165[27] , 
        \ScanLink105[23] , \wAIn2[3] , \wAMid3[24] , \wAMid3[17] , 
        \wAMid9[22] , \wAIn28[10] , \wAMid76[8] , \ScanLink110[17] , 
        \wBIn81[9] , \wBMid81[25] , \ScanLink146[16] , \ScanLink133[26] , 
        \wBIn84[31] , \wBIn84[28] , \wAIn85[10] , \wRegInA39[26] , 
        \wRegInA121[9] , \ScanLink91[4] , \wAIn90[24] , \wRegInB63[3] , 
        \wBMid103[29] , \wBMid120[18] , \wRegInA59[22] , \wBMid103[30] , 
        \wBIn116[7] , \wRegInB89[15] , \wRegInB31[21] , \wRegInB44[11] , 
        \ScanLink203[9] , \wRegInA94[26] , \wRegInB60[0] , \ScanLink92[7] , 
        \wAIn28[0] , \wBIn29[28] , \wRegInB12[10] , \wRegInB67[20] , 
        \wRegInB72[14] , \wBIn115[4] , \wBIn29[31] , \wAIn48[14] , 
        \wRegInB51[25] , \wBMid39[11] , \wAMid68[4] , \wAIn120[17] , 
        \wRegInB24[15] , \wRegInA81[12] , \ScanLink73[10] , \ScanLink25[11] , 
        \wBMid10[15] , \wAIn14[20] , \wBMid59[15] , \wAIn103[26] , 
        \wAIn116[12] , \ScanLink50[21] , \ScanLink40[1] , \ScanLink218[10] , 
        \ScanLink30[25] , \ScanLink45[15] , \ScanLink13[14] , \wAIn61[10] , 
        \ScanLink208[2] , \ScanLink66[24] , \wBIn15[18] , \wBMid17[0] , 
        \wAIn22[25] , \wBIn36[29] , \wAIn37[11] , \wAIn42[21] , 
        \ScanLink56[5] , \wRegInB78[21] , \wBIn43[19] , \wAIn57[15] , 
        \wBIn60[31] , \wBIn120[28] , \wRegInB18[25] , \ScanLink168[7] , 
        \wBIn60[28] , \wAMid121[1] , \wBIn36[30] , \wAIn74[24] , \wBIn103[19] , 
        \wBIn120[31] , \wBMid26[10] , \ScanLink231[14] , \ScanLink194[13] , 
        \wBIn46[8] , \wBMid53[20] , \wRegInB76[4] , \ScanLink244[24] , 
        \ScanLink19[21] , \wBMid70[11] , \ScanLink212[25] , \ScanLink84[3] , 
        \wBMid65[25] , \wBIn89[1] , \ScanLink207[11] , \ScanLink175[8] , 
        \wRegInA16[1] , \wAIn7[13] , \wBMid33[24] , \wBIn103[0] , 
        \wAIn109[13] , \wBMid46[14] , \ScanLink224[20] , \ScanLink181[27] , 
        \ScanLink79[25] , \ScanLink251[10] , \wBMid14[3] , \wBIn100[3] , 
        \wRegInA5[7] , \wRegInA6[4] , \wRegInB75[7] , \ScanLink139[13] , 
        \ScanLink87[0] , \ScanLink48[9] , \ScanLink9[5] , \ScanLink97[10] , 
        \ScanLink82[24] , \wRegInA15[2] , \ScanLink159[17] , \wAMid126[28] , 
        \wRegInA26[27] , \ScanLink55[6] , \wRegInA53[17] , \wRegInB83[20] , 
        \wRegInB68[8] , \wRegInA70[26] , \wRegInA10[22] , \wAIn20[8] , 
        \wBIn58[4] , \wAMid105[19] , \wAMid126[31] , \wRegInA65[12] , 
        \wRegInA33[13] , \wRegInB96[14] , \wAMid122[2] , \wRegInA46[23] , 
        \wAIn7[20] , \wBMid10[26] , \wBMid65[16] , \wAIn109[20] , 
        \wRegInA110[31] , \wBMid46[27] , \ScanLink207[22] , \ScanLink251[23] , 
        \wAMid8[31] , \wAMid8[28] , \wAIn14[13] , \wAIn22[16] , \wBMid26[23] , 
        \wBMid33[17] , \wRegInA110[28] , \wBMid53[13] , \wRegInB12[0] , 
        \ScanLink244[17] , \ScanLink224[13] , \ScanLink181[14] , 
        \ScanLink79[16] , \ScanLink19[12] , \ScanLink231[27] , 
        \ScanLink194[20] , \wBMid70[22] , \wAIn95[9] , \ScanLink212[16] , 
        \wRegInA72[5] , \wAIn57[26] , \ScanLink32[1] , \wAIn74[17] , 
        \wRegInB18[16] , \wRegInB101[8] , \wAMid19[7] , \wAIn37[22] , 
        \wAIn61[23] , \wBMid73[4] , \wRegInB78[12] , \wAIn42[12] , \wAIn59[3] , 
        \wAMid59[19] , \wAIn88[6] , \wBMid70[7] , \wAMid81[30] , 
        \wRegInA10[11] , \wRegInA65[21] , \wRegInA33[20] , \wRegInA46[10] , 
        \wRegInB96[27] , \ScanLink31[2] , \wRegInA53[24] , \wRegInA26[14] , 
        \wRegInB83[13] , \wAMid81[29] , \wRegInA70[15] , \wAIn110[8] , 
        \wRegInB11[3] , \ScanLink82[17] , \ScanLink159[24] , \wRegInA71[6] , 
        \ScanLink139[20] , \ScanLink97[23] , \wBMid9[10] , \wAMid65[1] , 
        \wAIn117[18] , \wAMid11[20] , \wAIn25[5] , \wBIn92[0] , \wBIn118[1] , 
        \wAMid32[11] , \wAMid47[21] , \wBIn48[26] , \wAMid64[10] , 
        \ScanLink213[3] , \wBIn108[26] , \wAIn1[0] , \wAIn26[6] , 
        \wAMid27[25] , \wBIn28[22] , \wBIn40[6] , \wAMid71[24] , 
        \wRegInA80[18] , \wBIn43[5] , \wAMid52[15] , \ScanLink173[6] , 
        \wBIn90[16] , \ScanLink0[10] , \wBMid117[17] , \wBMid121[12] , 
        \wRegInA58[28] , \wRegInB73[9] , \ScanLink210[0] , \ScanLink170[5] , 
        \wBIn85[22] , \wBMid102[23] , \wRegInA58[31] , \wBIn91[3] , 
        \wRegInB2[11] , \wRegInA3[9] , \wRegInB103[21] , \ScanLink171[19] , 
        \ScanLink152[31] , \ScanLink152[28] , \ScanLink104[29] , 
        \ScanLink53[8] , \wRegInB120[10] , \ScanLink127[18] , 
        \ScanLink104[30] , \wAMid66[2] , \wRegInB116[15] , \wRegInA4[14] , 
        \wBIn0[30] , \wRegInA0[25] , \wRegInA0[16] , \wBMid9[23] , 
        \wAMid11[13] , \wBIn24[2] , \wAMid27[16] , \wBIn28[11] , \wAMid52[26] , 
        \wAMid71[17] , \ScanLink29[0] , \wAMid47[12] , \ScanLink117[2] , 
        \wBIn48[15] , \wAIn29[30] , \wAIn29[29] , \wAMid32[22] , \wAIn115[5] , 
        \wRegInB13[29] , \wAMid64[23] , \wAIn93[7] , \wRegInB66[19] , 
        \wRegInB45[31] , \wBMid68[5] , \wBIn108[15] , \wRegInB13[30] , 
        \wRegInB30[18] , \wRegInB45[28] , \wRegInB107[6] , \ScanLink219[30] , 
        \ScanLink219[29] , \wAMid26[0] , \wBIn27[1] , \wBMid38[31] , 
        \ScanLink72[30] , \wBMid38[28] , \wAIn41[1] , \ScanLink51[18] , 
        \ScanLink24[28] , \wRegInA69[4] , \ScanLink72[29] , \wAIn42[2] , 
        \wBMid76[9] , \wBMid95[31] , \wRegInA4[27] , \wRegInB116[26] , 
        \ScanLink24[31] , \wRegInB104[5] , \wBMid95[28] , \wRegInB103[12] , 
        \ScanLink89[28] , \wRegInB2[22] , \wRegInB120[23] , \ScanLink89[31] , 
        \wAIn84[29] , \wBIn85[11] , \wBMid102[10] , \wBMid121[21] , 
        \wBIn90[25] , \ScanLink0[23] , \wBMid117[24] , \wAIn66[4] , 
        \wAIn84[30] , \wAIn90[4] , \wAIn116[6] , \ScanLink114[1] , 
        \wRegInA77[8] , \wBMid116[2] , \wRegInA81[8] , \wRegInB112[17] , 
        \wBMid4[4] , \wRegInB120[3] , \wAMid5[3] , \wBMid7[7] , \wAMid15[22] , 
        \wAMid23[27] , \wAMid75[26] , \wAIn80[18] , \wBIn81[20] , \wBMid80[9] , 
        \wBMid91[19] , \wRegInB6[13] , \wRegInB107[23] , \wBMid125[10] , 
        \wRegInB124[12] , \ScanLink130[7] , \wBMid106[21] , \wBIn94[14] , 
        \wBMid113[15] , \wBIn119[10] , \wRegInB99[30] , \ScanLink250[2] , 
        \ScanLink4[12] , \wRegInB99[29] , \wAMid36[13] , \wAMid56[17] , 
        \wBIn59[10] , \wAIn78[8] , \ScanLink133[4] , \wBIn39[14] , 
        \wAMid43[23] , \wRegInB62[28] , \wAIn58[28] , \wRegInB17[18] , 
        \wRegInB34[30] , \wAMid25[3] , \wAIn58[31] , \wAMid60[12] , 
        \wRegInB41[19] , \ScanLink253[1] , \wRegInB62[31] , \wBMid115[1] , 
        \wRegInB30[8] , \wRegInB34[29] , \wBMid49[30] , \wAIn65[7] , 
        \wBMid49[29] , \ScanLink55[29] , \ScanLink20[19] , \ScanLink10[9] , 
        \ScanLink55[30] , \wBIn67[3] , \wAMid90[2] , \wBIn94[27] , 
        \wBMid113[26] , \wRegInB123[0] , \ScanLink76[18] , \ScanLink4[21] , 
        \wBMid125[23] , \wRegInA29[29] , \ScanLink154[3] , \wRegInA29[30] , 
        \wRegInA115[5] , \ScanLink234[6] , \wAMid42[4] , \wBIn81[13] , 
        \wRegInB98[6] , \wBMid106[12] , \wRegInB107[10] , \ScanLink100[18] , 
        \ScanLink123[30] , \wRegInB6[20] , \ScanLink175[28] , \wRegInB112[24] , 
        \wRegInB124[21] , \ScanLink186[5] , \ScanLink229[9] , 
        \ScanLink175[31] , \ScanLink156[19] , \ScanLink123[29] , \wBMid1[9] , 
        \wAIn3[11] , \wAMid6[0] , \wAMid15[11] , \wBMid28[7] , \wBMid35[8] , 
        \wAMid103[9] , \wRegInB85[9] , \ScanLink185[6] , \wRegInA29[6] , 
        \wAMid36[20] , \wAMid41[7] , \wRegInB9[3] , \wAMid43[10] , 
        \wAIn113[30] , \wAIn113[29] , \wRegInB49[3] , \ScanLink157[0] , 
        \wBIn64[0] , \ScanLink198[9] , \wBIn39[27] , \wAMid60[21] , 
        \wBIn121[8] , \wRegInA34[9] , \wAMid93[1] , \wBIn119[23] , 
        \wRegInA84[29] , \wAMid7[15] , \wBMid14[17] , \wBIn18[6] , 
        \wAMid23[14] , \wAMid56[24] , \wBIn59[23] , \wAMid75[15] , 
        \ScanLink237[5] , \wRegInA84[30] , \ScanLink69[2] , \wRegInA116[6] , 
        \wBMid54[1] , \wRegInA14[20] , \wRegInA37[11] , \wRegInA61[10] , 
        \wRegInB92[16] , \wAMid85[18] , \wRegInA22[25] , \wRegInA42[21] , 
        \wRegInA87[6] , \ScanLink15[4] , \wRegInA57[15] , \wRegInB87[22] , 
        \wRegInA74[24] , \wBMid86[7] , \wRegInB35[5] , \wRegInA55[0] , 
        \ScanLink136[9] , \ScanLink86[26] , \ScanLink128[25] , 
        \wRegInB119[31] , \wRegInB119[28] , \ScanLink148[21] , 
        \ScanLink93[12] , \wBMid61[27] , \wRegInA56[3] , \ScanLink203[13] , 
        \wBMid37[26] , \wBMid42[16] , \wBMid85[4] , \wRegInA114[19] , 
        \ScanLink220[22] , \ScanLink185[25] , \wBIn8[2] , \wBMid22[12] , 
        \ScanLink255[12] , \ScanLink235[16] , \ScanLink190[11] , 
        \ScanLink68[13] , \wAIn53[17] , \wBMid57[22] , \ScanLink240[26] , 
        \wBMid74[13] , \wAIn118[25] , \wRegInB36[6] , \ScanLink216[27] , 
        \wAIn26[27] , \ScanLink128[5] , \wBMid57[2] , \wAIn63[9] , 
        \wAIn70[26] , \wRegInB69[17] , \wRegInA84[5] , \wAIn65[12] , 
        \ScanLink248[0] , \wAMid2[23] , \wAMid2[10] , \wAIn3[22] , 
        \wAMid7[26] , \wAIn10[22] , \wAIn10[11] , \wAIn19[1] , \wAMid28[18] , 
        \wAIn33[13] , \wAIn46[23] , \ScanLink16[7] , \wBIn124[5] , 
        \ScanLink148[12] , \wRegInA31[4] , \wBMid30[5] , \wAMid59[5] , 
        \ScanLink93[21] , \wAMid106[4] , \wRegInA22[16] , \wRegInB51[1] , 
        \ScanLink232[8] , \ScanLink86[15] , \wRegInA57[26] , \ScanLink128[16] , 
        \wRegInB87[11] , \wRegInA74[17] , \wBMid33[6] , \wAMid101[31] , 
        \wBMid118[19] , \wRegInA61[23] , \wAMid101[28] , \wAMid122[19] , 
        \wRegInB83[7] , \wRegInA14[13] , \wRegInA42[12] , \ScanLink71[0] , 
        \wRegInA37[22] , \wRegInB92[25] , \wBIn11[30] , \wAIn26[14] , 
        \wAIn33[20] , \wAMid47[9] , \wAMid88[0] , \wAIn65[21] , \wAIn46[10] , 
        \wAMid105[7] , \ScanLink183[8] , \wBIn11[29] , \wBIn32[18] , 
        \wBIn47[28] , \wRegInB69[24] , \ScanLink72[3] , \wAIn53[24] , 
        \wBIn107[31] , \wBIn124[19] , \wBMid22[21] , \wBIn47[31] , 
        \wAIn70[15] , \wBMid57[11] , \wBIn64[19] , \wBIn107[28] , 
        \wRegInB80[4] , \ScanLink240[15] , \ScanLink235[25] , 
        \ScanLink190[22] , \ScanLink68[20] , \wBMid74[20] , \wAIn118[16] , 
        \wAMid118[8] , \ScanLink216[14] , \wBIn127[6] , \wRegInA32[7] , 
        \wBMid14[24] , \wBMid61[14] , \wBMid42[25] , \wRegInA110[8] , 
        \ScanLink203[20] , \wBMid3[31] , \wAIn15[27] , \wBMid37[15] , 
        \wRegInB52[2] , \ScanLink255[21] , \wAIn60[17] , \ScanLink220[11] , 
        \ScanLink185[16] , \ScanLink218[5] , \wAIn23[22] , \wAIn36[16] , 
        \wAIn43[26] , \ScanLink46[2] , \wRegInB79[26] , \wAMid38[29] , 
        \wAIn56[12] , \wBIn84[9] , \wRegInB19[22] , \ScanLink178[0] , 
        \wBMid27[17] , \wAMid38[30] , \wAIn75[23] , \wAMid73[8] , 
        \wRegInA104[28] , \ScanLink230[13] , \ScanLink195[14] , \wBMid52[27] , 
        \ScanLink245[23] , \wRegInB66[3] , \ScanLink18[26] , \wBMid3[28] , 
        \wBMid71[16] , \wRegInA104[31] , \ScanLink213[22] , \ScanLink94[4] , 
        \wRegInA124[9] , \wRegInA127[19] , \wBMid11[12] , \wBMid64[22] , 
        \wBIn99[6] , \ScanLink206[16] , \wBIn113[7] , \wAIn6[14] , \wAIn9[5] , 
        \wBMid32[23] , \wAIn108[14] , \ScanLink78[22] , \wBMid47[13] , 
        \ScanLink225[27] , \ScanLink180[20] , \wBIn48[3] , \wAMid95[29] , 
        \wBIn110[4] , \wRegInB8[30] , \wRegInB65[0] , \ScanLink250[17] , 
        \ScanLink206[9] , \ScanLink138[14] , \ScanLink97[7] , \ScanLink96[17] , 
        \wRegInB8[29] , \wRegInB109[19] , \ScanLink83[23] , \ScanLink158[10] , 
        \wRegInA11[25] , \wRegInA27[20] , \wRegInB82[27] , \ScanLink45[1] , 
        \wRegInA52[10] , \wRegInA71[21] , \wRegInA32[14] , \wRegInA64[15] , 
        \wRegInB97[13] , \wAMid95[30] , \wRegInA47[24] , \wAIn6[27] , 
        \wBMid11[21] , \wBMid64[11] , \wAIn108[27] , \wBMid47[20] , 
        \ScanLink206[25] , \wBMid8[24] , \wBMid8[17] , \wAIn15[14] , 
        \wBIn22[30] , \wAIn23[11] , \wBMid27[24] , \wBMid32[10] , 
        \ScanLink250[24] , \ScanLink78[11] , \wBMid52[14] , \ScanLink245[10] , 
        \ScanLink225[14] , \ScanLink180[13] , \ScanLink230[20] , 
        \ScanLink195[27] , \ScanLink18[15] , \wBMid71[25] , \wRegInA62[2] , 
        \ScanLink213[11] , \wAIn56[21] , \ScanLink22[6] , \wBMid63[3] , 
        \wAIn75[10] , \wRegInB19[11] , \wBIn22[29] , \wAIn60[24] , 
        \wBIn74[28] , \wBIn117[19] , \wRegInB79[15] , \wBIn31[8] , 
        \wAIn36[25] , \wAIn43[15] , \wAIn57[8] , \wBIn74[31] , \wBIn57[19] , 
        \wAIn98[1] , \wBMid60[0] , \wBMid108[31] , \wRegInA11[16] , 
        \wRegInA64[26] , \wRegInA32[27] , \wRegInA47[17] , \ScanLink21[5] , 
        \wRegInA52[23] , \wRegInB97[20] , \wAMid111[19] , \wRegInA27[13] , 
        \wRegInB82[14] , \wRegInA71[12] , \wBMid108[28] , \ScanLink158[23] , 
        \ScanLink83[10] , \wAIn49[4] , \wRegInA61[1] , \ScanLink102[8] , 
        \ScanLink138[27] , \wBMid59[18] , \ScanLink96[24] , \ScanLink30[31] , 
        \ScanLink1[0] , \ScanLink13[19] , \wAMid75[6] , \ScanLink66[29] , 
        \wAMid10[27] , \wAMid33[16] , \wAIn35[2] , \wBIn82[7] , 
        \ScanLink30[28] , \wBIn108[6] , \ScanLink66[30] , \ScanLink45[18] , 
        \wAMid46[26] , \wBIn49[21] , \wRegInA122[7] , \wAMid10[14] , 
        \wAMid26[22] , \wBIn50[1] , \wAMid65[17] , \ScanLink203[4] , 
        \wAMid68[9] , \wBIn109[21] , \wRegInB24[18] , \wRegInB51[28] , 
        \wAMid70[23] , \wRegInB72[19] , \wRegInB51[31] , \wAMid26[11] , 
        \wBIn29[25] , \wAIn36[1] , \wAIn48[19] , \wBIn115[9] , 
        \ScanLink163[1] , \wBIn53[2] , \wAMid53[12] , \wBIn91[11] , 
        \wBMid116[10] , \wRegInA121[4] , \ScanLink200[7] , \ScanLink1[17] , 
        \ScanLink91[9] , \ScanLink160[2] , \wBIn81[4] , \wBIn84[25] , 
        \wAIn90[30] , \wBMid103[24] , \wBMid120[15] , \wRegInB89[18] , 
        \wAIn90[29] , \wRegInB3[16] , \wRegInB102[26] , \ScanLink2[3] , 
        \wRegInB121[17] , \wAMid53[21] , \wAMid70[10] , \wAMid76[5] , 
        \wBMid81[28] , \wRegInB117[12] , \wBMid81[31] , \wRegInA5[13] , 
        \ScanLink39[7] , \wBIn29[16] , \wAMid33[25] , \wBIn34[5] , 
        \wAMid46[15] , \wBIn49[12] , \ScanLink107[5] , \wAIn105[2] , 
        \wAMid65[24] , \wAIn83[0] , \wBMid78[2] , \wBIn109[12] , 
        \wRegInA94[18] , \wRegInB19[6] , \wRegInB117[1] , \ScanLink24[8] , 
        \wAMid11[2] , \wAIn51[6] , \wAIn103[18] , \wAIn120[30] , 
        \wRegInA79[3] , \wBMid121[0] , \wAIn120[29] , \ScanLink146[28] , 
        \ScanLink133[18] , \ScanLink110[30] , \wBIn0[29] , \wRegInA5[20] , 
        \wRegInB117[21] , \ScanLink110[29] , \ScanLink165[19] , 
        \ScanLink146[31] , \wBIn0[7] , \wBIn4[18] , \wAMid12[1] , 
        \wBMid122[3] , \wRegInB114[2] , \wRegInB102[15] , \wBIn37[6] , 
        \wAIn52[5] , \wRegInB3[25] , \wRegInB121[24] , \ScanLink119[9] , 
        \wBIn84[16] , \wBMid103[17] , \wBMid120[26] , \wBIn91[22] , 
        \wBMid116[23] , \ScanLink1[24] , \wBMid42[8] , \wAIn76[3] , 
        \wAIn80[3] , \wAIn106[1] , \wRegInA39[18] , \ScanLink104[6] , 
        \ScanLink161[31] , \ScanLink142[19] , \wBMid106[5] , \ScanLink161[28] , 
        \ScanLink137[29] , \wAMid36[7] , \wRegInB113[10] , \ScanLink137[30] , 
        \ScanLink114[18] , \wRegInA1[11] , \wRegInB7[14] , \wRegInB106[24] , 
        \wRegInB125[15] , \wRegInA0[31] , \wRegInA0[28] , \wAIn2[25] , 
        \wAIn2[16] , \wBIn3[4] , \wBIn10[3] , \wBIn13[0] , \wAIn122[7] , 
        \ScanLink120[0] , \wBMid124[17] , \wAMid74[21] , \wBIn80[27] , 
        \wRegInA43[9] , \wBIn95[13] , \wBMid107[26] , \wBMid112[12] , 
        \ScanLink5[15] , \wBIn118[17] , \wBMid118[9] , \wRegInA48[19] , 
        \ScanLink240[5] , \wAIn121[4] , \wBIn6[9] , \wAIn9[30] , \wAMid14[25] , 
        \wAMid22[20] , \wAMid37[14] , \wBIn38[13] , \wAMid57[10] , 
        \ScanLink123[3] , \wBIn58[17] , \wAMid42[24] , \wRegInA90[30] , 
        \wAMid35[4] , \wAMid61[15] , \ScanLink243[6] , \wBMid105[6] , 
        \wRegInA90[29] , \wAIn75[0] , \wAIn9[29] , \wAIn107[29] , 
        \wAIn124[18] , \wAIn11[4] , \wAIn12[7] , \wAMid52[3] , \wBIn77[4] , 
        \wAMid80[5] , \wBIn95[20] , \wAIn107[30] , \wBMid112[21] , 
        \ScanLink5[26] , \wRegInB7[8] , \wBIn80[14] , \wAIn94[18] , 
        \wBMid124[24] , \ScanLink144[4] , \wRegInB47[8] , \wRegInB88[1] , 
        \wRegInA105[2] , \ScanLink224[1] , \wBMid107[15] , \wRegInB106[17] , 
        \wRegInB7[27] , \wRegInB125[26] , \ScanLink196[2] , \wBIn69[8] , 
        \wBMid85[19] , \ScanLink67[9] , \wRegInA1[22] , \wRegInB113[23] , 
        \ScanLink209[18] , \ScanLink195[1] , \ScanLink99[19] , \wAMid14[16] , 
        \wBMid28[19] , \wAMid51[0] , \wRegInA39[1] , \ScanLink62[18] , 
        \ScanLink41[30] , \wAMid37[27] , \wBIn38[20] , \wAMid42[17] , 
        \wRegInB59[4] , \ScanLink147[7] , \ScanLink41[29] , \ScanLink17[28] , 
        \ScanLink34[19] , \ScanLink17[31] , \wBIn74[7] , \wBMid38[0] , 
        \wAMid61[26] , \wAMid83[6] , \wAMid22[13] , \wAIn39[18] , 
        \wAMid57[23] , \wAMid74[12] , \wBIn118[24] , \wRegInB20[29] , 
        \ScanLink227[2] , \wRegInB20[30] , \wRegInB55[19] , \wRegInB76[31] , 
        \ScanLink79[5] , \wBIn58[24] , \wRegInB76[28] , \wRegInA106[1] , 
        \wAMid30[9] , \wBMid44[6] , \wRegInA15[27] , \wRegInA60[17] , 
        \wBMid59[9] , \wBMid96[0] , \wAMid115[31] , \wAMid115[28] , 
        \wRegInA23[22] , \wRegInA36[16] , \wRegInA43[26] , \wRegInA58[8] , 
        \wRegInB93[11] , \wRegInA97[1] , \wRegInB86[25] , \wRegInA56[12] , 
        \wRegInA75[23] , \ScanLink87[21] , \wAMid6[12] , \wBMid15[10] , 
        \wAIn124[9] , \ScanLink129[22] , \wRegInB25[2] , \wRegInA45[7] , 
        \ScanLink149[26] , \ScanLink92[15] , \wBMid60[20] , \ScanLink202[14] , 
        \wRegInA46[4] , \wBMid36[21] , \wBMid43[11] , \wBMid95[3] , 
        \ScanLink221[25] , \ScanLink184[22] , \ScanLink254[15] , \wAMid6[21] , 
        \wBMid7[19] , \wAIn11[25] , \wBMid23[15] , \ScanLink245[8] , 
        \ScanLink234[11] , \ScanLink191[16] , \wAIn27[20] , \wAIn52[10] , 
        \wBMid56[25] , \wRegInB26[1] , \ScanLink241[21] , \ScanLink69[14] , 
        \wBMid75[14] , \wAIn119[22] , \ScanLink217[20] , \ScanLink138[2] , 
        \wBMid47[5] , \wRegInB68[10] , \wRegInA94[2] , \wBIn53[31] , 
        \wAIn71[21] , \wBMid103[8] , \wBIn113[28] , \wAIn64[15] , \wBIn70[19] , 
        \wAIn11[16] , \wAIn14[9] , \wBIn26[18] , \wAIn32[14] , \wAIn47[24] , 
        \wBIn53[28] , \wBIn113[31] , \wAMid49[2] , \wRegInA21[3] , 
        \ScanLink149[15] , \ScanLink92[26] , \wAMid116[3] , \wRegInB1[6] , 
        \wRegInA23[11] , \wRegInB41[6] , \ScanLink87[12] , \wRegInA56[21] , 
        \ScanLink129[11] , \wRegInB86[16] , \wBMid20[2] , \wAMid91[18] , 
        \wRegInA75[10] , \wRegInA15[14] , \wRegInA60[24] , \wRegInB93[0] , 
        \wRegInA36[25] , \wRegInA43[15] , \ScanLink61[7] , \wRegInB93[22] , 
        \wBMid23[26] , \wBMid23[1] , \wAIn27[13] , \wAIn32[27] , \wAIn64[26] , 
        \wAMid98[7] , \wAIn47[17] , \wAMid115[0] , \wAMid49[31] , 
        \wAMid49[28] , \wRegInB68[23] , \ScanLink62[4] , \wAIn52[23] , 
        \wBMid56[16] , \wAIn71[12] , \wRegInB90[3] , \ScanLink241[12] , 
        \wAMid85[8] , \wRegInB2[5] , \ScanLink234[22] , \ScanLink191[25] , 
        \wAIn119[11] , \wRegInA100[19] , \wRegInA123[31] , \ScanLink69[27] , 
        \ScanLink141[9] , \wBIn72[9] , \wBMid75[27] , \wRegInA22[0] , 
        \wRegInA123[28] , \ScanLink217[13] , \wBMid15[23] , \wBMid60[13] , 
        \wBMid43[22] , \ScanLink202[27] , \ScanLink254[26] , \wAIn8[10] , 
        \wAMid23[19] , \wBMid36[12] , \wAMid56[29] , \wAIn58[16] , 
        \wRegInB34[17] , \wRegInB42[5] , \ScanLink221[16] , \ScanLink184[11] , 
        \wRegInB41[27] , \wRegInA91[10] , \wBIn121[5] , \wRegInB17[26] , 
        \ScanLink198[4] , \wRegInA34[4] , \wRegInB62[16] , \wRegInB77[22] , 
        \wBMid35[5] , \wAIn38[12] , \wAMid56[30] , \wAMid75[18] , 
        \wRegInB21[23] , \wRegInA84[24] , \wRegInB54[13] , \ScanLink237[8] , 
        \wRegInB54[1] , \ScanLink76[26] , \wBMid49[17] , \wAIn125[21] , 
        \wBMid29[13] , \wBIn79[2] , \ScanLink55[17] , \wAMid103[4] , 
        \ScanLink208[12] , \wAIn106[10] , \ScanLink20[27] , \wAIn113[24] , 
        \ScanLink74[0] , \ScanLink40[23] , \ScanLink35[13] , \wBMid36[6] , 
        \wBMid91[27] , \wRegInB86[7] , \ScanLink63[12] , \ScanLink16[22] , 
        \ScanLink186[8] , \wAMid100[7] , \ScanLink149[1] , \ScanLink123[24] , 
        \ScanLink156[14] , \wAMid42[9] , \ScanLink100[15] , \wRegInB112[29] , 
        \ScanLink229[4] , \ScanLink175[25] , \ScanLink115[21] , \wBIn5[21] , 
        \wRegInB85[4] , \ScanLink160[11] , \ScanLink98[13] , \wBMid84[13] , 
        \wRegInB112[30] , \ScanLink136[10] , \wBIn5[12] , \wAIn8[23] , 
        \wBMid29[20] , \wBMid51[1] , \wAIn80[26] , \wBIn122[6] , 
        \wRegInB99[17] , \wRegInA108[7] , \ScanLink143[20] , \ScanLink77[3] , 
        \wRegInA37[7] , \wRegInA49[20] , \wAIn95[12] , \wAIn113[17] , 
        \wRegInA29[24] , \wRegInB57[2] , \wRegInA115[8] , \wRegInA82[6] , 
        \ScanLink35[20] , \ScanLink40[10] , \ScanLink16[11] , \wBMid49[24] , 
        \ScanLink63[21] , \wAIn38[21] , \wAIn106[23] , \wAIn125[12] , 
        \ScanLink76[15] , \ScanLink20[14] , \wRegInB77[11] , \ScanLink208[21] , 
        \ScanLink55[24] , \ScanLink10[4] , \ScanLink133[9] , \wAMid38[1] , 
        \wAIn78[5] , \wRegInA50[0] , \wBMid83[7] , \wBMid108[3] , 
        \wRegInB54[20] , \wBIn39[19] , \wRegInB21[10] , \wRegInA84[17] , 
        \wRegInB30[5] , \wRegInB34[24] , \wRegInB41[14] , \wRegInA91[23] , 
        \wAIn58[25] , \wRegInB62[25] , \wAIn80[15] , \wBMid80[4] , 
        \wRegInB17[15] , \wBIn94[19] , \wAIn95[21] , \wRegInA29[17] , 
        \wRegInA49[13] , \wRegInA53[3] , \wRegInB99[24] , \wBMid113[18] , 
        \wRegInB33[6] , \ScanLink160[22] , \wBMid52[2] , \ScanLink98[20] , 
        \wAIn66[9] , \wRegInA81[5] , \ScanLink143[13] , \ScanLink115[12] , 
        \ScanLink136[23] , \wBMid84[20] , \ScanLink13[7] , \wAMid0[3] , 
        \wBMid4[9] , \wBMid91[14] , \ScanLink156[27] , \ScanLink175[16] , 
        \ScanLink123[17] , \ScanLink100[26] , \wBMid6[13] , \wBIn62[3] , 
        \ScanLink151[3] , \wBMid42[28] , \wAMid95[2] , \wAMid118[5] , 
        \ScanLink235[31] , \wRegInA122[22] , \ScanLink216[19] , 
        \ScanLink240[18] , \ScanLink235[28] , \wRegInA101[13] , \wBIn1[23] , 
        \wBMid1[4] , \wAMid3[0] , \wBIn11[24] , \wBMid14[30] , \wBMid37[18] , 
        \ScanLink231[6] , \wRegInA114[27] , \wBMid14[29] , \wBMid42[31] , 
        \wBMid61[19] , \wBIn27[21] , \wRegInA110[5] , \ScanLink183[5] , 
        \wAMid28[26] , \wAMid47[4] , \wBIn52[11] , \wBIn71[20] , \wBIn112[11] , 
        \wAIn26[19] , \wBIn32[15] , \wAIn53[30] , \wBIn64[14] , 
        \wRegInB69[30] , \wAIn70[18] , \wBIn107[25] , \wRegInB80[9] , 
        \wBMid30[8] , \wBIn47[25] , \wAMid48[22] , \wAIn53[29] , 
        \wRegInB69[29] , \wBIn124[14] , \wAMid44[7] , \wAMid85[26] , 
        \wAMid59[8] , \wAMid90[12] , \wAMid101[25] , \wAMid106[9] , 
        \wAMid114[11] , \ScanLink180[6] , \wRegInB92[28] , \wBMid118[14] , 
        \wAMid122[14] , \wRegInB92[31] , \wBIn61[0] , \wAMid96[1] , 
        \wRegInB119[16] , \wBIn124[8] , \wRegInA31[9] , \ScanLink152[0] , 
        \wRegInA113[6] , \ScanLink232[5] , \ScanLink86[18] , \wBIn11[17] , 
        \wAMid23[0] , \wBIn64[27] , \wBMid113[2] , \wBMid98[6] , \wBIn107[16] , 
        \wBIn27[12] , \wBIn32[26] , \wBIn47[16] , \wAMid48[11] , \wBIn124[27] , 
        \ScanLink128[8] , \wBIn52[22] , \wAIn63[4] , \wRegInA84[8] , 
        \wAMid28[15] , \wBIn71[13] , \wBIn112[22] , \wBMid2[22] , \wBMid2[11] , 
        \wBMid2[7] , \wBMid6[20] , \wAMid7[18] , \wBMid85[9] , 
        \wRegInA114[14] , \wRegInB125[3] , \ScanLink185[31] , 
        \ScanLink185[28] , \ScanLink135[7] , \wAIn118[28] , \wRegInA99[7] , 
        \wRegInA122[11] , \wAMid20[3] , \wBMid49[3] , \wAIn118[31] , 
        \wRegInA101[20] , \ScanLink255[2] , \ScanLink136[4] , 
        \ScanLink128[31] , \ScanLink128[28] , \wAIn60[7] , \wAMid101[16] , 
        \wRegInB35[8] , \wRegInB119[25] , \ScanLink256[1] , \wAMid90[21] , 
        \wBMid110[1] , \wAMid122[27] , \wRegInA48[2] , \wBMid118[27] , 
        \wRegInA22[31] , \wRegInB28[7] , \wRegInA74[29] , \wRegInB126[0] , 
        \wAMid3[30] , \wBIn15[26] , \wBIn21[2] , \wAMid85[15] , \wAMid114[22] , 
        \wRegInA22[28] , \ScanLink15[9] , \wRegInB9[10] , \wRegInA57[18] , 
        \wRegInA74[30] , \ScanLink159[29] , \wRegInB108[20] , 
        \ScanLink159[30] , \wAIn44[1] , \wAMid81[24] , \wAMid94[10] , 
        \wAIn96[7] , \wAIn110[5] , \ScanLink112[2] , \wAMid105[27] , 
        \wBMid109[22] , \wAMid126[16] , \wRegInA53[30] , \wRegInB102[6] , 
        \wRegInA70[18] , \wRegInA26[19] , \wRegInA53[29] , \wAMid110[13] , 
        \wBIn23[23] , \wBIn36[17] , \wAMid39[10] , \wBIn60[16] , \wBIn103[27] , 
        \wRegInB101[5] , \wBIn43[27] , \wBIn120[16] , \wAIn47[2] , 
        \wBIn56[13] , \wAMid59[14] , \wBMid73[9] , \wBIn75[22] , \wBIn116[13] , 
        \wAMid3[29] , \wRegInA110[25] , \ScanLink181[19] , \wBIn22[1] , 
        \ScanLink111[1] , \wAIn7[3] , \wAIn20[5] , \wBIn58[9] , \wAMid81[17] , 
        \wAIn95[4] , \wAIn113[6] , \wRegInA72[8] , \wBMid109[11] , 
        \wRegInB68[5] , \wRegInA105[11] , \wRegInA126[20] , \wBIn97[0] , 
        \wAMid105[14] , \wAMid110[20] , \wRegInB96[19] , \wBIn45[6] , 
        \wAMid60[1] , \wAMid94[23] , \wAMid126[25] , \wRegInB9[23] , 
        \ScanLink216[3] , \ScanLink176[6] , \ScanLink48[4] , \ScanLink9[8] , 
        \wRegInB108[13] , \ScanLink82[30] , \wRegInA126[13] , 
        \ScanLink212[28] , \ScanLink82[29] , \ScanLink244[30] , \wAIn4[0] , 
        \wBMid10[18] , \wBMid33[29] , \wRegInB76[9] , \wRegInA105[22] , 
        \ScanLink231[19] , \ScanLink215[0] , \ScanLink212[31] , 
        \ScanLink244[29] , \wRegInA110[16] , \wBMid46[19] , \ScanLink79[28] , 
        \wBMid65[31] , \wRegInA6[9] , \wBIn23[10] , \wBMid33[30] , \wBIn46[5] , 
        \wBIn56[20] , \wBMid65[28] , \ScanLink175[5] , \ScanLink79[31] , 
        \ScanLink99[1] , \wAMid59[27] , \ScanLink56[8] , \wBIn60[25] , 
        \wAIn74[29] , \wBIn75[11] , \wBIn116[20] , \wRegInB18[31] , 
        \wBIn15[15] , \wBIn103[14] , \wAIn22[31] , \wAMid63[2] , \wAIn22[28] , 
        \wBIn43[14] , \wAIn57[18] , \wAIn74[30] , \wBIn94[3] , \wBIn120[25] , 
        \wRegInB18[28] , \wAIn23[6] , \wBIn36[24] , \wAMid39[23] , 
        \wAIn84[24] , \wAIn90[9] , \wAIn91[10] , \wRegInB17[0] , 
        \wRegInB119[7] , \wRegInA38[12] , \wRegInA58[16] , \wRegInB88[21] , 
        \wRegInA77[5] , \wBIn90[31] , \wBMid117[30] , \wBIn90[28] , 
        \wBMid117[29] , \wRegInB104[8] , \ScanLink164[13] , \ScanLink111[23] , 
        \wBIn1[10] , \wAMid8[16] , \wBIn39[0] , \wBMid38[25] , \wBMid58[21] , 
        \wBMid76[4] , \wBMid80[11] , \ScanLink132[12] , \wBMid95[25] , 
        \ScanLink147[22] , \ScanLink37[1] , \ScanLink152[16] , 
        \ScanLink127[26] , \ScanLink109[3] , \wAIn117[26] , \ScanLink219[24] , 
        \ScanLink171[27] , \ScanLink104[17] , \ScanLink89[25] , 
        \ScanLink44[21] , \ScanLink34[2] , \ScanLink67[10] , \ScanLink31[11] , 
        \ScanLink72[24] , \ScanLink12[20] , \wBMid75[7] , \wAIn121[23] , 
        \ScanLink51[15] , \wAIn108[7] , \wAIn29[24] , \wBIn48[18] , 
        \wAIn49[20] , \wAIn102[12] , \wRegInA69[9] , \ScanLink24[25] , 
        \wBMid68[8] , \wRegInB14[3] , \wRegInB25[21] , \wRegInB73[20] , 
        \wRegInA80[26] , \wRegInB50[11] , \wBIn108[18] , \wRegInB30[15] , 
        \wRegInB45[25] , \wRegInA95[12] , \wAIn115[8] , \wRegInB13[24] , 
        \wBMid95[16] , \wRegInB66[14] , \wRegInA74[6] , \ScanLink152[25] , 
        \ScanLink53[5] , \ScanLink171[14] , \ScanLink127[15] , 
        \ScanLink89[16] , \ScanLink164[20] , \ScanLink104[24] , \wBMid12[0] , 
        \wAMid27[28] , \wAIn29[17] , \wBIn43[8] , \wBMid80[22] , \wAMid124[1] , 
        \wRegInA4[19] , \wRegInB116[18] , \ScanLink111[10] , \ScanLink147[11] , 
        \ScanLink132[21] , \wAIn84[17] , \wRegInA38[21] , \ScanLink81[3] , 
        \wAIn91[23] , \wRegInB73[4] , \wRegInA3[4] , \wRegInA58[25] , 
        \ScanLink170[8] , \wBIn106[0] , \wRegInA13[1] , \wRegInB88[12] , 
        \wRegInB30[26] , \wRegInB45[16] , \wRegInB70[7] , \wRegInA95[21] , 
        \ScanLink82[0] , \wRegInB13[17] , \wRegInB66[27] , \wRegInB73[13] , 
        \wRegInA10[2] , \wAMid27[31] , \wAIn38[7] , \wAMid52[18] , 
        \wBIn105[3] , \wAIn49[13] , \wAMid71[30] , \wRegInB50[22] , 
        \wAMid78[3] , \wRegInA0[21] , \wRegInA0[12] , \wRegInA0[7] , 
        \wRegInB25[12] , \wRegInA80[15] , \wAIn3[26] , \wAIn3[15] , 
        \wBMid6[30] , \wBMid6[29] , \wBIn8[6] , \wAMid8[25] , \wBMid38[16] , 
        \wAMid71[29] , \wAIn121[10] , \ScanLink72[17] , \ScanLink24[16] , 
        \wAIn10[26] , \wBMid11[3] , \wAIn25[8] , \wAIn102[21] , 
        \ScanLink50[6] , \wAIn117[15] , \ScanLink51[26] , \ScanLink219[17] , 
        \ScanLink31[22] , \ScanLink44[12] , \wAIn33[17] , \wAIn46[27] , 
        \wBMid58[12] , \ScanLink67[23] , \ScanLink12[13] , \ScanLink16[3] , 
        \wAIn65[16] , \ScanLink248[4] , \wAMid23[9] , \wBMid57[6] , 
        \wAIn70[22] , \wAMid48[18] , \wAIn53[13] , \wAIn26[23] , 
        \ScanLink128[1] , \wAIn118[21] , \wRegInB69[13] , \wRegInA84[1] , 
        \wRegInA101[30] , \ScanLink216[23] , \wRegInA122[18] , \wBMid22[16] , 
        \wBMid74[17] , \wRegInA101[29] , \ScanLink235[12] , \ScanLink190[15] , 
        \wBMid57[26] , \wRegInB36[2] , \ScanLink240[22] , \ScanLink68[17] , 
        \wBMid37[22] , \wBMid42[12] , \wBMid85[0] , \ScanLink220[26] , 
        \ScanLink185[21] , \ScanLink255[16] , \wAMid7[11] , \wBMid14[13] , 
        \wBMid61[23] , \ScanLink203[17] , \wRegInA56[7] , \wBIn18[2] , 
        \wBMid86[3] , \wRegInB35[1] , \ScanLink256[8] , \wRegInA55[4] , 
        \ScanLink148[25] , \ScanLink93[16] , \ScanLink128[21] , 
        \wRegInA22[21] , \wRegInA74[20] , \wRegInB126[9] , \ScanLink86[22] , 
        \ScanLink15[0] , \wRegInA37[15] , \wRegInA57[11] , \wRegInB87[26] , 
        \wRegInB92[12] , \wBMid42[21] , \wBMid54[5] , \wAMid90[31] , 
        \wRegInA87[2] , \wRegInA14[24] , \wRegInA42[25] , \wAMid90[28] , 
        \wBMid110[8] , \wRegInA61[14] , \ScanLink255[25] , \wAMid3[9] , 
        \wAMid7[22] , \wBMid37[11] , \wRegInB52[6] , \ScanLink220[15] , 
        \ScanLink185[12] , \wAIn10[15] , \wBMid14[20] , \wBMid61[10] , 
        \wBMid22[25] , \wBMid57[15] , \wBMid74[24] , \wAIn118[12] , 
        \ScanLink203[24] , \wBIn127[2] , \ScanLink216[10] , \wRegInA32[3] , 
        \ScanLink240[11] , \ScanLink235[21] , \ScanLink190[26] , \wAIn26[10] , 
        \wAIn70[11] , \ScanLink68[24] , \wRegInB80[0] , \wBIn27[28] , 
        \wAIn53[20] , \wRegInB69[20] , \ScanLink72[7] , \wAIn33[24] , 
        \wAIn46[14] , \wAMid105[3] , \wBIn52[18] , \wBIn71[30] , \wBIn27[31] , 
        \wBMid30[1] , \wBMid33[2] , \wAIn65[25] , \wBIn71[29] , \wAMid88[4] , 
        \wBIn112[18] , \wRegInA14[17] , \wRegInA37[26] , \wRegInA42[16] , 
        \wRegInB92[21] , \ScanLink71[4] , \wRegInA61[27] , \wRegInB83[3] , 
        \wAMid106[0] , \wRegInA22[12] , \wRegInA57[22] , \wRegInA74[13] , 
        \wRegInB87[15] , \wAMid114[18] , \ScanLink128[12] , \ScanLink86[11] , 
        \wBMid4[0] , \wBMid7[3] , \wAIn19[5] , \wAMid59[1] , \wRegInB51[5] , 
        \ScanLink93[25] , \wBIn61[9] , \wAMid96[8] , \ScanLink148[16] , 
        \wBIn124[1] , \ScanLink152[9] , \wRegInA31[0] , \wAMid15[26] , 
        \wAMid25[7] , \wBMid29[30] , \wRegInB123[4] , \ScanLink208[31] , 
        \ScanLink208[28] , \ScanLink63[31] , \ScanLink35[29] , \wBMid51[8] , 
        \wAIn65[3] , \ScanLink40[19] , \wBMid115[5] , \ScanLink35[30] , 
        \ScanLink16[18] , \wBMid29[29] , \ScanLink63[28] , \wAMid23[23] , 
        \wAMid36[17] , \wBIn39[10] , \wAMid60[16] , \ScanLink253[5] , 
        \wAMid43[27] , \wRegInB54[30] , \wRegInB77[18] , \wAIn38[31] , 
        \wAIn38[28] , \wAMid56[13] , \wRegInA50[9] , \ScanLink133[0] , 
        \wBIn59[14] , \wRegInB54[29] , \wAMid38[8] , \wBIn119[14] , 
        \wRegInB21[19] , \wAMid75[22] , \wBIn81[24] , \wBIn94[10] , 
        \wBMid113[11] , \ScanLink4[16] , \ScanLink250[6] , \wAIn95[31] , 
        \wAIn95[28] , \wBMid106[25] , \wBMid125[14] , \ScanLink130[3] , 
        \wRegInB6[17] , \wRegInB120[7] , \wRegInB124[16] , \wAMid26[4] , 
        \wBMid84[30] , \wBMid116[6] , \wRegInB107[27] , \wRegInB112[13] , 
        \ScanLink98[29] , \wAMid6[4] , \wAMid23[10] , \wAMid56[20] , 
        \wAIn66[0] , \ScanLink98[30] , \wBMid84[29] , \ScanLink69[6] , 
        \wBIn59[27] , \wRegInA116[2] , \wBIn119[27] , \wAIn8[19] , 
        \wAMid15[15] , \wBMid28[3] , \wAMid60[25] , \wAMid75[11] , 
        \ScanLink237[1] , \wRegInB54[8] , \wRegInA91[19] , \wAMid36[24] , 
        \wBIn39[23] , \wAMid43[14] , \wAMid93[5] , \ScanLink157[4] , 
        \wBIn64[4] , \wRegInB9[7] , \wRegInB49[7] , \ScanLink74[9] , 
        \wAMid41[3] , \wAIn125[28] , \wAIn106[19] , \ScanLink185[2] , 
        \wAIn125[31] , \wRegInA29[2] , \wRegInB112[20] , \ScanLink115[28] , 
        \wAIn1[4] , \wBIn5[31] , \wBIn5[28] , \ScanLink160[18] , 
        \ScanLink143[30] , \ScanLink143[29] , \ScanLink136[19] , 
        \ScanLink115[31] , \wAMid5[7] , \wAMid42[0] , \wRegInB6[24] , 
        \wRegInB107[14] , \wRegInB124[25] , \ScanLink186[1] , \ScanLink149[8] , 
        \ScanLink234[2] , \wBIn67[7] , \wBIn81[17] , \wRegInB98[2] , 
        \wBMid106[16] , \wBMid125[27] , \wRegInA115[1] , \wAMid90[6] , 
        \wBIn94[23] , \wBMid113[22] , \wRegInA49[29] , \ScanLink154[7] , 
        \ScanLink4[25] , \wRegInA49[30] , \wBIn1[19] , \wBMid12[9] , 
        \ScanLink164[29] , \wAIn26[2] , \wAMid66[6] , \wRegInB116[11] , 
        \ScanLink111[19] , \ScanLink132[31] , \wBIn91[7] , \wRegInA4[10] , 
        \ScanLink164[30] , \ScanLink147[18] , \wAMid124[8] , \ScanLink132[28] , 
        \wAMid27[21] , \wBIn40[2] , \wBIn43[1] , \wBIn85[26] , \wBMid102[27] , 
        \wRegInB2[15] , \wRegInB103[25] , \wRegInB120[14] , \ScanLink170[1] , 
        \wBIn90[12] , \wBIn106[9] , \wBMid121[16] , \wRegInA13[8] , 
        \wRegInA38[28] , \wBMid117[13] , \wRegInA38[31] , \ScanLink210[4] , 
        \ScanLink0[14] , \wBIn28[26] , \wAMid52[11] , \ScanLink173[2] , 
        \wAIn2[7] , \wBMid9[14] , \wAMid11[24] , \wAMid71[20] , \wAMid32[15] , 
        \wAMid64[14] , \ScanLink213[7] , \wBIn108[22] , \wRegInA95[28] , 
        \ScanLink82[9] , \wAMid47[25] , \wBIn48[22] , \wRegInA95[31] , 
        \wAIn25[1] , \wBIn92[4] , \wBIn118[5] , \wBMid9[27] , \wBIn27[5] , 
        \wAMid65[5] , \wAIn102[31] , \wAIn121[19] , \wAIn102[28] , \wBIn39[9] , 
        \wAIn42[6] , \wBIn85[15] , \wAIn90[0] , \wAIn116[2] , \ScanLink114[5] , 
        \wBIn90[21] , \wAIn91[19] , \wBMid117[20] , \wRegInB88[31] , 
        \ScanLink0[27] , \wBMid102[14] , \wRegInB17[9] , \wBMid121[25] , 
        \wRegInB88[28] , \wRegInB2[26] , \wRegInB120[27] , \wBMid80[18] , 
        \wRegInA4[23] , \wRegInB103[16] , \wRegInB116[22] , \wRegInB104[1] , 
        \ScanLink37[8] , \wAIn41[5] , \wBMid58[31] , \wRegInA69[0] , 
        \ScanLink44[28] , \ScanLink12[30] , \wAMid11[17] , \wBMid58[28] , 
        \wRegInB107[2] , \ScanLink67[19] , \ScanLink44[31] , \ScanLink31[18] , 
        \ScanLink12[29] , \wAMid64[27] , \wBMid68[1] , \wBIn108[11] , 
        \wBIn24[6] , \wAMid47[16] , \wBIn48[11] , \ScanLink117[6] , 
        \wAMid27[12] , \wAMid32[26] , \wAIn115[1] , \wAIn49[29] , 
        \wAMid52[22] , \wAIn93[3] , \wRegInB25[31] , \ScanLink29[4] , 
        \wRegInB73[29] , \wBIn28[15] , \wRegInB25[28] , \wBIn0[20] , 
        \wBMid2[18] , \wAMid3[13] , \wAIn7[17] , \wBMid14[7] , \wAIn49[30] , 
        \wBIn58[0] , \wAMid71[13] , \wBIn97[9] , \wRegInB50[18] , 
        \wRegInB73[30] , \wRegInA33[17] , \wRegInB96[10] , \wAMid122[6] , 
        \wRegInA46[27] , \wBMid33[20] , \wAMid60[8] , \wRegInA10[26] , 
        \wRegInA65[16] , \wBIn100[7] , \wBMid109[18] , \wAMid110[30] , 
        \wRegInA70[22] , \wAMid110[29] , \wRegInA26[23] , \ScanLink55[2] , 
        \wRegInB83[24] , \wRegInA15[6] , \wRegInA53[13] , \ScanLink159[13] , 
        \wRegInA5[3] , \ScanLink82[20] , \wRegInB75[3] , \ScanLink139[17] , 
        \ScanLink97[14] , \ScanLink9[1] , \ScanLink87[4] , \ScanLink79[21] , 
        \wBMid46[10] , \ScanLink224[24] , \ScanLink181[23] , \wBMid10[11] , 
        \wRegInA6[0] , \ScanLink251[14] , \wBMid65[21] , \wBIn89[5] , 
        \ScanLink207[15] , \wRegInA16[5] , \wBIn103[4] , \wAIn4[9] , 
        \wBMid17[4] , \wBMid26[14] , \wBMid70[15] , \wAIn109[17] , 
        \ScanLink212[21] , \ScanLink84[7] , \ScanLink231[10] , 
        \ScanLink215[9] , \ScanLink194[17] , \wBMid53[24] , \ScanLink244[20] , 
        \wAIn74[20] , \wRegInB76[0] , \ScanLink19[25] , \wAIn14[24] , 
        \wAIn22[21] , \wAIn57[11] , \wRegInB18[21] , \ScanLink168[3] , 
        \wBIn23[19] , \wAIn37[15] , \wAIn42[25] , \wBIn56[29] , \wBIn116[30] , 
        \wAMid121[5] , \ScanLink99[8] , \ScanLink56[1] , \wRegInB78[25] , 
        \wBIn56[30] , \wAIn61[14] , \wBIn116[29] , \ScanLink208[6] , 
        \wBIn75[18] , \wAIn14[17] , \wAMid19[3] , \ScanLink97[27] , 
        \wAIn37[26] , \wAIn44[8] , \wAIn59[7] , \wRegInA71[2] , 
        \ScanLink139[24] , \wBMid70[3] , \wRegInB9[19] , \ScanLink159[20] , 
        \wRegInB11[7] , \wRegInB108[30] , \wRegInB108[29] , \ScanLink82[13] , 
        \wRegInA70[11] , \wRegInA26[10] , \wRegInA53[20] , \wRegInB83[17] , 
        \wAMid94[19] , \wRegInA33[24] , \wRegInA46[14] , \wRegInB96[23] , 
        \ScanLink31[6] , \wRegInA10[15] , \wRegInA65[25] , \wRegInB78[16] , 
        \wAIn42[16] , \wBMid73[0] , \wAIn88[2] , \wAIn22[12] , \wAIn61[27] , 
        \wAIn74[13] , \wAMid39[19] , \ScanLink32[5] , \wAIn57[22] , 
        \wBMid70[26] , \wRegInB18[12] , \ScanLink111[8] , \wAMid3[20] , 
        \wAIn7[24] , \wBIn22[8] , \wBMid26[27] , \wBMid53[17] , \wRegInA72[1] , 
        \wRegInA126[29] , \ScanLink212[12] , \ScanLink244[13] , 
        \wRegInA126[30] , \ScanLink231[23] , \ScanLink19[16] , 
        \ScanLink194[24] , \wBMid46[23] , \wRegInA105[18] , \wBMid33[13] , 
        \wRegInB12[4] , \ScanLink251[27] , \ScanLink79[12] , \ScanLink224[17] , 
        \ScanLink181[10] , \wAMid9[15] , \wBMid10[22] , \wBMid65[12] , 
        \wAIn109[24] , \wAMid26[18] , \wAIn28[27] , \wRegInB12[27] , 
        \ScanLink207[26] , \wAIn48[23] , \wAMid53[31] , \wAMid70[19] , 
        \wAIn83[9] , \wRegInB24[22] , \wRegInB31[16] , \wRegInA64[5] , 
        \wRegInB67[17] , \wRegInA94[11] , \wRegInB44[26] , \wRegInA81[25] , 
        \wRegInB51[12] , \wAMid53[28] , \wRegInB72[23] , \wBIn29[3] , 
        \ScanLink50[16] , \wAIn118[4] , \wAMid12[8] , \wBMid39[26] , 
        \wAIn103[11] , \ScanLink25[26] , \ScanLink73[27] , \wBMid59[22] , 
        \wBMid65[4] , \wAIn120[20] , \wBMid121[9] , \wRegInB117[8] , 
        \ScanLink66[13] , \wBMid66[7] , \wAIn116[25] , \ScanLink218[27] , 
        \ScanLink13[23] , \ScanLink45[22] , \ScanLink24[1] , \ScanLink30[12] , 
        \ScanLink105[14] , \wBMid81[12] , \wBMid94[26] , \ScanLink170[24] , 
        \ScanLink88[26] , \wRegInB117[31] , \ScanLink153[15] , 
        \ScanLink126[25] , \ScanLink119[0] , \ScanLink133[11] , \wRegInA5[30] , 
        \ScanLink27[2] , \wRegInA5[29] , \wRegInB117[28] , \ScanLink146[21] , 
        \ScanLink110[20] , \ScanLink165[10] , \wBIn0[13] , \wAMid9[26] , 
        \wBMid59[11] , \wAIn85[27] , \wAIn90[13] , \wAIn106[8] , 
        \wRegInA39[11] , \wRegInA59[15] , \wRegInA67[6] , \wRegInB89[22] , 
        \wRegInB109[4] , \wAIn116[16] , \ScanLink66[20] , \ScanLink13[10] , 
        \ScanLink218[14] , \ScanLink30[21] , \ScanLink45[11] , 
        \ScanLink25[15] , \wAIn28[14] , \wAIn28[4] , \wBMid39[15] , 
        \wAIn103[22] , \ScanLink40[5] , \wAIn120[13] , \ScanLink50[25] , 
        \ScanLink73[14] , \wBIn50[8] , \wAMid68[0] , \wRegInB51[21] , 
        \ScanLink1[9] , \wRegInB24[11] , \wRegInA81[16] , \wBIn115[0] , 
        \wRegInB72[10] , \ScanLink163[8] , \wAIn48[10] , \ScanLink92[3] , 
        \wAIn36[8] , \wBIn49[31] , \wBIn49[28] , \wRegInB67[24] , 
        \wBIn109[31] , \wRegInB12[14] , \wRegInB44[15] , \wAIn85[14] , 
        \wAIn90[20] , \wBIn109[28] , \wRegInB60[4] , \wRegInA94[22] , 
        \wBIn116[3] , \wRegInB31[25] , \wRegInA59[26] , \wRegInB89[11] , 
        \wBIn91[18] , \wBMid116[19] , \wRegInA39[22] , \wRegInB63[7] , 
        \ScanLink91[0] , \ScanLink146[12] , \wBMid81[21] , \ScanLink133[22] , 
        \ScanLink165[23] , \wAMid2[19] , \wBMid3[12] , \wBIn32[2] , 
        \wBMid94[15] , \ScanLink170[17] , \ScanLink110[13] , \ScanLink88[15] , 
        \ScanLink153[26] , \ScanLink105[27] , \ScanLink43[6] , 
        \wRegInA104[12] , \ScanLink245[19] , \ScanLink126[16] , 
        \ScanLink230[29] , \ScanLink101[2] , \wBMid11[31] , \wBMid11[28] , 
        \wBMid47[30] , \wBMid64[18] , \wAIn85[7] , \wAIn103[5] , 
        \ScanLink230[30] , \ScanLink213[18] , \wRegInA127[23] , \wBMid32[19] , 
        \wBMid47[29] , \ScanLink78[18] , \wBIn14[25] , \wAMid17[5] , 
        \wBIn117[10] , \wRegInA111[26] , \wBIn22[20] , \wBIn74[21] , 
        \wAIn23[18] , \wBIn37[14] , \wAMid38[13] , \wAIn57[1] , \wBIn57[10] , 
        \wAMid58[17] , \wAIn98[8] , \wBIn42[24] , \wAIn56[28] , \wBIn121[15] , 
        \wRegInB19[18] , \wBIn14[16] , \wAMid14[6] , \wAIn54[2] , \wAIn56[31] , 
        \wBIn61[15] , \wAIn75[19] , \wRegInB111[6] , \wBIn102[24] , 
        \wAMid111[10] , \wBMid60[9] , \wBMid124[4] , \wAMid80[27] , 
        \wBMid108[21] , \wBIn31[1] , \wAMid95[13] , \wAMid104[24] , 
        \wRegInB97[30] , \wRegInB112[5] , \wRegInB97[29] , \wAIn33[5] , 
        \wBIn37[27] , \wAMid38[20] , \wBIn42[17] , \wAIn86[4] , \wAIn100[6] , 
        \ScanLink102[1] , \wRegInB8[13] , \wRegInA61[8] , \wRegInB109[23] , 
        \ScanLink83[19] , \wBIn84[0] , \wBIn121[26] , \ScanLink178[9] , 
        \wBIn61[26] , \wBIn102[17] , \wBIn22[13] , \wBIn57[23] , \wAMid73[1] , 
        \wBIn74[12] , \wBIn117[23] , \ScanLink89[2] , \ScanLink7[7] , 
        \wAMid58[24] , \wBIn56[6] , \ScanLink180[30] , \ScanLink165[6] , 
        \wBMid3[21] , \wRegInA104[21] , \wRegInA111[15] , \ScanLink205[3] , 
        \ScanLink180[29] , \wRegInA127[10] , \wBMid19[2] , \wRegInB109[10] , 
        \wRegInA124[0] , \wAIn30[6] , \wBIn55[5] , \wRegInB8[20] , 
        \ScanLink166[5] , \wAMid70[2] , \wAMid95[20] , \wRegInA8[6] , 
        \wRegInB65[9] , \wRegInA127[3] , \ScanLink158[19] , \ScanLink58[7] , 
        \ScanLink206[0] , \wBIn87[3] , \wAMid104[17] , \wAMid80[14] , 
        \wBMid108[12] , \wAMid111[23] , \wRegInA18[3] , \wRegInA27[29] , 
        \ScanLink45[8] , \wRegInA27[30] , \wRegInA52[19] , \wRegInA71[31] , 
        \wRegInA71[28] , \wRegInB78[6] , \ScanLink4[4] , \wBIn0[22] , 
        \wBIn4[22] , \wBIn5[3] , \wBIn6[0] , \wAMid6[31] , \wAMid6[28] , 
        \wBIn10[27] , \wAIn14[0] , \wBIn71[3] , \wRegInA103[5] , 
        \ScanLink222[6] , \ScanLink129[18] , \wAMid86[2] , \wRegInB118[15] , 
        \ScanLink142[3] , \wAMid91[11] , \wAMid100[26] , \wBMid119[17] , 
        \wAMid123[17] , \wRegInB93[9] , \wAMid115[12] , \wRegInA23[18] , 
        \wRegInA56[28] , \ScanLink190[5] , \wBIn33[16] , \wAMid54[4] , 
        \wAMid84[25] , \wRegInA56[31] , \wRegInA75[19] , \wBIn46[26] , 
        \wAMid49[21] , \wBIn125[17] , \wAIn17[3] , \wBMid23[8] , \wBIn65[17] , 
        \wBIn106[26] , \wBIn26[22] , \wAMid57[7] , \wBIn70[23] , \wBIn113[12] , 
        \ScanLink193[6] , \wAMid29[25] , \wBIn53[12] , \wAMid115[9] , 
        \wRegInA100[6] , \wBMid7[10] , \wBIn72[0] , \wAMid85[1] , 
        \wRegInA115[24] , \ScanLink221[5] , \ScanLink184[18] , \wAIn119[18] , 
        \wRegInA100[10] , \ScanLink141[0] , \wAMid30[0] , \wAMid84[16] , 
        \wAMid108[6] , \wAMid115[21] , \wRegInA22[9] , \wRegInA123[21] , 
        \wRegInB38[4] , \wAMid91[22] , \wBMid100[2] , \wAMid123[24] , 
        \wBMid119[24] , \wBMid59[0] , \wAIn70[4] , \wAMid100[15] , 
        \wRegInB93[18] , \wBMid96[9] , \wRegInA58[1] , \wRegInA97[8] , 
        \wRegInB118[26] , \ScanLink18[5] , \ScanLink246[2] , \ScanLink87[28] , 
        \wBMid7[23] , \wBIn15[7] , \wAIn124[0] , \ScanLink126[7] , 
        \wRegInB26[8] , \wRegInA100[23] , \ScanLink245[1] , \ScanLink234[18] , 
        \ScanLink217[30] , \ScanLink87[31] , \ScanLink241[28] , 
        \wRegInA123[12] , \ScanLink217[29] , \ScanLink241[31] , \wBIn16[4] , 
        \wBMid15[19] , \wAIn127[3] , \wBMid36[31] , \wAMid8[2] , \wBIn10[14] , 
        \wBIn26[11] , \wBMid36[28] , \wBMid60[29] , \ScanLink125[4] , 
        \wRegInA89[4] , \wRegInA115[17] , \wBMid43[18] , \wBIn53[21] , 
        \wBMid60[30] , \wBIn70[10] , \wBIn113[21] , \wAIn27[30] , \wAIn27[29] , 
        \wAMid29[16] , \wBIn46[15] , \wAMid49[12] , \wAIn71[31] , \wAIn52[19] , 
        \wBIn125[24] , \wBIn33[25] , \wBIn65[24] , \wAIn71[28] , \wAIn73[7] , 
        \wRegInB68[19] , \wBMid103[1] , \wBMid88[5] , \wBIn106[15] , 
        \wAMid33[3] , \wAIn81[25] , \wAIn94[11] , \wRegInA28[27] , 
        \wRegInB88[8] , \ScanLink224[8] , \wRegInB47[1] , \wBMid85[10] , 
        \wBIn95[30] , \wBIn95[29] , \wBMid112[28] , \wRegInB7[1] , 
        \wRegInB98[14] , \wBMid112[31] , \wRegInA27[4] , \wRegInA48[23] , 
        \ScanLink137[13] , \wRegInA118[4] , \ScanLink142[23] , \ScanLink67[0] , 
        \ScanLink239[7] , \ScanLink114[22] , \wRegInB95[7] , \ScanLink161[12] , 
        \ScanLink99[10] , \wBIn4[11] , \wAIn9[13] , \wBMid25[6] , \wBMid26[5] , 
        \wBMid28[10] , \wBMid90[24] , \ScanLink174[26] , \ScanLink101[16] , 
        \wAMid110[4] , \ScanLink159[2] , \ScanLink122[27] , \ScanLink157[17] , 
        \wBIn69[1] , \wAIn112[27] , \wRegInB96[4] , \ScanLink62[11] , 
        \ScanLink17[21] , \ScanLink64[3] , \ScanLink41[20] , \ScanLink54[14] , 
        \ScanLink34[10] , \wAIn107[13] , \wAMid113[7] , \ScanLink209[11] , 
        \ScanLink195[8] , \wRegInA39[8] , \ScanLink21[24] , \ScanLink77[25] , 
        \wBMid48[14] , \wAMid51[9] , \wAIn124[22] , \wBIn38[30] , \wBIn38[29] , 
        \wAIn39[11] , \wRegInB20[20] , \wRegInB44[2] , \wRegInB55[10] , 
        \wRegInA85[27] , \wRegInB76[21] , \wRegInA106[8] , \wAIn59[15] , 
        \wRegInB16[25] , \ScanLink188[7] , \wBMid38[9] , \wRegInA24[7] , 
        \wRegInB63[15] , \wRegInB35[14] , \wRegInA90[13] , \wRegInB4[2] , 
        \wBMid85[23] , \wBMid90[17] , \wRegInB40[24] , \ScanLink174[15] , 
        \ScanLink157[24] , \ScanLink101[25] , \wRegInA91[6] , 
        \ScanLink142[10] , \ScanLink122[14] , \ScanLink137[20] , 
        \ScanLink161[21] , \wAIn9[20] , \wBMid9[5] , \wBMid42[1] , 
        \ScanLink99[23] , \wAIn81[16] , \wRegInA1[18] , \wRegInB113[19] , 
        \ScanLink114[11] , \wRegInB23[5] , \wBIn13[9] , \wRegInA48[10] , 
        \wRegInB98[27] , \ScanLink120[9] , \wAMid22[30] , \wAIn59[26] , 
        \wBMid90[7] , \wRegInA28[14] , \wRegInA43[0] , \wAIn94[22] , 
        \wRegInB63[26] , \wBMid118[0] , \wRegInB16[16] , \wRegInB20[6] , 
        \wRegInB40[17] , \wRegInB35[27] , \wRegInA90[20] , \wRegInB55[23] , 
        \wAMid22[29] , \wAMid28[2] , \wBMid93[4] , \wAIn39[22] , \wAMid74[28] , 
        \wRegInB20[13] , \wRegInA85[14] , \wRegInB76[12] , \wBMid48[27] , 
        \wAMid57[19] , \wRegInA40[3] , \wAIn68[6] , \wAMid74[31] , 
        \wAIn107[20] , \ScanLink21[17] , \ScanLink209[22] , \ScanLink54[27] , 
        \wBMid28[23] , \wBMid41[2] , \wAIn124[11] , \ScanLink77[16] , 
        \ScanLink17[12] , \wAIn75[9] , \wAIn112[14] , \ScanLink62[22] , 
        \ScanLink34[23] , \wAIn80[8] , \wAIn85[25] , \wAIn90[11] , 
        \wRegInA59[17] , \wRegInA92[5] , \ScanLink41[13] , \wRegInB89[20] , 
        \wRegInB109[6] , \wBIn91[29] , \wBMid116[28] , \wBIn91[30] , 
        \wBMid116[31] , \wRegInA67[4] , \wBMid81[10] , \wRegInA39[13] , 
        \ScanLink146[23] , \ScanLink133[13] , \ScanLink27[0] , 
        \ScanLink165[12] , \wBIn0[11] , \wAMid9[17] , \wBMid59[20] , 
        \wBMid66[5] , \wBMid122[8] , \wRegInB114[9] , \ScanLink170[26] , 
        \ScanLink110[22] , \ScanLink88[24] , \wBMid94[24] , \ScanLink153[17] , 
        \ScanLink105[16] , \ScanLink126[27] , \ScanLink119[2] , 
        \ScanLink13[21] , \wAIn116[27] , \ScanLink66[11] , \ScanLink218[25] , 
        \ScanLink30[10] , \ScanLink24[3] , \ScanLink45[20] , \ScanLink25[24] , 
        \wAMid11[9] , \wBIn29[1] , \wAIn103[13] , \wAIn118[6] , \wRegInA79[8] , 
        \ScanLink50[14] , \wAIn28[25] , \wBMid39[24] , \wAIn120[22] , 
        \wAIn48[21] , \wBMid65[6] , \ScanLink73[25] , \wRegInB24[20] , 
        \wRegInB51[10] , \wRegInA81[27] , \wRegInB72[21] , \wBIn49[19] , 
        \wRegInA64[7] , \wRegInB67[15] , \wBMid78[9] , \wAIn105[9] , 
        \wBIn109[19] , \wRegInB12[25] , \wRegInB44[24] , \wRegInB31[14] , 
        \wRegInA94[13] , \wBMid81[23] , \wBMid94[17] , \ScanLink170[15] , 
        \ScanLink105[25] , \ScanLink2[8] , \ScanLink88[17] , \ScanLink153[24] , 
        \ScanLink126[14] , \ScanLink43[4] , \ScanLink133[20] , \wRegInA5[18] , 
        \wRegInB117[19] , \ScanLink146[10] , \ScanLink110[11] , 
        \ScanLink165[21] , \wAMid2[31] , \wAMid2[28] , \wAMid9[24] , 
        \wAMid26[30] , \wAIn28[16] , \wBIn53[9] , \wAIn85[16] , \wRegInB63[5] , 
        \wBIn116[1] , \wRegInA39[20] , \wRegInB89[13] , \ScanLink91[2] , 
        \wRegInA59[24] , \ScanLink160[9] , \wAIn90[22] , \wRegInB12[16] , 
        \wAMid68[2] , \wRegInB24[13] , \wRegInB31[27] , \wRegInB67[26] , 
        \ScanLink92[1] , \wRegInB44[17] , \wRegInB60[6] , \wRegInA94[20] , 
        \wRegInA81[14] , \wAMid70[28] , \wRegInB51[23] , \wAMid26[29] , 
        \wAIn28[6] , \wAIn48[12] , \wAMid70[31] , \wBIn115[2] , \wAMid53[19] , 
        \wRegInB72[12] , \ScanLink50[27] , \wBIn14[27] , \wAMid14[4] , 
        \wBIn31[3] , \wAIn35[9] , \wBMid39[17] , \wAIn103[20] , 
        \ScanLink25[17] , \ScanLink40[7] , \wBMid59[13] , \wAIn120[11] , 
        \ScanLink73[16] , \ScanLink66[22] , \ScanLink13[12] , 
        \ScanLink218[16] , \wAIn86[6] , \wAIn116[14] , \ScanLink45[13] , 
        \wRegInB8[11] , \wRegInB109[21] , \ScanLink30[23] , \ScanLink158[31] , 
        \ScanLink158[28] , \wAIn100[4] , \wAIn54[0] , \wAMid95[11] , 
        \wRegInB112[7] , \ScanLink102[3] , \wAMid104[26] , \wRegInA27[18] , 
        \wAMid111[12] , \wRegInA52[28] , \wBIn37[16] , \wBIn42[26] , 
        \wAMid80[25] , \wBMid124[6] , \wRegInA71[19] , \wRegInA52[31] , 
        \wBMid108[23] , \wBIn121[17] , \wAMid38[11] , \wBIn61[17] , 
        \wRegInB111[4] , \wBIn102[26] , \wAMid17[7] , \wBIn74[23] , 
        \wBIn117[12] , \wBIn22[22] , \wAIn57[3] , \wBMid63[8] , \wBIn57[12] , 
        \wAMid58[15] , \wRegInA111[24] , \ScanLink180[18] , \wBMid3[10] , 
        \wAIn85[5] , \wRegInA62[9] , \wRegInA104[10] , \wRegInA127[21] , 
        \wAIn103[7] , \ScanLink101[0] , \wBIn32[0] , \wAMid111[21] , 
        \wRegInB78[4] , \ScanLink4[6] , \wRegInA0[23] , \wRegInA0[10] , 
        \wAMid0[8] , \wAIn3[17] , \wBIn4[20] , \wBMid3[23] , \wBMid19[0] , 
        \wAIn30[4] , \wAMid70[0] , \wAMid80[16] , \wAMid95[22] , 
        \wBMid108[10] , \wRegInA8[4] , \wBIn48[8] , \wBIn87[1] , 
        \wRegInA18[1] , \wAMid104[15] , \wRegInB97[18] , \wRegInB109[12] , 
        \wRegInA127[1] , \ScanLink206[2] , \ScanLink58[5] , \ScanLink83[28] , 
        \wBIn55[7] , \wRegInB8[22] , \ScanLink166[7] , \ScanLink83[31] , 
        \wRegInB66[8] , \ScanLink245[28] , \wRegInA104[23] , \ScanLink230[18] , 
        \ScanLink213[30] , \ScanLink205[1] , \wRegInA124[2] , 
        \ScanLink245[31] , \wBIn5[1] , \wAMid6[19] , \wBMid7[12] , 
        \wBMid11[19] , \wBMid32[31] , \wBIn56[4] , \wBMid64[29] , 
        \wRegInA127[12] , \ScanLink213[29] , \ScanLink78[30] , \wBIn14[14] , 
        \wBIn22[11] , \wBMid32[28] , \wBMid47[18] , \wBMid64[30] , 
        \ScanLink165[4] , \ScanLink78[29] , \wBIn74[10] , \wBIn117[21] , 
        \wRegInA111[17] , \ScanLink7[5] , \wAIn23[30] , \wAIn23[29] , 
        \wBIn37[25] , \wBIn57[21] , \wAMid58[26] , \ScanLink89[0] , 
        \ScanLink46[9] , \wAMid38[22] , \wAIn33[7] , \wBIn42[15] , 
        \wAIn56[19] , \wAIn75[31] , \wAMid73[3] , \wBIn84[2] , \wBIn121[24] , 
        \wRegInB19[29] , \wBIn61[24] , \wAIn75[28] , \wAMid85[3] , 
        \wBIn102[15] , \wRegInB19[30] , \wAMid108[4] , \wRegInA100[12] , 
        \ScanLink234[29] , \ScanLink241[19] , \ScanLink217[18] , 
        \wRegInA123[23] , \ScanLink234[30] , \ScanLink141[2] , \wBIn10[25] , 
        \wBMid15[31] , \wBMid15[28] , \wBIn72[2] , \wRegInA100[4] , 
        \wBMid43[30] , \wBMid60[18] , \wAIn17[1] , \wBMid36[19] , 
        \wRegInA115[26] , \wBMid43[29] , \wAMid57[5] , \wBIn113[10] , 
        \ScanLink221[7] , \wBIn70[21] , \wBIn26[20] , \wAMid29[27] , 
        \wBIn53[10] , \wAIn27[18] , \wBIn46[24] , \ScanLink193[4] , 
        \wAMid49[23] , \wAIn52[28] , \wBIn125[15] , \wBIn33[14] , \wAIn52[31] , 
        \wAIn71[19] , \wRegInB68[28] , \wBIn65[15] , \wBIn106[24] , 
        \wRegInB90[8] , \wBIn10[16] , \wAIn14[2] , \wAMid116[8] , 
        \wRegInB68[31] , \wBMid20[9] , \wAMid54[6] , \wAMid115[10] , 
        \ScanLink190[7] , \wBIn33[27] , \wAMid49[9] , \wBIn71[1] , 
        \wAMid84[27] , \wAMid91[13] , \wBMid119[15] , \wAMid123[15] , 
        \wRegInB93[30] , \wAMid100[24] , \wRegInA21[8] , \wRegInB93[29] , 
        \wRegInB118[17] , \ScanLink142[1] , \wAMid86[0] , \wRegInA103[7] , 
        \ScanLink222[4] , \ScanLink87[19] , \wBIn46[17] , \wAIn73[5] , 
        \wRegInA94[9] , \wAMid49[10] , \wBIn125[26] , \ScanLink138[9] , 
        \wBIn26[13] , \wAMid29[14] , \wAMid33[1] , \wBIn65[26] , \wBIn70[12] , 
        \wBMid88[7] , \wBMid103[3] , \wBIn106[17] , \wBIn113[23] , 
        \wBIn53[23] , \wBIn16[6] , \wRegInA89[6] , \wAIn127[1] , 
        \ScanLink125[6] , \wBIn6[2] , \wBMid7[21] , \wBMid95[8] , 
        \wRegInA115[15] , \ScanLink184[30] , \wAIn119[30] , \ScanLink184[29] , 
        \wAIn119[29] , \wRegInA100[21] , \ScanLink245[3] , \wBMid59[2] , 
        \wRegInA123[10] , \ScanLink129[30] , \ScanLink126[5] , \wAIn9[11] , 
        \wBIn15[5] , \wAMid22[18] , \wAMid30[2] , \wAMid91[20] , 
        \wBMid119[26] , \wAIn124[2] , \ScanLink129[29] , \wRegInB25[9] , 
        \ScanLink18[7] , \wRegInB118[24] , \ScanLink246[0] , \wAIn39[13] , 
        \wAMid57[31] , \wAIn59[17] , \wAIn70[6] , \wBMid100[0] , 
        \wAMid123[26] , \wAMid84[14] , \wAMid100[17] , \wRegInA58[3] , 
        \wAMid115[23] , \wRegInA23[29] , \wRegInA56[19] , \wRegInA75[31] , 
        \wRegInB38[6] , \wRegInA75[28] , \wRegInA23[30] , \wRegInA24[5] , 
        \wRegInB63[17] , \wRegInB4[0] , \wRegInB16[27] , \ScanLink188[5] , 
        \wRegInB20[22] , \wRegInB35[16] , \wRegInB40[26] , \wRegInB44[0] , 
        \wRegInA90[11] , \wRegInB55[12] , \wRegInA85[25] , \wAMid74[19] , 
        \ScanLink227[9] , \wRegInB76[23] , \wBMid48[16] , \wAMid57[28] , 
        \wBIn69[3] , \wAIn107[11] , \wAMid113[5] , \ScanLink21[26] , 
        \ScanLink209[13] , \ScanLink54[16] , \wBMid25[4] , \wAIn124[20] , 
        \ScanLink77[27] , \wBMid26[7] , \wBMid28[12] , \wRegInB96[6] , 
        \ScanLink17[23] , \ScanLink62[13] , \wAMid52[8] , \wAIn112[25] , 
        \ScanLink64[1] , \ScanLink34[12] , \ScanLink41[22] , \ScanLink174[24] , 
        \wBMid85[12] , \wBMid90[26] , \wAMid110[6] , \ScanLink157[15] , 
        \ScanLink101[14] , \wRegInA1[30] , \wRegInB113[31] , \wRegInA118[6] , 
        \ScanLink196[9] , \ScanLink159[0] , \ScanLink142[21] , 
        \ScanLink122[25] , \ScanLink137[11] , \ScanLink67[2] , \wRegInB95[5] , 
        \ScanLink161[10] , \wBIn4[13] , \wAMid8[0] , \wRegInA1[29] , 
        \wRegInB113[28] , \ScanLink99[12] , \ScanLink239[5] , 
        \ScanLink114[20] , \wAIn9[22] , \wBMid28[21] , \wAIn81[27] , 
        \wAIn94[13] , \wRegInB7[3] , \wRegInA27[6] , \wRegInA28[25] , 
        \wRegInA48[21] , \wRegInB98[16] , \wRegInA105[9] , \wRegInB47[3] , 
        \ScanLink62[20] , \wBMid41[0] , \wBMid48[25] , \wAIn107[22] , 
        \wAIn112[16] , \wRegInA92[7] , \ScanLink41[11] , \ScanLink17[10] , 
        \ScanLink209[20] , \ScanLink54[25] , \ScanLink34[21] , 
        \ScanLink21[15] , \ScanLink77[14] , \wAIn124[13] , \wBIn10[8] , 
        \wAMid28[0] , \wRegInB20[11] , \wRegInA85[16] , \wAIn68[4] , 
        \wBMid93[6] , \wBMid118[2] , \wRegInB55[21] , \wRegInA40[1] , 
        \wRegInB76[10] , \wBMid9[7] , \wBIn38[18] , \wAIn39[20] , \wAIn59[24] , 
        \ScanLink123[8] , \wRegInB16[14] , \wBMid90[5] , \wRegInB20[4] , 
        \wRegInB35[25] , \wRegInB63[24] , \wRegInA90[22] , \wRegInA28[16] , 
        \wRegInB40[15] , \wRegInA43[2] , \wAIn94[20] , \wRegInB23[7] , 
        \wBMid42[3] , \wAIn76[8] , \wAIn81[14] , \wBIn95[18] , \wBMid112[19] , 
        \wRegInA48[12] , \wRegInB98[25] , \wRegInA91[4] , \wBMid85[21] , 
        \ScanLink137[22] , \ScanLink161[23] , \ScanLink142[12] , 
        \ScanLink114[13] , \ScanLink99[21] , \wBIn18[0] , \wBMid90[15] , 
        \ScanLink174[17] , \ScanLink101[27] , \wRegInA42[27] , \wRegInA87[0] , 
        \ScanLink157[26] , \ScanLink122[16] , \wRegInA48[9] , \wAMid20[8] , 
        \wRegInA37[17] , \wRegInB92[10] , \wBMid42[10] , \wBMid49[8] , 
        \wBMid54[7] , \wRegInA61[16] , \wBMid86[1] , \wAMid114[30] , 
        \wRegInA14[26] , \wRegInA74[22] , \wAMid114[29] , \wRegInA22[23] , 
        \wRegInA57[13] , \wRegInB87[24] , \ScanLink15[2] , \wRegInA55[6] , 
        \ScanLink128[23] , \ScanLink86[20] , \wRegInB35[3] , \ScanLink148[27] , 
        \ScanLink93[14] , \wBMid6[18] , \wAMid7[13] , \wBMid37[20] , 
        \ScanLink255[14] , \wBMid85[2] , \ScanLink220[24] , \ScanLink185[23] , 
        \wBIn8[4] , \wBMid14[11] , \wBMid61[21] , \wRegInA56[5] , 
        \wBMid22[14] , \wBMid57[24] , \wBMid74[15] , \wAIn118[23] , 
        \ScanLink203[15] , \ScanLink240[20] , \ScanLink216[21] , 
        \wRegInB36[0] , \ScanLink255[9] , \ScanLink235[10] , \ScanLink190[17] , 
        \ScanLink68[15] , \wAIn26[21] , \wBMid57[4] , \wAIn70[20] , 
        \wBMid113[9] , \wAIn53[11] , \wRegInB69[11] , \wRegInA84[3] , 
        \ScanLink128[3] , \wAIn10[24] , \wBIn27[19] , \wAIn33[15] , 
        \wAIn46[25] , \wBIn112[30] , \wBIn52[29] , \ScanLink16[1] , 
        \wAIn10[17] , \wAIn19[7] , \wBIn52[30] , \wAIn65[14] , \wBIn71[18] , 
        \wBIn112[29] , \wRegInB125[8] , \ScanLink248[6] , \wAMid59[3] , 
        \wBIn124[3] , \wRegInA31[2] , \ScanLink93[27] , \wBMid30[3] , 
        \wRegInB51[7] , \ScanLink148[14] , \ScanLink128[10] , \wRegInA74[11] , 
        \ScanLink86[13] , \wAIn33[26] , \wAIn46[16] , \wAMid90[19] , 
        \wAMid106[2] , \wRegInA22[10] , \wRegInB87[17] , \wRegInA14[15] , 
        \wRegInA37[24] , \wRegInA57[20] , \wRegInA42[14] , \wRegInB92[23] , 
        \ScanLink71[6] , \wRegInB83[1] , \wAMid105[1] , \wRegInA61[25] , 
        \wBMid33[0] , \wAIn65[27] , \wAMid88[6] , \wAIn26[12] , \wAMid48[30] , 
        \wAMid48[29] , \wAIn53[22] , \wAIn70[13] , \wRegInB80[2] , 
        \ScanLink72[5] , \wBIn62[8] , \wAIn118[10] , \wBIn127[0] , 
        \wRegInA32[1] , \wRegInB69[22] , \ScanLink216[12] , \wRegInA122[29] , 
        \ScanLink151[8] , \wBMid22[27] , \wBMid74[26] , \wAMid95[9] , 
        \ScanLink235[23] , \ScanLink190[24] , \wRegInA101[18] , 
        \wRegInA122[30] , \ScanLink68[26] , \wBMid37[13] , \wBMid57[17] , 
        \ScanLink240[13] , \wRegInB52[4] , \wBMid42[23] , \ScanLink220[17] , 
        \ScanLink185[10] , \wAIn3[24] , \wAMid7[20] , \wBMid14[22] , 
        \ScanLink255[27] , \wBMid61[12] , \ScanLink203[26] , \wRegInB112[11] , 
        \ScanLink136[31] , \ScanLink115[19] , \wBIn5[19] , \wAMid26[6] , 
        \ScanLink160[29] , \wBMid4[2] , \wBMid52[9] , \wAIn66[2] , 
        \wBMid116[4] , \ScanLink136[28] , \wRegInB6[15] , \ScanLink160[30] , 
        \ScanLink143[18] , \wRegInB107[25] , \wRegInB120[5] , \wRegInB124[14] , 
        \wAMid5[5] , \wAIn8[31] , \wAIn8[28] , \wBMid7[1] , \wAMid15[24] , 
        \wAMid23[21] , \wAMid56[11] , \wBIn59[16] , \wBIn81[26] , 
        \wBMid106[27] , \wBIn94[12] , \wBMid125[16] , \wRegInA53[8] , 
        \ScanLink130[1] , \wRegInA49[18] , \wBMid113[13] , \ScanLink250[4] , 
        \ScanLink4[14] , \ScanLink133[2] , \wAMid60[14] , \wAMid75[20] , 
        \wBIn119[16] , \wBMid108[8] , \wRegInA91[28] , \ScanLink253[7] , 
        \wAMid25[5] , \wAMid36[15] , \wAMid43[25] , \wRegInA91[31] , 
        \wBIn39[12] , \wAIn65[1] , \wBMid115[7] , \wAIn106[31] , 
        \wRegInB123[6] , \wAIn106[28] , \wAIn125[19] , \wBIn67[5] , 
        \wBIn81[15] , \wAMid90[4] , \wBIn94[21] , \ScanLink154[5] , 
        \wBMid113[20] , \ScanLink4[27] , \wBMid106[14] , \wRegInB98[0] , 
        \wAIn95[19] , \wRegInB57[9] , \ScanLink234[0] , \wAMid42[2] , 
        \wBMid125[25] , \wRegInA115[3] , \wRegInB6[26] , \wRegInB124[27] , 
        \ScanLink186[3] , \wRegInB107[16] , \wRegInB112[22] , \ScanLink98[18] , 
        \wAIn2[5] , \wAMid6[6] , \wAMid15[17] , \wBMid29[18] , \wAMid41[1] , 
        \wBMid84[18] , \wRegInB9[5] , \ScanLink77[8] , \wBIn79[9] , 
        \wRegInA29[0] , \wRegInB49[5] , \ScanLink208[19] , \ScanLink185[0] , 
        \ScanLink40[28] , \ScanLink35[18] , \ScanLink16[30] , \ScanLink16[29] , 
        \wAMid93[7] , \ScanLink63[19] , \ScanLink40[31] , \wAMid23[12] , 
        \wBMid28[1] , \wAMid60[27] , \wAMid36[26] , \wBIn39[21] , 
        \wAMid43[16] , \wBIn64[6] , \ScanLink157[6] , \wRegInB77[29] , 
        \wRegInA116[0] , \wAIn38[19] , \wAMid56[22] , \wBIn59[25] , 
        \wRegInB21[31] , \ScanLink69[4] , \wRegInB54[18] , \wRegInB77[30] , 
        \wBMid9[16] , \wAIn25[3] , \wAMid75[13] , \wBIn119[25] , 
        \wRegInB21[28] , \wBIn118[7] , \ScanLink237[3] , \ScanLink44[19] , 
        \wBIn92[6] , \ScanLink67[31] , \ScanLink31[29] , \wBMid11[8] , 
        \wAMid65[7] , \ScanLink67[28] , \wBMid58[19] , \ScanLink12[18] , 
        \wAMid11[26] , \wAMid64[16] , \ScanLink31[30] , \wBIn108[20] , 
        \ScanLink213[5] , \wAMid27[23] , \wBIn28[24] , \wAMid32[17] , 
        \wAMid47[27] , \wBIn48[20] , \wBIn40[0] , \wAIn49[18] , \wAMid52[13] , 
        \wBIn105[8] , \wRegInA10[9] , \wRegInB50[30] , \wRegInB73[18] , 
        \ScanLink173[0] , \wAMid78[8] , \wAIn1[6] , \wBIn43[3] , \wAMid71[22] , 
        \wRegInB25[19] , \wBIn85[24] , \wBIn90[10] , \wBMid117[11] , 
        \wRegInB50[29] , \ScanLink81[8] , \ScanLink0[16] , \wAIn91[28] , 
        \ScanLink210[6] , \wBMid102[25] , \wBMid121[14] , \wRegInB88[19] , 
        \ScanLink170[3] , \wAMid66[4] , \wBMid80[30] , \wAIn91[31] , 
        \wRegInB2[17] , \wRegInA4[12] , \wRegInB103[27] , \wRegInB120[16] , 
        \wRegInB116[13] , \wAIn26[0] , \wAMid27[10] , \wBIn28[17] , 
        \wBMid80[29] , \wBIn91[5] , \wAMid52[20] , \ScanLink29[6] , 
        \wRegInB14[8] , \wRegInA0[19] , \wBIn1[31] , \wBIn1[28] , \wBMid9[25] , 
        \wAMid11[15] , \wAMid71[11] , \wBIn24[4] , \wAMid32[24] , 
        \wAMid64[25] , \wBMid68[3] , \wBIn108[13] , \wRegInA95[19] , 
        \wAMid47[14] , \wAIn93[1] , \wBIn48[13] , \wAIn115[3] , 
        \ScanLink117[4] , \wAIn41[7] , \wAIn121[28] , \wRegInB107[0] , 
        \ScanLink34[9] , \wAIn102[19] , \wAIn121[31] , \wRegInA69[2] , 
        \wRegInB104[3] , \ScanLink164[18] , \ScanLink147[30] , \wRegInA4[21] , 
        \wRegInB116[20] , \ScanLink111[28] , \ScanLink147[29] , \wBMid2[30] , 
        \wBMid2[29] , \wAIn14[26] , \wBIn27[7] , \wAIn42[4] , 
        \ScanLink132[19] , \ScanLink111[31] , \wBIn85[17] , \wRegInB2[24] , 
        \wRegInB103[14] , \wRegInB120[25] , \ScanLink109[8] , \wAIn90[2] , 
        \wBMid102[16] , \wBMid121[27] , \wAIn116[0] , \wAIn37[17] , 
        \wBIn90[23] , \wBMid117[22] , \wRegInA38[19] , \ScanLink114[7] , 
        \ScanLink0[25] , \wRegInB78[27] , \wAIn42[27] , \ScanLink56[3] , 
        \wBMid17[6] , \wAMid39[31] , \wAIn61[16] , \ScanLink208[4] , 
        \wAMid63[9] , \wAIn22[23] , \wAIn74[22] , \wAMid39[28] , \wAIn57[13] , 
        \wAMid121[7] , \wBMid70[17] , \wBIn94[8] , \wRegInB18[23] , 
        \ScanLink168[1] , \wRegInA105[30] , \wRegInA126[18] , 
        \ScanLink212[23] , \ScanLink84[5] , \ScanLink244[22] , \wAMid3[22] , 
        \wAMid3[11] , \wAIn7[15] , \wBMid26[16] , \wBMid53[26] , 
        \wRegInB76[2] , \ScanLink19[27] , \ScanLink231[12] , \ScanLink194[15] , 
        \wBMid46[12] , \wRegInA105[29] , \wRegInA6[2] , \ScanLink251[16] , 
        \wBMid33[22] , \ScanLink224[26] , \ScanLink79[23] , \ScanLink181[21] , 
        \wAIn7[26] , \wAIn7[8] , \wBMid10[13] , \wBMid65[23] , \wBIn103[6] , 
        \wAIn109[15] , \wRegInA16[7] , \wBIn58[2] , \wBIn89[7] , \wAMid94[31] , 
        \wBIn100[5] , \wRegInB75[1] , \ScanLink207[17] , \ScanLink9[3] , 
        \ScanLink216[8] , \ScanLink97[16] , \ScanLink139[15] , \ScanLink87[6] , 
        \wAMid122[4] , \wRegInA5[1] , \wRegInB9[28] , \wRegInA15[4] , 
        \ScanLink159[11] , \wRegInB9[31] , \ScanLink82[22] , \wRegInA26[21] , 
        \wRegInA53[11] , \wRegInA70[20] , \wRegInB108[18] , \wRegInB83[26] , 
        \ScanLink55[0] , \wRegInA46[25] , \wAMid94[28] , \wRegInA33[15] , 
        \wRegInB96[12] , \wRegInA65[14] , \wBMid14[5] , \wRegInA10[24] , 
        \wBMid33[11] , \wBMid46[21] , \wRegInB12[6] , \ScanLink79[10] , 
        \ScanLink224[15] , \ScanLink181[12] , \ScanLink251[25] , \wBMid10[20] , 
        \wBMid65[10] , \ScanLink207[24] , \wBIn5[23] , \wAIn14[15] , 
        \wAIn22[10] , \wBMid26[25] , \wBMid70[24] , \wAIn109[26] , 
        \wRegInA72[3] , \ScanLink212[10] , \ScanLink231[21] , 
        \ScanLink194[26] , \wBMid53[15] , \ScanLink244[11] , \ScanLink19[14] , 
        \wAIn57[20] , \wAIn74[11] , \wRegInB18[10] , \ScanLink32[7] , 
        \wBIn23[28] , \wAIn37[24] , \wAIn42[14] , \wAIn47[9] , \wBIn56[18] , 
        \wAIn88[0] , \wBIn75[30] , \wRegInB78[14] , \wAIn61[25] , 
        \wBIn116[18] , \wBIn75[29] , \wAMid19[1] , \wBIn23[31] , \wBMid73[2] , 
        \wBMid70[1] , \wRegInA10[17] , \wRegInA33[26] , \wRegInA46[16] , 
        \wRegInB96[21] , \ScanLink31[4] , \wRegInA65[27] , \wBMid109[30] , 
        \wBMid109[29] , \wRegInA70[13] , \wAMid110[18] , \wRegInA26[12] , 
        \wRegInB83[15] , \wRegInA53[22] , \wRegInB11[5] , \ScanLink159[22] , 
        \ScanLink82[11] , \wBIn21[9] , \wAIn59[5] , \wRegInA71[0] , 
        \ScanLink139[26] , \ScanLink97[25] , \wAIn80[24] , \wBIn94[31] , 
        \wAIn95[10] , \wRegInB57[0] , \wRegInB98[9] , \ScanLink112[9] , 
        \wBMid113[30] , \wRegInA29[26] , \ScanLink234[9] , \wRegInA37[5] , 
        \wBIn94[28] , \wBMid113[29] , \wBIn122[4] , \wRegInA49[22] , 
        \wRegInB99[15] , \wRegInB85[6] , \ScanLink160[13] , \wAIn8[12] , 
        \wBMid29[11] , \wBMid36[4] , \wBMid84[11] , \wRegInA108[5] , 
        \ScanLink229[6] , \ScanLink115[23] , \ScanLink98[11] , 
        \ScanLink143[22] , \ScanLink136[12] , \ScanLink77[1] , \wBMid91[25] , 
        \wAMid100[5] , \ScanLink156[16] , \ScanLink175[27] , \ScanLink149[3] , 
        \ScanLink123[26] , \wAIn113[26] , \ScanLink100[17] , \wRegInB86[5] , 
        \ScanLink74[2] , \ScanLink35[11] , \ScanLink40[21] , \ScanLink16[20] , 
        \ScanLink63[10] , \wBMid49[15] , \wBMid28[8] , \wBMid35[7] , 
        \wAMid41[8] , \wAIn125[23] , \ScanLink76[24] , \wAIn38[10] , 
        \wBIn79[0] , \wAMid103[6] , \ScanLink20[25] , \wAIn106[12] , 
        \wRegInA29[9] , \ScanLink208[10] , \ScanLink185[9] , \ScanLink55[15] , 
        \wRegInB77[20] , \wRegInA116[9] , \wBIn39[31] , \wRegInB21[21] , 
        \wRegInB54[11] , \wRegInB54[3] , \wRegInA84[26] , \wRegInB41[25] , 
        \wBIn39[28] , \wRegInB34[15] , \wRegInA91[12] , \wAIn58[14] , 
        \wBIn121[7] , \wRegInA34[6] , \wRegInB62[14] , \wBMid91[16] , 
        \wRegInB17[24] , \ScanLink198[6] , \wRegInB112[18] , \ScanLink175[14] , 
        \ScanLink156[25] , \ScanLink123[15] , \ScanLink13[5] , 
        \ScanLink100[24] , \ScanLink115[10] , \wAMid0[1] , \wAMid3[2] , 
        \wBIn5[10] , \wBMid52[0] , \ScanLink160[20] , \ScanLink98[22] , 
        \wAIn8[21] , \wBMid7[8] , \wAMid23[31] , \wAMid23[28] , \wAMid56[18] , 
        \wAIn58[27] , \wAIn80[17] , \wBMid84[22] , \wRegInA81[7] , 
        \ScanLink136[21] , \wRegInB33[4] , \wRegInA49[11] , \wRegInB99[26] , 
        \ScanLink143[11] , \wBMid80[6] , \wAIn95[23] , \wRegInA29[15] , 
        \wRegInB30[7] , \wRegInA53[1] , \ScanLink130[8] , \wRegInB34[26] , 
        \wRegInA91[21] , \wRegInB41[16] , \wAMid75[30] , \wAIn78[7] , 
        \wRegInB17[17] , \wRegInA50[2] , \wRegInB62[27] , \wRegInB77[13] , 
        \wAIn38[23] , \wAMid38[3] , \wRegInB21[12] , \wRegInA84[15] , 
        \wAMid75[29] , \wBMid83[5] , \wBMid108[1] , \wRegInB54[22] , 
        \wBMid49[26] , \ScanLink76[17] , \wAIn125[10] , \wBMid29[22] , 
        \wAIn65[8] , \wAIn106[21] , \ScanLink208[23] , \ScanLink55[26] , 
        \ScanLink20[16] , \ScanLink10[6] , \ScanLink40[12] , \wAIn113[15] , 
        \wRegInA82[4] , \ScanLink63[23] , \ScanLink35[22] , \wBMid51[3] , 
        \wRegInA113[4] , \ScanLink128[19] , \ScanLink16[13] , \ScanLink232[7] , 
        \wAMid7[30] , \wBIn11[26] , \wAMid44[5] , \wBIn61[2] , \wAMid96[3] , 
        \wRegInB119[14] , \wAMid90[10] , \wAMid101[27] , \ScanLink152[2] , 
        \wBMid118[16] , \wAMid122[16] , \wRegInB83[8] , \wBIn64[16] , 
        \wAMid85[24] , \wRegInA57[30] , \wRegInA74[18] , \wAMid114[13] , 
        \wRegInA22[19] , \wRegInA57[29] , \ScanLink180[4] , \wBIn107[27] , 
        \wBIn27[23] , \wAMid28[24] , \wBIn32[17] , \wBIn47[27] , \wAMid48[20] , 
        \wBIn124[16] , \wBIn52[13] , \wAMid105[8] , \wBMid33[9] , \wAMid47[6] , 
        \wBIn112[13] , \ScanLink183[7] , \wBIn71[22] , \wRegInA114[25] , 
        \ScanLink185[19] , \wBMid1[6] , \wBMid2[5] , \wBMid6[11] , 
        \wAMid7[29] , \wRegInA110[7] , \ScanLink231[4] , \wAIn118[19] , 
        \wAMid118[7] , \wBIn127[9] , \wRegInA122[20] , \wRegInA32[8] , 
        \ScanLink151[1] , \wBIn62[1] , \wAMid85[17] , \wAMid95[0] , 
        \wRegInB28[5] , \wRegInA101[11] , \wRegInB126[2] , \wBMid6[22] , 
        \wBIn18[9] , \wAIn60[5] , \wAMid114[20] , \wAMid101[14] , 
        \wRegInA48[0] , \wRegInA87[9] , \wRegInB92[19] , \wAMid20[1] , 
        \wAMid90[23] , \wBMid118[25] , \wBMid49[1] , \wBMid86[8] , 
        \wBMid110[3] , \wAMid122[25] , \wRegInB119[27] , \ScanLink256[3] , 
        \ScanLink136[6] , \ScanLink86[30] , \ScanLink86[29] , 
        \ScanLink240[30] , \wBMid14[18] , \wBMid37[30] , \wBMid37[29] , 
        \wBMid42[19] , \wBMid61[31] , \wRegInB36[9] , \wRegInA122[13] , 
        \ScanLink216[28] , \ScanLink240[29] , \wRegInA101[22] , 
        \ScanLink255[0] , \ScanLink235[19] , \ScanLink216[31] , \wBMid61[28] , 
        \wRegInA114[16] , \wRegInA99[5] , \wBIn27[10] , \wAMid28[17] , 
        \ScanLink135[5] , \wBIn52[20] , \ScanLink16[8] , \wBMid2[20] , 
        \wBMid2[13] , \wBIn11[15] , \wBIn71[11] , \wBIn112[20] , 
        \wRegInB125[1] , \wAMid23[2] , \wAIn26[31] , \wAIn26[28] , 
        \wBIn32[24] , \wBIn64[25] , \wAIn70[29] , \wBMid113[0] , \wBMid98[4] , 
        \wBIn107[14] , \wBIn47[14] , \wAIn53[18] , \wAIn63[6] , 
        \wRegInB69[18] , \wAMid48[13] , \wAIn70[30] , \wAIn95[6] , 
        \wBIn124[25] , \wRegInA126[22] , \ScanLink231[31] , \ScanLink212[19] , 
        \wAIn113[4] , \ScanLink111[3] , \wAMid3[18] , \wAIn4[2] , 
        \wBMid10[30] , \wBIn22[3] , \wRegInA105[13] , \ScanLink231[28] , 
        \wRegInA110[27] , \ScanLink244[18] , \wBMid10[29] , \wBMid33[18] , 
        \ScanLink79[19] , \wBMid46[28] , \wBIn15[24] , \wBIn23[21] , 
        \wAIn47[0] , \wBMid46[31] , \wBMid65[19] , \wBIn56[11] , \wAMid59[16] , 
        \wAIn88[9] , \wAIn57[30] , \wBIn60[14] , \wAIn74[18] , \wBIn75[20] , 
        \wBIn116[11] , \wRegInB101[7] , \wBIn103[25] , \wBIn15[17] , 
        \wAMid19[8] , \wAIn22[19] , \wBIn43[25] , \wAIn57[29] , \wBIn120[14] , 
        \wRegInB18[19] , \wBIn36[15] , \wAMid39[12] , \wAIn44[3] , 
        \wBMid70[8] , \wAMid81[26] , \wBMid109[20] , \wAMid110[11] , 
        \wAMid94[12] , \wAMid105[25] , \wAMid126[14] , \wRegInB96[28] , 
        \wRegInB96[31] , \wRegInB102[4] , \wBIn21[0] , \wAIn96[5] , 
        \wAIn110[7] , \wRegInA71[9] , \wAMid63[0] , \wRegInB9[12] , 
        \ScanLink112[0] , \wRegInB108[22] , \ScanLink82[18] , \wBIn60[27] , 
        \wBIn103[16] , \wAIn23[4] , \wBIn36[26] , \wAMid39[21] , \wBIn23[12] , 
        \wBIn43[16] , \wBIn94[1] , \wBIn120[27] , \ScanLink168[8] , 
        \wBIn56[22] , \wAMid59[25] , \ScanLink99[3] , \wBIn75[13] , 
        \wBIn116[22] , \wRegInA110[14] , \ScanLink181[28] , \wBIn46[7] , 
        \ScanLink181[31] , \ScanLink175[7] , \wAIn7[1] , \wAIn20[7] , 
        \wBIn45[4] , \wRegInB9[21] , \wRegInA105[20] , \wRegInA126[11] , 
        \ScanLink215[2] , \ScanLink176[4] , \ScanLink159[18] , \wRegInA5[8] , 
        \wRegInB75[8] , \wRegInB108[11] , \ScanLink216[1] , \ScanLink48[6] , 
        \wAMid60[3] , \wAMid94[21] , \wBIn97[2] , \wAMid105[16] , 
        \wAMid126[27] , \wAMid27[19] , \wAIn29[26] , \wAMid81[15] , 
        \wRegInB68[7] , \wRegInA70[29] , \wBMid109[13] , \wAMid110[22] , 
        \wRegInA26[31] , \wRegInA26[28] , \wRegInA53[18] , \wRegInA70[30] , 
        \ScanLink55[9] , \wRegInB30[17] , \wRegInB45[27] , \wRegInA95[10] , 
        \wAIn93[8] , \wRegInB66[16] , \wRegInB13[26] , \wRegInA74[4] , 
        \wRegInB73[22] , \wAIn49[22] , \wAMid52[29] , \wRegInB14[1] , 
        \wRegInB50[13] , \wRegInB25[23] , \wRegInA80[24] , \wRegInA0[5] , 
        \wBIn1[21] , \wAMid8[14] , \wBMid38[27] , \wAMid52[30] , \wAMid71[18] , 
        \wAIn121[21] , \wBMid75[5] , \ScanLink72[26] , \ScanLink24[27] , 
        \wBIn39[2] , \wAIn102[10] , \wAIn108[5] , \ScanLink51[17] , 
        \wBMid58[23] , \wAIn117[24] , \wRegInB107[9] , \ScanLink219[26] , 
        \ScanLink34[0] , \ScanLink31[13] , \ScanLink44[23] , \ScanLink12[22] , 
        \wBMid76[6] , \wBMid95[27] , \ScanLink152[14] , \ScanLink67[12] , 
        \ScanLink171[25] , \ScanLink127[24] , \ScanLink109[1] , 
        \ScanLink89[27] , \ScanLink164[11] , \ScanLink104[15] , \wAMid8[27] , 
        \wBMid11[1] , \wBMid80[13] , \wRegInA4[31] , \wRegInA4[28] , 
        \wRegInB116[29] , \ScanLink111[21] , \wRegInB116[30] , 
        \ScanLink147[20] , \ScanLink132[10] , \ScanLink37[3] , \wAIn84[26] , 
        \wAIn116[9] , \wRegInA77[7] , \wRegInA38[10] , \wAIn91[12] , 
        \wAIn117[17] , \wRegInB17[2] , \wRegInB119[5] , \wRegInA58[14] , 
        \wRegInB88[23] , \ScanLink219[15] , \ScanLink44[10] , \ScanLink67[21] , 
        \ScanLink31[20] , \wBMid38[14] , \wBMid58[10] , \ScanLink12[11] , 
        \wAIn121[12] , \ScanLink72[15] , \ScanLink51[24] , \wAIn38[5] , 
        \wAIn49[11] , \wAIn102[23] , \ScanLink24[14] , \wBIn105[1] , 
        \ScanLink50[4] , \wRegInA10[0] , \wBIn40[9] , \wRegInB73[11] , 
        \wAMid78[1] , \wRegInB25[10] , \ScanLink173[9] , \wRegInA80[17] , 
        \wBIn1[12] , \wBMid12[2] , \wAIn29[15] , \wBIn48[30] , \wRegInB50[20] , 
        \wBIn48[29] , \wBIn108[29] , \wRegInB70[5] , \wRegInA95[23] , 
        \wRegInB30[24] , \wRegInB45[14] , \wBIn108[30] , \wRegInB13[15] , 
        \wAIn84[15] , \wAIn91[21] , \wRegInA3[6] , \wRegInB66[25] , 
        \ScanLink82[2] , \wBIn106[2] , \wRegInB88[10] , \wRegInA13[3] , 
        \wRegInA38[23] , \wRegInA58[27] , \wRegInB73[6] , \ScanLink81[1] , 
        \wBIn90[19] , \wBMid117[18] , \ScanLink164[22] , \ScanLink111[12] , 
        \wAIn26[9] , \wAMid124[3] , \ScanLink132[23] , \wBIn48[1] , 
        \wAMid70[9] , \wBMid80[20] , \wBMid95[14] , \ScanLink147[13] , 
        \ScanLink171[16] , \ScanLink152[27] , \ScanLink127[17] , 
        \ScanLink53[7] , \ScanLink104[26] , \ScanLink89[14] , \wBIn87[8] , 
        \wRegInA11[27] , \wRegInA64[17] , \wRegInA18[8] , \wRegInA47[26] , 
        \wBMid108[19] , \wAMid111[28] , \wRegInA27[22] , \wRegInA32[16] , 
        \wRegInB97[11] , \wRegInA52[12] , \wRegInB82[25] , \ScanLink45[3] , 
        \wRegInA71[23] , \wBIn0[18] , \wAMid2[21] , \wAMid2[12] , \wBMid19[9] , 
        \wAMid111[31] , \ScanLink83[21] , \wBIn110[6] , \wRegInB65[2] , 
        \wRegInA127[8] , \ScanLink158[12] , \ScanLink138[16] , \ScanLink97[5] , 
        \ScanLink96[15] , \wBMid3[19] , \wAIn6[16] , \wBMid11[10] , 
        \wBMid64[20] , \wBIn113[5] , \wAIn108[16] , \wBMid47[11] , \wBIn99[4] , 
        \ScanLink206[14] , \ScanLink250[15] , \wAIn9[7] , \wBMid32[21] , 
        \ScanLink225[25] , \ScanLink180[22] , \ScanLink78[20] , \wAIn15[25] , 
        \wAIn23[20] , \wBMid27[15] , \wBMid52[25] , \wRegInB66[1] , 
        \ScanLink245[21] , \ScanLink18[24] , \ScanLink230[11] , 
        \ScanLink205[8] , \ScanLink195[16] , \wBMid71[14] , \ScanLink213[20] , 
        \ScanLink94[6] , \wAIn56[10] , \wAIn75[21] , \wRegInB19[20] , 
        \ScanLink178[2] , \wAIn15[16] , \wBIn22[18] , \wBIn57[31] , 
        \wBIn74[19] , \wBIn117[28] , \ScanLink218[7] , \wAIn60[15] , 
        \wRegInB79[24] , \wAIn36[14] , \wAIn43[24] , \wBIn117[31] , 
        \ScanLink89[9] , \wAIn49[6] , \wBIn57[28] , \wRegInA61[3] , 
        \ScanLink138[25] , \ScanLink46[0] , \wAIn54[9] , \wRegInB8[18] , 
        \wRegInB109[28] , \ScanLink96[26] , \ScanLink83[12] , \wRegInA27[11] , 
        \wRegInB109[31] , \ScanLink158[21] , \wRegInB82[16] , \wAIn60[26] , 
        \wBMid60[2] , \wRegInA52[21] , \wAMid95[18] , \wRegInA11[14] , 
        \wRegInA71[10] , \wRegInA32[25] , \wRegInA64[24] , \wRegInB97[22] , 
        \wRegInA47[15] , \ScanLink21[7] , \wAIn23[13] , \wAIn36[27] , 
        \wAIn43[17] , \wBMid63[1] , \wAIn98[3] , \wRegInB79[17] , 
        \wAMid38[18] , \wAIn56[23] , \wRegInB19[13] , \ScanLink22[4] , 
        \wBMid27[26] , \wAIn75[12] , \wRegInA104[19] , \ScanLink230[22] , 
        \ScanLink195[25] , \wBIn32[9] , \wBMid52[16] , \wRegInA127[31] , 
        \ScanLink245[12] , \ScanLink18[17] , \wRegInA62[0] , \ScanLink213[13] , 
        \wRegInA127[28] , \ScanLink101[9] , \wBMid71[27] , \wBMid11[23] , 
        \wBMid64[13] , \ScanLink206[27] , \wAIn6[25] , \wBMid32[12] , 
        \wAIn108[25] , \wBMid47[22] , \ScanLink225[16] , \ScanLink180[11] , 
        \ScanLink78[13] , \ScanLink250[26] , \wAIn36[3] , \wAMid76[7] , 
        \wBIn81[6] , \ScanLink133[29] , \wRegInA5[11] , \wRegInB117[10] , 
        \ScanLink165[31] , \ScanLink146[19] , \ScanLink133[30] , 
        \ScanLink110[18] , \ScanLink165[28] , \wBIn0[5] , \wBIn3[6] , 
        \wBMid8[26] , \wBMid8[15] , \wAMid10[25] , \wAMid26[20] , \wBIn29[27] , 
        \wBIn50[3] , \wBIn53[0] , \wBIn116[8] , \wRegInB3[14] , 
        \wRegInB102[24] , \ScanLink2[1] , \wRegInB121[15] , \wBMid120[17] , 
        \ScanLink160[0] , \wAMid53[10] , \wAMid70[21] , \wBIn84[27] , 
        \wBIn91[13] , \wBMid103[26] , \wBMid116[12] , \wRegInA39[30] , 
        \ScanLink1[15] , \wRegInA39[29] , \wRegInA121[6] , \ScanLink200[5] , 
        \ScanLink163[3] , \wAMid33[14] , \wAMid46[24] , \wBIn49[23] , 
        \wRegInA94[30] , \wRegInA122[5] , \wAMid65[15] , \ScanLink92[8] , 
        \wBIn109[23] , \wRegInA94[29] , \ScanLink203[6] , \wAIn35[0] , 
        \wAMid75[4] , \wBIn108[4] , \wBIn82[5] , \wAMid11[0] , \wAMid12[3] , 
        \wBIn37[4] , \wAIn80[1] , \wBIn91[20] , \wAIn103[30] , \wAIn103[29] , 
        \ScanLink1[2] , \wBMid116[21] , \wAIn120[18] , \ScanLink1[26] , 
        \wAIn106[3] , \wBIn84[14] , \wBMid120[24] , \ScanLink104[4] , 
        \wRegInB89[29] , \wAIn90[18] , \wBMid103[15] , \wRegInB89[30] , 
        \wBIn29[8] , \wAIn51[4] , \wAIn52[7] , \wBMid122[1] , \wRegInB102[17] , 
        \wBMid81[19] , \wRegInB3[27] , \wRegInB121[26] , \wRegInA5[22] , 
        \wRegInB114[0] , \ScanLink27[9] , \wRegInB117[23] , \wRegInA79[1] , 
        \wBMid59[29] , \wBMid121[2] , \wRegInB19[4] , \wRegInB117[3] , 
        \ScanLink66[18] , \ScanLink13[28] , \ScanLink45[30] , \ScanLink30[19] , 
        \wBIn10[1] , \wAMid10[16] , \wAMid33[27] , \wBMid59[30] , 
        \ScanLink45[29] , \ScanLink13[31] , \wBIn34[7] , \wAMid46[17] , 
        \wAIn83[2] , \wBIn49[10] , \wAIn105[0] , \ScanLink107[7] , 
        \wAMid14[27] , \wAMid26[13] , \wBIn29[14] , \wAIn48[31] , 
        \wAMid65[26] , \wBMid78[0] , \wBIn109[10] , \wRegInB24[29] , 
        \wRegInB51[19] , \wRegInB72[31] , \wAMid70[12] , \wRegInB72[28] , 
        \wBMid28[31] , \wBMid28[28] , \wAMid35[6] , \wAIn48[28] , 
        \wRegInB24[30] , \ScanLink39[5] , \wAMid53[23] , \ScanLink209[30] , 
        \ScanLink209[29] , \wBMid41[9] , \ScanLink62[29] , \wAIn75[2] , 
        \wBMid105[4] , \ScanLink34[31] , \ScanLink17[19] , \ScanLink41[18] , 
        \wAMid37[16] , \wAMid42[26] , \ScanLink62[30] , \ScanLink34[28] , 
        \wBIn38[11] , \wAMid61[17] , \ScanLink243[4] , \wAMid28[9] , 
        \wAIn39[30] , \wAMid74[23] , \wBIn118[15] , \wRegInB20[18] , 
        \wRegInB55[28] , \wAMid57[12] , \wBIn58[15] , \wRegInA40[8] , 
        \wRegInB55[31] , \wAMid22[22] , \wAIn39[29] , \wAIn121[6] , 
        \wRegInB76[19] , \ScanLink123[1] , \wBIn95[11] , \wBMid112[10] , 
        \ScanLink240[7] , \ScanLink5[17] , \ScanLink120[2] , \wAIn1[2] , 
        \wAIn2[27] , \wAIn2[14] , \wBIn4[30] , \wAIn9[18] , \wAIn11[6] , 
        \wBIn13[2] , \wAIn94[30] , \wAMid14[14] , \wAMid22[11] , \wAMid36[5] , 
        \wAIn76[1] , \wBIn80[25] , \wAIn94[29] , \wAIn122[5] , \wBMid124[15] , 
        \wBMid107[24] , \wRegInB7[16] , \wRegInB106[26] , \wRegInB125[17] , 
        \wBMid85[28] , \wRegInA1[13] , \wRegInB113[12] , \ScanLink99[31] , 
        \wAMid74[10] , \wBMid85[31] , \wBMid106[7] , \ScanLink99[28] , 
        \wBIn118[26] , \wRegInB44[9] , \wRegInA106[3] , \ScanLink227[0] , 
        \wAMid37[25] , \wAMid57[21] , \wBIn58[26] , \ScanLink79[7] , 
        \wBIn38[22] , \wAMid42[15] , \wBIn74[5] , \ScanLink147[5] , 
        \wRegInB4[9] , \wBMid38[2] , \wAMid61[24] , \wAMid83[4] , 
        \wRegInA90[18] , \wRegInB59[6] , \ScanLink64[8] , \wAMid51[2] , 
        \wAIn107[18] , \wAIn124[30] , \wRegInA39[3] , \ScanLink195[3] , 
        \wAIn124[29] , \ScanLink142[28] , \wBIn4[29] , \ScanLink161[19] , 
        \ScanLink142[31] , \ScanLink137[18] , \ScanLink114[30] , \wBIn5[8] , 
        \wAMid6[10] , \wBMid7[31] , \wAMid8[9] , \wRegInB113[21] , 
        \ScanLink114[29] , \wAIn11[27] , \wAIn12[5] , \wAMid52[1] , 
        \wRegInA1[20] , \wRegInB106[15] , \wBIn77[6] , \wBIn80[16] , 
        \wBMid107[17] , \wBMid124[26] , \wRegInB7[25] , \wRegInA105[0] , 
        \wRegInB125[24] , \ScanLink196[0] , \ScanLink159[9] , \wRegInB88[3] , 
        \wAMid80[7] , \wBIn95[22] , \ScanLink224[3] , \wBMid112[23] , 
        \wRegInA48[31] , \ScanLink5[24] , \wRegInA48[28] , \ScanLink144[6] , 
        \wAIn27[22] , \wAIn32[16] , \wAIn64[17] , \wAIn47[26] , \wAMid33[8] , 
        \wAMid49[19] , \wRegInB68[12] , \wRegInA94[0] , \wAIn52[12] , 
        \ScanLink138[0] , \wBMid47[7] , \wAIn71[23] , \ScanLink241[23] , 
        \wBMid7[28] , \wBMid23[17] , \wBMid56[27] , \wRegInB26[3] , 
        \ScanLink234[13] , \ScanLink191[14] , \ScanLink69[16] , \wAIn119[20] , 
        \wRegInA100[28] , \wBMid75[16] , \wRegInA100[31] , \wRegInA123[19] , 
        \ScanLink217[22] , \wBMid15[12] , \wBMid60[22] , \wRegInA46[6] , 
        \wAIn127[8] , \wBMid43[13] , \ScanLink202[16] , \wAMid6[23] , 
        \wBMid15[21] , \wBMid36[23] , \ScanLink254[17] , \wBMid44[4] , 
        \wAMid91[29] , \wBMid95[1] , \wBMid96[2] , \wRegInB25[0] , 
        \ScanLink221[27] , \ScanLink184[20] , \ScanLink149[24] , 
        \ScanLink246[9] , \ScanLink92[17] , \ScanLink87[23] , \wRegInA23[20] , 
        \wRegInA45[5] , \wRegInA56[10] , \ScanLink129[20] , \wRegInA75[21] , 
        \wRegInB86[27] , \wBMid100[9] , \wRegInA60[15] , \wAMid91[30] , 
        \wRegInA15[25] , \wRegInA36[14] , \wRegInA43[24] , \wRegInA97[3] , 
        \wRegInB93[13] , \wBMid60[11] , \ScanLink202[25] , \wBMid36[10] , 
        \wRegInB42[7] , \wBMid43[20] , \ScanLink221[14] , \ScanLink184[13] , 
        \wAMid3[26] , \wAMid3[15] , \wAIn11[14] , \wBMid23[24] , \wRegInB2[7] , 
        \ScanLink254[24] , \ScanLink234[20] , \ScanLink191[27] , 
        \ScanLink69[25] , \wBMid23[3] , \wBIn26[30] , \wAIn27[11] , 
        \wAIn52[21] , \wBMid56[14] , \ScanLink241[10] , \wBMid75[25] , 
        \wAIn119[13] , \wRegInA22[2] , \ScanLink217[11] , \ScanLink62[6] , 
        \wAIn64[24] , \wAIn71[10] , \wRegInB68[21] , \wAMid98[5] , 
        \wRegInB90[1] , \wBIn113[19] , \wBIn70[28] , \wBMid14[1] , \wAIn17[8] , 
        \wBMid20[0] , \wBIn26[29] , \wAIn32[25] , \wAIn47[15] , \wBIn53[19] , 
        \wAMid115[2] , \wBIn70[31] , \wAMid115[19] , \wRegInA15[16] , 
        \wRegInB93[2] , \wRegInA23[13] , \wRegInA36[27] , \wRegInA60[26] , 
        \wRegInB93[20] , \wRegInA43[17] , \ScanLink61[5] , \wRegInB86[14] , 
        \wAMid116[1] , \wRegInA56[23] , \wRegInA75[12] , \wAMid49[0] , 
        \wBIn71[8] , \wRegInA21[1] , \wRegInB41[4] , \ScanLink129[13] , 
        \ScanLink87[10] , \ScanLink149[17] , \ScanLink142[8] , \wAMid86[9] , 
        \wRegInB1[4] , \wRegInA65[10] , \ScanLink92[24] , \wBIn45[9] , 
        \wBIn58[6] , \wAMid122[0] , \wRegInA10[20] , \wRegInA46[21] , 
        \wAMid81[18] , \wRegInA26[25] , \wRegInA33[11] , \wRegInA53[15] , 
        \wRegInB96[16] , \wRegInB83[22] , \wRegInA70[24] , \ScanLink55[4] , 
        \wBIn100[1] , \wRegInA5[5] , \ScanLink82[26] , \wRegInA15[0] , 
        \ScanLink159[15] , \ScanLink176[9] , \wBIn103[2] , \wRegInB75[5] , 
        \ScanLink139[11] , \ScanLink87[2] , \ScanLink97[12] , \ScanLink9[7] , 
        \wAIn7[11] , \wBMid10[17] , \wBMid65[27] , \wRegInA16[3] , 
        \wAIn109[11] , \wBMid46[16] , \wBIn89[3] , \ScanLink207[13] , 
        \wRegInA6[6] , \wBMid10[24] , \wAIn14[22] , \wBMid17[2] , \wAIn22[27] , 
        \wBMid26[12] , \wBMid33[26] , \wRegInA110[19] , \ScanLink251[12] , 
        \ScanLink79[27] , \wBMid53[22] , \ScanLink244[26] , \ScanLink224[22] , 
        \ScanLink181[25] , \wRegInB76[6] , \ScanLink231[16] , 
        \ScanLink194[11] , \ScanLink19[23] , \wBMid70[13] , \ScanLink212[27] , 
        \ScanLink84[1] , \wAIn23[9] , \wAMid121[3] , \wAIn57[17] , 
        \wAIn74[26] , \wRegInB18[27] , \ScanLink168[5] , \wAIn14[11] , 
        \wAMid19[5] , \wAIn37[13] , \wAMid59[31] , \wAIn61[12] , 
        \ScanLink208[0] , \wRegInB78[23] , \wAIn42[23] , \wAIn59[1] , 
        \wAMid59[28] , \wAIn96[8] , \wRegInA71[4] , \ScanLink56[7] , 
        \ScanLink139[22] , \wAIn61[21] , \wBMid70[5] , \wRegInB11[1] , 
        \ScanLink97[21] , \wRegInA26[16] , \wRegInB83[11] , \ScanLink159[26] , 
        \ScanLink82[15] , \wRegInA53[26] , \wRegInA70[17] , \wAMid105[31] , 
        \wAMid126[19] , \wAMid105[28] , \wRegInA10[13] , \wRegInB102[9] , 
        \wRegInA65[23] , \wRegInA33[22] , \wRegInA46[12] , \wRegInB96[25] , 
        \ScanLink31[0] , \wBMid73[6] , \wBIn15[30] , \wAIn22[14] , 
        \wBIn36[18] , \wAIn37[20] , \wAIn42[10] , \wAIn88[4] , \wRegInB78[10] , 
        \wBIn43[28] , \wAIn57[24] , \wBIn103[31] , \wBIn120[19] , 
        \wRegInB18[14] , \ScanLink32[3] , \wBIn15[29] , \wBIn43[31] , 
        \wBIn60[19] , \wAIn74[15] , \wBIn103[28] , \wBMid26[21] , 
        \ScanLink231[25] , \ScanLink194[22] , \wBMid53[11] , \ScanLink244[15] , 
        \wBMid70[20] , \wAIn113[9] , \wRegInA72[7] , \ScanLink212[14] , 
        \ScanLink19[10] , \wBMid65[14] , \ScanLink207[20] , \wAIn7[22] , 
        \wBMid33[15] , \wAIn109[22] , \wRegInB12[2] , \ScanLink79[14] , 
        \wBMid46[25] , \ScanLink224[11] , \ScanLink181[16] , \wAIn26[4] , 
        \ScanLink251[21] , \wAMid66[0] , \wBIn91[1] , \wRegInA4[16] , 
        \wRegInB116[17] , \wBIn43[7] , \wBMid95[19] , \wRegInB2[13] , 
        \wRegInB103[23] , \ScanLink89[19] , \wRegInB120[12] , \ScanLink170[7] , 
        \wAIn84[18] , \wBIn85[20] , \wBMid121[10] , \wBIn90[14] , 
        \wBMid102[21] , \wBMid117[15] , \ScanLink0[12] , \ScanLink210[2] , 
        \wRegInA0[8] , \wAMid71[26] , \wAIn2[1] , \wAMid11[22] , \wAMid27[27] , 
        \wAIn38[8] , \wAMid52[17] , \wBIn40[4] , \ScanLink173[4] , 
        \wBIn28[20] , \wAIn29[18] , \wAMid32[13] , \wAMid47[23] , \wBIn48[24] , 
        \wRegInB13[18] , \wRegInB30[30] , \wAMid64[12] , \wRegInB66[28] , 
        \wBIn108[24] , \wRegInB30[29] , \wRegInB70[8] , \ScanLink213[1] , 
        \wAMid65[3] , \wRegInB45[19] , \wRegInB66[31] , \wAMid8[19] , 
        \wBMid9[12] , \wAIn25[7] , \wBIn118[3] , \ScanLink219[18] , 
        \wBIn92[2] , \wBIn27[3] , \wBMid38[19] , \ScanLink51[29] , 
        \ScanLink50[9] , \ScanLink24[19] , \wAIn90[6] , \wBIn90[27] , 
        \wBMid117[26] , \ScanLink72[18] , \ScanLink51[30] , \ScanLink0[21] , 
        \wAIn116[4] , \wAIn42[0] , \wBIn85[13] , \wBMid121[23] , 
        \wRegInA58[19] , \ScanLink114[3] , \wBMid102[12] , \wRegInB103[10] , 
        \wRegInB119[8] , \ScanLink171[28] , \ScanLink127[30] , 
        \ScanLink104[18] , \ScanLink171[31] , \wRegInB2[20] , 
        \ScanLink152[19] , \wRegInA4[25] , \wRegInB104[7] , \wRegInB120[21] , 
        \ScanLink127[29] , \wRegInB116[24] , \wBMid9[21] , \wAIn41[3] , 
        \wBMid75[8] , \wAIn108[8] , \wRegInA69[6] , \wAIn117[30] , 
        \wAIn117[29] , \wRegInB107[4] , \wAMid11[11] , \wBIn24[0] , 
        \wAMid32[20] , \wAMid47[10] , \wBIn48[17] , \wAIn93[5] , 
        \wRegInA74[9] , \wAIn115[7] , \ScanLink117[0] , \wAMid64[21] , 
        \wBMid68[7] , \wBIn108[17] , \wRegInA80[29] , \wBIn0[8] , 
        \wRegInA0[27] , \wRegInA0[14] , \wBMid4[6] , \wBMid7[5] , 
        \wAMid27[14] , \wAMid71[15] , \wBIn28[13] , \wAMid52[24] , 
        \wRegInA80[30] , \ScanLink29[2] , \wAMid15[20] , \wAMid25[1] , 
        \wRegInB123[2] , \wAMid36[11] , \wBIn39[16] , \wAMid43[21] , 
        \wAIn65[5] , \wBMid115[3] , \wRegInA82[9] , \wAIn113[18] , 
        \wAMid60[10] , \ScanLink253[3] , \wAMid23[25] , \wAMid56[15] , 
        \wAMid75[24] , \wBIn119[12] , \wRegInA84[18] , \wBMid83[8] , 
        \wBIn59[12] , \ScanLink133[6] , \wBIn81[22] , \wBIn94[16] , 
        \wRegInB33[9] , \ScanLink4[10] , \wBMid106[23] , \wBMid113[17] , 
        \wBMid125[12] , \wRegInA29[18] , \ScanLink250[0] , \ScanLink130[5] , 
        \wRegInB107[21] , \wRegInB120[1] , \ScanLink100[29] , \wAIn66[6] , 
        \wRegInB6[11] , \ScanLink175[19] , \ScanLink156[31] , \wRegInB124[10] , 
        \ScanLink123[18] , \ScanLink100[30] , \ScanLink156[28] , 
        \ScanLink13[8] , \wRegInB112[15] , \wAMid6[2] , \wAMid26[2] , 
        \wBMid116[0] , \wAMid15[13] , \wAMid23[16] , \wAMid75[17] , 
        \wBIn119[21] , \wRegInA116[4] , \ScanLink237[7] , \wAMid36[22] , 
        \wBIn39[25] , \wAMid56[26] , \ScanLink69[0] , \wBIn59[21] , 
        \wAMid43[12] , \wRegInB41[31] , \wRegInB62[19] , \wAIn58[19] , 
        \ScanLink157[2] , \wBIn64[2] , \wRegInB17[29] , \wBMid28[5] , 
        \wAMid60[23] , \wAMid93[3] , \wRegInB41[28] , \wRegInB17[30] , 
        \wAMid41[5] , \wBMid49[18] , \wRegInA29[4] , \wRegInB34[18] , 
        \wRegInB49[1] , \wRegInB86[8] , \ScanLink20[28] , \ScanLink185[4] , 
        \ScanLink76[30] , \ScanLink55[18] , \wRegInB9[1] , \ScanLink20[31] , 
        \wRegInA108[8] , \ScanLink76[29] , \wRegInB112[26] , \wAIn3[20] , 
        \wAIn3[13] , \wAMid5[1] , \wBMid36[9] , \wAMid42[6] , \wBIn81[11] , 
        \wBMid91[31] , \wBMid91[28] , \wAMid100[8] , \wRegInB107[12] , 
        \wBMid106[10] , \wBMid125[21] , \wRegInB6[22] , \wRegInA115[7] , 
        \wRegInB124[23] , \ScanLink186[7] , \wRegInB98[4] , \ScanLink234[4] , 
        \wAMid7[17] , \wBIn8[0] , \wAIn10[20] , \wBIn67[1] , \wAIn80[30] , 
        \wAIn80[29] , \wAMid90[0] , \wBIn94[25] , \ScanLink4[23] , 
        \wBMid113[24] , \wBIn122[9] , \wRegInA37[8] , \wRegInB99[18] , 
        \ScanLink154[1] , \wAIn26[25] , \wAIn33[11] , \wAIn65[10] , 
        \ScanLink248[2] , \wAIn46[21] , \ScanLink16[5] , \wBIn32[29] , 
        \wBIn47[19] , \wRegInB69[15] , \wRegInA84[7] , \wAIn53[15] , 
        \wBIn64[31] , \wBIn124[28] , \ScanLink128[7] , \wBIn11[18] , 
        \wBMid22[10] , \wBIn32[30] , \wBMid57[20] , \wBMid57[0] , \wBIn64[28] , 
        \wAIn70[24] , \wBMid98[9] , \wBIn107[19] , \wBIn124[31] , 
        \wRegInB36[4] , \ScanLink240[24] , \ScanLink235[14] , 
        \ScanLink190[13] , \wBMid74[11] , \wAIn118[27] , \ScanLink68[11] , 
        \ScanLink216[25] , \wBMid14[15] , \wBMid61[25] , \wRegInA56[1] , 
        \wRegInA99[8] , \wBMid42[14] , \ScanLink203[11] , \ScanLink135[8] , 
        \ScanLink255[10] , \wBMid2[8] , \wBMid37[24] , \wBMid85[6] , 
        \wBMid86[5] , \wRegInB35[7] , \ScanLink220[20] , \ScanLink185[27] , 
        \ScanLink148[23] , \ScanLink93[10] , \ScanLink86[24] , \wRegInA22[27] , 
        \wRegInA55[2] , \wRegInA57[17] , \ScanLink128[27] , \wRegInB87[20] , 
        \wRegInB28[8] , \wRegInA74[26] , \ScanLink15[6] , \wAMid7[24] , 
        \wBMid14[26] , \wBIn18[4] , \wBMid54[3] , \wBMid118[28] , 
        \wAMid122[28] , \wRegInA61[12] , \wRegInA14[22] , \wAIn60[8] , 
        \wBMid118[31] , \wRegInA87[4] , \wAMid101[19] , \wRegInA42[23] , 
        \wAMid122[31] , \wRegInA37[13] , \wRegInB92[14] , \wRegInA114[31] , 
        \wBMid61[16] , \ScanLink203[22] , \wBMid37[17] , \wBMid42[27] , 
        \wRegInB52[0] , \wRegInA114[28] , \ScanLink220[13] , \ScanLink185[14] , 
        \ScanLink255[23] , \wBIn4[24] , \wAIn10[13] , \wBMid22[23] , 
        \ScanLink235[27] , \ScanLink231[9] , \ScanLink190[20] , \wAIn26[16] , 
        \wAIn53[26] , \wBMid57[13] , \ScanLink240[17] , \ScanLink68[22] , 
        \wBMid74[22] , \wAIn118[14] , \wBIn127[4] , \wRegInA32[5] , 
        \ScanLink216[16] , \ScanLink72[1] , \wAMid28[30] , \wAIn65[23] , 
        \wAIn70[17] , \wRegInB69[26] , \wAMid88[2] , \wRegInB80[6] , 
        \wAIn19[3] , \wAMid28[29] , \wAIn33[22] , \wBMid33[4] , \wAIn46[12] , 
        \wAMid105[5] , \wBMid30[7] , \wAMid44[8] , \wAMid85[30] , 
        \wAMid106[6] , \wRegInA14[11] , \wRegInB83[5] , \wRegInA22[14] , 
        \wRegInA37[20] , \wRegInA61[21] , \wRegInA42[10] , \wRegInB92[27] , 
        \ScanLink71[2] , \wRegInB87[13] , \wRegInA57[24] , \ScanLink180[9] , 
        \wAMid85[29] , \wRegInA74[15] , \wBIn124[7] , \wRegInA31[6] , 
        \wRegInB51[3] , \wRegInA113[9] , \ScanLink128[14] , \ScanLink86[17] , 
        \wAMid59[7] , \ScanLink148[10] , \wAIn81[23] , \wAIn94[17] , 
        \wRegInB47[7] , \wRegInB119[19] , \ScanLink93[23] , \wRegInA27[2] , 
        \wRegInA28[21] , \ScanLink5[30] , \wRegInA48[25] , \wRegInB98[12] , 
        \ScanLink5[29] , \wRegInB7[7] , \wRegInB95[1] , \ScanLink161[14] , 
        \wBIn4[17] , \wAMid8[4] , \ScanLink239[1] , \ScanLink99[16] , 
        \ScanLink114[24] , \wAIn9[15] , \wAIn12[8] , \wBMid85[16] , 
        \wRegInA118[2] , \ScanLink142[25] , \ScanLink137[15] , \ScanLink67[6] , 
        \wBMid26[3] , \wBMid90[22] , \wAMid110[2] , \ScanLink157[11] , 
        \wRegInB7[28] , \wRegInB7[31] , \wRegInB125[29] , \ScanLink174[20] , 
        \ScanLink159[4] , \ScanLink122[21] , \wBMid28[16] , \wAIn112[21] , 
        \wRegInB106[18] , \ScanLink101[10] , \wRegInB125[30] , \wRegInB96[2] , 
        \ScanLink64[5] , \ScanLink34[16] , \ScanLink41[26] , \ScanLink17[27] , 
        \wBMid48[12] , \ScanLink62[17] , \wAMid14[19] , \wBMid25[0] , 
        \wAIn124[24] , \ScanLink77[23] , \wAMid37[31] , \wAIn39[17] , 
        \wBIn69[7] , \wAIn107[15] , \wAMid113[1] , \ScanLink21[22] , 
        \ScanLink209[17] , \ScanLink54[12] , \wRegInB76[27] , \wRegInB20[26] , 
        \wRegInB44[4] , \wRegInB55[16] , \wRegInA85[21] , \wAMid83[9] , 
        \wRegInB4[4] , \wAMid36[8] , \wAMid37[28] , \wAMid61[29] , 
        \wRegInB40[22] , \wRegInB35[12] , \wRegInA90[15] , \wAMid42[18] , 
        \wAIn59[13] , \wRegInA24[1] , \wRegInB63[13] , \wAMid61[30] , 
        \ScanLink147[8] , \wBIn74[8] , \wBMid90[11] , \wRegInB16[23] , 
        \ScanLink188[1] , \ScanLink174[13] , \ScanLink157[22] , 
        \ScanLink122[12] , \ScanLink101[23] , \ScanLink114[17] , \wBMid42[7] , 
        \ScanLink161[27] , \ScanLink99[25] , \wBMid9[3] , \wBMid85[25] , 
        \wRegInA91[0] , \ScanLink137[26] , \wRegInB23[3] , \wRegInA48[16] , 
        \wRegInB98[21] , \ScanLink142[16] , \wBIn80[28] , \wAIn81[10] , 
        \wBMid90[1] , \wAIn94[24] , \wBMid107[29] , \wRegInA28[12] , 
        \wRegInA43[6] , \wAIn2[19] , \wBIn6[6] , \wBMid7[16] , \wAIn9[26] , 
        \wAMid28[4] , \wAIn39[24] , \wBIn58[18] , \wAIn59[20] , \wBIn80[31] , 
        \wBMid107[30] , \wAIn122[8] , \wBMid124[18] , \wRegInB20[0] , 
        \wRegInB35[21] , \wRegInB40[11] , \wRegInA90[26] , \ScanLink243[9] , 
        \wAIn68[0] , \wRegInB16[10] , \wRegInA40[5] , \wRegInB63[20] , 
        \wRegInB76[14] , \wBIn118[18] , \wRegInA85[12] , \wRegInB20[15] , 
        \wBMid48[21] , \wBMid93[2] , \wBMid118[6] , \wRegInB55[25] , 
        \ScanLink77[10] , \wAIn124[17] , \wBIn10[21] , \wAIn14[6] , 
        \wBMid28[25] , \wAIn107[26] , \ScanLink209[24] , \ScanLink54[21] , 
        \ScanLink21[11] , \wAIn112[12] , \wRegInA92[3] , \ScanLink41[15] , 
        \ScanLink34[25] , \wBMid41[4] , \wBMid105[9] , \ScanLink62[24] , 
        \wAMid54[2] , \wBIn71[5] , \wAMid86[4] , \wRegInB1[9] , \wRegInB41[9] , 
        \wRegInA103[3] , \ScanLink17[14] , \wRegInB118[13] , \ScanLink222[0] , 
        \ScanLink92[29] , \wAMid91[17] , \wAMid100[20] , \ScanLink142[5] , 
        \ScanLink92[30] , \wAMid123[11] , \ScanLink61[8] , \wBMid119[11] , 
        \wAMid84[23] , \wAMid115[14] , \wRegInB86[19] , \wBIn65[11] , 
        \ScanLink190[3] , \wBIn106[20] , \wAIn11[19] , \wAIn17[5] , 
        \wBIn33[10] , \wBIn46[20] , \wAMid49[27] , \wBIn125[11] , \wBIn26[24] , 
        \wAIn47[18] , \wBIn53[14] , \wAIn64[30] , \wAMid29[23] , \wAIn32[28] , 
        \wAMid57[1] , \wBIn70[25] , \wAMid98[8] , \wBIn113[14] , 
        \ScanLink193[0] , \wAIn64[29] , \wBMid23[30] , \wAIn32[31] , 
        \wAMid108[0] , \wRegInA100[0] , \wRegInA115[22] , \ScanLink254[29] , 
        \ScanLink221[19] , \ScanLink221[3] , \ScanLink202[31] , 
        \ScanLink254[30] , \ScanLink202[28] , \ScanLink69[31] , 
        \wRegInA123[27] , \ScanLink141[6] , \wBMid23[29] , \wBIn72[6] , 
        \wBMid75[28] , \wAMid85[7] , \ScanLink69[28] , \wAMid30[6] , 
        \wBMid56[19] , \wBMid75[31] , \wRegInA100[16] , \wAIn70[2] , 
        \wAMid84[10] , \wRegInB38[2] , \wAMid115[27] , \wAMid91[24] , 
        \wAMid100[13] , \wRegInA43[29] , \wRegInA58[7] , \wRegInA15[31] , 
        \wRegInA36[19] , \wBMid119[22] , \wRegInA60[18] , \wBMid44[9] , 
        \wAMid123[22] , \wRegInA43[30] , \wBMid100[4] , \wRegInA15[28] , 
        \wRegInA45[8] , \wRegInB118[20] , \ScanLink149[30] , \ScanLink246[4] , 
        \ScanLink149[29] , \ScanLink18[3] , \ScanLink126[1] , \wBMid7[25] , 
        \wBIn15[1] , \wBMid59[6] , \wAIn124[6] , \wRegInA100[25] , 
        \wRegInA123[14] , \ScanLink245[7] , \ScanLink191[19] , \wBMid3[27] , 
        \wBMid3[14] , \wBIn5[5] , \wBIn16[2] , \wRegInA89[2] , 
        \wRegInA115[11] , \wAIn127[5] , \ScanLink125[2] , \wBIn10[12] , 
        \wBIn26[17] , \wAMid29[10] , \wAMid33[5] , \wBIn53[27] , \wBIn70[16] , 
        \wBIn113[27] , \wBIn33[23] , \wBIn65[22] , \wBMid88[3] , \wBMid103[7] , 
        \wBIn106[13] , \wBIn46[13] , \wAMid49[14] , \wAIn73[1] , \wAIn85[1] , 
        \wBIn125[22] , \wRegInA127[25] , \ScanLink195[31] , \ScanLink101[4] , 
        \wAIn6[31] , \wAIn6[28] , \wBIn32[4] , \wAIn103[3] , \wAIn108[31] , 
        \wRegInA104[14] , \ScanLink195[28] , \wRegInA111[20] , \wAIn108[28] , 
        \wBIn14[23] , \wAMid17[3] , \wBIn22[26] , \wAIn57[7] , \wBIn57[16] , 
        \wAMid58[11] , \wBIn117[16] , \wBIn61[13] , \wBIn74[27] , 
        \wRegInB111[0] , \wBIn102[22] , \wBIn14[10] , \wAMid14[0] , 
        \wBIn37[12] , \wAMid38[15] , \wBIn42[22] , \wBIn121[13] , 
        \ScanLink22[9] , \wBIn31[7] , \wAIn54[4] , \wAMid80[21] , 
        \wBMid108[27] , \wBMid124[2] , \wAMid111[16] , \wAIn86[2] , 
        \wAMid95[15] , \wAMid104[22] , \wRegInA11[19] , \wRegInA32[28] , 
        \wRegInA47[18] , \wRegInA64[30] , \wRegInA32[31] , \wRegInB112[3] , 
        \wRegInA64[29] , \ScanLink138[31] , \ScanLink138[28] , \wAIn100[0] , 
        \wRegInB8[15] , \ScanLink102[7] , \wRegInB109[25] , \wAIn15[31] , 
        \wAIn33[3] , \wBIn37[21] , \wAMid38[26] , \wBIn61[20] , \wAMid73[7] , 
        \wBIn102[11] , \wAIn36[19] , \wBIn42[11] , \wBIn84[6] , \wBIn121[20] , 
        \wRegInB79[29] , \wAIn15[28] , \wBIn22[15] , \wAIn43[29] , 
        \wBIn57[25] , \ScanLink89[4] , \wAMid58[22] , \wRegInB79[30] , 
        \wAIn43[30] , \wAIn60[18] , \wBIn117[25] , \ScanLink7[1] , 
        \wBMid52[31] , \wBIn56[0] , \wBIn74[14] , \wBIn113[8] , 
        \wRegInA111[13] , \ScanLink250[18] , \ScanLink225[28] , \wBIn99[9] , 
        \ScanLink206[19] , \ScanLink165[0] , \ScanLink225[31] , 
        \ScanLink18[30] , \wBMid71[19] , \wBMid19[4] , \wBMid27[18] , 
        \wBMid52[28] , \wRegInA124[6] , \wRegInA127[16] , \ScanLink18[29] , 
        \wRegInA104[27] , \ScanLink205[5] , \wBIn55[3] , \wRegInB8[26] , 
        \ScanLink166[3] , \wRegInB109[16] , \wAIn30[0] , \wRegInA127[5] , 
        \ScanLink206[6] , \ScanLink96[18] , \ScanLink97[8] , \ScanLink58[1] , 
        \wAMid70[4] , \wBIn87[5] , \wRegInA18[5] , \wAMid95[26] , 
        \wAMid104[11] , \wRegInA8[0] , \wBMid108[14] , \wRegInB78[0] , 
        \ScanLink4[2] , \wBIn0[26] , \wAMid9[13] , \wAIn28[21] , \wAMid80[12] , 
        \wAMid111[25] , \wRegInB82[31] , \wRegInB82[28] , \wRegInB31[10] , 
        \wRegInB44[20] , \wRegInA94[17] , \wBIn29[19] , \wRegInB12[21] , 
        \wRegInA64[3] , \wRegInB67[11] , \wRegInB72[25] , \wBMid39[20] , 
        \wAIn48[25] , \ScanLink39[8] , \wAIn120[26] , \wRegInB24[24] , 
        \wRegInB51[14] , \wRegInA81[23] , \ScanLink73[21] , \wAIn51[9] , 
        \wBMid65[2] , \ScanLink25[20] , \wBIn29[5] , \wAIn103[17] , 
        \wAIn118[2] , \ScanLink50[10] , \wBMid59[24] , \wAIn116[23] , 
        \wRegInB19[9] , \ScanLink218[21] , \ScanLink30[14] , \ScanLink24[7] , 
        \ScanLink45[24] , \wBMid66[1] , \wBMid94[20] , \ScanLink153[13] , 
        \ScanLink66[15] , \ScanLink13[25] , \ScanLink170[22] , 
        \ScanLink126[23] , \ScanLink119[6] , \ScanLink88[20] , 
        \ScanLink165[16] , \ScanLink105[12] , \wBIn0[15] , \wBMid8[18] , 
        \wBIn37[9] , \wBMid81[14] , \ScanLink146[27] , \ScanLink110[26] , 
        \ScanLink133[17] , \ScanLink27[4] , \wRegInA67[0] , \wBIn84[19] , 
        \wAIn85[21] , \wRegInA39[17] , \ScanLink104[9] , \wAIn90[15] , 
        \wBMid120[30] , \wBMid103[18] , \wRegInB109[2] , \wBIn108[9] , 
        \wBMid120[29] , \wRegInA59[13] , \wRegInB89[24] , \ScanLink218[12] , 
        \wAIn116[10] , \ScanLink45[17] , \ScanLink30[27] , \wAMid9[20] , 
        \wBMid39[13] , \wBMid59[17] , \wAMid75[9] , \wBIn82[8] , 
        \ScanLink66[26] , \ScanLink73[12] , \ScanLink13[16] , \wAIn120[15] , 
        \ScanLink50[23] , \wAMid10[31] , \wAMid10[28] , \wAIn28[2] , 
        \wAIn48[16] , \wAIn103[24] , \ScanLink40[3] , \ScanLink25[13] , 
        \wBIn115[6] , \wAMid46[30] , \wAMid68[6] , \wRegInB24[17] , 
        \wRegInB72[16] , \wRegInA81[10] , \wRegInB51[27] , \wAMid65[18] , 
        \wRegInB31[23] , \wRegInB60[2] , \wRegInA94[24] , \wAMid46[29] , 
        \wRegInB44[13] , \wRegInB12[12] , \wRegInA122[8] , \wAIn28[12] , 
        \wAMid33[19] , \ScanLink92[5] , \wAIn85[12] , \wAIn90[26] , 
        \wRegInB67[22] , \wBIn116[5] , \wRegInB89[17] , \wRegInA39[24] , 
        \wRegInA59[20] , \wRegInB63[1] , \ScanLink91[6] , \ScanLink200[8] , 
        \ScanLink1[18] , \ScanLink165[25] , \ScanLink110[15] , \wBIn0[1] , 
        \wAIn2[23] , \wAIn2[10] , \wBIn15[8] , \wBMid44[0] , \wBMid81[27] , 
        \ScanLink133[24] , \wBMid94[13] , \ScanLink146[14] , \wRegInB3[19] , 
        \wRegInA15[21] , \wRegInA36[10] , \wRegInA43[20] , \wRegInA97[7] , 
        \wRegInB102[30] , \wRegInB121[18] , \ScanLink126[10] , 
        \wRegInB102[29] , \ScanLink153[20] , \ScanLink43[0] , 
        \ScanLink170[11] , \ScanLink105[21] , \ScanLink88[13] , 
        \wRegInB93[17] , \wRegInA60[11] , \wAMid84[19] , \wRegInA75[25] , 
        \wRegInA23[24] , \wRegInA56[14] , \wRegInA45[1] , \wRegInB86[23] , 
        \ScanLink129[24] , \ScanLink126[8] , \wBMid43[17] , \wBMid96[6] , 
        \ScanLink87[27] , \wRegInB25[4] , \wRegInB118[30] , \wRegInB118[29] , 
        \ScanLink92[13] , \ScanLink149[20] , \ScanLink254[13] , \wAMid6[14] , 
        \wBMid36[27] , \wRegInA115[18] , \wBMid95[5] , \ScanLink221[23] , 
        \ScanLink184[24] , \wBIn10[31] , \wBIn10[28] , \wAIn11[23] , 
        \wBMid15[16] , \wBMid60[26] , \wRegInA46[2] , \wBMid23[13] , 
        \wBMid56[23] , \wBMid75[12] , \wAIn119[24] , \ScanLink202[12] , 
        \wRegInB26[7] , \ScanLink241[27] , \ScanLink217[26] , 
        \ScanLink234[17] , \ScanLink191[10] , \wAIn27[26] , \wBMid47[3] , 
        \ScanLink69[12] , \wAIn71[27] , \wAMid29[19] , \wAIn52[16] , 
        \wAIn73[8] , \wRegInB68[16] , \wRegInA94[4] , \ScanLink138[4] , 
        \wAIn32[12] , \wAIn47[22] , \wAIn11[10] , \wBMid20[4] , \wAMid49[4] , 
        \wAIn64[13] , \wRegInB1[0] , \wRegInA21[5] , \ScanLink92[20] , 
        \wRegInB41[0] , \ScanLink149[13] , \ScanLink129[17] , \ScanLink222[9] , 
        \ScanLink87[14] , \wAIn32[21] , \wAIn47[11] , \wAMid100[30] , 
        \wAMid100[29] , \wAMid116[5] , \wRegInA23[17] , \wRegInA75[16] , 
        \wRegInB86[10] , \wRegInA56[27] , \wAMid123[18] , \wRegInA36[23] , 
        \wRegInB93[24] , \wRegInA43[13] , \ScanLink61[1] , \wRegInB93[6] , 
        \wAMid115[6] , \wBMid119[18] , \wRegInA15[12] , \wRegInA60[22] , 
        \ScanLink193[9] , \wAMid57[8] , \wAIn64[20] , \wAMid98[1] , 
        \wBMid23[7] , \wBIn46[30] , \wBIn65[18] , \wAIn71[14] , \wBIn106[29] , 
        \wRegInB90[5] , \wBIn33[19] , \wBIn46[29] , \wAIn52[25] , 
        \wBIn106[30] , \wBIn125[18] , \ScanLink62[2] , \wBMid23[20] , 
        \wAIn27[15] , \wBMid75[21] , \wAMid108[9] , \wRegInB68[25] , 
        \wAIn119[17] , \wRegInA22[6] , \ScanLink217[15] , \wRegInB2[3] , 
        \ScanLink234[24] , \ScanLink191[23] , \wBMid36[14] , \wBMid56[10] , 
        \ScanLink241[14] , \ScanLink69[21] , \wBMid43[24] , \wRegInB42[3] , 
        \ScanLink221[10] , \ScanLink184[17] , \ScanLink254[20] , \wAMid6[27] , 
        \wBMid15[25] , \wRegInA100[9] , \wBMid60[15] , \ScanLink202[21] , 
        \wAMid36[1] , \wRegInA1[17] , \wRegInB113[16] , \wAIn76[5] , 
        \wBMid106[3] , \wBIn80[21] , \wBMid90[18] , \wRegInA91[9] , 
        \wBMid90[8] , \wRegInB7[12] , \wRegInB106[22] , \wRegInB125[13] , 
        \wBMid107[20] , \ScanLink120[6] , \wRegInA0[1] , \wBIn1[25] , 
        \wAMid2[25] , \wAMid2[16] , \wBIn3[2] , \wBIn10[5] , \wBIn13[6] , 
        \wBMid124[11] , \wAMid57[16] , \wAIn81[19] , \wBIn95[15] , 
        \wAIn122[1] , \wRegInB98[31] , \wRegInB98[28] , \ScanLink5[13] , 
        \wBMid112[14] , \ScanLink240[3] , \wBIn58[11] , \wAIn68[9] , 
        \wAIn121[2] , \ScanLink123[5] , \wAIn6[12] , \wBMid8[22] , 
        \wBMid8[11] , \wAMid9[30] , \wAIn11[2] , \wAIn12[1] , \wAMid14[23] , 
        \wAMid22[26] , \wAIn59[30] , \wAMid61[13] , \wAMid74[27] , 
        \wBIn118[11] , \wRegInB20[9] , \wRegInB35[28] , \ScanLink243[0] , 
        \wAMid35[2] , \wAMid37[12] , \wBIn38[15] , \wAMid42[22] , \wAIn59[29] , 
        \wRegInB40[18] , \wRegInB63[30] , \wRegInB16[19] , \wRegInB35[31] , 
        \wAIn75[6] , \wRegInB63[29] , \wBMid48[31] , \wBMid48[28] , 
        \wBMid105[0] , \ScanLink77[19] , \ScanLink54[31] , \ScanLink54[28] , 
        \ScanLink21[18] , \wBIn77[2] , \wBIn80[12] , \wAMid80[3] , 
        \wBIn95[26] , \ScanLink144[2] , \ScanLink5[20] , \wBMid112[27] , 
        \wBMid107[13] , \wRegInB88[7] , \wBMid124[22] , \wRegInA28[31] , 
        \wRegInA105[4] , \ScanLink224[7] , \wRegInA28[28] , \ScanLink174[30] , 
        \ScanLink157[18] , \wBMid25[9] , \wAMid51[6] , \wAMid52[5] , 
        \wRegInB7[21] , \wRegInB125[20] , \ScanLink196[4] , \ScanLink122[28] , 
        \wRegInA1[24] , \wRegInB95[8] , \wRegInB106[11] , \ScanLink174[29] , 
        \ScanLink122[31] , \ScanLink101[19] , \wRegInB113[25] , 
        \ScanLink239[8] , \wAMid113[8] , \wAMid14[10] , \wAMid83[0] , 
        \wAIn112[31] , \wAIn112[28] , \wRegInA39[7] , \ScanLink195[7] , 
        \wRegInB59[2] , \wAMid22[15] , \wAMid37[21] , \wBIn38[26] , 
        \wBMid38[6] , \wAMid61[20] , \wAMid42[11] , \wRegInA24[8] , 
        \wBIn74[1] , \ScanLink188[8] , \ScanLink147[1] , \wRegInA106[7] , 
        \wAMid57[25] , \wRegInA85[31] , \ScanLink79[3] , \wBIn58[22] , 
        \wAMid74[14] , \wBIn118[22] , \wRegInA85[28] , \ScanLink227[4] , 
        \ScanLink1[6] , \wAMid9[29] , \wAIn35[4] , \wBIn108[0] , \wBIn82[1] , 
        \wAIn116[19] , \wAMid10[21] , \wAMid65[11] , \wAMid75[0] , 
        \wBIn109[27] , \ScanLink203[2] , \wAMid10[12] , \wAMid26[24] , 
        \wAMid33[10] , \wAMid46[20] , \wBIn49[27] , \wRegInA122[1] , 
        \wBIn50[7] , \wAMid53[14] , \ScanLink163[7] , \wAMid26[17] , 
        \wBIn29[23] , \wAIn36[7] , \wBIn53[4] , \wAMid70[25] , \wRegInA81[19] , 
        \wBIn84[23] , \wBIn91[17] , \wBMid116[16] , \wRegInB63[8] , 
        \wRegInA121[2] , \wRegInA59[30] , \ScanLink200[1] , \ScanLink1[11] , 
        \wBMid103[22] , \wRegInA59[29] , \ScanLink160[4] , \wAMid76[3] , 
        \wBMid120[13] , \wRegInB3[10] , \wRegInA5[15] , \wRegInB102[20] , 
        \wRegInB121[11] , \ScanLink105[31] , \ScanLink153[29] , 
        \ScanLink126[19] , \ScanLink43[9] , \ScanLink105[28] , \ScanLink2[5] , 
        \wRegInB117[14] , \ScanLink170[18] , \ScanLink153[30] , \wBIn81[2] , 
        \wAIn28[31] , \wBIn29[10] , \wAMid53[27] , \ScanLink39[1] , 
        \wAMid70[16] , \wAIn28[28] , \wAMid65[22] , \wRegInB44[29] , 
        \wBMid78[4] , \wBIn109[14] , \wRegInB12[31] , \wRegInB31[19] , 
        \wAMid33[23] , \wBIn34[3] , \wAMid46[13] , \wBIn49[14] , \wAIn83[6] , 
        \wRegInB44[30] , \wRegInB67[18] , \wAIn105[4] , \wRegInB12[28] , 
        \ScanLink107[3] , \wAMid11[4] , \wRegInB19[0] , \wRegInB117[7] , 
        \ScanLink218[28] , \ScanLink218[31] , \ScanLink25[30] , \wAMid12[7] , 
        \wBMid39[30] , \wBMid39[29] , \wAIn51[0] , \wBMid121[6] , 
        \ScanLink73[28] , \ScanLink25[29] , \wRegInA79[5] , \ScanLink50[19] , 
        \wAIn52[3] , \wRegInA5[26] , \wRegInB114[4] , \ScanLink73[31] , 
        \wRegInB117[27] , \ScanLink88[30] , \wBMid94[29] , \wRegInB3[23] , 
        \wRegInB121[22] , \wBIn14[19] , \wAIn15[21] , \wAIn36[10] , 
        \wBIn37[0] , \wBMid66[8] , \ScanLink88[29] , \wAIn80[5] , \wBIn84[10] , 
        \wBMid94[30] , \wBMid122[5] , \wRegInB102[13] , \wAIn85[31] , 
        \wBMid103[11] , \wBMid120[20] , \wAIn106[7] , \wRegInA67[9] , 
        \wAIn85[28] , \ScanLink104[0] , \wBIn91[24] , \wBMid116[25] , 
        \wRegInB79[20] , \ScanLink1[22] , \wAIn43[20] , \ScanLink46[4] , 
        \ScanLink7[8] , \wAIn60[11] , \ScanLink218[3] , \wAIn23[24] , 
        \wBIn37[31] , \wBIn61[29] , \wAIn75[25] , \wBIn102[18] , \wBIn121[30] , 
        \wBMid27[11] , \wBIn37[28] , \wBIn42[18] , \wBMid52[21] , \wAIn56[14] , 
        \wBIn61[30] , \wBMid71[10] , \wBIn121[29] , \wRegInB19[24] , 
        \ScanLink178[6] , \ScanLink245[25] , \ScanLink213[24] , 
        \ScanLink94[2] , \wRegInB66[5] , \ScanLink230[15] , \ScanLink18[20] , 
        \ScanLink195[12] , \wBMid47[15] , \wAIn9[3] , \wBMid32[25] , 
        \ScanLink250[11] , \ScanLink78[24] , \ScanLink225[21] , 
        \ScanLink180[26] , \wBIn113[1] , \wAIn6[21] , \wBMid11[14] , 
        \wBMid64[24] , \wAIn108[12] , \wAIn30[9] , \wBIn56[9] , \wBIn99[0] , 
        \wBIn110[2] , \wRegInB65[6] , \ScanLink206[10] , \ScanLink165[9] , 
        \ScanLink138[12] , \ScanLink96[11] , \ScanLink58[8] , \ScanLink97[1] , 
        \wRegInA27[26] , \wRegInA52[16] , \wRegInA71[27] , \wRegInB78[9] , 
        \ScanLink158[16] , \ScanLink83[25] , \wRegInB82[21] , \ScanLink45[7] , 
        \wBMid32[16] , \wBIn48[5] , \wAMid104[18] , \wRegInA47[22] , 
        \wRegInA8[9] , \wRegInA32[12] , \wRegInB97[15] , \wRegInA11[23] , 
        \wRegInA64[13] , \ScanLink78[17] , \wBMid47[26] , \wRegInA111[29] , 
        \ScanLink225[12] , \ScanLink180[15] , \wBMid11[27] , \ScanLink250[22] , 
        \wBMid64[17] , \wRegInA111[30] , \ScanLink206[23] , \wAMid14[9] , 
        \wAIn15[12] , \wAIn23[17] , \wBMid27[22] , \wBMid71[23] , \wAIn85[8] , 
        \wAIn108[21] , \ScanLink213[17] , \wRegInA62[4] , \ScanLink230[26] , 
        \ScanLink195[21] , \wBMid52[12] , \ScanLink245[16] , \wAIn56[27] , 
        \wAIn75[16] , \wRegInB111[9] , \ScanLink18[13] , \wRegInB19[17] , 
        \ScanLink22[0] , \wAIn36[23] , \wAIn43[13] , \wAMid58[18] , 
        \wAIn98[7] , \wRegInB79[13] , \wAIn60[22] , \wBMid63[5] , 
        \wRegInA11[10] , \wRegInA32[21] , \wRegInB97[26] , \wRegInA47[11] , 
        \ScanLink21[3] , \wRegInA64[20] , \wAIn49[2] , \wBMid60[6] , 
        \wRegInA71[14] , \wAMid80[31] , \wAMid80[28] , \wRegInA27[15] , 
        \wRegInA52[25] , \wRegInB82[12] , \wRegInA61[7] , \ScanLink158[25] , 
        \ScanLink96[22] , \ScanLink83[16] , \ScanLink138[21] , \wBMid80[17] , 
        \wAIn84[22] , \wAIn91[16] , \wAIn100[9] , \wRegInA58[10] , 
        \wRegInB88[27] , \wRegInB119[1] , \wRegInB17[6] , \ScanLink0[28] , 
        \wRegInA38[14] , \wRegInA77[3] , \ScanLink0[31] , \ScanLink147[24] , 
        \ScanLink132[14] , \ScanLink37[7] , \ScanLink164[15] , \wBIn1[16] , 
        \wAMid8[10] , \wBMid9[31] , \wAIn42[9] , \wBMid76[2] , \wRegInB2[30] , 
        \ScanLink171[21] , \ScanLink111[25] , \ScanLink89[23] , 
        \wRegInB103[19] , \wRegInB120[31] , \ScanLink104[11] , 
        \ScanLink152[10] , \wBMid58[27] , \wBMid95[23] , \wRegInB2[29] , 
        \wRegInB120[28] , \ScanLink127[20] , \ScanLink109[5] , 
        \ScanLink12[26] , \wBMid9[28] , \wAIn117[20] , \ScanLink67[16] , 
        \ScanLink31[17] , \ScanLink219[22] , \ScanLink34[4] , \ScanLink44[27] , 
        \ScanLink24[23] , \wAMid11[18] , \wBIn24[9] , \wAIn29[22] , 
        \wAMid32[29] , \wBIn39[6] , \wAIn102[14] , \wAIn108[1] , 
        \ScanLink51[13] , \wBMid38[23] , \wAIn121[25] , \ScanLink72[22] , 
        \wAIn49[26] , \wBMid75[1] , \wRegInB14[5] , \wRegInB50[17] , 
        \wRegInB25[27] , \wRegInB73[26] , \wRegInA80[20] , \wAMid47[19] , 
        \wAMid64[31] , \wRegInB66[12] , \wRegInA74[0] , \ScanLink117[9] , 
        \wAMid32[30] , \wRegInB13[22] , \wBMid12[6] , \wAMid64[28] , 
        \wRegInB45[23] , \wAMid66[9] , \wBMid80[24] , \wBMid95[10] , 
        \wRegInB30[13] , \wRegInA95[14] , \ScanLink171[12] , \ScanLink104[22] , 
        \ScanLink89[10] , \wAMid124[7] , \ScanLink152[23] , \ScanLink127[13] , 
        \ScanLink53[3] , \ScanLink132[27] , \wBIn91[8] , \ScanLink147[17] , 
        \ScanLink111[16] , \ScanLink164[26] , \wAIn29[11] , \wAIn84[11] , 
        \wRegInB73[2] , \wBIn85[30] , \wBMid102[31] , \wBIn106[6] , 
        \wRegInA38[27] , \wRegInB88[14] , \ScanLink81[5] , \wRegInA13[7] , 
        \wRegInA58[23] , \wBIn85[29] , \wBMid102[28] , \wBMid121[19] , 
        \wRegInA3[2] , \wAIn91[25] , \wRegInB13[11] , \wAMid78[5] , 
        \wRegInB25[14] , \wRegInB30[20] , \wRegInB66[21] , \ScanLink82[6] , 
        \wRegInA95[27] , \wRegInB45[10] , \wRegInB70[1] , \ScanLink213[8] , 
        \wRegInA80[13] , \wAMid0[5] , \wAIn2[8] , \wAMid8[23] , \wBIn28[30] , 
        \wRegInB50[24] , \wBIn28[29] , \wAIn38[1] , \wAIn49[15] , \wBIn105[5] , 
        \wRegInA10[4] , \wRegInB73[15] , \ScanLink51[20] , \wBMid11[5] , 
        \wBMid38[10] , \wAIn102[27] , \ScanLink50[0] , \ScanLink24[10] , 
        \ScanLink72[11] , \wAIn121[16] , \ScanLink67[25] , \wAIn3[30] , 
        \wBMid2[24] , \wBMid2[17] , \wAIn14[18] , \wBIn15[20] , \wBIn21[4] , 
        \wAIn59[8] , \wBMid58[14] , \wAIn96[1] , \wAIn117[13] , 
        \ScanLink219[11] , \ScanLink12[15] , \ScanLink44[14] , \wRegInB9[16] , 
        \wRegInB11[8] , \ScanLink31[24] , \wRegInB108[26] , \wAIn110[3] , 
        \wBIn36[11] , \wAMid39[16] , \wBIn43[21] , \wAIn44[7] , \wAMid94[16] , 
        \wAMid126[10] , \ScanLink112[4] , \ScanLink97[31] , \ScanLink97[28] , 
        \wRegInB102[0] , \wAMid105[21] , \wRegInB83[18] , \ScanLink31[9] , 
        \wAMid81[22] , \wBMid109[24] , \wAMid110[15] , \wBIn120[10] , 
        \wBIn60[10] , \wRegInB101[3] , \wBIn103[21] , \wAIn61[28] , 
        \wBIn75[24] , \wBIn116[15] , \wBIn23[25] , \wAIn37[30] , \wAIn42[19] , 
        \wAIn47[4] , \wBIn56[15] , \wAMid59[12] , \wAIn61[31] , 
        \wRegInB78[19] , \wBMid26[31] , \wBMid26[28] , \wAIn37[29] , 
        \wRegInA110[23] , \ScanLink251[31] , \ScanLink207[29] , 
        \ScanLink251[28] , \ScanLink224[18] , \ScanLink207[30] , \wBMid53[18] , 
        \wBMid70[30] , \wRegInA105[17] , \ScanLink19[19] , \wRegInA126[26] , 
        \wBMid70[29] , \wAIn95[2] , \ScanLink111[7] , \wAIn7[5] , \wBIn22[7] , 
        \wAIn113[0] , \wAMid60[7] , \wAMid81[11] , \wBMid109[17] , 
        \wAMid110[26] , \wRegInB68[3] , \wAMid94[25] , \wRegInA65[19] , 
        \wAMid126[23] , \wRegInA46[31] , \wBMid14[8] , \wRegInA10[29] , 
        \wAIn20[3] , \wBIn45[0] , \wBIn97[6] , \wAMid122[9] , \wRegInA46[28] , 
        \wBIn100[8] , \wAMid105[12] , \wRegInA10[30] , \wRegInA33[18] , 
        \wRegInA15[9] , \wRegInB108[15] , \ScanLink216[5] , \ScanLink139[18] , 
        \ScanLink48[2] , \wRegInB9[25] , \ScanLink176[0] , \wRegInA105[24] , 
        \ScanLink215[6] , \ScanLink194[18] , \wAIn4[6] , \wAIn7[18] , 
        \wBIn46[3] , \wAIn109[18] , \wRegInA126[15] , \ScanLink84[8] , 
        \ScanLink175[3] , \wBIn15[13] , \wAIn23[0] , \wBIn23[16] , 
        \wBIn75[17] , \wBIn116[26] , \wRegInA110[10] , \ScanLink208[9] , 
        \wBIn36[22] , \wAMid39[25] , \wBIn56[26] , \ScanLink99[7] , 
        \wAMid59[21] , \wBIn43[12] , \wBIn94[5] , \wBIn120[23] , \wBIn60[23] , 
        \wAMid63[4] , \wBIn103[12] , \wBMid6[15] , \wAMid95[4] , \wAMid118[3] , 
        \wRegInA101[15] , \ScanLink190[29] , \ScanLink190[30] , 
        \wRegInA122[24] , \ScanLink151[5] , \wBIn62[5] , \wRegInA110[3] , 
        \wRegInB52[9] , \wRegInA114[21] , \wBMid1[2] , \wAIn3[29] , 
        \ScanLink231[0] , \wAMid3[6] , \wBIn11[22] , \wBIn27[27] , 
        \wAMid47[2] , \wBIn71[26] , \wBIn112[17] , \wBIn52[17] , \wAMid28[20] , 
        \wBIn32[13] , \wBIn47[23] , \wAMid48[24] , \ScanLink183[3] , 
        \wBIn124[12] , \wBIn64[12] , \ScanLink72[8] , \wBIn107[23] , 
        \wAMid44[1] , \wAMid114[17] , \ScanLink180[0] , \wBIn61[6] , 
        \wAMid85[20] , \wAMid90[14] , \wAMid122[12] , \wRegInA14[18] , 
        \wRegInA37[30] , \wAMid101[23] , \wBMid118[12] , \wRegInA61[28] , 
        \wRegInA37[29] , \wRegInA42[19] , \wRegInA61[31] , \ScanLink148[19] , 
        \wAMid96[7] , \wRegInB119[10] , \ScanLink152[6] , \ScanLink232[3] , 
        \wBIn8[9] , \wBIn32[20] , \wRegInA113[0] , \wBIn47[10] , \wAMid48[17] , 
        \wAIn63[2] , \wBIn11[11] , \wAMid23[6] , \wBIn124[21] , \wBMid57[9] , 
        \wBIn64[21] , \wBMid98[0] , \wBMid113[4] , \wBIn107[10] , \wBMid2[1] , 
        \wBMid6[26] , \wAIn10[30] , \wAIn10[29] , \wRegInB125[5] , 
        \wBIn27[14] , \wAIn33[18] , \wAIn46[31] , \wAIn65[19] , \wBIn112[24] , 
        \wBIn71[15] , \wBMid22[19] , \wAMid28[13] , \wAIn46[28] , \wBIn52[24] , 
        \wBMid57[29] , \wRegInA56[8] , \wRegInA99[1] , \wRegInA114[12] , 
        \ScanLink255[19] , \ScanLink220[30] , \ScanLink203[18] , 
        \ScanLink135[1] , \ScanLink220[29] , \wRegInA101[26] , 
        \ScanLink255[4] , \ScanLink68[18] , \wBMid57[30] , \wAMid20[5] , 
        \wBMid49[5] , \wBMid74[18] , \wRegInA122[17] , \wAMid90[27] , 
        \wRegInB119[23] , \ScanLink136[2] , \ScanLink93[19] , \ScanLink256[7] , 
        \wBMid118[21] , \wAIn60[1] , \wBMid110[7] , \wAMid122[21] , 
        \wAMid85[13] , \wAMid101[10] , \wRegInA48[4] , \wAMid114[24] , 
        \wRegInB87[29] , \wRegInB28[1] , \wRegInB126[6] , \wBIn5[27] , 
        \wAIn8[16] , \wAIn38[14] , \wAIn58[10] , \wBIn121[3] , \wRegInA34[2] , 
        \wRegInB87[30] , \wRegInB62[10] , \wBIn59[31] , \wBIn119[28] , 
        \wRegInB17[20] , \wRegInB34[11] , \wRegInB41[21] , \ScanLink198[2] , 
        \wRegInA91[16] , \wRegInB54[15] , \wRegInB54[7] , \wRegInB21[25] , 
        \wRegInA84[22] , \wRegInB77[24] , \wBMid49[11] , \wBIn59[28] , 
        \wBIn119[31] , \ScanLink69[9] , \wBIn79[4] , \wAMid103[2] , 
        \ScanLink20[21] , \wAIn106[16] , \ScanLink208[14] , \ScanLink55[11] , 
        \wRegInB9[8] , \wBMid29[15] , \wBMid35[3] , \wAIn125[27] , 
        \ScanLink76[20] , \wRegInB49[8] , \wRegInB86[1] , \ScanLink16[24] , 
        \wBMid36[0] , \wAIn113[22] , \ScanLink63[14] , \ScanLink175[23] , 
        \ScanLink74[6] , \ScanLink35[15] , \ScanLink40[25] , \wBMid84[15] , 
        \wBMid91[21] , \wAMid100[1] , \ScanLink156[12] , \ScanLink100[13] , 
        \wRegInA108[1] , \ScanLink149[7] , \ScanLink123[22] , 
        \ScanLink143[26] , \ScanLink136[16] , \ScanLink77[5] , \wRegInB85[2] , 
        \ScanLink160[17] , \wBIn5[14] , \wAMid5[8] , \wBIn67[8] , \wAIn80[20] , 
        \ScanLink229[2] , \ScanLink98[15] , \ScanLink115[27] , \wAMid90[9] , 
        \wBIn122[0] , \wRegInA37[1] , \wRegInA49[26] , \wBIn81[18] , 
        \wAIn95[14] , \wBMid125[28] , \wRegInB99[11] , \ScanLink154[8] , 
        \wRegInA29[22] , \wRegInB57[4] , \wBMid125[31] , \wBMid106[19] , 
        \wAIn8[25] , \wAMid25[8] , \wBMid29[26] , \wBMid49[22] , \wBMid51[7] , 
        \ScanLink63[27] , \wAIn106[25] , \wAIn113[11] , \wRegInA82[0] , 
        \ScanLink40[16] , \ScanLink16[17] , \ScanLink208[27] , 
        \ScanLink55[22] , \ScanLink35[26] , \ScanLink20[12] , \ScanLink76[13] , 
        \ScanLink10[2] , \wAIn125[14] , \wAMid15[30] , \wAIn38[27] , 
        \wAMid38[7] , \wRegInB21[16] , \wRegInA84[11] , \wAIn78[3] , 
        \wBMid83[1] , \wBMid108[5] , \wRegInB54[26] , \wRegInA50[6] , 
        \wRegInB77[17] , \wAMid43[28] , \wAIn58[23] , \wRegInB17[13] , 
        \wAMid15[29] , \wAMid36[18] , \wAMid43[31] , \wRegInB62[23] , 
        \wAMid60[19] , \wRegInB30[3] , \wRegInB34[22] , \wRegInA91[25] , 
        \wBMid52[4] , \wAIn80[13] , \wBMid80[2] , \wRegInA29[11] , 
        \wRegInB41[12] , \wRegInA53[5] , \wAIn95[27] , \wRegInB33[0] , 
        \wBMid84[26] , \wRegInA49[15] , \wRegInB99[22] , \ScanLink250[9] , 
        \ScanLink4[19] , \wRegInA81[3] , \ScanLink136[25] , \wBMid116[9] , 
        \ScanLink160[24] , \ScanLink143[15] , \ScanLink115[14] , 
        \ScanLink98[26] , \wBMid91[12] , \wRegInB6[18] , \wRegInB107[28] , 
        \wRegInB120[8] , \ScanLink100[20] , \ScanLink175[10] , 
        \wRegInB107[31] , \wRegInB124[19] , \ScanLink123[11] , 
        \ScanLink156[21] , \ScanLink13[1] ;
    BubbleSort_Node_WIDTH32 BSN1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn0[31] , 
        \wAIn0[30] , \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , \wAIn0[26] , 
        \wAIn0[25] , \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , \wAIn0[21] , 
        \wAIn0[20] , \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , \wAIn0[16] , 
        \wAIn0[15] , \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , \wAIn0[11] , 
        \wAIn0[10] , \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , \wAIn0[6] , 
        \wAIn0[5] , \wAIn0[4] , \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , \wAIn0[0] 
        }), .BIn({\wBIn0[31] , \wBIn0[30] , \wBIn0[29] , \wBIn0[28] , 
        \wBIn0[27] , \wBIn0[26] , \wBIn0[25] , \wBIn0[24] , \wBIn0[23] , 
        \wBIn0[22] , \wBIn0[21] , \wBIn0[20] , \wBIn0[19] , \wBIn0[18] , 
        \wBIn0[17] , \wBIn0[16] , \wBIn0[15] , \wBIn0[14] , \wBIn0[13] , 
        \wBIn0[12] , \wBIn0[11] , \wBIn0[10] , \wBIn0[9] , \wBIn0[8] , 
        \wBIn0[7] , \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , \wBIn0[3] , \wBIn0[2] , 
        \wBIn0[1] , \wBIn0[0] }), .HiOut({\wRegInA0[31] , \wRegInA0[30] , 
        \wRegInA0[29] , \wRegInA0[28] , \wRegInA0[27] , \wRegInA0[26] , 
        \wRegInA0[25] , \wRegInA0[24] , \wRegInA0[23] , \wRegInA0[22] , 
        \wRegInA0[21] , \wRegInA0[20] , \wRegInA0[19] , \wRegInA0[18] , 
        \wRegInA0[17] , \wRegInA0[16] , \wRegInA0[15] , \wRegInA0[14] , 
        \wRegInA0[13] , \wRegInA0[12] , \wRegInA0[11] , \wRegInA0[10] , 
        \wRegInA0[9] , \wRegInA0[8] , \wRegInA0[7] , \wRegInA0[6] , 
        \wRegInA0[5] , \wRegInA0[4] , \wRegInA0[3] , \wRegInA0[2] , 
        \wRegInA0[1] , \wRegInA0[0] }), .LoOut({\wAMid0[31] , \wAMid0[30] , 
        \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , \wAMid0[25] , 
        \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , \wAMid0[20] , 
        \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , \wAMid0[15] , 
        \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , \wAMid0[10] , 
        \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , \wAMid0[5] , 
        \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , \wAMid0[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn2[31] , 
        \wAIn2[30] , \wAIn2[29] , \wAIn2[28] , \wAIn2[27] , \wAIn2[26] , 
        \wAIn2[25] , \wAIn2[24] , \wAIn2[23] , \wAIn2[22] , \wAIn2[21] , 
        \wAIn2[20] , \wAIn2[19] , \wAIn2[18] , \wAIn2[17] , \wAIn2[16] , 
        \wAIn2[15] , \wAIn2[14] , \wAIn2[13] , \wAIn2[12] , \wAIn2[11] , 
        \wAIn2[10] , \wAIn2[9] , \wAIn2[8] , \wAIn2[7] , \wAIn2[6] , 
        \wAIn2[5] , \wAIn2[4] , \wAIn2[3] , \wAIn2[2] , \wAIn2[1] , \wAIn2[0] 
        }), .BIn({\wBIn2[31] , \wBIn2[30] , \wBIn2[29] , \wBIn2[28] , 
        \wBIn2[27] , \wBIn2[26] , \wBIn2[25] , \wBIn2[24] , \wBIn2[23] , 
        \wBIn2[22] , \wBIn2[21] , \wBIn2[20] , \wBIn2[19] , \wBIn2[18] , 
        \wBIn2[17] , \wBIn2[16] , \wBIn2[15] , \wBIn2[14] , \wBIn2[13] , 
        \wBIn2[12] , \wBIn2[11] , \wBIn2[10] , \wBIn2[9] , \wBIn2[8] , 
        \wBIn2[7] , \wBIn2[6] , \wBIn2[5] , \wBIn2[4] , \wBIn2[3] , \wBIn2[2] , 
        \wBIn2[1] , \wBIn2[0] }), .HiOut({\wBMid1[31] , \wBMid1[30] , 
        \wBMid1[29] , \wBMid1[28] , \wBMid1[27] , \wBMid1[26] , \wBMid1[25] , 
        \wBMid1[24] , \wBMid1[23] , \wBMid1[22] , \wBMid1[21] , \wBMid1[20] , 
        \wBMid1[19] , \wBMid1[18] , \wBMid1[17] , \wBMid1[16] , \wBMid1[15] , 
        \wBMid1[14] , \wBMid1[13] , \wBMid1[12] , \wBMid1[11] , \wBMid1[10] , 
        \wBMid1[9] , \wBMid1[8] , \wBMid1[7] , \wBMid1[6] , \wBMid1[5] , 
        \wBMid1[4] , \wBMid1[3] , \wBMid1[2] , \wBMid1[1] , \wBMid1[0] }), 
        .LoOut({\wAMid2[31] , \wAMid2[30] , \wAMid2[29] , \wAMid2[28] , 
        \wAMid2[27] , \wAMid2[26] , \wAMid2[25] , \wAMid2[24] , \wAMid2[23] , 
        \wAMid2[22] , \wAMid2[21] , \wAMid2[20] , \wAMid2[19] , \wAMid2[18] , 
        \wAMid2[17] , \wAMid2[16] , \wAMid2[15] , \wAMid2[14] , \wAMid2[13] , 
        \wAMid2[12] , \wAMid2[11] , \wAMid2[10] , \wAMid2[9] , \wAMid2[8] , 
        \wAMid2[7] , \wAMid2[6] , \wAMid2[5] , \wAMid2[4] , \wAMid2[3] , 
        \wAMid2[2] , \wAMid2[1] , \wAMid2[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn3[31] , 
        \wAIn3[30] , \wAIn3[29] , \wAIn3[28] , \wAIn3[27] , \wAIn3[26] , 
        \wAIn3[25] , \wAIn3[24] , \wAIn3[23] , \wAIn3[22] , \wAIn3[21] , 
        \wAIn3[20] , \wAIn3[19] , \wAIn3[18] , \wAIn3[17] , \wAIn3[16] , 
        \wAIn3[15] , \wAIn3[14] , \wAIn3[13] , \wAIn3[12] , \wAIn3[11] , 
        \wAIn3[10] , \wAIn3[9] , \wAIn3[8] , \wAIn3[7] , \wAIn3[6] , 
        \wAIn3[5] , \wAIn3[4] , \wAIn3[3] , \wAIn3[2] , \wAIn3[1] , \wAIn3[0] 
        }), .BIn({\wBIn3[31] , \wBIn3[30] , \wBIn3[29] , \wBIn3[28] , 
        \wBIn3[27] , \wBIn3[26] , \wBIn3[25] , \wBIn3[24] , \wBIn3[23] , 
        \wBIn3[22] , \wBIn3[21] , \wBIn3[20] , \wBIn3[19] , \wBIn3[18] , 
        \wBIn3[17] , \wBIn3[16] , \wBIn3[15] , \wBIn3[14] , \wBIn3[13] , 
        \wBIn3[12] , \wBIn3[11] , \wBIn3[10] , \wBIn3[9] , \wBIn3[8] , 
        \wBIn3[7] , \wBIn3[6] , \wBIn3[5] , \wBIn3[4] , \wBIn3[3] , \wBIn3[2] , 
        \wBIn3[1] , \wBIn3[0] }), .HiOut({\wBMid2[31] , \wBMid2[30] , 
        \wBMid2[29] , \wBMid2[28] , \wBMid2[27] , \wBMid2[26] , \wBMid2[25] , 
        \wBMid2[24] , \wBMid2[23] , \wBMid2[22] , \wBMid2[21] , \wBMid2[20] , 
        \wBMid2[19] , \wBMid2[18] , \wBMid2[17] , \wBMid2[16] , \wBMid2[15] , 
        \wBMid2[14] , \wBMid2[13] , \wBMid2[12] , \wBMid2[11] , \wBMid2[10] , 
        \wBMid2[9] , \wBMid2[8] , \wBMid2[7] , \wBMid2[6] , \wBMid2[5] , 
        \wBMid2[4] , \wBMid2[3] , \wBMid2[2] , \wBMid2[1] , \wBMid2[0] }), 
        .LoOut({\wAMid3[31] , \wAMid3[30] , \wAMid3[29] , \wAMid3[28] , 
        \wAMid3[27] , \wAMid3[26] , \wAMid3[25] , \wAMid3[24] , \wAMid3[23] , 
        \wAMid3[22] , \wAMid3[21] , \wAMid3[20] , \wAMid3[19] , \wAMid3[18] , 
        \wAMid3[17] , \wAMid3[16] , \wAMid3[15] , \wAMid3[14] , \wAMid3[13] , 
        \wAMid3[12] , \wAMid3[11] , \wAMid3[10] , \wAMid3[9] , \wAMid3[8] , 
        \wAMid3[7] , \wAMid3[6] , \wAMid3[5] , \wAMid3[4] , \wAMid3[3] , 
        \wAMid3[2] , \wAMid3[1] , \wAMid3[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn4[31] , 
        \wAIn4[30] , \wAIn4[29] , \wAIn4[28] , \wAIn4[27] , \wAIn4[26] , 
        \wAIn4[25] , \wAIn4[24] , \wAIn4[23] , \wAIn4[22] , \wAIn4[21] , 
        \wAIn4[20] , \wAIn4[19] , \wAIn4[18] , \wAIn4[17] , \wAIn4[16] , 
        \wAIn4[15] , \wAIn4[14] , \wAIn4[13] , \wAIn4[12] , \wAIn4[11] , 
        \wAIn4[10] , \wAIn4[9] , \wAIn4[8] , \wAIn4[7] , \wAIn4[6] , 
        \wAIn4[5] , \wAIn4[4] , \wAIn4[3] , \wAIn4[2] , \wAIn4[1] , \wAIn4[0] 
        }), .BIn({\wBIn4[31] , \wBIn4[30] , \wBIn4[29] , \wBIn4[28] , 
        \wBIn4[27] , \wBIn4[26] , \wBIn4[25] , \wBIn4[24] , \wBIn4[23] , 
        \wBIn4[22] , \wBIn4[21] , \wBIn4[20] , \wBIn4[19] , \wBIn4[18] , 
        \wBIn4[17] , \wBIn4[16] , \wBIn4[15] , \wBIn4[14] , \wBIn4[13] , 
        \wBIn4[12] , \wBIn4[11] , \wBIn4[10] , \wBIn4[9] , \wBIn4[8] , 
        \wBIn4[7] , \wBIn4[6] , \wBIn4[5] , \wBIn4[4] , \wBIn4[3] , \wBIn4[2] , 
        \wBIn4[1] , \wBIn4[0] }), .HiOut({\wBMid3[31] , \wBMid3[30] , 
        \wBMid3[29] , \wBMid3[28] , \wBMid3[27] , \wBMid3[26] , \wBMid3[25] , 
        \wBMid3[24] , \wBMid3[23] , \wBMid3[22] , \wBMid3[21] , \wBMid3[20] , 
        \wBMid3[19] , \wBMid3[18] , \wBMid3[17] , \wBMid3[16] , \wBMid3[15] , 
        \wBMid3[14] , \wBMid3[13] , \wBMid3[12] , \wBMid3[11] , \wBMid3[10] , 
        \wBMid3[9] , \wBMid3[8] , \wBMid3[7] , \wBMid3[6] , \wBMid3[5] , 
        \wBMid3[4] , \wBMid3[3] , \wBMid3[2] , \wBMid3[1] , \wBMid3[0] }), 
        .LoOut({\wAMid4[31] , \wAMid4[30] , \wAMid4[29] , \wAMid4[28] , 
        \wAMid4[27] , \wAMid4[26] , \wAMid4[25] , \wAMid4[24] , \wAMid4[23] , 
        \wAMid4[22] , \wAMid4[21] , \wAMid4[20] , \wAMid4[19] , \wAMid4[18] , 
        \wAMid4[17] , \wAMid4[16] , \wAMid4[15] , \wAMid4[14] , \wAMid4[13] , 
        \wAMid4[12] , \wAMid4[11] , \wAMid4[10] , \wAMid4[9] , \wAMid4[8] , 
        \wAMid4[7] , \wAMid4[6] , \wAMid4[5] , \wAMid4[4] , \wAMid4[3] , 
        \wAMid4[2] , \wAMid4[1] , \wAMid4[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn82[31] , \wAIn82[30] , \wAIn82[29] , \wAIn82[28] , \wAIn82[27] , 
        \wAIn82[26] , \wAIn82[25] , \wAIn82[24] , \wAIn82[23] , \wAIn82[22] , 
        \wAIn82[21] , \wAIn82[20] , \wAIn82[19] , \wAIn82[18] , \wAIn82[17] , 
        \wAIn82[16] , \wAIn82[15] , \wAIn82[14] , \wAIn82[13] , \wAIn82[12] , 
        \wAIn82[11] , \wAIn82[10] , \wAIn82[9] , \wAIn82[8] , \wAIn82[7] , 
        \wAIn82[6] , \wAIn82[5] , \wAIn82[4] , \wAIn82[3] , \wAIn82[2] , 
        \wAIn82[1] , \wAIn82[0] }), .BIn({\wBIn82[31] , \wBIn82[30] , 
        \wBIn82[29] , \wBIn82[28] , \wBIn82[27] , \wBIn82[26] , \wBIn82[25] , 
        \wBIn82[24] , \wBIn82[23] , \wBIn82[22] , \wBIn82[21] , \wBIn82[20] , 
        \wBIn82[19] , \wBIn82[18] , \wBIn82[17] , \wBIn82[16] , \wBIn82[15] , 
        \wBIn82[14] , \wBIn82[13] , \wBIn82[12] , \wBIn82[11] , \wBIn82[10] , 
        \wBIn82[9] , \wBIn82[8] , \wBIn82[7] , \wBIn82[6] , \wBIn82[5] , 
        \wBIn82[4] , \wBIn82[3] , \wBIn82[2] , \wBIn82[1] , \wBIn82[0] }), 
        .HiOut({\wBMid81[31] , \wBMid81[30] , \wBMid81[29] , \wBMid81[28] , 
        \wBMid81[27] , \wBMid81[26] , \wBMid81[25] , \wBMid81[24] , 
        \wBMid81[23] , \wBMid81[22] , \wBMid81[21] , \wBMid81[20] , 
        \wBMid81[19] , \wBMid81[18] , \wBMid81[17] , \wBMid81[16] , 
        \wBMid81[15] , \wBMid81[14] , \wBMid81[13] , \wBMid81[12] , 
        \wBMid81[11] , \wBMid81[10] , \wBMid81[9] , \wBMid81[8] , \wBMid81[7] , 
        \wBMid81[6] , \wBMid81[5] , \wBMid81[4] , \wBMid81[3] , \wBMid81[2] , 
        \wBMid81[1] , \wBMid81[0] }), .LoOut({\wAMid82[31] , \wAMid82[30] , 
        \wAMid82[29] , \wAMid82[28] , \wAMid82[27] , \wAMid82[26] , 
        \wAMid82[25] , \wAMid82[24] , \wAMid82[23] , \wAMid82[22] , 
        \wAMid82[21] , \wAMid82[20] , \wAMid82[19] , \wAMid82[18] , 
        \wAMid82[17] , \wAMid82[16] , \wAMid82[15] , \wAMid82[14] , 
        \wAMid82[13] , \wAMid82[12] , \wAMid82[11] , \wAMid82[10] , 
        \wAMid82[9] , \wAMid82[8] , \wAMid82[7] , \wAMid82[6] , \wAMid82[5] , 
        \wAMid82[4] , \wAMid82[3] , \wAMid82[2] , \wAMid82[1] , \wAMid82[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid39[31] , \wAMid39[30] , \wAMid39[29] , \wAMid39[28] , 
        \wAMid39[27] , \wAMid39[26] , \wAMid39[25] , \wAMid39[24] , 
        \wAMid39[23] , \wAMid39[22] , \wAMid39[21] , \wAMid39[20] , 
        \wAMid39[19] , \wAMid39[18] , \wAMid39[17] , \wAMid39[16] , 
        \wAMid39[15] , \wAMid39[14] , \wAMid39[13] , \wAMid39[12] , 
        \wAMid39[11] , \wAMid39[10] , \wAMid39[9] , \wAMid39[8] , \wAMid39[7] , 
        \wAMid39[6] , \wAMid39[5] , \wAMid39[4] , \wAMid39[3] , \wAMid39[2] , 
        \wAMid39[1] , \wAMid39[0] }), .BIn({\wBMid39[31] , \wBMid39[30] , 
        \wBMid39[29] , \wBMid39[28] , \wBMid39[27] , \wBMid39[26] , 
        \wBMid39[25] , \wBMid39[24] , \wBMid39[23] , \wBMid39[22] , 
        \wBMid39[21] , \wBMid39[20] , \wBMid39[19] , \wBMid39[18] , 
        \wBMid39[17] , \wBMid39[16] , \wBMid39[15] , \wBMid39[14] , 
        \wBMid39[13] , \wBMid39[12] , \wBMid39[11] , \wBMid39[10] , 
        \wBMid39[9] , \wBMid39[8] , \wBMid39[7] , \wBMid39[6] , \wBMid39[5] , 
        \wBMid39[4] , \wBMid39[3] , \wBMid39[2] , \wBMid39[1] , \wBMid39[0] }), 
        .HiOut({\wRegInB39[31] , \wRegInB39[30] , \wRegInB39[29] , 
        \wRegInB39[28] , \wRegInB39[27] , \wRegInB39[26] , \wRegInB39[25] , 
        \wRegInB39[24] , \wRegInB39[23] , \wRegInB39[22] , \wRegInB39[21] , 
        \wRegInB39[20] , \wRegInB39[19] , \wRegInB39[18] , \wRegInB39[17] , 
        \wRegInB39[16] , \wRegInB39[15] , \wRegInB39[14] , \wRegInB39[13] , 
        \wRegInB39[12] , \wRegInB39[11] , \wRegInB39[10] , \wRegInB39[9] , 
        \wRegInB39[8] , \wRegInB39[7] , \wRegInB39[6] , \wRegInB39[5] , 
        \wRegInB39[4] , \wRegInB39[3] , \wRegInB39[2] , \wRegInB39[1] , 
        \wRegInB39[0] }), .LoOut({\wRegInA40[31] , \wRegInA40[30] , 
        \wRegInA40[29] , \wRegInA40[28] , \wRegInA40[27] , \wRegInA40[26] , 
        \wRegInA40[25] , \wRegInA40[24] , \wRegInA40[23] , \wRegInA40[22] , 
        \wRegInA40[21] , \wRegInA40[20] , \wRegInA40[19] , \wRegInA40[18] , 
        \wRegInA40[17] , \wRegInA40[16] , \wRegInA40[15] , \wRegInA40[14] , 
        \wRegInA40[13] , \wRegInA40[12] , \wRegInA40[11] , \wRegInA40[10] , 
        \wRegInA40[9] , \wRegInA40[8] , \wRegInA40[7] , \wRegInA40[6] , 
        \wRegInA40[5] , \wRegInA40[4] , \wRegInA40[3] , \wRegInA40[2] , 
        \wRegInA40[1] , \wRegInA40[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_187 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink188[31] , \ScanLink188[30] , \ScanLink188[29] , 
        \ScanLink188[28] , \ScanLink188[27] , \ScanLink188[26] , 
        \ScanLink188[25] , \ScanLink188[24] , \ScanLink188[23] , 
        \ScanLink188[22] , \ScanLink188[21] , \ScanLink188[20] , 
        \ScanLink188[19] , \ScanLink188[18] , \ScanLink188[17] , 
        \ScanLink188[16] , \ScanLink188[15] , \ScanLink188[14] , 
        \ScanLink188[13] , \ScanLink188[12] , \ScanLink188[11] , 
        \ScanLink188[10] , \ScanLink188[9] , \ScanLink188[8] , 
        \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , \ScanLink188[4] , 
        \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , \ScanLink188[0] 
        }), .ScanOut({\ScanLink187[31] , \ScanLink187[30] , \ScanLink187[29] , 
        \ScanLink187[28] , \ScanLink187[27] , \ScanLink187[26] , 
        \ScanLink187[25] , \ScanLink187[24] , \ScanLink187[23] , 
        \ScanLink187[22] , \ScanLink187[21] , \ScanLink187[20] , 
        \ScanLink187[19] , \ScanLink187[18] , \ScanLink187[17] , 
        \ScanLink187[16] , \ScanLink187[15] , \ScanLink187[14] , 
        \ScanLink187[13] , \ScanLink187[12] , \ScanLink187[11] , 
        \ScanLink187[10] , \ScanLink187[9] , \ScanLink187[8] , 
        \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , \ScanLink187[4] , 
        \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , \ScanLink187[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA34[31] , \wRegInA34[30] , \wRegInA34[29] , 
        \wRegInA34[28] , \wRegInA34[27] , \wRegInA34[26] , \wRegInA34[25] , 
        \wRegInA34[24] , \wRegInA34[23] , \wRegInA34[22] , \wRegInA34[21] , 
        \wRegInA34[20] , \wRegInA34[19] , \wRegInA34[18] , \wRegInA34[17] , 
        \wRegInA34[16] , \wRegInA34[15] , \wRegInA34[14] , \wRegInA34[13] , 
        \wRegInA34[12] , \wRegInA34[11] , \wRegInA34[10] , \wRegInA34[9] , 
        \wRegInA34[8] , \wRegInA34[7] , \wRegInA34[6] , \wRegInA34[5] , 
        \wRegInA34[4] , \wRegInA34[3] , \wRegInA34[2] , \wRegInA34[1] , 
        \wRegInA34[0] }), .Out({\wAIn34[31] , \wAIn34[30] , \wAIn34[29] , 
        \wAIn34[28] , \wAIn34[27] , \wAIn34[26] , \wAIn34[25] , \wAIn34[24] , 
        \wAIn34[23] , \wAIn34[22] , \wAIn34[21] , \wAIn34[20] , \wAIn34[19] , 
        \wAIn34[18] , \wAIn34[17] , \wAIn34[16] , \wAIn34[15] , \wAIn34[14] , 
        \wAIn34[13] , \wAIn34[12] , \wAIn34[11] , \wAIn34[10] , \wAIn34[9] , 
        \wAIn34[8] , \wAIn34[7] , \wAIn34[6] , \wAIn34[5] , \wAIn34[4] , 
        \wAIn34[3] , \wAIn34[2] , \wAIn34[1] , \wAIn34[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn12[31] , \wAIn12[30] , \wAIn12[29] , \wAIn12[28] , \wAIn12[27] , 
        \wAIn12[26] , \wAIn12[25] , \wAIn12[24] , \wAIn12[23] , \wAIn12[22] , 
        \wAIn12[21] , \wAIn12[20] , \wAIn12[19] , \wAIn12[18] , \wAIn12[17] , 
        \wAIn12[16] , \wAIn12[15] , \wAIn12[14] , \wAIn12[13] , \wAIn12[12] , 
        \wAIn12[11] , \wAIn12[10] , \wAIn12[9] , \wAIn12[8] , \wAIn12[7] , 
        \wAIn12[6] , \wAIn12[5] , \wAIn12[4] , \wAIn12[3] , \wAIn12[2] , 
        \wAIn12[1] , \wAIn12[0] }), .BIn({\wBIn12[31] , \wBIn12[30] , 
        \wBIn12[29] , \wBIn12[28] , \wBIn12[27] , \wBIn12[26] , \wBIn12[25] , 
        \wBIn12[24] , \wBIn12[23] , \wBIn12[22] , \wBIn12[21] , \wBIn12[20] , 
        \wBIn12[19] , \wBIn12[18] , \wBIn12[17] , \wBIn12[16] , \wBIn12[15] , 
        \wBIn12[14] , \wBIn12[13] , \wBIn12[12] , \wBIn12[11] , \wBIn12[10] , 
        \wBIn12[9] , \wBIn12[8] , \wBIn12[7] , \wBIn12[6] , \wBIn12[5] , 
        \wBIn12[4] , \wBIn12[3] , \wBIn12[2] , \wBIn12[1] , \wBIn12[0] }), 
        .HiOut({\wBMid11[31] , \wBMid11[30] , \wBMid11[29] , \wBMid11[28] , 
        \wBMid11[27] , \wBMid11[26] , \wBMid11[25] , \wBMid11[24] , 
        \wBMid11[23] , \wBMid11[22] , \wBMid11[21] , \wBMid11[20] , 
        \wBMid11[19] , \wBMid11[18] , \wBMid11[17] , \wBMid11[16] , 
        \wBMid11[15] , \wBMid11[14] , \wBMid11[13] , \wBMid11[12] , 
        \wBMid11[11] , \wBMid11[10] , \wBMid11[9] , \wBMid11[8] , \wBMid11[7] , 
        \wBMid11[6] , \wBMid11[5] , \wBMid11[4] , \wBMid11[3] , \wBMid11[2] , 
        \wBMid11[1] , \wBMid11[0] }), .LoOut({\wAMid12[31] , \wAMid12[30] , 
        \wAMid12[29] , \wAMid12[28] , \wAMid12[27] , \wAMid12[26] , 
        \wAMid12[25] , \wAMid12[24] , \wAMid12[23] , \wAMid12[22] , 
        \wAMid12[21] , \wAMid12[20] , \wAMid12[19] , \wAMid12[18] , 
        \wAMid12[17] , \wAMid12[16] , \wAMid12[15] , \wAMid12[14] , 
        \wAMid12[13] , \wAMid12[12] , \wAMid12[11] , \wAMid12[10] , 
        \wAMid12[9] , \wAMid12[8] , \wAMid12[7] , \wAMid12[6] , \wAMid12[5] , 
        \wAMid12[4] , \wAMid12[3] , \wAMid12[2] , \wAMid12[1] , \wAMid12[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn35[31] , \wAIn35[30] , \wAIn35[29] , \wAIn35[28] , \wAIn35[27] , 
        \wAIn35[26] , \wAIn35[25] , \wAIn35[24] , \wAIn35[23] , \wAIn35[22] , 
        \wAIn35[21] , \wAIn35[20] , \wAIn35[19] , \wAIn35[18] , \wAIn35[17] , 
        \wAIn35[16] , \wAIn35[15] , \wAIn35[14] , \wAIn35[13] , \wAIn35[12] , 
        \wAIn35[11] , \wAIn35[10] , \wAIn35[9] , \wAIn35[8] , \wAIn35[7] , 
        \wAIn35[6] , \wAIn35[5] , \wAIn35[4] , \wAIn35[3] , \wAIn35[2] , 
        \wAIn35[1] , \wAIn35[0] }), .BIn({\wBIn35[31] , \wBIn35[30] , 
        \wBIn35[29] , \wBIn35[28] , \wBIn35[27] , \wBIn35[26] , \wBIn35[25] , 
        \wBIn35[24] , \wBIn35[23] , \wBIn35[22] , \wBIn35[21] , \wBIn35[20] , 
        \wBIn35[19] , \wBIn35[18] , \wBIn35[17] , \wBIn35[16] , \wBIn35[15] , 
        \wBIn35[14] , \wBIn35[13] , \wBIn35[12] , \wBIn35[11] , \wBIn35[10] , 
        \wBIn35[9] , \wBIn35[8] , \wBIn35[7] , \wBIn35[6] , \wBIn35[5] , 
        \wBIn35[4] , \wBIn35[3] , \wBIn35[2] , \wBIn35[1] , \wBIn35[0] }), 
        .HiOut({\wBMid34[31] , \wBMid34[30] , \wBMid34[29] , \wBMid34[28] , 
        \wBMid34[27] , \wBMid34[26] , \wBMid34[25] , \wBMid34[24] , 
        \wBMid34[23] , \wBMid34[22] , \wBMid34[21] , \wBMid34[20] , 
        \wBMid34[19] , \wBMid34[18] , \wBMid34[17] , \wBMid34[16] , 
        \wBMid34[15] , \wBMid34[14] , \wBMid34[13] , \wBMid34[12] , 
        \wBMid34[11] , \wBMid34[10] , \wBMid34[9] , \wBMid34[8] , \wBMid34[7] , 
        \wBMid34[6] , \wBMid34[5] , \wBMid34[4] , \wBMid34[3] , \wBMid34[2] , 
        \wBMid34[1] , \wBMid34[0] }), .LoOut({\wAMid35[31] , \wAMid35[30] , 
        \wAMid35[29] , \wAMid35[28] , \wAMid35[27] , \wAMid35[26] , 
        \wAMid35[25] , \wAMid35[24] , \wAMid35[23] , \wAMid35[22] , 
        \wAMid35[21] , \wAMid35[20] , \wAMid35[19] , \wAMid35[18] , 
        \wAMid35[17] , \wAMid35[16] , \wAMid35[15] , \wAMid35[14] , 
        \wAMid35[13] , \wAMid35[12] , \wAMid35[11] , \wAMid35[10] , 
        \wAMid35[9] , \wAMid35[8] , \wAMid35[7] , \wAMid35[6] , \wAMid35[5] , 
        \wAMid35[4] , \wAMid35[3] , \wAMid35[2] , \wAMid35[1] , \wAMid35[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn40[31] , \wAIn40[30] , \wAIn40[29] , \wAIn40[28] , \wAIn40[27] , 
        \wAIn40[26] , \wAIn40[25] , \wAIn40[24] , \wAIn40[23] , \wAIn40[22] , 
        \wAIn40[21] , \wAIn40[20] , \wAIn40[19] , \wAIn40[18] , \wAIn40[17] , 
        \wAIn40[16] , \wAIn40[15] , \wAIn40[14] , \wAIn40[13] , \wAIn40[12] , 
        \wAIn40[11] , \wAIn40[10] , \wAIn40[9] , \wAIn40[8] , \wAIn40[7] , 
        \wAIn40[6] , \wAIn40[5] , \wAIn40[4] , \wAIn40[3] , \wAIn40[2] , 
        \wAIn40[1] , \wAIn40[0] }), .BIn({\wBIn40[31] , \wBIn40[30] , 
        \wBIn40[29] , \wBIn40[28] , \wBIn40[27] , \wBIn40[26] , \wBIn40[25] , 
        \wBIn40[24] , \wBIn40[23] , \wBIn40[22] , \wBIn40[21] , \wBIn40[20] , 
        \wBIn40[19] , \wBIn40[18] , \wBIn40[17] , \wBIn40[16] , \wBIn40[15] , 
        \wBIn40[14] , \wBIn40[13] , \wBIn40[12] , \wBIn40[11] , \wBIn40[10] , 
        \wBIn40[9] , \wBIn40[8] , \wBIn40[7] , \wBIn40[6] , \wBIn40[5] , 
        \wBIn40[4] , \wBIn40[3] , \wBIn40[2] , \wBIn40[1] , \wBIn40[0] }), 
        .HiOut({\wBMid39[31] , \wBMid39[30] , \wBMid39[29] , \wBMid39[28] , 
        \wBMid39[27] , \wBMid39[26] , \wBMid39[25] , \wBMid39[24] , 
        \wBMid39[23] , \wBMid39[22] , \wBMid39[21] , \wBMid39[20] , 
        \wBMid39[19] , \wBMid39[18] , \wBMid39[17] , \wBMid39[16] , 
        \wBMid39[15] , \wBMid39[14] , \wBMid39[13] , \wBMid39[12] , 
        \wBMid39[11] , \wBMid39[10] , \wBMid39[9] , \wBMid39[8] , \wBMid39[7] , 
        \wBMid39[6] , \wBMid39[5] , \wBMid39[4] , \wBMid39[3] , \wBMid39[2] , 
        \wBMid39[1] , \wBMid39[0] }), .LoOut({\wAMid40[31] , \wAMid40[30] , 
        \wAMid40[29] , \wAMid40[28] , \wAMid40[27] , \wAMid40[26] , 
        \wAMid40[25] , \wAMid40[24] , \wAMid40[23] , \wAMid40[22] , 
        \wAMid40[21] , \wAMid40[20] , \wAMid40[19] , \wAMid40[18] , 
        \wAMid40[17] , \wAMid40[16] , \wAMid40[15] , \wAMid40[14] , 
        \wAMid40[13] , \wAMid40[12] , \wAMid40[11] , \wAMid40[10] , 
        \wAMid40[9] , \wAMid40[8] , \wAMid40[7] , \wAMid40[6] , \wAMid40[5] , 
        \wAMid40[4] , \wAMid40[3] , \wAMid40[2] , \wAMid40[1] , \wAMid40[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid70[31] , \wAMid70[30] , \wAMid70[29] , \wAMid70[28] , 
        \wAMid70[27] , \wAMid70[26] , \wAMid70[25] , \wAMid70[24] , 
        \wAMid70[23] , \wAMid70[22] , \wAMid70[21] , \wAMid70[20] , 
        \wAMid70[19] , \wAMid70[18] , \wAMid70[17] , \wAMid70[16] , 
        \wAMid70[15] , \wAMid70[14] , \wAMid70[13] , \wAMid70[12] , 
        \wAMid70[11] , \wAMid70[10] , \wAMid70[9] , \wAMid70[8] , \wAMid70[7] , 
        \wAMid70[6] , \wAMid70[5] , \wAMid70[4] , \wAMid70[3] , \wAMid70[2] , 
        \wAMid70[1] , \wAMid70[0] }), .BIn({\wBMid70[31] , \wBMid70[30] , 
        \wBMid70[29] , \wBMid70[28] , \wBMid70[27] , \wBMid70[26] , 
        \wBMid70[25] , \wBMid70[24] , \wBMid70[23] , \wBMid70[22] , 
        \wBMid70[21] , \wBMid70[20] , \wBMid70[19] , \wBMid70[18] , 
        \wBMid70[17] , \wBMid70[16] , \wBMid70[15] , \wBMid70[14] , 
        \wBMid70[13] , \wBMid70[12] , \wBMid70[11] , \wBMid70[10] , 
        \wBMid70[9] , \wBMid70[8] , \wBMid70[7] , \wBMid70[6] , \wBMid70[5] , 
        \wBMid70[4] , \wBMid70[3] , \wBMid70[2] , \wBMid70[1] , \wBMid70[0] }), 
        .HiOut({\wRegInB70[31] , \wRegInB70[30] , \wRegInB70[29] , 
        \wRegInB70[28] , \wRegInB70[27] , \wRegInB70[26] , \wRegInB70[25] , 
        \wRegInB70[24] , \wRegInB70[23] , \wRegInB70[22] , \wRegInB70[21] , 
        \wRegInB70[20] , \wRegInB70[19] , \wRegInB70[18] , \wRegInB70[17] , 
        \wRegInB70[16] , \wRegInB70[15] , \wRegInB70[14] , \wRegInB70[13] , 
        \wRegInB70[12] , \wRegInB70[11] , \wRegInB70[10] , \wRegInB70[9] , 
        \wRegInB70[8] , \wRegInB70[7] , \wRegInB70[6] , \wRegInB70[5] , 
        \wRegInB70[4] , \wRegInB70[3] , \wRegInB70[2] , \wRegInB70[1] , 
        \wRegInB70[0] }), .LoOut({\wRegInA71[31] , \wRegInA71[30] , 
        \wRegInA71[29] , \wRegInA71[28] , \wRegInA71[27] , \wRegInA71[26] , 
        \wRegInA71[25] , \wRegInA71[24] , \wRegInA71[23] , \wRegInA71[22] , 
        \wRegInA71[21] , \wRegInA71[20] , \wRegInA71[19] , \wRegInA71[18] , 
        \wRegInA71[17] , \wRegInA71[16] , \wRegInA71[15] , \wRegInA71[14] , 
        \wRegInA71[13] , \wRegInA71[12] , \wRegInA71[11] , \wRegInA71[10] , 
        \wRegInA71[9] , \wRegInA71[8] , \wRegInA71[7] , \wRegInA71[6] , 
        \wRegInA71[5] , \wRegInA71[4] , \wRegInA71[3] , \wRegInA71[2] , 
        \wRegInA71[1] , \wRegInA71[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid95[31] , \wAMid95[30] , \wAMid95[29] , \wAMid95[28] , 
        \wAMid95[27] , \wAMid95[26] , \wAMid95[25] , \wAMid95[24] , 
        \wAMid95[23] , \wAMid95[22] , \wAMid95[21] , \wAMid95[20] , 
        \wAMid95[19] , \wAMid95[18] , \wAMid95[17] , \wAMid95[16] , 
        \wAMid95[15] , \wAMid95[14] , \wAMid95[13] , \wAMid95[12] , 
        \wAMid95[11] , \wAMid95[10] , \wAMid95[9] , \wAMid95[8] , \wAMid95[7] , 
        \wAMid95[6] , \wAMid95[5] , \wAMid95[4] , \wAMid95[3] , \wAMid95[2] , 
        \wAMid95[1] , \wAMid95[0] }), .BIn({\wBMid95[31] , \wBMid95[30] , 
        \wBMid95[29] , \wBMid95[28] , \wBMid95[27] , \wBMid95[26] , 
        \wBMid95[25] , \wBMid95[24] , \wBMid95[23] , \wBMid95[22] , 
        \wBMid95[21] , \wBMid95[20] , \wBMid95[19] , \wBMid95[18] , 
        \wBMid95[17] , \wBMid95[16] , \wBMid95[15] , \wBMid95[14] , 
        \wBMid95[13] , \wBMid95[12] , \wBMid95[11] , \wBMid95[10] , 
        \wBMid95[9] , \wBMid95[8] , \wBMid95[7] , \wBMid95[6] , \wBMid95[5] , 
        \wBMid95[4] , \wBMid95[3] , \wBMid95[2] , \wBMid95[1] , \wBMid95[0] }), 
        .HiOut({\wRegInB95[31] , \wRegInB95[30] , \wRegInB95[29] , 
        \wRegInB95[28] , \wRegInB95[27] , \wRegInB95[26] , \wRegInB95[25] , 
        \wRegInB95[24] , \wRegInB95[23] , \wRegInB95[22] , \wRegInB95[21] , 
        \wRegInB95[20] , \wRegInB95[19] , \wRegInB95[18] , \wRegInB95[17] , 
        \wRegInB95[16] , \wRegInB95[15] , \wRegInB95[14] , \wRegInB95[13] , 
        \wRegInB95[12] , \wRegInB95[11] , \wRegInB95[10] , \wRegInB95[9] , 
        \wRegInB95[8] , \wRegInB95[7] , \wRegInB95[6] , \wRegInB95[5] , 
        \wRegInB95[4] , \wRegInB95[3] , \wRegInB95[2] , \wRegInB95[1] , 
        \wRegInB95[0] }), .LoOut({\wRegInA96[31] , \wRegInA96[30] , 
        \wRegInA96[29] , \wRegInA96[28] , \wRegInA96[27] , \wRegInA96[26] , 
        \wRegInA96[25] , \wRegInA96[24] , \wRegInA96[23] , \wRegInA96[22] , 
        \wRegInA96[21] , \wRegInA96[20] , \wRegInA96[19] , \wRegInA96[18] , 
        \wRegInA96[17] , \wRegInA96[16] , \wRegInA96[15] , \wRegInA96[14] , 
        \wRegInA96[13] , \wRegInA96[12] , \wRegInA96[11] , \wRegInA96[10] , 
        \wRegInA96[9] , \wRegInA96[8] , \wRegInA96[7] , \wRegInA96[6] , 
        \wRegInA96[5] , \wRegInA96[4] , \wRegInA96[3] , \wRegInA96[2] , 
        \wRegInA96[1] , \wRegInA96[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_145 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink146[31] , \ScanLink146[30] , \ScanLink146[29] , 
        \ScanLink146[28] , \ScanLink146[27] , \ScanLink146[26] , 
        \ScanLink146[25] , \ScanLink146[24] , \ScanLink146[23] , 
        \ScanLink146[22] , \ScanLink146[21] , \ScanLink146[20] , 
        \ScanLink146[19] , \ScanLink146[18] , \ScanLink146[17] , 
        \ScanLink146[16] , \ScanLink146[15] , \ScanLink146[14] , 
        \ScanLink146[13] , \ScanLink146[12] , \ScanLink146[11] , 
        \ScanLink146[10] , \ScanLink146[9] , \ScanLink146[8] , 
        \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , \ScanLink146[4] , 
        \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , \ScanLink146[0] 
        }), .ScanOut({\ScanLink145[31] , \ScanLink145[30] , \ScanLink145[29] , 
        \ScanLink145[28] , \ScanLink145[27] , \ScanLink145[26] , 
        \ScanLink145[25] , \ScanLink145[24] , \ScanLink145[23] , 
        \ScanLink145[22] , \ScanLink145[21] , \ScanLink145[20] , 
        \ScanLink145[19] , \ScanLink145[18] , \ScanLink145[17] , 
        \ScanLink145[16] , \ScanLink145[15] , \ScanLink145[14] , 
        \ScanLink145[13] , \ScanLink145[12] , \ScanLink145[11] , 
        \ScanLink145[10] , \ScanLink145[9] , \ScanLink145[8] , 
        \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , \ScanLink145[4] , 
        \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , \ScanLink145[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA55[31] , \wRegInA55[30] , \wRegInA55[29] , 
        \wRegInA55[28] , \wRegInA55[27] , \wRegInA55[26] , \wRegInA55[25] , 
        \wRegInA55[24] , \wRegInA55[23] , \wRegInA55[22] , \wRegInA55[21] , 
        \wRegInA55[20] , \wRegInA55[19] , \wRegInA55[18] , \wRegInA55[17] , 
        \wRegInA55[16] , \wRegInA55[15] , \wRegInA55[14] , \wRegInA55[13] , 
        \wRegInA55[12] , \wRegInA55[11] , \wRegInA55[10] , \wRegInA55[9] , 
        \wRegInA55[8] , \wRegInA55[7] , \wRegInA55[6] , \wRegInA55[5] , 
        \wRegInA55[4] , \wRegInA55[3] , \wRegInA55[2] , \wRegInA55[1] , 
        \wRegInA55[0] }), .Out({\wAIn55[31] , \wAIn55[30] , \wAIn55[29] , 
        \wAIn55[28] , \wAIn55[27] , \wAIn55[26] , \wAIn55[25] , \wAIn55[24] , 
        \wAIn55[23] , \wAIn55[22] , \wAIn55[21] , \wAIn55[20] , \wAIn55[19] , 
        \wAIn55[18] , \wAIn55[17] , \wAIn55[16] , \wAIn55[15] , \wAIn55[14] , 
        \wAIn55[13] , \wAIn55[12] , \wAIn55[11] , \wAIn55[10] , \wAIn55[9] , 
        \wAIn55[8] , \wAIn55[7] , \wAIn55[6] , \wAIn55[5] , \wAIn55[4] , 
        \wAIn55[3] , \wAIn55[2] , \wAIn55[1] , \wAIn55[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_15 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[31] , \ScanLink16[30] , \ScanLink16[29] , 
        \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , \ScanLink16[25] , 
        \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , \ScanLink16[21] , 
        \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , \ScanLink16[17] , 
        \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , \ScanLink16[13] , 
        \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , \ScanLink16[9] , 
        \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA120[31] , \wRegInA120[30] , 
        \wRegInA120[29] , \wRegInA120[28] , \wRegInA120[27] , \wRegInA120[26] , 
        \wRegInA120[25] , \wRegInA120[24] , \wRegInA120[23] , \wRegInA120[22] , 
        \wRegInA120[21] , \wRegInA120[20] , \wRegInA120[19] , \wRegInA120[18] , 
        \wRegInA120[17] , \wRegInA120[16] , \wRegInA120[15] , \wRegInA120[14] , 
        \wRegInA120[13] , \wRegInA120[12] , \wRegInA120[11] , \wRegInA120[10] , 
        \wRegInA120[9] , \wRegInA120[8] , \wRegInA120[7] , \wRegInA120[6] , 
        \wRegInA120[5] , \wRegInA120[4] , \wRegInA120[3] , \wRegInA120[2] , 
        \wRegInA120[1] , \wRegInA120[0] }), .Out({\wAIn120[31] , \wAIn120[30] , 
        \wAIn120[29] , \wAIn120[28] , \wAIn120[27] , \wAIn120[26] , 
        \wAIn120[25] , \wAIn120[24] , \wAIn120[23] , \wAIn120[22] , 
        \wAIn120[21] , \wAIn120[20] , \wAIn120[19] , \wAIn120[18] , 
        \wAIn120[17] , \wAIn120[16] , \wAIn120[15] , \wAIn120[14] , 
        \wAIn120[13] , \wAIn120[12] , \wAIn120[11] , \wAIn120[10] , 
        \wAIn120[9] , \wAIn120[8] , \wAIn120[7] , \wAIn120[6] , \wAIn120[5] , 
        \wAIn120[4] , \wAIn120[3] , \wAIn120[2] , \wAIn120[1] , \wAIn120[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn67[31] , \wAIn67[30] , \wAIn67[29] , \wAIn67[28] , \wAIn67[27] , 
        \wAIn67[26] , \wAIn67[25] , \wAIn67[24] , \wAIn67[23] , \wAIn67[22] , 
        \wAIn67[21] , \wAIn67[20] , \wAIn67[19] , \wAIn67[18] , \wAIn67[17] , 
        \wAIn67[16] , \wAIn67[15] , \wAIn67[14] , \wAIn67[13] , \wAIn67[12] , 
        \wAIn67[11] , \wAIn67[10] , \wAIn67[9] , \wAIn67[8] , \wAIn67[7] , 
        \wAIn67[6] , \wAIn67[5] , \wAIn67[4] , \wAIn67[3] , \wAIn67[2] , 
        \wAIn67[1] , \wAIn67[0] }), .BIn({\wBIn67[31] , \wBIn67[30] , 
        \wBIn67[29] , \wBIn67[28] , \wBIn67[27] , \wBIn67[26] , \wBIn67[25] , 
        \wBIn67[24] , \wBIn67[23] , \wBIn67[22] , \wBIn67[21] , \wBIn67[20] , 
        \wBIn67[19] , \wBIn67[18] , \wBIn67[17] , \wBIn67[16] , \wBIn67[15] , 
        \wBIn67[14] , \wBIn67[13] , \wBIn67[12] , \wBIn67[11] , \wBIn67[10] , 
        \wBIn67[9] , \wBIn67[8] , \wBIn67[7] , \wBIn67[6] , \wBIn67[5] , 
        \wBIn67[4] , \wBIn67[3] , \wBIn67[2] , \wBIn67[1] , \wBIn67[0] }), 
        .HiOut({\wBMid66[31] , \wBMid66[30] , \wBMid66[29] , \wBMid66[28] , 
        \wBMid66[27] , \wBMid66[26] , \wBMid66[25] , \wBMid66[24] , 
        \wBMid66[23] , \wBMid66[22] , \wBMid66[21] , \wBMid66[20] , 
        \wBMid66[19] , \wBMid66[18] , \wBMid66[17] , \wBMid66[16] , 
        \wBMid66[15] , \wBMid66[14] , \wBMid66[13] , \wBMid66[12] , 
        \wBMid66[11] , \wBMid66[10] , \wBMid66[9] , \wBMid66[8] , \wBMid66[7] , 
        \wBMid66[6] , \wBMid66[5] , \wBMid66[4] , \wBMid66[3] , \wBMid66[2] , 
        \wBMid66[1] , \wBMid66[0] }), .LoOut({\wAMid67[31] , \wAMid67[30] , 
        \wAMid67[29] , \wAMid67[28] , \wAMid67[27] , \wAMid67[26] , 
        \wAMid67[25] , \wAMid67[24] , \wAMid67[23] , \wAMid67[22] , 
        \wAMid67[21] , \wAMid67[20] , \wAMid67[19] , \wAMid67[18] , 
        \wAMid67[17] , \wAMid67[16] , \wAMid67[15] , \wAMid67[14] , 
        \wAMid67[13] , \wAMid67[12] , \wAMid67[11] , \wAMid67[10] , 
        \wAMid67[9] , \wAMid67[8] , \wAMid67[7] , \wAMid67[6] , \wAMid67[5] , 
        \wAMid67[4] , \wAMid67[3] , \wAMid67[2] , \wAMid67[1] , \wAMid67[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn117[31] , \wAIn117[30] , \wAIn117[29] , \wAIn117[28] , 
        \wAIn117[27] , \wAIn117[26] , \wAIn117[25] , \wAIn117[24] , 
        \wAIn117[23] , \wAIn117[22] , \wAIn117[21] , \wAIn117[20] , 
        \wAIn117[19] , \wAIn117[18] , \wAIn117[17] , \wAIn117[16] , 
        \wAIn117[15] , \wAIn117[14] , \wAIn117[13] , \wAIn117[12] , 
        \wAIn117[11] , \wAIn117[10] , \wAIn117[9] , \wAIn117[8] , \wAIn117[7] , 
        \wAIn117[6] , \wAIn117[5] , \wAIn117[4] , \wAIn117[3] , \wAIn117[2] , 
        \wAIn117[1] , \wAIn117[0] }), .BIn({\wBIn117[31] , \wBIn117[30] , 
        \wBIn117[29] , \wBIn117[28] , \wBIn117[27] , \wBIn117[26] , 
        \wBIn117[25] , \wBIn117[24] , \wBIn117[23] , \wBIn117[22] , 
        \wBIn117[21] , \wBIn117[20] , \wBIn117[19] , \wBIn117[18] , 
        \wBIn117[17] , \wBIn117[16] , \wBIn117[15] , \wBIn117[14] , 
        \wBIn117[13] , \wBIn117[12] , \wBIn117[11] , \wBIn117[10] , 
        \wBIn117[9] , \wBIn117[8] , \wBIn117[7] , \wBIn117[6] , \wBIn117[5] , 
        \wBIn117[4] , \wBIn117[3] , \wBIn117[2] , \wBIn117[1] , \wBIn117[0] }), 
        .HiOut({\wBMid116[31] , \wBMid116[30] , \wBMid116[29] , \wBMid116[28] , 
        \wBMid116[27] , \wBMid116[26] , \wBMid116[25] , \wBMid116[24] , 
        \wBMid116[23] , \wBMid116[22] , \wBMid116[21] , \wBMid116[20] , 
        \wBMid116[19] , \wBMid116[18] , \wBMid116[17] , \wBMid116[16] , 
        \wBMid116[15] , \wBMid116[14] , \wBMid116[13] , \wBMid116[12] , 
        \wBMid116[11] , \wBMid116[10] , \wBMid116[9] , \wBMid116[8] , 
        \wBMid116[7] , \wBMid116[6] , \wBMid116[5] , \wBMid116[4] , 
        \wBMid116[3] , \wBMid116[2] , \wBMid116[1] , \wBMid116[0] }), .LoOut({
        \wAMid117[31] , \wAMid117[30] , \wAMid117[29] , \wAMid117[28] , 
        \wAMid117[27] , \wAMid117[26] , \wAMid117[25] , \wAMid117[24] , 
        \wAMid117[23] , \wAMid117[22] , \wAMid117[21] , \wAMid117[20] , 
        \wAMid117[19] , \wAMid117[18] , \wAMid117[17] , \wAMid117[16] , 
        \wAMid117[15] , \wAMid117[14] , \wAMid117[13] , \wAMid117[12] , 
        \wAMid117[11] , \wAMid117[10] , \wAMid117[9] , \wAMid117[8] , 
        \wAMid117[7] , \wAMid117[6] , \wAMid117[5] , \wAMid117[4] , 
        \wAMid117[3] , \wAMid117[2] , \wAMid117[1] , \wAMid117[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_252 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink253[31] , \ScanLink253[30] , \ScanLink253[29] , 
        \ScanLink253[28] , \ScanLink253[27] , \ScanLink253[26] , 
        \ScanLink253[25] , \ScanLink253[24] , \ScanLink253[23] , 
        \ScanLink253[22] , \ScanLink253[21] , \ScanLink253[20] , 
        \ScanLink253[19] , \ScanLink253[18] , \ScanLink253[17] , 
        \ScanLink253[16] , \ScanLink253[15] , \ScanLink253[14] , 
        \ScanLink253[13] , \ScanLink253[12] , \ScanLink253[11] , 
        \ScanLink253[10] , \ScanLink253[9] , \ScanLink253[8] , 
        \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , \ScanLink253[4] , 
        \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , \ScanLink253[0] 
        }), .ScanOut({\ScanLink252[31] , \ScanLink252[30] , \ScanLink252[29] , 
        \ScanLink252[28] , \ScanLink252[27] , \ScanLink252[26] , 
        \ScanLink252[25] , \ScanLink252[24] , \ScanLink252[23] , 
        \ScanLink252[22] , \ScanLink252[21] , \ScanLink252[20] , 
        \ScanLink252[19] , \ScanLink252[18] , \ScanLink252[17] , 
        \ScanLink252[16] , \ScanLink252[15] , \ScanLink252[14] , 
        \ScanLink252[13] , \ScanLink252[12] , \ScanLink252[11] , 
        \ScanLink252[10] , \ScanLink252[9] , \ScanLink252[8] , 
        \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , \ScanLink252[4] , 
        \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , \ScanLink252[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB1[31] , \wRegInB1[30] , \wRegInB1[29] , \wRegInB1[28] , 
        \wRegInB1[27] , \wRegInB1[26] , \wRegInB1[25] , \wRegInB1[24] , 
        \wRegInB1[23] , \wRegInB1[22] , \wRegInB1[21] , \wRegInB1[20] , 
        \wRegInB1[19] , \wRegInB1[18] , \wRegInB1[17] , \wRegInB1[16] , 
        \wRegInB1[15] , \wRegInB1[14] , \wRegInB1[13] , \wRegInB1[12] , 
        \wRegInB1[11] , \wRegInB1[10] , \wRegInB1[9] , \wRegInB1[8] , 
        \wRegInB1[7] , \wRegInB1[6] , \wRegInB1[5] , \wRegInB1[4] , 
        \wRegInB1[3] , \wRegInB1[2] , \wRegInB1[1] , \wRegInB1[0] }), .Out({
        \wBIn1[31] , \wBIn1[30] , \wBIn1[29] , \wBIn1[28] , \wBIn1[27] , 
        \wBIn1[26] , \wBIn1[25] , \wBIn1[24] , \wBIn1[23] , \wBIn1[22] , 
        \wBIn1[21] , \wBIn1[20] , \wBIn1[19] , \wBIn1[18] , \wBIn1[17] , 
        \wBIn1[16] , \wBIn1[15] , \wBIn1[14] , \wBIn1[13] , \wBIn1[12] , 
        \wBIn1[11] , \wBIn1[10] , \wBIn1[9] , \wBIn1[8] , \wBIn1[7] , 
        \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , \wBIn1[3] , \wBIn1[2] , \wBIn1[1] , 
        \wBIn1[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid57[31] , \wAMid57[30] , \wAMid57[29] , \wAMid57[28] , 
        \wAMid57[27] , \wAMid57[26] , \wAMid57[25] , \wAMid57[24] , 
        \wAMid57[23] , \wAMid57[22] , \wAMid57[21] , \wAMid57[20] , 
        \wAMid57[19] , \wAMid57[18] , \wAMid57[17] , \wAMid57[16] , 
        \wAMid57[15] , \wAMid57[14] , \wAMid57[13] , \wAMid57[12] , 
        \wAMid57[11] , \wAMid57[10] , \wAMid57[9] , \wAMid57[8] , \wAMid57[7] , 
        \wAMid57[6] , \wAMid57[5] , \wAMid57[4] , \wAMid57[3] , \wAMid57[2] , 
        \wAMid57[1] , \wAMid57[0] }), .BIn({\wBMid57[31] , \wBMid57[30] , 
        \wBMid57[29] , \wBMid57[28] , \wBMid57[27] , \wBMid57[26] , 
        \wBMid57[25] , \wBMid57[24] , \wBMid57[23] , \wBMid57[22] , 
        \wBMid57[21] , \wBMid57[20] , \wBMid57[19] , \wBMid57[18] , 
        \wBMid57[17] , \wBMid57[16] , \wBMid57[15] , \wBMid57[14] , 
        \wBMid57[13] , \wBMid57[12] , \wBMid57[11] , \wBMid57[10] , 
        \wBMid57[9] , \wBMid57[8] , \wBMid57[7] , \wBMid57[6] , \wBMid57[5] , 
        \wBMid57[4] , \wBMid57[3] , \wBMid57[2] , \wBMid57[1] , \wBMid57[0] }), 
        .HiOut({\wRegInB57[31] , \wRegInB57[30] , \wRegInB57[29] , 
        \wRegInB57[28] , \wRegInB57[27] , \wRegInB57[26] , \wRegInB57[25] , 
        \wRegInB57[24] , \wRegInB57[23] , \wRegInB57[22] , \wRegInB57[21] , 
        \wRegInB57[20] , \wRegInB57[19] , \wRegInB57[18] , \wRegInB57[17] , 
        \wRegInB57[16] , \wRegInB57[15] , \wRegInB57[14] , \wRegInB57[13] , 
        \wRegInB57[12] , \wRegInB57[11] , \wRegInB57[10] , \wRegInB57[9] , 
        \wRegInB57[8] , \wRegInB57[7] , \wRegInB57[6] , \wRegInB57[5] , 
        \wRegInB57[4] , \wRegInB57[3] , \wRegInB57[2] , \wRegInB57[1] , 
        \wRegInB57[0] }), .LoOut({\wRegInA58[31] , \wRegInA58[30] , 
        \wRegInA58[29] , \wRegInA58[28] , \wRegInA58[27] , \wRegInA58[26] , 
        \wRegInA58[25] , \wRegInA58[24] , \wRegInA58[23] , \wRegInA58[22] , 
        \wRegInA58[21] , \wRegInA58[20] , \wRegInA58[19] , \wRegInA58[18] , 
        \wRegInA58[17] , \wRegInA58[16] , \wRegInA58[15] , \wRegInA58[14] , 
        \wRegInA58[13] , \wRegInA58[12] , \wRegInA58[11] , \wRegInA58[10] , 
        \wRegInA58[9] , \wRegInA58[8] , \wRegInA58[7] , \wRegInA58[6] , 
        \wRegInA58[5] , \wRegInA58[4] , \wRegInA58[3] , \wRegInA58[2] , 
        \wRegInA58[1] , \wRegInA58[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_162 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink163[31] , \ScanLink163[30] , \ScanLink163[29] , 
        \ScanLink163[28] , \ScanLink163[27] , \ScanLink163[26] , 
        \ScanLink163[25] , \ScanLink163[24] , \ScanLink163[23] , 
        \ScanLink163[22] , \ScanLink163[21] , \ScanLink163[20] , 
        \ScanLink163[19] , \ScanLink163[18] , \ScanLink163[17] , 
        \ScanLink163[16] , \ScanLink163[15] , \ScanLink163[14] , 
        \ScanLink163[13] , \ScanLink163[12] , \ScanLink163[11] , 
        \ScanLink163[10] , \ScanLink163[9] , \ScanLink163[8] , 
        \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , \ScanLink163[4] , 
        \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , \ScanLink163[0] 
        }), .ScanOut({\ScanLink162[31] , \ScanLink162[30] , \ScanLink162[29] , 
        \ScanLink162[28] , \ScanLink162[27] , \ScanLink162[26] , 
        \ScanLink162[25] , \ScanLink162[24] , \ScanLink162[23] , 
        \ScanLink162[22] , \ScanLink162[21] , \ScanLink162[20] , 
        \ScanLink162[19] , \ScanLink162[18] , \ScanLink162[17] , 
        \ScanLink162[16] , \ScanLink162[15] , \ScanLink162[14] , 
        \ScanLink162[13] , \ScanLink162[12] , \ScanLink162[11] , 
        \ScanLink162[10] , \ScanLink162[9] , \ScanLink162[8] , 
        \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , \ScanLink162[4] , 
        \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , \ScanLink162[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB46[31] , \wRegInB46[30] , \wRegInB46[29] , 
        \wRegInB46[28] , \wRegInB46[27] , \wRegInB46[26] , \wRegInB46[25] , 
        \wRegInB46[24] , \wRegInB46[23] , \wRegInB46[22] , \wRegInB46[21] , 
        \wRegInB46[20] , \wRegInB46[19] , \wRegInB46[18] , \wRegInB46[17] , 
        \wRegInB46[16] , \wRegInB46[15] , \wRegInB46[14] , \wRegInB46[13] , 
        \wRegInB46[12] , \wRegInB46[11] , \wRegInB46[10] , \wRegInB46[9] , 
        \wRegInB46[8] , \wRegInB46[7] , \wRegInB46[6] , \wRegInB46[5] , 
        \wRegInB46[4] , \wRegInB46[3] , \wRegInB46[2] , \wRegInB46[1] , 
        \wRegInB46[0] }), .Out({\wBIn46[31] , \wBIn46[30] , \wBIn46[29] , 
        \wBIn46[28] , \wBIn46[27] , \wBIn46[26] , \wBIn46[25] , \wBIn46[24] , 
        \wBIn46[23] , \wBIn46[22] , \wBIn46[21] , \wBIn46[20] , \wBIn46[19] , 
        \wBIn46[18] , \wBIn46[17] , \wBIn46[16] , \wBIn46[15] , \wBIn46[14] , 
        \wBIn46[13] , \wBIn46[12] , \wBIn46[11] , \wBIn46[10] , \wBIn46[9] , 
        \wBIn46[8] , \wBIn46[7] , \wBIn46[6] , \wBIn46[5] , \wBIn46[4] , 
        \wBIn46[3] , \wBIn46[2] , \wBIn46[1] , \wBIn46[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_32 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink33[31] , \ScanLink33[30] , \ScanLink33[29] , 
        \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , \ScanLink33[25] , 
        \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , \ScanLink33[21] , 
        \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , \ScanLink33[17] , 
        \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , \ScanLink33[13] , 
        \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , \ScanLink33[9] , 
        \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , \ScanLink33[5] , 
        \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , \ScanLink33[1] , 
        \ScanLink33[0] }), .ScanOut({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB111[31] , \wRegInB111[30] , 
        \wRegInB111[29] , \wRegInB111[28] , \wRegInB111[27] , \wRegInB111[26] , 
        \wRegInB111[25] , \wRegInB111[24] , \wRegInB111[23] , \wRegInB111[22] , 
        \wRegInB111[21] , \wRegInB111[20] , \wRegInB111[19] , \wRegInB111[18] , 
        \wRegInB111[17] , \wRegInB111[16] , \wRegInB111[15] , \wRegInB111[14] , 
        \wRegInB111[13] , \wRegInB111[12] , \wRegInB111[11] , \wRegInB111[10] , 
        \wRegInB111[9] , \wRegInB111[8] , \wRegInB111[7] , \wRegInB111[6] , 
        \wRegInB111[5] , \wRegInB111[4] , \wRegInB111[3] , \wRegInB111[2] , 
        \wRegInB111[1] , \wRegInB111[0] }), .Out({\wBIn111[31] , \wBIn111[30] , 
        \wBIn111[29] , \wBIn111[28] , \wBIn111[27] , \wBIn111[26] , 
        \wBIn111[25] , \wBIn111[24] , \wBIn111[23] , \wBIn111[22] , 
        \wBIn111[21] , \wBIn111[20] , \wBIn111[19] , \wBIn111[18] , 
        \wBIn111[17] , \wBIn111[16] , \wBIn111[15] , \wBIn111[14] , 
        \wBIn111[13] , \wBIn111[12] , \wBIn111[11] , \wBIn111[10] , 
        \wBIn111[9] , \wBIn111[8] , \wBIn111[7] , \wBIn111[6] , \wBIn111[5] , 
        \wBIn111[4] , \wBIn111[3] , \wBIn111[2] , \wBIn111[1] , \wBIn111[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn99[31] , \wAIn99[30] , \wAIn99[29] , \wAIn99[28] , \wAIn99[27] , 
        \wAIn99[26] , \wAIn99[25] , \wAIn99[24] , \wAIn99[23] , \wAIn99[22] , 
        \wAIn99[21] , \wAIn99[20] , \wAIn99[19] , \wAIn99[18] , \wAIn99[17] , 
        \wAIn99[16] , \wAIn99[15] , \wAIn99[14] , \wAIn99[13] , \wAIn99[12] , 
        \wAIn99[11] , \wAIn99[10] , \wAIn99[9] , \wAIn99[8] , \wAIn99[7] , 
        \wAIn99[6] , \wAIn99[5] , \wAIn99[4] , \wAIn99[3] , \wAIn99[2] , 
        \wAIn99[1] , \wAIn99[0] }), .BIn({\wBIn99[31] , \wBIn99[30] , 
        \wBIn99[29] , \wBIn99[28] , \wBIn99[27] , \wBIn99[26] , \wBIn99[25] , 
        \wBIn99[24] , \wBIn99[23] , \wBIn99[22] , \wBIn99[21] , \wBIn99[20] , 
        \wBIn99[19] , \wBIn99[18] , \wBIn99[17] , \wBIn99[16] , \wBIn99[15] , 
        \wBIn99[14] , \wBIn99[13] , \wBIn99[12] , \wBIn99[11] , \wBIn99[10] , 
        \wBIn99[9] , \wBIn99[8] , \wBIn99[7] , \wBIn99[6] , \wBIn99[5] , 
        \wBIn99[4] , \wBIn99[3] , \wBIn99[2] , \wBIn99[1] , \wBIn99[0] }), 
        .HiOut({\wBMid98[31] , \wBMid98[30] , \wBMid98[29] , \wBMid98[28] , 
        \wBMid98[27] , \wBMid98[26] , \wBMid98[25] , \wBMid98[24] , 
        \wBMid98[23] , \wBMid98[22] , \wBMid98[21] , \wBMid98[20] , 
        \wBMid98[19] , \wBMid98[18] , \wBMid98[17] , \wBMid98[16] , 
        \wBMid98[15] , \wBMid98[14] , \wBMid98[13] , \wBMid98[12] , 
        \wBMid98[11] , \wBMid98[10] , \wBMid98[9] , \wBMid98[8] , \wBMid98[7] , 
        \wBMid98[6] , \wBMid98[5] , \wBMid98[4] , \wBMid98[3] , \wBMid98[2] , 
        \wBMid98[1] , \wBMid98[0] }), .LoOut({\wAMid99[31] , \wAMid99[30] , 
        \wAMid99[29] , \wAMid99[28] , \wAMid99[27] , \wAMid99[26] , 
        \wAMid99[25] , \wAMid99[24] , \wAMid99[23] , \wAMid99[22] , 
        \wAMid99[21] , \wAMid99[20] , \wAMid99[19] , \wAMid99[18] , 
        \wAMid99[17] , \wAMid99[16] , \wAMid99[15] , \wAMid99[14] , 
        \wAMid99[13] , \wAMid99[12] , \wAMid99[11] , \wAMid99[10] , 
        \wAMid99[9] , \wAMid99[8] , \wAMid99[7] , \wAMid99[6] , \wAMid99[5] , 
        \wAMid99[4] , \wAMid99[3] , \wAMid99[2] , \wAMid99[1] , \wAMid99[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid106[31] , \wAMid106[30] , \wAMid106[29] , \wAMid106[28] , 
        \wAMid106[27] , \wAMid106[26] , \wAMid106[25] , \wAMid106[24] , 
        \wAMid106[23] , \wAMid106[22] , \wAMid106[21] , \wAMid106[20] , 
        \wAMid106[19] , \wAMid106[18] , \wAMid106[17] , \wAMid106[16] , 
        \wAMid106[15] , \wAMid106[14] , \wAMid106[13] , \wAMid106[12] , 
        \wAMid106[11] , \wAMid106[10] , \wAMid106[9] , \wAMid106[8] , 
        \wAMid106[7] , \wAMid106[6] , \wAMid106[5] , \wAMid106[4] , 
        \wAMid106[3] , \wAMid106[2] , \wAMid106[1] , \wAMid106[0] }), .BIn({
        \wBMid106[31] , \wBMid106[30] , \wBMid106[29] , \wBMid106[28] , 
        \wBMid106[27] , \wBMid106[26] , \wBMid106[25] , \wBMid106[24] , 
        \wBMid106[23] , \wBMid106[22] , \wBMid106[21] , \wBMid106[20] , 
        \wBMid106[19] , \wBMid106[18] , \wBMid106[17] , \wBMid106[16] , 
        \wBMid106[15] , \wBMid106[14] , \wBMid106[13] , \wBMid106[12] , 
        \wBMid106[11] , \wBMid106[10] , \wBMid106[9] , \wBMid106[8] , 
        \wBMid106[7] , \wBMid106[6] , \wBMid106[5] , \wBMid106[4] , 
        \wBMid106[3] , \wBMid106[2] , \wBMid106[1] , \wBMid106[0] }), .HiOut({
        \wRegInB106[31] , \wRegInB106[30] , \wRegInB106[29] , \wRegInB106[28] , 
        \wRegInB106[27] , \wRegInB106[26] , \wRegInB106[25] , \wRegInB106[24] , 
        \wRegInB106[23] , \wRegInB106[22] , \wRegInB106[21] , \wRegInB106[20] , 
        \wRegInB106[19] , \wRegInB106[18] , \wRegInB106[17] , \wRegInB106[16] , 
        \wRegInB106[15] , \wRegInB106[14] , \wRegInB106[13] , \wRegInB106[12] , 
        \wRegInB106[11] , \wRegInB106[10] , \wRegInB106[9] , \wRegInB106[8] , 
        \wRegInB106[7] , \wRegInB106[6] , \wRegInB106[5] , \wRegInB106[4] , 
        \wRegInB106[3] , \wRegInB106[2] , \wRegInB106[1] , \wRegInB106[0] }), 
        .LoOut({\wRegInA107[31] , \wRegInA107[30] , \wRegInA107[29] , 
        \wRegInA107[28] , \wRegInA107[27] , \wRegInA107[26] , \wRegInA107[25] , 
        \wRegInA107[24] , \wRegInA107[23] , \wRegInA107[22] , \wRegInA107[21] , 
        \wRegInA107[20] , \wRegInA107[19] , \wRegInA107[18] , \wRegInA107[17] , 
        \wRegInA107[16] , \wRegInA107[15] , \wRegInA107[14] , \wRegInA107[13] , 
        \wRegInA107[12] , \wRegInA107[11] , \wRegInA107[10] , \wRegInA107[9] , 
        \wRegInA107[8] , \wRegInA107[7] , \wRegInA107[6] , \wRegInA107[5] , 
        \wRegInA107[4] , \wRegInA107[3] , \wRegInA107[2] , \wRegInA107[1] , 
        \wRegInA107[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid121[31] , \wAMid121[30] , \wAMid121[29] , \wAMid121[28] , 
        \wAMid121[27] , \wAMid121[26] , \wAMid121[25] , \wAMid121[24] , 
        \wAMid121[23] , \wAMid121[22] , \wAMid121[21] , \wAMid121[20] , 
        \wAMid121[19] , \wAMid121[18] , \wAMid121[17] , \wAMid121[16] , 
        \wAMid121[15] , \wAMid121[14] , \wAMid121[13] , \wAMid121[12] , 
        \wAMid121[11] , \wAMid121[10] , \wAMid121[9] , \wAMid121[8] , 
        \wAMid121[7] , \wAMid121[6] , \wAMid121[5] , \wAMid121[4] , 
        \wAMid121[3] , \wAMid121[2] , \wAMid121[1] , \wAMid121[0] }), .BIn({
        \wBMid121[31] , \wBMid121[30] , \wBMid121[29] , \wBMid121[28] , 
        \wBMid121[27] , \wBMid121[26] , \wBMid121[25] , \wBMid121[24] , 
        \wBMid121[23] , \wBMid121[22] , \wBMid121[21] , \wBMid121[20] , 
        \wBMid121[19] , \wBMid121[18] , \wBMid121[17] , \wBMid121[16] , 
        \wBMid121[15] , \wBMid121[14] , \wBMid121[13] , \wBMid121[12] , 
        \wBMid121[11] , \wBMid121[10] , \wBMid121[9] , \wBMid121[8] , 
        \wBMid121[7] , \wBMid121[6] , \wBMid121[5] , \wBMid121[4] , 
        \wBMid121[3] , \wBMid121[2] , \wBMid121[1] , \wBMid121[0] }), .HiOut({
        \wRegInB121[31] , \wRegInB121[30] , \wRegInB121[29] , \wRegInB121[28] , 
        \wRegInB121[27] , \wRegInB121[26] , \wRegInB121[25] , \wRegInB121[24] , 
        \wRegInB121[23] , \wRegInB121[22] , \wRegInB121[21] , \wRegInB121[20] , 
        \wRegInB121[19] , \wRegInB121[18] , \wRegInB121[17] , \wRegInB121[16] , 
        \wRegInB121[15] , \wRegInB121[14] , \wRegInB121[13] , \wRegInB121[12] , 
        \wRegInB121[11] , \wRegInB121[10] , \wRegInB121[9] , \wRegInB121[8] , 
        \wRegInB121[7] , \wRegInB121[6] , \wRegInB121[5] , \wRegInB121[4] , 
        \wRegInB121[3] , \wRegInB121[2] , \wRegInB121[1] , \wRegInB121[0] }), 
        .LoOut({\wRegInA122[31] , \wRegInA122[30] , \wRegInA122[29] , 
        \wRegInA122[28] , \wRegInA122[27] , \wRegInA122[26] , \wRegInA122[25] , 
        \wRegInA122[24] , \wRegInA122[23] , \wRegInA122[22] , \wRegInA122[21] , 
        \wRegInA122[20] , \wRegInA122[19] , \wRegInA122[18] , \wRegInA122[17] , 
        \wRegInA122[16] , \wRegInA122[15] , \wRegInA122[14] , \wRegInA122[13] , 
        \wRegInA122[12] , \wRegInA122[11] , \wRegInA122[10] , \wRegInA122[9] , 
        \wRegInA122[8] , \wRegInA122[7] , \wRegInA122[6] , \wRegInA122[5] , 
        \wRegInA122[4] , \wRegInA122[3] , \wRegInA122[2] , \wRegInA122[1] , 
        \wRegInA122[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_249 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink250[31] , \ScanLink250[30] , \ScanLink250[29] , 
        \ScanLink250[28] , \ScanLink250[27] , \ScanLink250[26] , 
        \ScanLink250[25] , \ScanLink250[24] , \ScanLink250[23] , 
        \ScanLink250[22] , \ScanLink250[21] , \ScanLink250[20] , 
        \ScanLink250[19] , \ScanLink250[18] , \ScanLink250[17] , 
        \ScanLink250[16] , \ScanLink250[15] , \ScanLink250[14] , 
        \ScanLink250[13] , \ScanLink250[12] , \ScanLink250[11] , 
        \ScanLink250[10] , \ScanLink250[9] , \ScanLink250[8] , 
        \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , \ScanLink250[4] , 
        \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , \ScanLink250[0] 
        }), .ScanOut({\ScanLink249[31] , \ScanLink249[30] , \ScanLink249[29] , 
        \ScanLink249[28] , \ScanLink249[27] , \ScanLink249[26] , 
        \ScanLink249[25] , \ScanLink249[24] , \ScanLink249[23] , 
        \ScanLink249[22] , \ScanLink249[21] , \ScanLink249[20] , 
        \ScanLink249[19] , \ScanLink249[18] , \ScanLink249[17] , 
        \ScanLink249[16] , \ScanLink249[15] , \ScanLink249[14] , 
        \ScanLink249[13] , \ScanLink249[12] , \ScanLink249[11] , 
        \ScanLink249[10] , \ScanLink249[9] , \ScanLink249[8] , 
        \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , \ScanLink249[4] , 
        \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , \ScanLink249[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA3[31] , \wRegInA3[30] , \wRegInA3[29] , \wRegInA3[28] , 
        \wRegInA3[27] , \wRegInA3[26] , \wRegInA3[25] , \wRegInA3[24] , 
        \wRegInA3[23] , \wRegInA3[22] , \wRegInA3[21] , \wRegInA3[20] , 
        \wRegInA3[19] , \wRegInA3[18] , \wRegInA3[17] , \wRegInA3[16] , 
        \wRegInA3[15] , \wRegInA3[14] , \wRegInA3[13] , \wRegInA3[12] , 
        \wRegInA3[11] , \wRegInA3[10] , \wRegInA3[9] , \wRegInA3[8] , 
        \wRegInA3[7] , \wRegInA3[6] , \wRegInA3[5] , \wRegInA3[4] , 
        \wRegInA3[3] , \wRegInA3[2] , \wRegInA3[1] , \wRegInA3[0] }), .Out({
        \wAIn3[31] , \wAIn3[30] , \wAIn3[29] , \wAIn3[28] , \wAIn3[27] , 
        \wAIn3[26] , \wAIn3[25] , \wAIn3[24] , \wAIn3[23] , \wAIn3[22] , 
        \wAIn3[21] , \wAIn3[20] , \wAIn3[19] , \wAIn3[18] , \wAIn3[17] , 
        \wAIn3[16] , \wAIn3[15] , \wAIn3[14] , \wAIn3[13] , \wAIn3[12] , 
        \wAIn3[11] , \wAIn3[10] , \wAIn3[9] , \wAIn3[8] , \wAIn3[7] , 
        \wAIn3[6] , \wAIn3[5] , \wAIn3[4] , \wAIn3[3] , \wAIn3[2] , \wAIn3[1] , 
        \wAIn3[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_179 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink180[31] , \ScanLink180[30] , \ScanLink180[29] , 
        \ScanLink180[28] , \ScanLink180[27] , \ScanLink180[26] , 
        \ScanLink180[25] , \ScanLink180[24] , \ScanLink180[23] , 
        \ScanLink180[22] , \ScanLink180[21] , \ScanLink180[20] , 
        \ScanLink180[19] , \ScanLink180[18] , \ScanLink180[17] , 
        \ScanLink180[16] , \ScanLink180[15] , \ScanLink180[14] , 
        \ScanLink180[13] , \ScanLink180[12] , \ScanLink180[11] , 
        \ScanLink180[10] , \ScanLink180[9] , \ScanLink180[8] , 
        \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , \ScanLink180[4] , 
        \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , \ScanLink180[0] 
        }), .ScanOut({\ScanLink179[31] , \ScanLink179[30] , \ScanLink179[29] , 
        \ScanLink179[28] , \ScanLink179[27] , \ScanLink179[26] , 
        \ScanLink179[25] , \ScanLink179[24] , \ScanLink179[23] , 
        \ScanLink179[22] , \ScanLink179[21] , \ScanLink179[20] , 
        \ScanLink179[19] , \ScanLink179[18] , \ScanLink179[17] , 
        \ScanLink179[16] , \ScanLink179[15] , \ScanLink179[14] , 
        \ScanLink179[13] , \ScanLink179[12] , \ScanLink179[11] , 
        \ScanLink179[10] , \ScanLink179[9] , \ScanLink179[8] , 
        \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , \ScanLink179[4] , 
        \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , \ScanLink179[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA38[31] , \wRegInA38[30] , \wRegInA38[29] , 
        \wRegInA38[28] , \wRegInA38[27] , \wRegInA38[26] , \wRegInA38[25] , 
        \wRegInA38[24] , \wRegInA38[23] , \wRegInA38[22] , \wRegInA38[21] , 
        \wRegInA38[20] , \wRegInA38[19] , \wRegInA38[18] , \wRegInA38[17] , 
        \wRegInA38[16] , \wRegInA38[15] , \wRegInA38[14] , \wRegInA38[13] , 
        \wRegInA38[12] , \wRegInA38[11] , \wRegInA38[10] , \wRegInA38[9] , 
        \wRegInA38[8] , \wRegInA38[7] , \wRegInA38[6] , \wRegInA38[5] , 
        \wRegInA38[4] , \wRegInA38[3] , \wRegInA38[2] , \wRegInA38[1] , 
        \wRegInA38[0] }), .Out({\wAIn38[31] , \wAIn38[30] , \wAIn38[29] , 
        \wAIn38[28] , \wAIn38[27] , \wAIn38[26] , \wAIn38[25] , \wAIn38[24] , 
        \wAIn38[23] , \wAIn38[22] , \wAIn38[21] , \wAIn38[20] , \wAIn38[19] , 
        \wAIn38[18] , \wAIn38[17] , \wAIn38[16] , \wAIn38[15] , \wAIn38[14] , 
        \wAIn38[13] , \wAIn38[12] , \wAIn38[11] , \wAIn38[10] , \wAIn38[9] , 
        \wAIn38[8] , \wAIn38[7] , \wAIn38[6] , \wAIn38[5] , \wAIn38[4] , 
        \wAIn38[3] , \wAIn38[2] , \wAIn38[1] , \wAIn38[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_29 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink30[31] , \ScanLink30[30] , \ScanLink30[29] , 
        \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , \ScanLink30[25] , 
        \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , \ScanLink30[21] , 
        \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , \ScanLink30[17] , 
        \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , \ScanLink30[13] , 
        \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , \ScanLink30[9] , 
        \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , \ScanLink30[5] , 
        \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , \ScanLink30[1] , 
        \ScanLink30[0] }), .ScanOut({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA113[31] , \wRegInA113[30] , 
        \wRegInA113[29] , \wRegInA113[28] , \wRegInA113[27] , \wRegInA113[26] , 
        \wRegInA113[25] , \wRegInA113[24] , \wRegInA113[23] , \wRegInA113[22] , 
        \wRegInA113[21] , \wRegInA113[20] , \wRegInA113[19] , \wRegInA113[18] , 
        \wRegInA113[17] , \wRegInA113[16] , \wRegInA113[15] , \wRegInA113[14] , 
        \wRegInA113[13] , \wRegInA113[12] , \wRegInA113[11] , \wRegInA113[10] , 
        \wRegInA113[9] , \wRegInA113[8] , \wRegInA113[7] , \wRegInA113[6] , 
        \wRegInA113[5] , \wRegInA113[4] , \wRegInA113[3] , \wRegInA113[2] , 
        \wRegInA113[1] , \wRegInA113[0] }), .Out({\wAIn113[31] , \wAIn113[30] , 
        \wAIn113[29] , \wAIn113[28] , \wAIn113[27] , \wAIn113[26] , 
        \wAIn113[25] , \wAIn113[24] , \wAIn113[23] , \wAIn113[22] , 
        \wAIn113[21] , \wAIn113[20] , \wAIn113[19] , \wAIn113[18] , 
        \wAIn113[17] , \wAIn113[16] , \wAIn113[15] , \wAIn113[14] , 
        \wAIn113[13] , \wAIn113[12] , \wAIn113[11] , \wAIn113[10] , 
        \wAIn113[9] , \wAIn113[8] , \wAIn113[7] , \wAIn113[6] , \wAIn113[5] , 
        \wAIn113[4] , \wAIn113[3] , \wAIn113[2] , \wAIn113[1] , \wAIn113[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_85 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink86[31] , \ScanLink86[30] , \ScanLink86[29] , 
        \ScanLink86[28] , \ScanLink86[27] , \ScanLink86[26] , \ScanLink86[25] , 
        \ScanLink86[24] , \ScanLink86[23] , \ScanLink86[22] , \ScanLink86[21] , 
        \ScanLink86[20] , \ScanLink86[19] , \ScanLink86[18] , \ScanLink86[17] , 
        \ScanLink86[16] , \ScanLink86[15] , \ScanLink86[14] , \ScanLink86[13] , 
        \ScanLink86[12] , \ScanLink86[11] , \ScanLink86[10] , \ScanLink86[9] , 
        \ScanLink86[8] , \ScanLink86[7] , \ScanLink86[6] , \ScanLink86[5] , 
        \ScanLink86[4] , \ScanLink86[3] , \ScanLink86[2] , \ScanLink86[1] , 
        \ScanLink86[0] }), .ScanOut({\ScanLink85[31] , \ScanLink85[30] , 
        \ScanLink85[29] , \ScanLink85[28] , \ScanLink85[27] , \ScanLink85[26] , 
        \ScanLink85[25] , \ScanLink85[24] , \ScanLink85[23] , \ScanLink85[22] , 
        \ScanLink85[21] , \ScanLink85[20] , \ScanLink85[19] , \ScanLink85[18] , 
        \ScanLink85[17] , \ScanLink85[16] , \ScanLink85[15] , \ScanLink85[14] , 
        \ScanLink85[13] , \ScanLink85[12] , \ScanLink85[11] , \ScanLink85[10] , 
        \ScanLink85[9] , \ScanLink85[8] , \ScanLink85[7] , \ScanLink85[6] , 
        \ScanLink85[5] , \ScanLink85[4] , \ScanLink85[3] , \ScanLink85[2] , 
        \ScanLink85[1] , \ScanLink85[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA85[31] , \wRegInA85[30] , 
        \wRegInA85[29] , \wRegInA85[28] , \wRegInA85[27] , \wRegInA85[26] , 
        \wRegInA85[25] , \wRegInA85[24] , \wRegInA85[23] , \wRegInA85[22] , 
        \wRegInA85[21] , \wRegInA85[20] , \wRegInA85[19] , \wRegInA85[18] , 
        \wRegInA85[17] , \wRegInA85[16] , \wRegInA85[15] , \wRegInA85[14] , 
        \wRegInA85[13] , \wRegInA85[12] , \wRegInA85[11] , \wRegInA85[10] , 
        \wRegInA85[9] , \wRegInA85[8] , \wRegInA85[7] , \wRegInA85[6] , 
        \wRegInA85[5] , \wRegInA85[4] , \wRegInA85[3] , \wRegInA85[2] , 
        \wRegInA85[1] , \wRegInA85[0] }), .Out({\wAIn85[31] , \wAIn85[30] , 
        \wAIn85[29] , \wAIn85[28] , \wAIn85[27] , \wAIn85[26] , \wAIn85[25] , 
        \wAIn85[24] , \wAIn85[23] , \wAIn85[22] , \wAIn85[21] , \wAIn85[20] , 
        \wAIn85[19] , \wAIn85[18] , \wAIn85[17] , \wAIn85[16] , \wAIn85[15] , 
        \wAIn85[14] , \wAIn85[13] , \wAIn85[12] , \wAIn85[11] , \wAIn85[10] , 
        \wAIn85[9] , \wAIn85[8] , \wAIn85[7] , \wAIn85[6] , \wAIn85[5] , 
        \wAIn85[4] , \wAIn85[3] , \wAIn85[2] , \wAIn85[1] , \wAIn85[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid8[31] , 
        \wAMid8[30] , \wAMid8[29] , \wAMid8[28] , \wAMid8[27] , \wAMid8[26] , 
        \wAMid8[25] , \wAMid8[24] , \wAMid8[23] , \wAMid8[22] , \wAMid8[21] , 
        \wAMid8[20] , \wAMid8[19] , \wAMid8[18] , \wAMid8[17] , \wAMid8[16] , 
        \wAMid8[15] , \wAMid8[14] , \wAMid8[13] , \wAMid8[12] , \wAMid8[11] , 
        \wAMid8[10] , \wAMid8[9] , \wAMid8[8] , \wAMid8[7] , \wAMid8[6] , 
        \wAMid8[5] , \wAMid8[4] , \wAMid8[3] , \wAMid8[2] , \wAMid8[1] , 
        \wAMid8[0] }), .BIn({\wBMid8[31] , \wBMid8[30] , \wBMid8[29] , 
        \wBMid8[28] , \wBMid8[27] , \wBMid8[26] , \wBMid8[25] , \wBMid8[24] , 
        \wBMid8[23] , \wBMid8[22] , \wBMid8[21] , \wBMid8[20] , \wBMid8[19] , 
        \wBMid8[18] , \wBMid8[17] , \wBMid8[16] , \wBMid8[15] , \wBMid8[14] , 
        \wBMid8[13] , \wBMid8[12] , \wBMid8[11] , \wBMid8[10] , \wBMid8[9] , 
        \wBMid8[8] , \wBMid8[7] , \wBMid8[6] , \wBMid8[5] , \wBMid8[4] , 
        \wBMid8[3] , \wBMid8[2] , \wBMid8[1] , \wBMid8[0] }), .HiOut({
        \wRegInB8[31] , \wRegInB8[30] , \wRegInB8[29] , \wRegInB8[28] , 
        \wRegInB8[27] , \wRegInB8[26] , \wRegInB8[25] , \wRegInB8[24] , 
        \wRegInB8[23] , \wRegInB8[22] , \wRegInB8[21] , \wRegInB8[20] , 
        \wRegInB8[19] , \wRegInB8[18] , \wRegInB8[17] , \wRegInB8[16] , 
        \wRegInB8[15] , \wRegInB8[14] , \wRegInB8[13] , \wRegInB8[12] , 
        \wRegInB8[11] , \wRegInB8[10] , \wRegInB8[9] , \wRegInB8[8] , 
        \wRegInB8[7] , \wRegInB8[6] , \wRegInB8[5] , \wRegInB8[4] , 
        \wRegInB8[3] , \wRegInB8[2] , \wRegInB8[1] , \wRegInB8[0] }), .LoOut({
        \wRegInA9[31] , \wRegInA9[30] , \wRegInA9[29] , \wRegInA9[28] , 
        \wRegInA9[27] , \wRegInA9[26] , \wRegInA9[25] , \wRegInA9[24] , 
        \wRegInA9[23] , \wRegInA9[22] , \wRegInA9[21] , \wRegInA9[20] , 
        \wRegInA9[19] , \wRegInA9[18] , \wRegInA9[17] , \wRegInA9[16] , 
        \wRegInA9[15] , \wRegInA9[14] , \wRegInA9[13] , \wRegInA9[12] , 
        \wRegInA9[11] , \wRegInA9[10] , \wRegInA9[9] , \wRegInA9[8] , 
        \wRegInA9[7] , \wRegInA9[6] , \wRegInA9[5] , \wRegInA9[4] , 
        \wRegInA9[3] , \wRegInA9[2] , \wRegInA9[1] , \wRegInA9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_200 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink201[31] , \ScanLink201[30] , \ScanLink201[29] , 
        \ScanLink201[28] , \ScanLink201[27] , \ScanLink201[26] , 
        \ScanLink201[25] , \ScanLink201[24] , \ScanLink201[23] , 
        \ScanLink201[22] , \ScanLink201[21] , \ScanLink201[20] , 
        \ScanLink201[19] , \ScanLink201[18] , \ScanLink201[17] , 
        \ScanLink201[16] , \ScanLink201[15] , \ScanLink201[14] , 
        \ScanLink201[13] , \ScanLink201[12] , \ScanLink201[11] , 
        \ScanLink201[10] , \ScanLink201[9] , \ScanLink201[8] , 
        \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , \ScanLink201[4] , 
        \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , \ScanLink201[0] 
        }), .ScanOut({\ScanLink200[31] , \ScanLink200[30] , \ScanLink200[29] , 
        \ScanLink200[28] , \ScanLink200[27] , \ScanLink200[26] , 
        \ScanLink200[25] , \ScanLink200[24] , \ScanLink200[23] , 
        \ScanLink200[22] , \ScanLink200[21] , \ScanLink200[20] , 
        \ScanLink200[19] , \ScanLink200[18] , \ScanLink200[17] , 
        \ScanLink200[16] , \ScanLink200[15] , \ScanLink200[14] , 
        \ScanLink200[13] , \ScanLink200[12] , \ScanLink200[11] , 
        \ScanLink200[10] , \ScanLink200[9] , \ScanLink200[8] , 
        \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , \ScanLink200[4] , 
        \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , \ScanLink200[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB27[31] , \wRegInB27[30] , \wRegInB27[29] , 
        \wRegInB27[28] , \wRegInB27[27] , \wRegInB27[26] , \wRegInB27[25] , 
        \wRegInB27[24] , \wRegInB27[23] , \wRegInB27[22] , \wRegInB27[21] , 
        \wRegInB27[20] , \wRegInB27[19] , \wRegInB27[18] , \wRegInB27[17] , 
        \wRegInB27[16] , \wRegInB27[15] , \wRegInB27[14] , \wRegInB27[13] , 
        \wRegInB27[12] , \wRegInB27[11] , \wRegInB27[10] , \wRegInB27[9] , 
        \wRegInB27[8] , \wRegInB27[7] , \wRegInB27[6] , \wRegInB27[5] , 
        \wRegInB27[4] , \wRegInB27[3] , \wRegInB27[2] , \wRegInB27[1] , 
        \wRegInB27[0] }), .Out({\wBIn27[31] , \wBIn27[30] , \wBIn27[29] , 
        \wBIn27[28] , \wBIn27[27] , \wBIn27[26] , \wBIn27[25] , \wBIn27[24] , 
        \wBIn27[23] , \wBIn27[22] , \wBIn27[21] , \wBIn27[20] , \wBIn27[19] , 
        \wBIn27[18] , \wBIn27[17] , \wBIn27[16] , \wBIn27[15] , \wBIn27[14] , 
        \wBIn27[13] , \wBIn27[12] , \wBIn27[11] , \wBIn27[10] , \wBIn27[9] , 
        \wBIn27[8] , \wBIn27[7] , \wBIn27[6] , \wBIn27[5] , \wBIn27[4] , 
        \wBIn27[3] , \wBIn27[2] , \wBIn27[1] , \wBIn27[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_4 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[31] , \ScanLink5[30] , \ScanLink5[29] , 
        \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , \ScanLink5[25] , 
        \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , \ScanLink5[21] , 
        \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , \ScanLink5[17] , 
        \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , \ScanLink5[13] , 
        \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , \ScanLink5[9] , 
        \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB125[31] , \wRegInB125[30] , 
        \wRegInB125[29] , \wRegInB125[28] , \wRegInB125[27] , \wRegInB125[26] , 
        \wRegInB125[25] , \wRegInB125[24] , \wRegInB125[23] , \wRegInB125[22] , 
        \wRegInB125[21] , \wRegInB125[20] , \wRegInB125[19] , \wRegInB125[18] , 
        \wRegInB125[17] , \wRegInB125[16] , \wRegInB125[15] , \wRegInB125[14] , 
        \wRegInB125[13] , \wRegInB125[12] , \wRegInB125[11] , \wRegInB125[10] , 
        \wRegInB125[9] , \wRegInB125[8] , \wRegInB125[7] , \wRegInB125[6] , 
        \wRegInB125[5] , \wRegInB125[4] , \wRegInB125[3] , \wRegInB125[2] , 
        \wRegInB125[1] , \wRegInB125[0] }), .Out({\wBIn125[31] , \wBIn125[30] , 
        \wBIn125[29] , \wBIn125[28] , \wBIn125[27] , \wBIn125[26] , 
        \wBIn125[25] , \wBIn125[24] , \wBIn125[23] , \wBIn125[22] , 
        \wBIn125[21] , \wBIn125[20] , \wBIn125[19] , \wBIn125[18] , 
        \wBIn125[17] , \wBIn125[16] , \wBIn125[15] , \wBIn125[14] , 
        \wBIn125[13] , \wBIn125[12] , \wBIn125[11] , \wBIn125[10] , 
        \wBIn125[9] , \wBIn125[8] , \wBIn125[7] , \wBIn125[6] , \wBIn125[5] , 
        \wBIn125[4] , \wBIn125[3] , \wBIn125[2] , \wBIn125[1] , \wBIn125[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_130 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink131[31] , \ScanLink131[30] , \ScanLink131[29] , 
        \ScanLink131[28] , \ScanLink131[27] , \ScanLink131[26] , 
        \ScanLink131[25] , \ScanLink131[24] , \ScanLink131[23] , 
        \ScanLink131[22] , \ScanLink131[21] , \ScanLink131[20] , 
        \ScanLink131[19] , \ScanLink131[18] , \ScanLink131[17] , 
        \ScanLink131[16] , \ScanLink131[15] , \ScanLink131[14] , 
        \ScanLink131[13] , \ScanLink131[12] , \ScanLink131[11] , 
        \ScanLink131[10] , \ScanLink131[9] , \ScanLink131[8] , 
        \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , \ScanLink131[4] , 
        \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , \ScanLink131[0] 
        }), .ScanOut({\ScanLink130[31] , \ScanLink130[30] , \ScanLink130[29] , 
        \ScanLink130[28] , \ScanLink130[27] , \ScanLink130[26] , 
        \ScanLink130[25] , \ScanLink130[24] , \ScanLink130[23] , 
        \ScanLink130[22] , \ScanLink130[21] , \ScanLink130[20] , 
        \ScanLink130[19] , \ScanLink130[18] , \ScanLink130[17] , 
        \ScanLink130[16] , \ScanLink130[15] , \ScanLink130[14] , 
        \ScanLink130[13] , \ScanLink130[12] , \ScanLink130[11] , 
        \ScanLink130[10] , \ScanLink130[9] , \ScanLink130[8] , 
        \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , \ScanLink130[4] , 
        \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , \ScanLink130[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB62[31] , \wRegInB62[30] , \wRegInB62[29] , 
        \wRegInB62[28] , \wRegInB62[27] , \wRegInB62[26] , \wRegInB62[25] , 
        \wRegInB62[24] , \wRegInB62[23] , \wRegInB62[22] , \wRegInB62[21] , 
        \wRegInB62[20] , \wRegInB62[19] , \wRegInB62[18] , \wRegInB62[17] , 
        \wRegInB62[16] , \wRegInB62[15] , \wRegInB62[14] , \wRegInB62[13] , 
        \wRegInB62[12] , \wRegInB62[11] , \wRegInB62[10] , \wRegInB62[9] , 
        \wRegInB62[8] , \wRegInB62[7] , \wRegInB62[6] , \wRegInB62[5] , 
        \wRegInB62[4] , \wRegInB62[3] , \wRegInB62[2] , \wRegInB62[1] , 
        \wRegInB62[0] }), .Out({\wBIn62[31] , \wBIn62[30] , \wBIn62[29] , 
        \wBIn62[28] , \wBIn62[27] , \wBIn62[26] , \wBIn62[25] , \wBIn62[24] , 
        \wBIn62[23] , \wBIn62[22] , \wBIn62[21] , \wBIn62[20] , \wBIn62[19] , 
        \wBIn62[18] , \wBIn62[17] , \wBIn62[16] , \wBIn62[15] , \wBIn62[14] , 
        \wBIn62[13] , \wBIn62[12] , \wBIn62[11] , \wBIn62[10] , \wBIn62[9] , 
        \wBIn62[8] , \wBIn62[7] , \wBIn62[6] , \wBIn62[5] , \wBIn62[4] , 
        \wBIn62[3] , \wBIn62[2] , \wBIn62[1] , \wBIn62[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_60 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink61[31] , \ScanLink61[30] , \ScanLink61[29] , 
        \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , \ScanLink61[25] , 
        \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , \ScanLink61[21] , 
        \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , \ScanLink61[17] , 
        \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , \ScanLink61[13] , 
        \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , \ScanLink61[9] , 
        \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , \ScanLink61[5] , 
        \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , \ScanLink61[1] , 
        \ScanLink61[0] }), .ScanOut({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB97[31] , \wRegInB97[30] , 
        \wRegInB97[29] , \wRegInB97[28] , \wRegInB97[27] , \wRegInB97[26] , 
        \wRegInB97[25] , \wRegInB97[24] , \wRegInB97[23] , \wRegInB97[22] , 
        \wRegInB97[21] , \wRegInB97[20] , \wRegInB97[19] , \wRegInB97[18] , 
        \wRegInB97[17] , \wRegInB97[16] , \wRegInB97[15] , \wRegInB97[14] , 
        \wRegInB97[13] , \wRegInB97[12] , \wRegInB97[11] , \wRegInB97[10] , 
        \wRegInB97[9] , \wRegInB97[8] , \wRegInB97[7] , \wRegInB97[6] , 
        \wRegInB97[5] , \wRegInB97[4] , \wRegInB97[3] , \wRegInB97[2] , 
        \wRegInB97[1] , \wRegInB97[0] }), .Out({\wBIn97[31] , \wBIn97[30] , 
        \wBIn97[29] , \wBIn97[28] , \wBIn97[27] , \wBIn97[26] , \wBIn97[25] , 
        \wBIn97[24] , \wBIn97[23] , \wBIn97[22] , \wBIn97[21] , \wBIn97[20] , 
        \wBIn97[19] , \wBIn97[18] , \wBIn97[17] , \wBIn97[16] , \wBIn97[15] , 
        \wBIn97[14] , \wBIn97[13] , \wBIn97[12] , \wBIn97[11] , \wBIn97[10] , 
        \wBIn97[9] , \wBIn97[8] , \wBIn97[7] , \wBIn97[6] , \wBIn97[5] , 
        \wBIn97[4] , \wBIn97[3] , \wBIn97[2] , \wBIn97[1] , \wBIn97[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn15[31] , \wAIn15[30] , \wAIn15[29] , \wAIn15[28] , \wAIn15[27] , 
        \wAIn15[26] , \wAIn15[25] , \wAIn15[24] , \wAIn15[23] , \wAIn15[22] , 
        \wAIn15[21] , \wAIn15[20] , \wAIn15[19] , \wAIn15[18] , \wAIn15[17] , 
        \wAIn15[16] , \wAIn15[15] , \wAIn15[14] , \wAIn15[13] , \wAIn15[12] , 
        \wAIn15[11] , \wAIn15[10] , \wAIn15[9] , \wAIn15[8] , \wAIn15[7] , 
        \wAIn15[6] , \wAIn15[5] , \wAIn15[4] , \wAIn15[3] , \wAIn15[2] , 
        \wAIn15[1] , \wAIn15[0] }), .BIn({\wBIn15[31] , \wBIn15[30] , 
        \wBIn15[29] , \wBIn15[28] , \wBIn15[27] , \wBIn15[26] , \wBIn15[25] , 
        \wBIn15[24] , \wBIn15[23] , \wBIn15[22] , \wBIn15[21] , \wBIn15[20] , 
        \wBIn15[19] , \wBIn15[18] , \wBIn15[17] , \wBIn15[16] , \wBIn15[15] , 
        \wBIn15[14] , \wBIn15[13] , \wBIn15[12] , \wBIn15[11] , \wBIn15[10] , 
        \wBIn15[9] , \wBIn15[8] , \wBIn15[7] , \wBIn15[6] , \wBIn15[5] , 
        \wBIn15[4] , \wBIn15[3] , \wBIn15[2] , \wBIn15[1] , \wBIn15[0] }), 
        .HiOut({\wBMid14[31] , \wBMid14[30] , \wBMid14[29] , \wBMid14[28] , 
        \wBMid14[27] , \wBMid14[26] , \wBMid14[25] , \wBMid14[24] , 
        \wBMid14[23] , \wBMid14[22] , \wBMid14[21] , \wBMid14[20] , 
        \wBMid14[19] , \wBMid14[18] , \wBMid14[17] , \wBMid14[16] , 
        \wBMid14[15] , \wBMid14[14] , \wBMid14[13] , \wBMid14[12] , 
        \wBMid14[11] , \wBMid14[10] , \wBMid14[9] , \wBMid14[8] , \wBMid14[7] , 
        \wBMid14[6] , \wBMid14[5] , \wBMid14[4] , \wBMid14[3] , \wBMid14[2] , 
        \wBMid14[1] , \wBMid14[0] }), .LoOut({\wAMid15[31] , \wAMid15[30] , 
        \wAMid15[29] , \wAMid15[28] , \wAMid15[27] , \wAMid15[26] , 
        \wAMid15[25] , \wAMid15[24] , \wAMid15[23] , \wAMid15[22] , 
        \wAMid15[21] , \wAMid15[20] , \wAMid15[19] , \wAMid15[18] , 
        \wAMid15[17] , \wAMid15[16] , \wAMid15[15] , \wAMid15[14] , 
        \wAMid15[13] , \wAMid15[12] , \wAMid15[11] , \wAMid15[10] , 
        \wAMid15[9] , \wAMid15[8] , \wAMid15[7] , \wAMid15[6] , \wAMid15[5] , 
        \wAMid15[4] , \wAMid15[3] , \wAMid15[2] , \wAMid15[1] , \wAMid15[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn20[31] , \wAIn20[30] , \wAIn20[29] , \wAIn20[28] , \wAIn20[27] , 
        \wAIn20[26] , \wAIn20[25] , \wAIn20[24] , \wAIn20[23] , \wAIn20[22] , 
        \wAIn20[21] , \wAIn20[20] , \wAIn20[19] , \wAIn20[18] , \wAIn20[17] , 
        \wAIn20[16] , \wAIn20[15] , \wAIn20[14] , \wAIn20[13] , \wAIn20[12] , 
        \wAIn20[11] , \wAIn20[10] , \wAIn20[9] , \wAIn20[8] , \wAIn20[7] , 
        \wAIn20[6] , \wAIn20[5] , \wAIn20[4] , \wAIn20[3] , \wAIn20[2] , 
        \wAIn20[1] , \wAIn20[0] }), .BIn({\wBIn20[31] , \wBIn20[30] , 
        \wBIn20[29] , \wBIn20[28] , \wBIn20[27] , \wBIn20[26] , \wBIn20[25] , 
        \wBIn20[24] , \wBIn20[23] , \wBIn20[22] , \wBIn20[21] , \wBIn20[20] , 
        \wBIn20[19] , \wBIn20[18] , \wBIn20[17] , \wBIn20[16] , \wBIn20[15] , 
        \wBIn20[14] , \wBIn20[13] , \wBIn20[12] , \wBIn20[11] , \wBIn20[10] , 
        \wBIn20[9] , \wBIn20[8] , \wBIn20[7] , \wBIn20[6] , \wBIn20[5] , 
        \wBIn20[4] , \wBIn20[3] , \wBIn20[2] , \wBIn20[1] , \wBIn20[0] }), 
        .HiOut({\wBMid19[31] , \wBMid19[30] , \wBMid19[29] , \wBMid19[28] , 
        \wBMid19[27] , \wBMid19[26] , \wBMid19[25] , \wBMid19[24] , 
        \wBMid19[23] , \wBMid19[22] , \wBMid19[21] , \wBMid19[20] , 
        \wBMid19[19] , \wBMid19[18] , \wBMid19[17] , \wBMid19[16] , 
        \wBMid19[15] , \wBMid19[14] , \wBMid19[13] , \wBMid19[12] , 
        \wBMid19[11] , \wBMid19[10] , \wBMid19[9] , \wBMid19[8] , \wBMid19[7] , 
        \wBMid19[6] , \wBMid19[5] , \wBMid19[4] , \wBMid19[3] , \wBMid19[2] , 
        \wBMid19[1] , \wBMid19[0] }), .LoOut({\wAMid20[31] , \wAMid20[30] , 
        \wAMid20[29] , \wAMid20[28] , \wAMid20[27] , \wAMid20[26] , 
        \wAMid20[25] , \wAMid20[24] , \wAMid20[23] , \wAMid20[22] , 
        \wAMid20[21] , \wAMid20[20] , \wAMid20[19] , \wAMid20[18] , 
        \wAMid20[17] , \wAMid20[16] , \wAMid20[15] , \wAMid20[14] , 
        \wAMid20[13] , \wAMid20[12] , \wAMid20[11] , \wAMid20[10] , 
        \wAMid20[9] , \wAMid20[8] , \wAMid20[7] , \wAMid20[6] , \wAMid20[5] , 
        \wAMid20[4] , \wAMid20[3] , \wAMid20[2] , \wAMid20[1] , \wAMid20[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn27[31] , \wAIn27[30] , \wAIn27[29] , \wAIn27[28] , \wAIn27[27] , 
        \wAIn27[26] , \wAIn27[25] , \wAIn27[24] , \wAIn27[23] , \wAIn27[22] , 
        \wAIn27[21] , \wAIn27[20] , \wAIn27[19] , \wAIn27[18] , \wAIn27[17] , 
        \wAIn27[16] , \wAIn27[15] , \wAIn27[14] , \wAIn27[13] , \wAIn27[12] , 
        \wAIn27[11] , \wAIn27[10] , \wAIn27[9] , \wAIn27[8] , \wAIn27[7] , 
        \wAIn27[6] , \wAIn27[5] , \wAIn27[4] , \wAIn27[3] , \wAIn27[2] , 
        \wAIn27[1] , \wAIn27[0] }), .BIn({\wBIn27[31] , \wBIn27[30] , 
        \wBIn27[29] , \wBIn27[28] , \wBIn27[27] , \wBIn27[26] , \wBIn27[25] , 
        \wBIn27[24] , \wBIn27[23] , \wBIn27[22] , \wBIn27[21] , \wBIn27[20] , 
        \wBIn27[19] , \wBIn27[18] , \wBIn27[17] , \wBIn27[16] , \wBIn27[15] , 
        \wBIn27[14] , \wBIn27[13] , \wBIn27[12] , \wBIn27[11] , \wBIn27[10] , 
        \wBIn27[9] , \wBIn27[8] , \wBIn27[7] , \wBIn27[6] , \wBIn27[5] , 
        \wBIn27[4] , \wBIn27[3] , \wBIn27[2] , \wBIn27[1] , \wBIn27[0] }), 
        .HiOut({\wBMid26[31] , \wBMid26[30] , \wBMid26[29] , \wBMid26[28] , 
        \wBMid26[27] , \wBMid26[26] , \wBMid26[25] , \wBMid26[24] , 
        \wBMid26[23] , \wBMid26[22] , \wBMid26[21] , \wBMid26[20] , 
        \wBMid26[19] , \wBMid26[18] , \wBMid26[17] , \wBMid26[16] , 
        \wBMid26[15] , \wBMid26[14] , \wBMid26[13] , \wBMid26[12] , 
        \wBMid26[11] , \wBMid26[10] , \wBMid26[9] , \wBMid26[8] , \wBMid26[7] , 
        \wBMid26[6] , \wBMid26[5] , \wBMid26[4] , \wBMid26[3] , \wBMid26[2] , 
        \wBMid26[1] , \wBMid26[0] }), .LoOut({\wAMid27[31] , \wAMid27[30] , 
        \wAMid27[29] , \wAMid27[28] , \wAMid27[27] , \wAMid27[26] , 
        \wAMid27[25] , \wAMid27[24] , \wAMid27[23] , \wAMid27[22] , 
        \wAMid27[21] , \wAMid27[20] , \wAMid27[19] , \wAMid27[18] , 
        \wAMid27[17] , \wAMid27[16] , \wAMid27[15] , \wAMid27[14] , 
        \wAMid27[13] , \wAMid27[12] , \wAMid27[11] , \wAMid27[10] , 
        \wAMid27[9] , \wAMid27[8] , \wAMid27[7] , \wAMid27[6] , \wAMid27[5] , 
        \wAMid27[4] , \wAMid27[3] , \wAMid27[2] , \wAMid27[1] , \wAMid27[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid22[31] , \wAMid22[30] , \wAMid22[29] , \wAMid22[28] , 
        \wAMid22[27] , \wAMid22[26] , \wAMid22[25] , \wAMid22[24] , 
        \wAMid22[23] , \wAMid22[22] , \wAMid22[21] , \wAMid22[20] , 
        \wAMid22[19] , \wAMid22[18] , \wAMid22[17] , \wAMid22[16] , 
        \wAMid22[15] , \wAMid22[14] , \wAMid22[13] , \wAMid22[12] , 
        \wAMid22[11] , \wAMid22[10] , \wAMid22[9] , \wAMid22[8] , \wAMid22[7] , 
        \wAMid22[6] , \wAMid22[5] , \wAMid22[4] , \wAMid22[3] , \wAMid22[2] , 
        \wAMid22[1] , \wAMid22[0] }), .BIn({\wBMid22[31] , \wBMid22[30] , 
        \wBMid22[29] , \wBMid22[28] , \wBMid22[27] , \wBMid22[26] , 
        \wBMid22[25] , \wBMid22[24] , \wBMid22[23] , \wBMid22[22] , 
        \wBMid22[21] , \wBMid22[20] , \wBMid22[19] , \wBMid22[18] , 
        \wBMid22[17] , \wBMid22[16] , \wBMid22[15] , \wBMid22[14] , 
        \wBMid22[13] , \wBMid22[12] , \wBMid22[11] , \wBMid22[10] , 
        \wBMid22[9] , \wBMid22[8] , \wBMid22[7] , \wBMid22[6] , \wBMid22[5] , 
        \wBMid22[4] , \wBMid22[3] , \wBMid22[2] , \wBMid22[1] , \wBMid22[0] }), 
        .HiOut({\wRegInB22[31] , \wRegInB22[30] , \wRegInB22[29] , 
        \wRegInB22[28] , \wRegInB22[27] , \wRegInB22[26] , \wRegInB22[25] , 
        \wRegInB22[24] , \wRegInB22[23] , \wRegInB22[22] , \wRegInB22[21] , 
        \wRegInB22[20] , \wRegInB22[19] , \wRegInB22[18] , \wRegInB22[17] , 
        \wRegInB22[16] , \wRegInB22[15] , \wRegInB22[14] , \wRegInB22[13] , 
        \wRegInB22[12] , \wRegInB22[11] , \wRegInB22[10] , \wRegInB22[9] , 
        \wRegInB22[8] , \wRegInB22[7] , \wRegInB22[6] , \wRegInB22[5] , 
        \wRegInB22[4] , \wRegInB22[3] , \wRegInB22[2] , \wRegInB22[1] , 
        \wRegInB22[0] }), .LoOut({\wRegInA23[31] , \wRegInA23[30] , 
        \wRegInA23[29] , \wRegInA23[28] , \wRegInA23[27] , \wRegInA23[26] , 
        \wRegInA23[25] , \wRegInA23[24] , \wRegInA23[23] , \wRegInA23[22] , 
        \wRegInA23[21] , \wRegInA23[20] , \wRegInA23[19] , \wRegInA23[18] , 
        \wRegInA23[17] , \wRegInA23[16] , \wRegInA23[15] , \wRegInA23[14] , 
        \wRegInA23[13] , \wRegInA23[12] , \wRegInA23[11] , \wRegInA23[10] , 
        \wRegInA23[9] , \wRegInA23[8] , \wRegInA23[7] , \wRegInA23[6] , 
        \wRegInA23[5] , \wRegInA23[4] , \wRegInA23[3] , \wRegInA23[2] , 
        \wRegInA23[1] , \wRegInA23[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_117 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink118[31] , \ScanLink118[30] , \ScanLink118[29] , 
        \ScanLink118[28] , \ScanLink118[27] , \ScanLink118[26] , 
        \ScanLink118[25] , \ScanLink118[24] , \ScanLink118[23] , 
        \ScanLink118[22] , \ScanLink118[21] , \ScanLink118[20] , 
        \ScanLink118[19] , \ScanLink118[18] , \ScanLink118[17] , 
        \ScanLink118[16] , \ScanLink118[15] , \ScanLink118[14] , 
        \ScanLink118[13] , \ScanLink118[12] , \ScanLink118[11] , 
        \ScanLink118[10] , \ScanLink118[9] , \ScanLink118[8] , 
        \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , \ScanLink118[4] , 
        \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , \ScanLink118[0] 
        }), .ScanOut({\ScanLink117[31] , \ScanLink117[30] , \ScanLink117[29] , 
        \ScanLink117[28] , \ScanLink117[27] , \ScanLink117[26] , 
        \ScanLink117[25] , \ScanLink117[24] , \ScanLink117[23] , 
        \ScanLink117[22] , \ScanLink117[21] , \ScanLink117[20] , 
        \ScanLink117[19] , \ScanLink117[18] , \ScanLink117[17] , 
        \ScanLink117[16] , \ScanLink117[15] , \ScanLink117[14] , 
        \ScanLink117[13] , \ScanLink117[12] , \ScanLink117[11] , 
        \ScanLink117[10] , \ScanLink117[9] , \ScanLink117[8] , 
        \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , \ScanLink117[4] , 
        \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , \ScanLink117[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA69[31] , \wRegInA69[30] , \wRegInA69[29] , 
        \wRegInA69[28] , \wRegInA69[27] , \wRegInA69[26] , \wRegInA69[25] , 
        \wRegInA69[24] , \wRegInA69[23] , \wRegInA69[22] , \wRegInA69[21] , 
        \wRegInA69[20] , \wRegInA69[19] , \wRegInA69[18] , \wRegInA69[17] , 
        \wRegInA69[16] , \wRegInA69[15] , \wRegInA69[14] , \wRegInA69[13] , 
        \wRegInA69[12] , \wRegInA69[11] , \wRegInA69[10] , \wRegInA69[9] , 
        \wRegInA69[8] , \wRegInA69[7] , \wRegInA69[6] , \wRegInA69[5] , 
        \wRegInA69[4] , \wRegInA69[3] , \wRegInA69[2] , \wRegInA69[1] , 
        \wRegInA69[0] }), .Out({\wAIn69[31] , \wAIn69[30] , \wAIn69[29] , 
        \wAIn69[28] , \wAIn69[27] , \wAIn69[26] , \wAIn69[25] , \wAIn69[24] , 
        \wAIn69[23] , \wAIn69[22] , \wAIn69[21] , \wAIn69[20] , \wAIn69[19] , 
        \wAIn69[18] , \wAIn69[17] , \wAIn69[16] , \wAIn69[15] , \wAIn69[14] , 
        \wAIn69[13] , \wAIn69[12] , \wAIn69[11] , \wAIn69[10] , \wAIn69[9] , 
        \wAIn69[8] , \wAIn69[7] , \wAIn69[6] , \wAIn69[5] , \wAIn69[4] , 
        \wAIn69[3] , \wAIn69[2] , \wAIn69[1] , \wAIn69[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_227 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink228[31] , \ScanLink228[30] , \ScanLink228[29] , 
        \ScanLink228[28] , \ScanLink228[27] , \ScanLink228[26] , 
        \ScanLink228[25] , \ScanLink228[24] , \ScanLink228[23] , 
        \ScanLink228[22] , \ScanLink228[21] , \ScanLink228[20] , 
        \ScanLink228[19] , \ScanLink228[18] , \ScanLink228[17] , 
        \ScanLink228[16] , \ScanLink228[15] , \ScanLink228[14] , 
        \ScanLink228[13] , \ScanLink228[12] , \ScanLink228[11] , 
        \ScanLink228[10] , \ScanLink228[9] , \ScanLink228[8] , 
        \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , \ScanLink228[4] , 
        \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , \ScanLink228[0] 
        }), .ScanOut({\ScanLink227[31] , \ScanLink227[30] , \ScanLink227[29] , 
        \ScanLink227[28] , \ScanLink227[27] , \ScanLink227[26] , 
        \ScanLink227[25] , \ScanLink227[24] , \ScanLink227[23] , 
        \ScanLink227[22] , \ScanLink227[21] , \ScanLink227[20] , 
        \ScanLink227[19] , \ScanLink227[18] , \ScanLink227[17] , 
        \ScanLink227[16] , \ScanLink227[15] , \ScanLink227[14] , 
        \ScanLink227[13] , \ScanLink227[12] , \ScanLink227[11] , 
        \ScanLink227[10] , \ScanLink227[9] , \ScanLink227[8] , 
        \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , \ScanLink227[4] , 
        \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , \ScanLink227[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA14[31] , \wRegInA14[30] , \wRegInA14[29] , 
        \wRegInA14[28] , \wRegInA14[27] , \wRegInA14[26] , \wRegInA14[25] , 
        \wRegInA14[24] , \wRegInA14[23] , \wRegInA14[22] , \wRegInA14[21] , 
        \wRegInA14[20] , \wRegInA14[19] , \wRegInA14[18] , \wRegInA14[17] , 
        \wRegInA14[16] , \wRegInA14[15] , \wRegInA14[14] , \wRegInA14[13] , 
        \wRegInA14[12] , \wRegInA14[11] , \wRegInA14[10] , \wRegInA14[9] , 
        \wRegInA14[8] , \wRegInA14[7] , \wRegInA14[6] , \wRegInA14[5] , 
        \wRegInA14[4] , \wRegInA14[3] , \wRegInA14[2] , \wRegInA14[1] , 
        \wRegInA14[0] }), .Out({\wAIn14[31] , \wAIn14[30] , \wAIn14[29] , 
        \wAIn14[28] , \wAIn14[27] , \wAIn14[26] , \wAIn14[25] , \wAIn14[24] , 
        \wAIn14[23] , \wAIn14[22] , \wAIn14[21] , \wAIn14[20] , \wAIn14[19] , 
        \wAIn14[18] , \wAIn14[17] , \wAIn14[16] , \wAIn14[15] , \wAIn14[14] , 
        \wAIn14[13] , \wAIn14[12] , \wAIn14[11] , \wAIn14[10] , \wAIn14[9] , 
        \wAIn14[8] , \wAIn14[7] , \wAIn14[6] , \wAIn14[5] , \wAIn14[4] , 
        \wAIn14[3] , \wAIn14[2] , \wAIn14[1] , \wAIn14[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_47 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink48[31] , \ScanLink48[30] , \ScanLink48[29] , 
        \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , \ScanLink48[25] , 
        \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , \ScanLink48[21] , 
        \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , \ScanLink48[17] , 
        \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , \ScanLink48[13] , 
        \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , \ScanLink48[9] , 
        \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , \ScanLink48[5] , 
        \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , \ScanLink48[1] , 
        \ScanLink48[0] }), .ScanOut({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA104[31] , \wRegInA104[30] , 
        \wRegInA104[29] , \wRegInA104[28] , \wRegInA104[27] , \wRegInA104[26] , 
        \wRegInA104[25] , \wRegInA104[24] , \wRegInA104[23] , \wRegInA104[22] , 
        \wRegInA104[21] , \wRegInA104[20] , \wRegInA104[19] , \wRegInA104[18] , 
        \wRegInA104[17] , \wRegInA104[16] , \wRegInA104[15] , \wRegInA104[14] , 
        \wRegInA104[13] , \wRegInA104[12] , \wRegInA104[11] , \wRegInA104[10] , 
        \wRegInA104[9] , \wRegInA104[8] , \wRegInA104[7] , \wRegInA104[6] , 
        \wRegInA104[5] , \wRegInA104[4] , \wRegInA104[3] , \wRegInA104[2] , 
        \wRegInA104[1] , \wRegInA104[0] }), .Out({\wAIn104[31] , \wAIn104[30] , 
        \wAIn104[29] , \wAIn104[28] , \wAIn104[27] , \wAIn104[26] , 
        \wAIn104[25] , \wAIn104[24] , \wAIn104[23] , \wAIn104[22] , 
        \wAIn104[21] , \wAIn104[20] , \wAIn104[19] , \wAIn104[18] , 
        \wAIn104[17] , \wAIn104[16] , \wAIn104[15] , \wAIn104[14] , 
        \wAIn104[13] , \wAIn104[12] , \wAIn104[11] , \wAIn104[10] , 
        \wAIn104[9] , \wAIn104[8] , \wAIn104[7] , \wAIn104[6] , \wAIn104[5] , 
        \wAIn104[4] , \wAIn104[3] , \wAIn104[2] , \wAIn104[1] , \wAIn104[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_212 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink213[31] , \ScanLink213[30] , \ScanLink213[29] , 
        \ScanLink213[28] , \ScanLink213[27] , \ScanLink213[26] , 
        \ScanLink213[25] , \ScanLink213[24] , \ScanLink213[23] , 
        \ScanLink213[22] , \ScanLink213[21] , \ScanLink213[20] , 
        \ScanLink213[19] , \ScanLink213[18] , \ScanLink213[17] , 
        \ScanLink213[16] , \ScanLink213[15] , \ScanLink213[14] , 
        \ScanLink213[13] , \ScanLink213[12] , \ScanLink213[11] , 
        \ScanLink213[10] , \ScanLink213[9] , \ScanLink213[8] , 
        \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , \ScanLink213[4] , 
        \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , \ScanLink213[0] 
        }), .ScanOut({\ScanLink212[31] , \ScanLink212[30] , \ScanLink212[29] , 
        \ScanLink212[28] , \ScanLink212[27] , \ScanLink212[26] , 
        \ScanLink212[25] , \ScanLink212[24] , \ScanLink212[23] , 
        \ScanLink212[22] , \ScanLink212[21] , \ScanLink212[20] , 
        \ScanLink212[19] , \ScanLink212[18] , \ScanLink212[17] , 
        \ScanLink212[16] , \ScanLink212[15] , \ScanLink212[14] , 
        \ScanLink212[13] , \ScanLink212[12] , \ScanLink212[11] , 
        \ScanLink212[10] , \ScanLink212[9] , \ScanLink212[8] , 
        \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , \ScanLink212[4] , 
        \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , \ScanLink212[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB21[31] , \wRegInB21[30] , \wRegInB21[29] , 
        \wRegInB21[28] , \wRegInB21[27] , \wRegInB21[26] , \wRegInB21[25] , 
        \wRegInB21[24] , \wRegInB21[23] , \wRegInB21[22] , \wRegInB21[21] , 
        \wRegInB21[20] , \wRegInB21[19] , \wRegInB21[18] , \wRegInB21[17] , 
        \wRegInB21[16] , \wRegInB21[15] , \wRegInB21[14] , \wRegInB21[13] , 
        \wRegInB21[12] , \wRegInB21[11] , \wRegInB21[10] , \wRegInB21[9] , 
        \wRegInB21[8] , \wRegInB21[7] , \wRegInB21[6] , \wRegInB21[5] , 
        \wRegInB21[4] , \wRegInB21[3] , \wRegInB21[2] , \wRegInB21[1] , 
        \wRegInB21[0] }), .Out({\wBIn21[31] , \wBIn21[30] , \wBIn21[29] , 
        \wBIn21[28] , \wBIn21[27] , \wBIn21[26] , \wBIn21[25] , \wBIn21[24] , 
        \wBIn21[23] , \wBIn21[22] , \wBIn21[21] , \wBIn21[20] , \wBIn21[19] , 
        \wBIn21[18] , \wBIn21[17] , \wBIn21[16] , \wBIn21[15] , \wBIn21[14] , 
        \wBIn21[13] , \wBIn21[12] , \wBIn21[11] , \wBIn21[10] , \wBIn21[9] , 
        \wBIn21[8] , \wBIn21[7] , \wBIn21[6] , \wBIn21[5] , \wBIn21[4] , 
        \wBIn21[3] , \wBIn21[2] , \wBIn21[1] , \wBIn21[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn49[31] , \wAIn49[30] , \wAIn49[29] , \wAIn49[28] , \wAIn49[27] , 
        \wAIn49[26] , \wAIn49[25] , \wAIn49[24] , \wAIn49[23] , \wAIn49[22] , 
        \wAIn49[21] , \wAIn49[20] , \wAIn49[19] , \wAIn49[18] , \wAIn49[17] , 
        \wAIn49[16] , \wAIn49[15] , \wAIn49[14] , \wAIn49[13] , \wAIn49[12] , 
        \wAIn49[11] , \wAIn49[10] , \wAIn49[9] , \wAIn49[8] , \wAIn49[7] , 
        \wAIn49[6] , \wAIn49[5] , \wAIn49[4] , \wAIn49[3] , \wAIn49[2] , 
        \wAIn49[1] , \wAIn49[0] }), .BIn({\wBIn49[31] , \wBIn49[30] , 
        \wBIn49[29] , \wBIn49[28] , \wBIn49[27] , \wBIn49[26] , \wBIn49[25] , 
        \wBIn49[24] , \wBIn49[23] , \wBIn49[22] , \wBIn49[21] , \wBIn49[20] , 
        \wBIn49[19] , \wBIn49[18] , \wBIn49[17] , \wBIn49[16] , \wBIn49[15] , 
        \wBIn49[14] , \wBIn49[13] , \wBIn49[12] , \wBIn49[11] , \wBIn49[10] , 
        \wBIn49[9] , \wBIn49[8] , \wBIn49[7] , \wBIn49[6] , \wBIn49[5] , 
        \wBIn49[4] , \wBIn49[3] , \wBIn49[2] , \wBIn49[1] , \wBIn49[0] }), 
        .HiOut({\wBMid48[31] , \wBMid48[30] , \wBMid48[29] , \wBMid48[28] , 
        \wBMid48[27] , \wBMid48[26] , \wBMid48[25] , \wBMid48[24] , 
        \wBMid48[23] , \wBMid48[22] , \wBMid48[21] , \wBMid48[20] , 
        \wBMid48[19] , \wBMid48[18] , \wBMid48[17] , \wBMid48[16] , 
        \wBMid48[15] , \wBMid48[14] , \wBMid48[13] , \wBMid48[12] , 
        \wBMid48[11] , \wBMid48[10] , \wBMid48[9] , \wBMid48[8] , \wBMid48[7] , 
        \wBMid48[6] , \wBMid48[5] , \wBMid48[4] , \wBMid48[3] , \wBMid48[2] , 
        \wBMid48[1] , \wBMid48[0] }), .LoOut({\wAMid49[31] , \wAMid49[30] , 
        \wAMid49[29] , \wAMid49[28] , \wAMid49[27] , \wAMid49[26] , 
        \wAMid49[25] , \wAMid49[24] , \wAMid49[23] , \wAMid49[22] , 
        \wAMid49[21] , \wAMid49[20] , \wAMid49[19] , \wAMid49[18] , 
        \wAMid49[17] , \wAMid49[16] , \wAMid49[15] , \wAMid49[14] , 
        \wAMid49[13] , \wAMid49[12] , \wAMid49[11] , \wAMid49[10] , 
        \wAMid49[9] , \wAMid49[8] , \wAMid49[7] , \wAMid49[6] , \wAMid49[5] , 
        \wAMid49[4] , \wAMid49[3] , \wAMid49[2] , \wAMid49[1] , \wAMid49[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid17[31] , \wAMid17[30] , \wAMid17[29] , \wAMid17[28] , 
        \wAMid17[27] , \wAMid17[26] , \wAMid17[25] , \wAMid17[24] , 
        \wAMid17[23] , \wAMid17[22] , \wAMid17[21] , \wAMid17[20] , 
        \wAMid17[19] , \wAMid17[18] , \wAMid17[17] , \wAMid17[16] , 
        \wAMid17[15] , \wAMid17[14] , \wAMid17[13] , \wAMid17[12] , 
        \wAMid17[11] , \wAMid17[10] , \wAMid17[9] , \wAMid17[8] , \wAMid17[7] , 
        \wAMid17[6] , \wAMid17[5] , \wAMid17[4] , \wAMid17[3] , \wAMid17[2] , 
        \wAMid17[1] , \wAMid17[0] }), .BIn({\wBMid17[31] , \wBMid17[30] , 
        \wBMid17[29] , \wBMid17[28] , \wBMid17[27] , \wBMid17[26] , 
        \wBMid17[25] , \wBMid17[24] , \wBMid17[23] , \wBMid17[22] , 
        \wBMid17[21] , \wBMid17[20] , \wBMid17[19] , \wBMid17[18] , 
        \wBMid17[17] , \wBMid17[16] , \wBMid17[15] , \wBMid17[14] , 
        \wBMid17[13] , \wBMid17[12] , \wBMid17[11] , \wBMid17[10] , 
        \wBMid17[9] , \wBMid17[8] , \wBMid17[7] , \wBMid17[6] , \wBMid17[5] , 
        \wBMid17[4] , \wBMid17[3] , \wBMid17[2] , \wBMid17[1] , \wBMid17[0] }), 
        .HiOut({\wRegInB17[31] , \wRegInB17[30] , \wRegInB17[29] , 
        \wRegInB17[28] , \wRegInB17[27] , \wRegInB17[26] , \wRegInB17[25] , 
        \wRegInB17[24] , \wRegInB17[23] , \wRegInB17[22] , \wRegInB17[21] , 
        \wRegInB17[20] , \wRegInB17[19] , \wRegInB17[18] , \wRegInB17[17] , 
        \wRegInB17[16] , \wRegInB17[15] , \wRegInB17[14] , \wRegInB17[13] , 
        \wRegInB17[12] , \wRegInB17[11] , \wRegInB17[10] , \wRegInB17[9] , 
        \wRegInB17[8] , \wRegInB17[7] , \wRegInB17[6] , \wRegInB17[5] , 
        \wRegInB17[4] , \wRegInB17[3] , \wRegInB17[2] , \wRegInB17[1] , 
        \wRegInB17[0] }), .LoOut({\wRegInA18[31] , \wRegInA18[30] , 
        \wRegInA18[29] , \wRegInA18[28] , \wRegInA18[27] , \wRegInA18[26] , 
        \wRegInA18[25] , \wRegInA18[24] , \wRegInA18[23] , \wRegInA18[22] , 
        \wRegInA18[21] , \wRegInA18[20] , \wRegInA18[19] , \wRegInA18[18] , 
        \wRegInA18[17] , \wRegInA18[16] , \wRegInA18[15] , \wRegInA18[14] , 
        \wRegInA18[13] , \wRegInA18[12] , \wRegInA18[11] , \wRegInA18[10] , 
        \wRegInA18[9] , \wRegInA18[8] , \wRegInA18[7] , \wRegInA18[6] , 
        \wRegInA18[5] , \wRegInA18[4] , \wRegInA18[3] , \wRegInA18[2] , 
        \wRegInA18[1] , \wRegInA18[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_72 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink73[31] , \ScanLink73[30] , \ScanLink73[29] , 
        \ScanLink73[28] , \ScanLink73[27] , \ScanLink73[26] , \ScanLink73[25] , 
        \ScanLink73[24] , \ScanLink73[23] , \ScanLink73[22] , \ScanLink73[21] , 
        \ScanLink73[20] , \ScanLink73[19] , \ScanLink73[18] , \ScanLink73[17] , 
        \ScanLink73[16] , \ScanLink73[15] , \ScanLink73[14] , \ScanLink73[13] , 
        \ScanLink73[12] , \ScanLink73[11] , \ScanLink73[10] , \ScanLink73[9] , 
        \ScanLink73[8] , \ScanLink73[7] , \ScanLink73[6] , \ScanLink73[5] , 
        \ScanLink73[4] , \ScanLink73[3] , \ScanLink73[2] , \ScanLink73[1] , 
        \ScanLink73[0] }), .ScanOut({\ScanLink72[31] , \ScanLink72[30] , 
        \ScanLink72[29] , \ScanLink72[28] , \ScanLink72[27] , \ScanLink72[26] , 
        \ScanLink72[25] , \ScanLink72[24] , \ScanLink72[23] , \ScanLink72[22] , 
        \ScanLink72[21] , \ScanLink72[20] , \ScanLink72[19] , \ScanLink72[18] , 
        \ScanLink72[17] , \ScanLink72[16] , \ScanLink72[15] , \ScanLink72[14] , 
        \ScanLink72[13] , \ScanLink72[12] , \ScanLink72[11] , \ScanLink72[10] , 
        \ScanLink72[9] , \ScanLink72[8] , \ScanLink72[7] , \ScanLink72[6] , 
        \ScanLink72[5] , \ScanLink72[4] , \ScanLink72[3] , \ScanLink72[2] , 
        \ScanLink72[1] , \ScanLink72[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB91[31] , \wRegInB91[30] , 
        \wRegInB91[29] , \wRegInB91[28] , \wRegInB91[27] , \wRegInB91[26] , 
        \wRegInB91[25] , \wRegInB91[24] , \wRegInB91[23] , \wRegInB91[22] , 
        \wRegInB91[21] , \wRegInB91[20] , \wRegInB91[19] , \wRegInB91[18] , 
        \wRegInB91[17] , \wRegInB91[16] , \wRegInB91[15] , \wRegInB91[14] , 
        \wRegInB91[13] , \wRegInB91[12] , \wRegInB91[11] , \wRegInB91[10] , 
        \wRegInB91[9] , \wRegInB91[8] , \wRegInB91[7] , \wRegInB91[6] , 
        \wRegInB91[5] , \wRegInB91[4] , \wRegInB91[3] , \wRegInB91[2] , 
        \wRegInB91[1] , \wRegInB91[0] }), .Out({\wBIn91[31] , \wBIn91[30] , 
        \wBIn91[29] , \wBIn91[28] , \wBIn91[27] , \wBIn91[26] , \wBIn91[25] , 
        \wBIn91[24] , \wBIn91[23] , \wBIn91[22] , \wBIn91[21] , \wBIn91[20] , 
        \wBIn91[19] , \wBIn91[18] , \wBIn91[17] , \wBIn91[16] , \wBIn91[15] , 
        \wBIn91[14] , \wBIn91[13] , \wBIn91[12] , \wBIn91[11] , \wBIn91[10] , 
        \wBIn91[9] , \wBIn91[8] , \wBIn91[7] , \wBIn91[6] , \wBIn91[5] , 
        \wBIn91[4] , \wBIn91[3] , \wBIn91[2] , \wBIn91[1] , \wBIn91[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid30[31] , \wAMid30[30] , \wAMid30[29] , \wAMid30[28] , 
        \wAMid30[27] , \wAMid30[26] , \wAMid30[25] , \wAMid30[24] , 
        \wAMid30[23] , \wAMid30[22] , \wAMid30[21] , \wAMid30[20] , 
        \wAMid30[19] , \wAMid30[18] , \wAMid30[17] , \wAMid30[16] , 
        \wAMid30[15] , \wAMid30[14] , \wAMid30[13] , \wAMid30[12] , 
        \wAMid30[11] , \wAMid30[10] , \wAMid30[9] , \wAMid30[8] , \wAMid30[7] , 
        \wAMid30[6] , \wAMid30[5] , \wAMid30[4] , \wAMid30[3] , \wAMid30[2] , 
        \wAMid30[1] , \wAMid30[0] }), .BIn({\wBMid30[31] , \wBMid30[30] , 
        \wBMid30[29] , \wBMid30[28] , \wBMid30[27] , \wBMid30[26] , 
        \wBMid30[25] , \wBMid30[24] , \wBMid30[23] , \wBMid30[22] , 
        \wBMid30[21] , \wBMid30[20] , \wBMid30[19] , \wBMid30[18] , 
        \wBMid30[17] , \wBMid30[16] , \wBMid30[15] , \wBMid30[14] , 
        \wBMid30[13] , \wBMid30[12] , \wBMid30[11] , \wBMid30[10] , 
        \wBMid30[9] , \wBMid30[8] , \wBMid30[7] , \wBMid30[6] , \wBMid30[5] , 
        \wBMid30[4] , \wBMid30[3] , \wBMid30[2] , \wBMid30[1] , \wBMid30[0] }), 
        .HiOut({\wRegInB30[31] , \wRegInB30[30] , \wRegInB30[29] , 
        \wRegInB30[28] , \wRegInB30[27] , \wRegInB30[26] , \wRegInB30[25] , 
        \wRegInB30[24] , \wRegInB30[23] , \wRegInB30[22] , \wRegInB30[21] , 
        \wRegInB30[20] , \wRegInB30[19] , \wRegInB30[18] , \wRegInB30[17] , 
        \wRegInB30[16] , \wRegInB30[15] , \wRegInB30[14] , \wRegInB30[13] , 
        \wRegInB30[12] , \wRegInB30[11] , \wRegInB30[10] , \wRegInB30[9] , 
        \wRegInB30[8] , \wRegInB30[7] , \wRegInB30[6] , \wRegInB30[5] , 
        \wRegInB30[4] , \wRegInB30[3] , \wRegInB30[2] , \wRegInB30[1] , 
        \wRegInB30[0] }), .LoOut({\wRegInA31[31] , \wRegInA31[30] , 
        \wRegInA31[29] , \wRegInA31[28] , \wRegInA31[27] , \wRegInA31[26] , 
        \wRegInA31[25] , \wRegInA31[24] , \wRegInA31[23] , \wRegInA31[22] , 
        \wRegInA31[21] , \wRegInA31[20] , \wRegInA31[19] , \wRegInA31[18] , 
        \wRegInA31[17] , \wRegInA31[16] , \wRegInA31[15] , \wRegInA31[14] , 
        \wRegInA31[13] , \wRegInA31[12] , \wRegInA31[11] , \wRegInA31[10] , 
        \wRegInA31[9] , \wRegInA31[8] , \wRegInA31[7] , \wRegInA31[6] , 
        \wRegInA31[5] , \wRegInA31[4] , \wRegInA31[3] , \wRegInA31[2] , 
        \wRegInA31[1] , \wRegInA31[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_122 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink123[31] , \ScanLink123[30] , \ScanLink123[29] , 
        \ScanLink123[28] , \ScanLink123[27] , \ScanLink123[26] , 
        \ScanLink123[25] , \ScanLink123[24] , \ScanLink123[23] , 
        \ScanLink123[22] , \ScanLink123[21] , \ScanLink123[20] , 
        \ScanLink123[19] , \ScanLink123[18] , \ScanLink123[17] , 
        \ScanLink123[16] , \ScanLink123[15] , \ScanLink123[14] , 
        \ScanLink123[13] , \ScanLink123[12] , \ScanLink123[11] , 
        \ScanLink123[10] , \ScanLink123[9] , \ScanLink123[8] , 
        \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , \ScanLink123[4] , 
        \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , \ScanLink123[0] 
        }), .ScanOut({\ScanLink122[31] , \ScanLink122[30] , \ScanLink122[29] , 
        \ScanLink122[28] , \ScanLink122[27] , \ScanLink122[26] , 
        \ScanLink122[25] , \ScanLink122[24] , \ScanLink122[23] , 
        \ScanLink122[22] , \ScanLink122[21] , \ScanLink122[20] , 
        \ScanLink122[19] , \ScanLink122[18] , \ScanLink122[17] , 
        \ScanLink122[16] , \ScanLink122[15] , \ScanLink122[14] , 
        \ScanLink122[13] , \ScanLink122[12] , \ScanLink122[11] , 
        \ScanLink122[10] , \ScanLink122[9] , \ScanLink122[8] , 
        \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , \ScanLink122[4] , 
        \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , \ScanLink122[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB66[31] , \wRegInB66[30] , \wRegInB66[29] , 
        \wRegInB66[28] , \wRegInB66[27] , \wRegInB66[26] , \wRegInB66[25] , 
        \wRegInB66[24] , \wRegInB66[23] , \wRegInB66[22] , \wRegInB66[21] , 
        \wRegInB66[20] , \wRegInB66[19] , \wRegInB66[18] , \wRegInB66[17] , 
        \wRegInB66[16] , \wRegInB66[15] , \wRegInB66[14] , \wRegInB66[13] , 
        \wRegInB66[12] , \wRegInB66[11] , \wRegInB66[10] , \wRegInB66[9] , 
        \wRegInB66[8] , \wRegInB66[7] , \wRegInB66[6] , \wRegInB66[5] , 
        \wRegInB66[4] , \wRegInB66[3] , \wRegInB66[2] , \wRegInB66[1] , 
        \wRegInB66[0] }), .Out({\wBIn66[31] , \wBIn66[30] , \wBIn66[29] , 
        \wBIn66[28] , \wBIn66[27] , \wBIn66[26] , \wBIn66[25] , \wBIn66[24] , 
        \wBIn66[23] , \wBIn66[22] , \wBIn66[21] , \wBIn66[20] , \wBIn66[19] , 
        \wBIn66[18] , \wBIn66[17] , \wBIn66[16] , \wBIn66[15] , \wBIn66[14] , 
        \wBIn66[13] , \wBIn66[12] , \wBIn66[11] , \wBIn66[10] , \wBIn66[9] , 
        \wBIn66[8] , \wBIn66[7] , \wBIn66[6] , \wBIn66[5] , \wBIn66[4] , 
        \wBIn66[3] , \wBIn66[2] , \wBIn66[1] , \wBIn66[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid114[31] , \wAMid114[30] , \wAMid114[29] , \wAMid114[28] , 
        \wAMid114[27] , \wAMid114[26] , \wAMid114[25] , \wAMid114[24] , 
        \wAMid114[23] , \wAMid114[22] , \wAMid114[21] , \wAMid114[20] , 
        \wAMid114[19] , \wAMid114[18] , \wAMid114[17] , \wAMid114[16] , 
        \wAMid114[15] , \wAMid114[14] , \wAMid114[13] , \wAMid114[12] , 
        \wAMid114[11] , \wAMid114[10] , \wAMid114[9] , \wAMid114[8] , 
        \wAMid114[7] , \wAMid114[6] , \wAMid114[5] , \wAMid114[4] , 
        \wAMid114[3] , \wAMid114[2] , \wAMid114[1] , \wAMid114[0] }), .BIn({
        \wBMid114[31] , \wBMid114[30] , \wBMid114[29] , \wBMid114[28] , 
        \wBMid114[27] , \wBMid114[26] , \wBMid114[25] , \wBMid114[24] , 
        \wBMid114[23] , \wBMid114[22] , \wBMid114[21] , \wBMid114[20] , 
        \wBMid114[19] , \wBMid114[18] , \wBMid114[17] , \wBMid114[16] , 
        \wBMid114[15] , \wBMid114[14] , \wBMid114[13] , \wBMid114[12] , 
        \wBMid114[11] , \wBMid114[10] , \wBMid114[9] , \wBMid114[8] , 
        \wBMid114[7] , \wBMid114[6] , \wBMid114[5] , \wBMid114[4] , 
        \wBMid114[3] , \wBMid114[2] , \wBMid114[1] , \wBMid114[0] }), .HiOut({
        \wRegInB114[31] , \wRegInB114[30] , \wRegInB114[29] , \wRegInB114[28] , 
        \wRegInB114[27] , \wRegInB114[26] , \wRegInB114[25] , \wRegInB114[24] , 
        \wRegInB114[23] , \wRegInB114[22] , \wRegInB114[21] , \wRegInB114[20] , 
        \wRegInB114[19] , \wRegInB114[18] , \wRegInB114[17] , \wRegInB114[16] , 
        \wRegInB114[15] , \wRegInB114[14] , \wRegInB114[13] , \wRegInB114[12] , 
        \wRegInB114[11] , \wRegInB114[10] , \wRegInB114[9] , \wRegInB114[8] , 
        \wRegInB114[7] , \wRegInB114[6] , \wRegInB114[5] , \wRegInB114[4] , 
        \wRegInB114[3] , \wRegInB114[2] , \wRegInB114[1] , \wRegInB114[0] }), 
        .LoOut({\wRegInA115[31] , \wRegInA115[30] , \wRegInA115[29] , 
        \wRegInA115[28] , \wRegInA115[27] , \wRegInA115[26] , \wRegInA115[25] , 
        \wRegInA115[24] , \wRegInA115[23] , \wRegInA115[22] , \wRegInA115[21] , 
        \wRegInA115[20] , \wRegInA115[19] , \wRegInA115[18] , \wRegInA115[17] , 
        \wRegInA115[16] , \wRegInA115[15] , \wRegInA115[14] , \wRegInA115[13] , 
        \wRegInA115[12] , \wRegInA115[11] , \wRegInA115[10] , \wRegInA115[9] , 
        \wRegInA115[8] , \wRegInA115[7] , \wRegInA115[6] , \wRegInA115[5] , 
        \wRegInA115[4] , \wRegInA115[3] , \wRegInA115[2] , \wRegInA115[1] , 
        \wRegInA115[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_235 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink236[31] , \ScanLink236[30] , \ScanLink236[29] , 
        \ScanLink236[28] , \ScanLink236[27] , \ScanLink236[26] , 
        \ScanLink236[25] , \ScanLink236[24] , \ScanLink236[23] , 
        \ScanLink236[22] , \ScanLink236[21] , \ScanLink236[20] , 
        \ScanLink236[19] , \ScanLink236[18] , \ScanLink236[17] , 
        \ScanLink236[16] , \ScanLink236[15] , \ScanLink236[14] , 
        \ScanLink236[13] , \ScanLink236[12] , \ScanLink236[11] , 
        \ScanLink236[10] , \ScanLink236[9] , \ScanLink236[8] , 
        \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , \ScanLink236[4] , 
        \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , \ScanLink236[0] 
        }), .ScanOut({\ScanLink235[31] , \ScanLink235[30] , \ScanLink235[29] , 
        \ScanLink235[28] , \ScanLink235[27] , \ScanLink235[26] , 
        \ScanLink235[25] , \ScanLink235[24] , \ScanLink235[23] , 
        \ScanLink235[22] , \ScanLink235[21] , \ScanLink235[20] , 
        \ScanLink235[19] , \ScanLink235[18] , \ScanLink235[17] , 
        \ScanLink235[16] , \ScanLink235[15] , \ScanLink235[14] , 
        \ScanLink235[13] , \ScanLink235[12] , \ScanLink235[11] , 
        \ScanLink235[10] , \ScanLink235[9] , \ScanLink235[8] , 
        \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , \ScanLink235[4] , 
        \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , \ScanLink235[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA10[31] , \wRegInA10[30] , \wRegInA10[29] , 
        \wRegInA10[28] , \wRegInA10[27] , \wRegInA10[26] , \wRegInA10[25] , 
        \wRegInA10[24] , \wRegInA10[23] , \wRegInA10[22] , \wRegInA10[21] , 
        \wRegInA10[20] , \wRegInA10[19] , \wRegInA10[18] , \wRegInA10[17] , 
        \wRegInA10[16] , \wRegInA10[15] , \wRegInA10[14] , \wRegInA10[13] , 
        \wRegInA10[12] , \wRegInA10[11] , \wRegInA10[10] , \wRegInA10[9] , 
        \wRegInA10[8] , \wRegInA10[7] , \wRegInA10[6] , \wRegInA10[5] , 
        \wRegInA10[4] , \wRegInA10[3] , \wRegInA10[2] , \wRegInA10[1] , 
        \wRegInA10[0] }), .Out({\wAIn10[31] , \wAIn10[30] , \wAIn10[29] , 
        \wAIn10[28] , \wAIn10[27] , \wAIn10[26] , \wAIn10[25] , \wAIn10[24] , 
        \wAIn10[23] , \wAIn10[22] , \wAIn10[21] , \wAIn10[20] , \wAIn10[19] , 
        \wAIn10[18] , \wAIn10[17] , \wAIn10[16] , \wAIn10[15] , \wAIn10[14] , 
        \wAIn10[13] , \wAIn10[12] , \wAIn10[11] , \wAIn10[10] , \wAIn10[9] , 
        \wAIn10[8] , \wAIn10[7] , \wAIn10[6] , \wAIn10[5] , \wAIn10[4] , 
        \wAIn10[3] , \wAIn10[2] , \wAIn10[1] , \wAIn10[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_105 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink106[31] , \ScanLink106[30] , \ScanLink106[29] , 
        \ScanLink106[28] , \ScanLink106[27] , \ScanLink106[26] , 
        \ScanLink106[25] , \ScanLink106[24] , \ScanLink106[23] , 
        \ScanLink106[22] , \ScanLink106[21] , \ScanLink106[20] , 
        \ScanLink106[19] , \ScanLink106[18] , \ScanLink106[17] , 
        \ScanLink106[16] , \ScanLink106[15] , \ScanLink106[14] , 
        \ScanLink106[13] , \ScanLink106[12] , \ScanLink106[11] , 
        \ScanLink106[10] , \ScanLink106[9] , \ScanLink106[8] , 
        \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , \ScanLink106[4] , 
        \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , \ScanLink106[0] 
        }), .ScanOut({\ScanLink105[31] , \ScanLink105[30] , \ScanLink105[29] , 
        \ScanLink105[28] , \ScanLink105[27] , \ScanLink105[26] , 
        \ScanLink105[25] , \ScanLink105[24] , \ScanLink105[23] , 
        \ScanLink105[22] , \ScanLink105[21] , \ScanLink105[20] , 
        \ScanLink105[19] , \ScanLink105[18] , \ScanLink105[17] , 
        \ScanLink105[16] , \ScanLink105[15] , \ScanLink105[14] , 
        \ScanLink105[13] , \ScanLink105[12] , \ScanLink105[11] , 
        \ScanLink105[10] , \ScanLink105[9] , \ScanLink105[8] , 
        \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , \ScanLink105[4] , 
        \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , \ScanLink105[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA75[31] , \wRegInA75[30] , \wRegInA75[29] , 
        \wRegInA75[28] , \wRegInA75[27] , \wRegInA75[26] , \wRegInA75[25] , 
        \wRegInA75[24] , \wRegInA75[23] , \wRegInA75[22] , \wRegInA75[21] , 
        \wRegInA75[20] , \wRegInA75[19] , \wRegInA75[18] , \wRegInA75[17] , 
        \wRegInA75[16] , \wRegInA75[15] , \wRegInA75[14] , \wRegInA75[13] , 
        \wRegInA75[12] , \wRegInA75[11] , \wRegInA75[10] , \wRegInA75[9] , 
        \wRegInA75[8] , \wRegInA75[7] , \wRegInA75[6] , \wRegInA75[5] , 
        \wRegInA75[4] , \wRegInA75[3] , \wRegInA75[2] , \wRegInA75[1] , 
        \wRegInA75[0] }), .Out({\wAIn75[31] , \wAIn75[30] , \wAIn75[29] , 
        \wAIn75[28] , \wAIn75[27] , \wAIn75[26] , \wAIn75[25] , \wAIn75[24] , 
        \wAIn75[23] , \wAIn75[22] , \wAIn75[21] , \wAIn75[20] , \wAIn75[19] , 
        \wAIn75[18] , \wAIn75[17] , \wAIn75[16] , \wAIn75[15] , \wAIn75[14] , 
        \wAIn75[13] , \wAIn75[12] , \wAIn75[11] , \wAIn75[10] , \wAIn75[9] , 
        \wAIn75[8] , \wAIn75[7] , \wAIn75[6] , \wAIn75[5] , \wAIn75[4] , 
        \wAIn75[3] , \wAIn75[2] , \wAIn75[1] , \wAIn75[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_55 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink56[31] , \ScanLink56[30] , \ScanLink56[29] , 
        \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , \ScanLink56[25] , 
        \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , \ScanLink56[21] , 
        \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , \ScanLink56[17] , 
        \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , \ScanLink56[13] , 
        \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , \ScanLink56[9] , 
        \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , \ScanLink56[5] , 
        \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , \ScanLink56[1] , 
        \ScanLink56[0] }), .ScanOut({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA100[31] , \wRegInA100[30] , 
        \wRegInA100[29] , \wRegInA100[28] , \wRegInA100[27] , \wRegInA100[26] , 
        \wRegInA100[25] , \wRegInA100[24] , \wRegInA100[23] , \wRegInA100[22] , 
        \wRegInA100[21] , \wRegInA100[20] , \wRegInA100[19] , \wRegInA100[18] , 
        \wRegInA100[17] , \wRegInA100[16] , \wRegInA100[15] , \wRegInA100[14] , 
        \wRegInA100[13] , \wRegInA100[12] , \wRegInA100[11] , \wRegInA100[10] , 
        \wRegInA100[9] , \wRegInA100[8] , \wRegInA100[7] , \wRegInA100[6] , 
        \wRegInA100[5] , \wRegInA100[4] , \wRegInA100[3] , \wRegInA100[2] , 
        \wRegInA100[1] , \wRegInA100[0] }), .Out({\wAIn100[31] , \wAIn100[30] , 
        \wAIn100[29] , \wAIn100[28] , \wAIn100[27] , \wAIn100[26] , 
        \wAIn100[25] , \wAIn100[24] , \wAIn100[23] , \wAIn100[22] , 
        \wAIn100[21] , \wAIn100[20] , \wAIn100[19] , \wAIn100[18] , 
        \wAIn100[17] , \wAIn100[16] , \wAIn100[15] , \wAIn100[14] , 
        \wAIn100[13] , \wAIn100[12] , \wAIn100[11] , \wAIn100[10] , 
        \wAIn100[9] , \wAIn100[8] , \wAIn100[7] , \wAIn100[6] , \wAIn100[5] , 
        \wAIn100[4] , \wAIn100[3] , \wAIn100[2] , \wAIn100[1] , \wAIn100[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_97 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink98[31] , \ScanLink98[30] , \ScanLink98[29] , 
        \ScanLink98[28] , \ScanLink98[27] , \ScanLink98[26] , \ScanLink98[25] , 
        \ScanLink98[24] , \ScanLink98[23] , \ScanLink98[22] , \ScanLink98[21] , 
        \ScanLink98[20] , \ScanLink98[19] , \ScanLink98[18] , \ScanLink98[17] , 
        \ScanLink98[16] , \ScanLink98[15] , \ScanLink98[14] , \ScanLink98[13] , 
        \ScanLink98[12] , \ScanLink98[11] , \ScanLink98[10] , \ScanLink98[9] , 
        \ScanLink98[8] , \ScanLink98[7] , \ScanLink98[6] , \ScanLink98[5] , 
        \ScanLink98[4] , \ScanLink98[3] , \ScanLink98[2] , \ScanLink98[1] , 
        \ScanLink98[0] }), .ScanOut({\ScanLink97[31] , \ScanLink97[30] , 
        \ScanLink97[29] , \ScanLink97[28] , \ScanLink97[27] , \ScanLink97[26] , 
        \ScanLink97[25] , \ScanLink97[24] , \ScanLink97[23] , \ScanLink97[22] , 
        \ScanLink97[21] , \ScanLink97[20] , \ScanLink97[19] , \ScanLink97[18] , 
        \ScanLink97[17] , \ScanLink97[16] , \ScanLink97[15] , \ScanLink97[14] , 
        \ScanLink97[13] , \ScanLink97[12] , \ScanLink97[11] , \ScanLink97[10] , 
        \ScanLink97[9] , \ScanLink97[8] , \ScanLink97[7] , \ScanLink97[6] , 
        \ScanLink97[5] , \ScanLink97[4] , \ScanLink97[3] , \ScanLink97[2] , 
        \ScanLink97[1] , \ScanLink97[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA79[31] , \wRegInA79[30] , 
        \wRegInA79[29] , \wRegInA79[28] , \wRegInA79[27] , \wRegInA79[26] , 
        \wRegInA79[25] , \wRegInA79[24] , \wRegInA79[23] , \wRegInA79[22] , 
        \wRegInA79[21] , \wRegInA79[20] , \wRegInA79[19] , \wRegInA79[18] , 
        \wRegInA79[17] , \wRegInA79[16] , \wRegInA79[15] , \wRegInA79[14] , 
        \wRegInA79[13] , \wRegInA79[12] , \wRegInA79[11] , \wRegInA79[10] , 
        \wRegInA79[9] , \wRegInA79[8] , \wRegInA79[7] , \wRegInA79[6] , 
        \wRegInA79[5] , \wRegInA79[4] , \wRegInA79[3] , \wRegInA79[2] , 
        \wRegInA79[1] , \wRegInA79[0] }), .Out({\wAIn79[31] , \wAIn79[30] , 
        \wAIn79[29] , \wAIn79[28] , \wAIn79[27] , \wAIn79[26] , \wAIn79[25] , 
        \wAIn79[24] , \wAIn79[23] , \wAIn79[22] , \wAIn79[21] , \wAIn79[20] , 
        \wAIn79[19] , \wAIn79[18] , \wAIn79[17] , \wAIn79[16] , \wAIn79[15] , 
        \wAIn79[14] , \wAIn79[13] , \wAIn79[12] , \wAIn79[11] , \wAIn79[10] , 
        \wAIn79[9] , \wAIn79[8] , \wAIn79[7] , \wAIn79[6] , \wAIn79[5] , 
        \wAIn79[4] , \wAIn79[3] , \wAIn79[2] , \wAIn79[1] , \wAIn79[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn52[31] , \wAIn52[30] , \wAIn52[29] , \wAIn52[28] , \wAIn52[27] , 
        \wAIn52[26] , \wAIn52[25] , \wAIn52[24] , \wAIn52[23] , \wAIn52[22] , 
        \wAIn52[21] , \wAIn52[20] , \wAIn52[19] , \wAIn52[18] , \wAIn52[17] , 
        \wAIn52[16] , \wAIn52[15] , \wAIn52[14] , \wAIn52[13] , \wAIn52[12] , 
        \wAIn52[11] , \wAIn52[10] , \wAIn52[9] , \wAIn52[8] , \wAIn52[7] , 
        \wAIn52[6] , \wAIn52[5] , \wAIn52[4] , \wAIn52[3] , \wAIn52[2] , 
        \wAIn52[1] , \wAIn52[0] }), .BIn({\wBIn52[31] , \wBIn52[30] , 
        \wBIn52[29] , \wBIn52[28] , \wBIn52[27] , \wBIn52[26] , \wBIn52[25] , 
        \wBIn52[24] , \wBIn52[23] , \wBIn52[22] , \wBIn52[21] , \wBIn52[20] , 
        \wBIn52[19] , \wBIn52[18] , \wBIn52[17] , \wBIn52[16] , \wBIn52[15] , 
        \wBIn52[14] , \wBIn52[13] , \wBIn52[12] , \wBIn52[11] , \wBIn52[10] , 
        \wBIn52[9] , \wBIn52[8] , \wBIn52[7] , \wBIn52[6] , \wBIn52[5] , 
        \wBIn52[4] , \wBIn52[3] , \wBIn52[2] , \wBIn52[1] , \wBIn52[0] }), 
        .HiOut({\wBMid51[31] , \wBMid51[30] , \wBMid51[29] , \wBMid51[28] , 
        \wBMid51[27] , \wBMid51[26] , \wBMid51[25] , \wBMid51[24] , 
        \wBMid51[23] , \wBMid51[22] , \wBMid51[21] , \wBMid51[20] , 
        \wBMid51[19] , \wBMid51[18] , \wBMid51[17] , \wBMid51[16] , 
        \wBMid51[15] , \wBMid51[14] , \wBMid51[13] , \wBMid51[12] , 
        \wBMid51[11] , \wBMid51[10] , \wBMid51[9] , \wBMid51[8] , \wBMid51[7] , 
        \wBMid51[6] , \wBMid51[5] , \wBMid51[4] , \wBMid51[3] , \wBMid51[2] , 
        \wBMid51[1] , \wBMid51[0] }), .LoOut({\wAMid52[31] , \wAMid52[30] , 
        \wAMid52[29] , \wAMid52[28] , \wAMid52[27] , \wAMid52[26] , 
        \wAMid52[25] , \wAMid52[24] , \wAMid52[23] , \wAMid52[22] , 
        \wAMid52[21] , \wAMid52[20] , \wAMid52[19] , \wAMid52[18] , 
        \wAMid52[17] , \wAMid52[16] , \wAMid52[15] , \wAMid52[14] , 
        \wAMid52[13] , \wAMid52[12] , \wAMid52[11] , \wAMid52[10] , 
        \wAMid52[9] , \wAMid52[8] , \wAMid52[7] , \wAMid52[6] , \wAMid52[5] , 
        \wAMid52[4] , \wAMid52[3] , \wAMid52[2] , \wAMid52[1] , \wAMid52[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid62[31] , \wAMid62[30] , \wAMid62[29] , \wAMid62[28] , 
        \wAMid62[27] , \wAMid62[26] , \wAMid62[25] , \wAMid62[24] , 
        \wAMid62[23] , \wAMid62[22] , \wAMid62[21] , \wAMid62[20] , 
        \wAMid62[19] , \wAMid62[18] , \wAMid62[17] , \wAMid62[16] , 
        \wAMid62[15] , \wAMid62[14] , \wAMid62[13] , \wAMid62[12] , 
        \wAMid62[11] , \wAMid62[10] , \wAMid62[9] , \wAMid62[8] , \wAMid62[7] , 
        \wAMid62[6] , \wAMid62[5] , \wAMid62[4] , \wAMid62[3] , \wAMid62[2] , 
        \wAMid62[1] , \wAMid62[0] }), .BIn({\wBMid62[31] , \wBMid62[30] , 
        \wBMid62[29] , \wBMid62[28] , \wBMid62[27] , \wBMid62[26] , 
        \wBMid62[25] , \wBMid62[24] , \wBMid62[23] , \wBMid62[22] , 
        \wBMid62[21] , \wBMid62[20] , \wBMid62[19] , \wBMid62[18] , 
        \wBMid62[17] , \wBMid62[16] , \wBMid62[15] , \wBMid62[14] , 
        \wBMid62[13] , \wBMid62[12] , \wBMid62[11] , \wBMid62[10] , 
        \wBMid62[9] , \wBMid62[8] , \wBMid62[7] , \wBMid62[6] , \wBMid62[5] , 
        \wBMid62[4] , \wBMid62[3] , \wBMid62[2] , \wBMid62[1] , \wBMid62[0] }), 
        .HiOut({\wRegInB62[31] , \wRegInB62[30] , \wRegInB62[29] , 
        \wRegInB62[28] , \wRegInB62[27] , \wRegInB62[26] , \wRegInB62[25] , 
        \wRegInB62[24] , \wRegInB62[23] , \wRegInB62[22] , \wRegInB62[21] , 
        \wRegInB62[20] , \wRegInB62[19] , \wRegInB62[18] , \wRegInB62[17] , 
        \wRegInB62[16] , \wRegInB62[15] , \wRegInB62[14] , \wRegInB62[13] , 
        \wRegInB62[12] , \wRegInB62[11] , \wRegInB62[10] , \wRegInB62[9] , 
        \wRegInB62[8] , \wRegInB62[7] , \wRegInB62[6] , \wRegInB62[5] , 
        \wRegInB62[4] , \wRegInB62[3] , \wRegInB62[2] , \wRegInB62[1] , 
        \wRegInB62[0] }), .LoOut({\wRegInA63[31] , \wRegInA63[30] , 
        \wRegInA63[29] , \wRegInA63[28] , \wRegInA63[27] , \wRegInA63[26] , 
        \wRegInA63[25] , \wRegInA63[24] , \wRegInA63[23] , \wRegInA63[22] , 
        \wRegInA63[21] , \wRegInA63[20] , \wRegInA63[19] , \wRegInA63[18] , 
        \wRegInA63[17] , \wRegInA63[16] , \wRegInA63[15] , \wRegInA63[14] , 
        \wRegInA63[13] , \wRegInA63[12] , \wRegInA63[11] , \wRegInA63[10] , 
        \wRegInA63[9] , \wRegInA63[8] , \wRegInA63[7] , \wRegInA63[6] , 
        \wRegInA63[5] , \wRegInA63[4] , \wRegInA63[3] , \wRegInA63[2] , 
        \wRegInA63[1] , \wRegInA63[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid79[31] , \wAMid79[30] , \wAMid79[29] , \wAMid79[28] , 
        \wAMid79[27] , \wAMid79[26] , \wAMid79[25] , \wAMid79[24] , 
        \wAMid79[23] , \wAMid79[22] , \wAMid79[21] , \wAMid79[20] , 
        \wAMid79[19] , \wAMid79[18] , \wAMid79[17] , \wAMid79[16] , 
        \wAMid79[15] , \wAMid79[14] , \wAMid79[13] , \wAMid79[12] , 
        \wAMid79[11] , \wAMid79[10] , \wAMid79[9] , \wAMid79[8] , \wAMid79[7] , 
        \wAMid79[6] , \wAMid79[5] , \wAMid79[4] , \wAMid79[3] , \wAMid79[2] , 
        \wAMid79[1] , \wAMid79[0] }), .BIn({\wBMid79[31] , \wBMid79[30] , 
        \wBMid79[29] , \wBMid79[28] , \wBMid79[27] , \wBMid79[26] , 
        \wBMid79[25] , \wBMid79[24] , \wBMid79[23] , \wBMid79[22] , 
        \wBMid79[21] , \wBMid79[20] , \wBMid79[19] , \wBMid79[18] , 
        \wBMid79[17] , \wBMid79[16] , \wBMid79[15] , \wBMid79[14] , 
        \wBMid79[13] , \wBMid79[12] , \wBMid79[11] , \wBMid79[10] , 
        \wBMid79[9] , \wBMid79[8] , \wBMid79[7] , \wBMid79[6] , \wBMid79[5] , 
        \wBMid79[4] , \wBMid79[3] , \wBMid79[2] , \wBMid79[1] , \wBMid79[0] }), 
        .HiOut({\wRegInB79[31] , \wRegInB79[30] , \wRegInB79[29] , 
        \wRegInB79[28] , \wRegInB79[27] , \wRegInB79[26] , \wRegInB79[25] , 
        \wRegInB79[24] , \wRegInB79[23] , \wRegInB79[22] , \wRegInB79[21] , 
        \wRegInB79[20] , \wRegInB79[19] , \wRegInB79[18] , \wRegInB79[17] , 
        \wRegInB79[16] , \wRegInB79[15] , \wRegInB79[14] , \wRegInB79[13] , 
        \wRegInB79[12] , \wRegInB79[11] , \wRegInB79[10] , \wRegInB79[9] , 
        \wRegInB79[8] , \wRegInB79[7] , \wRegInB79[6] , \wRegInB79[5] , 
        \wRegInB79[4] , \wRegInB79[3] , \wRegInB79[2] , \wRegInB79[1] , 
        \wRegInB79[0] }), .LoOut({\wRegInA80[31] , \wRegInA80[30] , 
        \wRegInA80[29] , \wRegInA80[28] , \wRegInA80[27] , \wRegInA80[26] , 
        \wRegInA80[25] , \wRegInA80[24] , \wRegInA80[23] , \wRegInA80[22] , 
        \wRegInA80[21] , \wRegInA80[20] , \wRegInA80[19] , \wRegInA80[18] , 
        \wRegInA80[17] , \wRegInA80[16] , \wRegInA80[15] , \wRegInA80[14] , 
        \wRegInA80[13] , \wRegInA80[12] , \wRegInA80[11] , \wRegInA80[10] , 
        \wRegInA80[9] , \wRegInA80[8] , \wRegInA80[7] , \wRegInA80[6] , 
        \wRegInA80[5] , \wRegInA80[4] , \wRegInA80[3] , \wRegInA80[2] , 
        \wRegInA80[1] , \wRegInA80[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_157 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink158[31] , \ScanLink158[30] , \ScanLink158[29] , 
        \ScanLink158[28] , \ScanLink158[27] , \ScanLink158[26] , 
        \ScanLink158[25] , \ScanLink158[24] , \ScanLink158[23] , 
        \ScanLink158[22] , \ScanLink158[21] , \ScanLink158[20] , 
        \ScanLink158[19] , \ScanLink158[18] , \ScanLink158[17] , 
        \ScanLink158[16] , \ScanLink158[15] , \ScanLink158[14] , 
        \ScanLink158[13] , \ScanLink158[12] , \ScanLink158[11] , 
        \ScanLink158[10] , \ScanLink158[9] , \ScanLink158[8] , 
        \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , \ScanLink158[4] , 
        \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , \ScanLink158[0] 
        }), .ScanOut({\ScanLink157[31] , \ScanLink157[30] , \ScanLink157[29] , 
        \ScanLink157[28] , \ScanLink157[27] , \ScanLink157[26] , 
        \ScanLink157[25] , \ScanLink157[24] , \ScanLink157[23] , 
        \ScanLink157[22] , \ScanLink157[21] , \ScanLink157[20] , 
        \ScanLink157[19] , \ScanLink157[18] , \ScanLink157[17] , 
        \ScanLink157[16] , \ScanLink157[15] , \ScanLink157[14] , 
        \ScanLink157[13] , \ScanLink157[12] , \ScanLink157[11] , 
        \ScanLink157[10] , \ScanLink157[9] , \ScanLink157[8] , 
        \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , \ScanLink157[4] , 
        \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , \ScanLink157[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA49[31] , \wRegInA49[30] , \wRegInA49[29] , 
        \wRegInA49[28] , \wRegInA49[27] , \wRegInA49[26] , \wRegInA49[25] , 
        \wRegInA49[24] , \wRegInA49[23] , \wRegInA49[22] , \wRegInA49[21] , 
        \wRegInA49[20] , \wRegInA49[19] , \wRegInA49[18] , \wRegInA49[17] , 
        \wRegInA49[16] , \wRegInA49[15] , \wRegInA49[14] , \wRegInA49[13] , 
        \wRegInA49[12] , \wRegInA49[11] , \wRegInA49[10] , \wRegInA49[9] , 
        \wRegInA49[8] , \wRegInA49[7] , \wRegInA49[6] , \wRegInA49[5] , 
        \wRegInA49[4] , \wRegInA49[3] , \wRegInA49[2] , \wRegInA49[1] , 
        \wRegInA49[0] }), .Out({\wAIn49[31] , \wAIn49[30] , \wAIn49[29] , 
        \wAIn49[28] , \wAIn49[27] , \wAIn49[26] , \wAIn49[25] , \wAIn49[24] , 
        \wAIn49[23] , \wAIn49[22] , \wAIn49[21] , \wAIn49[20] , \wAIn49[19] , 
        \wAIn49[18] , \wAIn49[17] , \wAIn49[16] , \wAIn49[15] , \wAIn49[14] , 
        \wAIn49[13] , \wAIn49[12] , \wAIn49[11] , \wAIn49[10] , \wAIn49[9] , 
        \wAIn49[8] , \wAIn49[7] , \wAIn49[6] , \wAIn49[5] , \wAIn49[4] , 
        \wAIn49[3] , \wAIn49[2] , \wAIn49[1] , \wAIn49[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn55[31] , \wAIn55[30] , \wAIn55[29] , \wAIn55[28] , \wAIn55[27] , 
        \wAIn55[26] , \wAIn55[25] , \wAIn55[24] , \wAIn55[23] , \wAIn55[22] , 
        \wAIn55[21] , \wAIn55[20] , \wAIn55[19] , \wAIn55[18] , \wAIn55[17] , 
        \wAIn55[16] , \wAIn55[15] , \wAIn55[14] , \wAIn55[13] , \wAIn55[12] , 
        \wAIn55[11] , \wAIn55[10] , \wAIn55[9] , \wAIn55[8] , \wAIn55[7] , 
        \wAIn55[6] , \wAIn55[5] , \wAIn55[4] , \wAIn55[3] , \wAIn55[2] , 
        \wAIn55[1] , \wAIn55[0] }), .BIn({\wBIn55[31] , \wBIn55[30] , 
        \wBIn55[29] , \wBIn55[28] , \wBIn55[27] , \wBIn55[26] , \wBIn55[25] , 
        \wBIn55[24] , \wBIn55[23] , \wBIn55[22] , \wBIn55[21] , \wBIn55[20] , 
        \wBIn55[19] , \wBIn55[18] , \wBIn55[17] , \wBIn55[16] , \wBIn55[15] , 
        \wBIn55[14] , \wBIn55[13] , \wBIn55[12] , \wBIn55[11] , \wBIn55[10] , 
        \wBIn55[9] , \wBIn55[8] , \wBIn55[7] , \wBIn55[6] , \wBIn55[5] , 
        \wBIn55[4] , \wBIn55[3] , \wBIn55[2] , \wBIn55[1] , \wBIn55[0] }), 
        .HiOut({\wBMid54[31] , \wBMid54[30] , \wBMid54[29] , \wBMid54[28] , 
        \wBMid54[27] , \wBMid54[26] , \wBMid54[25] , \wBMid54[24] , 
        \wBMid54[23] , \wBMid54[22] , \wBMid54[21] , \wBMid54[20] , 
        \wBMid54[19] , \wBMid54[18] , \wBMid54[17] , \wBMid54[16] , 
        \wBMid54[15] , \wBMid54[14] , \wBMid54[13] , \wBMid54[12] , 
        \wBMid54[11] , \wBMid54[10] , \wBMid54[9] , \wBMid54[8] , \wBMid54[7] , 
        \wBMid54[6] , \wBMid54[5] , \wBMid54[4] , \wBMid54[3] , \wBMid54[2] , 
        \wBMid54[1] , \wBMid54[0] }), .LoOut({\wAMid55[31] , \wAMid55[30] , 
        \wAMid55[29] , \wAMid55[28] , \wAMid55[27] , \wAMid55[26] , 
        \wAMid55[25] , \wAMid55[24] , \wAMid55[23] , \wAMid55[22] , 
        \wAMid55[21] , \wAMid55[20] , \wAMid55[19] , \wAMid55[18] , 
        \wAMid55[17] , \wAMid55[16] , \wAMid55[15] , \wAMid55[14] , 
        \wAMid55[13] , \wAMid55[12] , \wAMid55[11] , \wAMid55[10] , 
        \wAMid55[9] , \wAMid55[8] , \wAMid55[7] , \wAMid55[6] , \wAMid55[5] , 
        \wAMid55[4] , \wAMid55[3] , \wAMid55[2] , \wAMid55[1] , \wAMid55[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn72[31] , \wAIn72[30] , \wAIn72[29] , \wAIn72[28] , \wAIn72[27] , 
        \wAIn72[26] , \wAIn72[25] , \wAIn72[24] , \wAIn72[23] , \wAIn72[22] , 
        \wAIn72[21] , \wAIn72[20] , \wAIn72[19] , \wAIn72[18] , \wAIn72[17] , 
        \wAIn72[16] , \wAIn72[15] , \wAIn72[14] , \wAIn72[13] , \wAIn72[12] , 
        \wAIn72[11] , \wAIn72[10] , \wAIn72[9] , \wAIn72[8] , \wAIn72[7] , 
        \wAIn72[6] , \wAIn72[5] , \wAIn72[4] , \wAIn72[3] , \wAIn72[2] , 
        \wAIn72[1] , \wAIn72[0] }), .BIn({\wBIn72[31] , \wBIn72[30] , 
        \wBIn72[29] , \wBIn72[28] , \wBIn72[27] , \wBIn72[26] , \wBIn72[25] , 
        \wBIn72[24] , \wBIn72[23] , \wBIn72[22] , \wBIn72[21] , \wBIn72[20] , 
        \wBIn72[19] , \wBIn72[18] , \wBIn72[17] , \wBIn72[16] , \wBIn72[15] , 
        \wBIn72[14] , \wBIn72[13] , \wBIn72[12] , \wBIn72[11] , \wBIn72[10] , 
        \wBIn72[9] , \wBIn72[8] , \wBIn72[7] , \wBIn72[6] , \wBIn72[5] , 
        \wBIn72[4] , \wBIn72[3] , \wBIn72[2] , \wBIn72[1] , \wBIn72[0] }), 
        .HiOut({\wBMid71[31] , \wBMid71[30] , \wBMid71[29] , \wBMid71[28] , 
        \wBMid71[27] , \wBMid71[26] , \wBMid71[25] , \wBMid71[24] , 
        \wBMid71[23] , \wBMid71[22] , \wBMid71[21] , \wBMid71[20] , 
        \wBMid71[19] , \wBMid71[18] , \wBMid71[17] , \wBMid71[16] , 
        \wBMid71[15] , \wBMid71[14] , \wBMid71[13] , \wBMid71[12] , 
        \wBMid71[11] , \wBMid71[10] , \wBMid71[9] , \wBMid71[8] , \wBMid71[7] , 
        \wBMid71[6] , \wBMid71[5] , \wBMid71[4] , \wBMid71[3] , \wBMid71[2] , 
        \wBMid71[1] , \wBMid71[0] }), .LoOut({\wAMid72[31] , \wAMid72[30] , 
        \wAMid72[29] , \wAMid72[28] , \wAMid72[27] , \wAMid72[26] , 
        \wAMid72[25] , \wAMid72[24] , \wAMid72[23] , \wAMid72[22] , 
        \wAMid72[21] , \wAMid72[20] , \wAMid72[19] , \wAMid72[18] , 
        \wAMid72[17] , \wAMid72[16] , \wAMid72[15] , \wAMid72[14] , 
        \wAMid72[13] , \wAMid72[12] , \wAMid72[11] , \wAMid72[10] , 
        \wAMid72[9] , \wAMid72[8] , \wAMid72[7] , \wAMid72[6] , \wAMid72[5] , 
        \wAMid72[4] , \wAMid72[3] , \wAMid72[2] , \wAMid72[1] , \wAMid72[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn75[31] , \wAIn75[30] , \wAIn75[29] , \wAIn75[28] , \wAIn75[27] , 
        \wAIn75[26] , \wAIn75[25] , \wAIn75[24] , \wAIn75[23] , \wAIn75[22] , 
        \wAIn75[21] , \wAIn75[20] , \wAIn75[19] , \wAIn75[18] , \wAIn75[17] , 
        \wAIn75[16] , \wAIn75[15] , \wAIn75[14] , \wAIn75[13] , \wAIn75[12] , 
        \wAIn75[11] , \wAIn75[10] , \wAIn75[9] , \wAIn75[8] , \wAIn75[7] , 
        \wAIn75[6] , \wAIn75[5] , \wAIn75[4] , \wAIn75[3] , \wAIn75[2] , 
        \wAIn75[1] , \wAIn75[0] }), .BIn({\wBIn75[31] , \wBIn75[30] , 
        \wBIn75[29] , \wBIn75[28] , \wBIn75[27] , \wBIn75[26] , \wBIn75[25] , 
        \wBIn75[24] , \wBIn75[23] , \wBIn75[22] , \wBIn75[21] , \wBIn75[20] , 
        \wBIn75[19] , \wBIn75[18] , \wBIn75[17] , \wBIn75[16] , \wBIn75[15] , 
        \wBIn75[14] , \wBIn75[13] , \wBIn75[12] , \wBIn75[11] , \wBIn75[10] , 
        \wBIn75[9] , \wBIn75[8] , \wBIn75[7] , \wBIn75[6] , \wBIn75[5] , 
        \wBIn75[4] , \wBIn75[3] , \wBIn75[2] , \wBIn75[1] , \wBIn75[0] }), 
        .HiOut({\wBMid74[31] , \wBMid74[30] , \wBMid74[29] , \wBMid74[28] , 
        \wBMid74[27] , \wBMid74[26] , \wBMid74[25] , \wBMid74[24] , 
        \wBMid74[23] , \wBMid74[22] , \wBMid74[21] , \wBMid74[20] , 
        \wBMid74[19] , \wBMid74[18] , \wBMid74[17] , \wBMid74[16] , 
        \wBMid74[15] , \wBMid74[14] , \wBMid74[13] , \wBMid74[12] , 
        \wBMid74[11] , \wBMid74[10] , \wBMid74[9] , \wBMid74[8] , \wBMid74[7] , 
        \wBMid74[6] , \wBMid74[5] , \wBMid74[4] , \wBMid74[3] , \wBMid74[2] , 
        \wBMid74[1] , \wBMid74[0] }), .LoOut({\wAMid75[31] , \wAMid75[30] , 
        \wAMid75[29] , \wAMid75[28] , \wAMid75[27] , \wAMid75[26] , 
        \wAMid75[25] , \wAMid75[24] , \wAMid75[23] , \wAMid75[22] , 
        \wAMid75[21] , \wAMid75[20] , \wAMid75[19] , \wAMid75[18] , 
        \wAMid75[17] , \wAMid75[16] , \wAMid75[15] , \wAMid75[14] , 
        \wAMid75[13] , \wAMid75[12] , \wAMid75[11] , \wAMid75[10] , 
        \wAMid75[9] , \wAMid75[8] , \wAMid75[7] , \wAMid75[6] , \wAMid75[5] , 
        \wAMid75[4] , \wAMid75[3] , \wAMid75[2] , \wAMid75[1] , \wAMid75[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn105[31] , \wAIn105[30] , \wAIn105[29] , \wAIn105[28] , 
        \wAIn105[27] , \wAIn105[26] , \wAIn105[25] , \wAIn105[24] , 
        \wAIn105[23] , \wAIn105[22] , \wAIn105[21] , \wAIn105[20] , 
        \wAIn105[19] , \wAIn105[18] , \wAIn105[17] , \wAIn105[16] , 
        \wAIn105[15] , \wAIn105[14] , \wAIn105[13] , \wAIn105[12] , 
        \wAIn105[11] , \wAIn105[10] , \wAIn105[9] , \wAIn105[8] , \wAIn105[7] , 
        \wAIn105[6] , \wAIn105[5] , \wAIn105[4] , \wAIn105[3] , \wAIn105[2] , 
        \wAIn105[1] , \wAIn105[0] }), .BIn({\wBIn105[31] , \wBIn105[30] , 
        \wBIn105[29] , \wBIn105[28] , \wBIn105[27] , \wBIn105[26] , 
        \wBIn105[25] , \wBIn105[24] , \wBIn105[23] , \wBIn105[22] , 
        \wBIn105[21] , \wBIn105[20] , \wBIn105[19] , \wBIn105[18] , 
        \wBIn105[17] , \wBIn105[16] , \wBIn105[15] , \wBIn105[14] , 
        \wBIn105[13] , \wBIn105[12] , \wBIn105[11] , \wBIn105[10] , 
        \wBIn105[9] , \wBIn105[8] , \wBIn105[7] , \wBIn105[6] , \wBIn105[5] , 
        \wBIn105[4] , \wBIn105[3] , \wBIn105[2] , \wBIn105[1] , \wBIn105[0] }), 
        .HiOut({\wBMid104[31] , \wBMid104[30] , \wBMid104[29] , \wBMid104[28] , 
        \wBMid104[27] , \wBMid104[26] , \wBMid104[25] , \wBMid104[24] , 
        \wBMid104[23] , \wBMid104[22] , \wBMid104[21] , \wBMid104[20] , 
        \wBMid104[19] , \wBMid104[18] , \wBMid104[17] , \wBMid104[16] , 
        \wBMid104[15] , \wBMid104[14] , \wBMid104[13] , \wBMid104[12] , 
        \wBMid104[11] , \wBMid104[10] , \wBMid104[9] , \wBMid104[8] , 
        \wBMid104[7] , \wBMid104[6] , \wBMid104[5] , \wBMid104[4] , 
        \wBMid104[3] , \wBMid104[2] , \wBMid104[1] , \wBMid104[0] }), .LoOut({
        \wAMid105[31] , \wAMid105[30] , \wAMid105[29] , \wAMid105[28] , 
        \wAMid105[27] , \wAMid105[26] , \wAMid105[25] , \wAMid105[24] , 
        \wAMid105[23] , \wAMid105[22] , \wAMid105[21] , \wAMid105[20] , 
        \wAMid105[19] , \wAMid105[18] , \wAMid105[17] , \wAMid105[16] , 
        \wAMid105[15] , \wAMid105[14] , \wAMid105[13] , \wAMid105[12] , 
        \wAMid105[11] , \wAMid105[10] , \wAMid105[9] , \wAMid105[8] , 
        \wAMid105[7] , \wAMid105[6] , \wAMid105[5] , \wAMid105[4] , 
        \wAMid105[3] , \wAMid105[2] , \wAMid105[1] , \wAMid105[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn122[31] , \wAIn122[30] , \wAIn122[29] , \wAIn122[28] , 
        \wAIn122[27] , \wAIn122[26] , \wAIn122[25] , \wAIn122[24] , 
        \wAIn122[23] , \wAIn122[22] , \wAIn122[21] , \wAIn122[20] , 
        \wAIn122[19] , \wAIn122[18] , \wAIn122[17] , \wAIn122[16] , 
        \wAIn122[15] , \wAIn122[14] , \wAIn122[13] , \wAIn122[12] , 
        \wAIn122[11] , \wAIn122[10] , \wAIn122[9] , \wAIn122[8] , \wAIn122[7] , 
        \wAIn122[6] , \wAIn122[5] , \wAIn122[4] , \wAIn122[3] , \wAIn122[2] , 
        \wAIn122[1] , \wAIn122[0] }), .BIn({\wBIn122[31] , \wBIn122[30] , 
        \wBIn122[29] , \wBIn122[28] , \wBIn122[27] , \wBIn122[26] , 
        \wBIn122[25] , \wBIn122[24] , \wBIn122[23] , \wBIn122[22] , 
        \wBIn122[21] , \wBIn122[20] , \wBIn122[19] , \wBIn122[18] , 
        \wBIn122[17] , \wBIn122[16] , \wBIn122[15] , \wBIn122[14] , 
        \wBIn122[13] , \wBIn122[12] , \wBIn122[11] , \wBIn122[10] , 
        \wBIn122[9] , \wBIn122[8] , \wBIn122[7] , \wBIn122[6] , \wBIn122[5] , 
        \wBIn122[4] , \wBIn122[3] , \wBIn122[2] , \wBIn122[1] , \wBIn122[0] }), 
        .HiOut({\wBMid121[31] , \wBMid121[30] , \wBMid121[29] , \wBMid121[28] , 
        \wBMid121[27] , \wBMid121[26] , \wBMid121[25] , \wBMid121[24] , 
        \wBMid121[23] , \wBMid121[22] , \wBMid121[21] , \wBMid121[20] , 
        \wBMid121[19] , \wBMid121[18] , \wBMid121[17] , \wBMid121[16] , 
        \wBMid121[15] , \wBMid121[14] , \wBMid121[13] , \wBMid121[12] , 
        \wBMid121[11] , \wBMid121[10] , \wBMid121[9] , \wBMid121[8] , 
        \wBMid121[7] , \wBMid121[6] , \wBMid121[5] , \wBMid121[4] , 
        \wBMid121[3] , \wBMid121[2] , \wBMid121[1] , \wBMid121[0] }), .LoOut({
        \wAMid122[31] , \wAMid122[30] , \wAMid122[29] , \wAMid122[28] , 
        \wAMid122[27] , \wAMid122[26] , \wAMid122[25] , \wAMid122[24] , 
        \wAMid122[23] , \wAMid122[22] , \wAMid122[21] , \wAMid122[20] , 
        \wAMid122[19] , \wAMid122[18] , \wAMid122[17] , \wAMid122[16] , 
        \wAMid122[15] , \wAMid122[14] , \wAMid122[13] , \wAMid122[12] , 
        \wAMid122[11] , \wAMid122[10] , \wAMid122[9] , \wAMid122[8] , 
        \wAMid122[7] , \wAMid122[6] , \wAMid122[5] , \wAMid122[4] , 
        \wAMid122[3] , \wAMid122[2] , \wAMid122[1] , \wAMid122[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_240 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink241[31] , \ScanLink241[30] , \ScanLink241[29] , 
        \ScanLink241[28] , \ScanLink241[27] , \ScanLink241[26] , 
        \ScanLink241[25] , \ScanLink241[24] , \ScanLink241[23] , 
        \ScanLink241[22] , \ScanLink241[21] , \ScanLink241[20] , 
        \ScanLink241[19] , \ScanLink241[18] , \ScanLink241[17] , 
        \ScanLink241[16] , \ScanLink241[15] , \ScanLink241[14] , 
        \ScanLink241[13] , \ScanLink241[12] , \ScanLink241[11] , 
        \ScanLink241[10] , \ScanLink241[9] , \ScanLink241[8] , 
        \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , \ScanLink241[4] , 
        \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , \ScanLink241[0] 
        }), .ScanOut({\ScanLink240[31] , \ScanLink240[30] , \ScanLink240[29] , 
        \ScanLink240[28] , \ScanLink240[27] , \ScanLink240[26] , 
        \ScanLink240[25] , \ScanLink240[24] , \ScanLink240[23] , 
        \ScanLink240[22] , \ScanLink240[21] , \ScanLink240[20] , 
        \ScanLink240[19] , \ScanLink240[18] , \ScanLink240[17] , 
        \ScanLink240[16] , \ScanLink240[15] , \ScanLink240[14] , 
        \ScanLink240[13] , \ScanLink240[12] , \ScanLink240[11] , 
        \ScanLink240[10] , \ScanLink240[9] , \ScanLink240[8] , 
        \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , \ScanLink240[4] , 
        \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , \ScanLink240[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB7[31] , \wRegInB7[30] , \wRegInB7[29] , \wRegInB7[28] , 
        \wRegInB7[27] , \wRegInB7[26] , \wRegInB7[25] , \wRegInB7[24] , 
        \wRegInB7[23] , \wRegInB7[22] , \wRegInB7[21] , \wRegInB7[20] , 
        \wRegInB7[19] , \wRegInB7[18] , \wRegInB7[17] , \wRegInB7[16] , 
        \wRegInB7[15] , \wRegInB7[14] , \wRegInB7[13] , \wRegInB7[12] , 
        \wRegInB7[11] , \wRegInB7[10] , \wRegInB7[9] , \wRegInB7[8] , 
        \wRegInB7[7] , \wRegInB7[6] , \wRegInB7[5] , \wRegInB7[4] , 
        \wRegInB7[3] , \wRegInB7[2] , \wRegInB7[1] , \wRegInB7[0] }), .Out({
        \wBIn7[31] , \wBIn7[30] , \wBIn7[29] , \wBIn7[28] , \wBIn7[27] , 
        \wBIn7[26] , \wBIn7[25] , \wBIn7[24] , \wBIn7[23] , \wBIn7[22] , 
        \wBIn7[21] , \wBIn7[20] , \wBIn7[19] , \wBIn7[18] , \wBIn7[17] , 
        \wBIn7[16] , \wBIn7[15] , \wBIn7[14] , \wBIn7[13] , \wBIn7[12] , 
        \wBIn7[11] , \wBIn7[10] , \wBIn7[9] , \wBIn7[8] , \wBIn7[7] , 
        \wBIn7[6] , \wBIn7[5] , \wBIn7[4] , \wBIn7[3] , \wBIn7[2] , \wBIn7[1] , 
        \wBIn7[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid45[31] , \wAMid45[30] , \wAMid45[29] , \wAMid45[28] , 
        \wAMid45[27] , \wAMid45[26] , \wAMid45[25] , \wAMid45[24] , 
        \wAMid45[23] , \wAMid45[22] , \wAMid45[21] , \wAMid45[20] , 
        \wAMid45[19] , \wAMid45[18] , \wAMid45[17] , \wAMid45[16] , 
        \wAMid45[15] , \wAMid45[14] , \wAMid45[13] , \wAMid45[12] , 
        \wAMid45[11] , \wAMid45[10] , \wAMid45[9] , \wAMid45[8] , \wAMid45[7] , 
        \wAMid45[6] , \wAMid45[5] , \wAMid45[4] , \wAMid45[3] , \wAMid45[2] , 
        \wAMid45[1] , \wAMid45[0] }), .BIn({\wBMid45[31] , \wBMid45[30] , 
        \wBMid45[29] , \wBMid45[28] , \wBMid45[27] , \wBMid45[26] , 
        \wBMid45[25] , \wBMid45[24] , \wBMid45[23] , \wBMid45[22] , 
        \wBMid45[21] , \wBMid45[20] , \wBMid45[19] , \wBMid45[18] , 
        \wBMid45[17] , \wBMid45[16] , \wBMid45[15] , \wBMid45[14] , 
        \wBMid45[13] , \wBMid45[12] , \wBMid45[11] , \wBMid45[10] , 
        \wBMid45[9] , \wBMid45[8] , \wBMid45[7] , \wBMid45[6] , \wBMid45[5] , 
        \wBMid45[4] , \wBMid45[3] , \wBMid45[2] , \wBMid45[1] , \wBMid45[0] }), 
        .HiOut({\wRegInB45[31] , \wRegInB45[30] , \wRegInB45[29] , 
        \wRegInB45[28] , \wRegInB45[27] , \wRegInB45[26] , \wRegInB45[25] , 
        \wRegInB45[24] , \wRegInB45[23] , \wRegInB45[22] , \wRegInB45[21] , 
        \wRegInB45[20] , \wRegInB45[19] , \wRegInB45[18] , \wRegInB45[17] , 
        \wRegInB45[16] , \wRegInB45[15] , \wRegInB45[14] , \wRegInB45[13] , 
        \wRegInB45[12] , \wRegInB45[11] , \wRegInB45[10] , \wRegInB45[9] , 
        \wRegInB45[8] , \wRegInB45[7] , \wRegInB45[6] , \wRegInB45[5] , 
        \wRegInB45[4] , \wRegInB45[3] , \wRegInB45[2] , \wRegInB45[1] , 
        \wRegInB45[0] }), .LoOut({\wRegInA46[31] , \wRegInA46[30] , 
        \wRegInA46[29] , \wRegInA46[28] , \wRegInA46[27] , \wRegInA46[26] , 
        \wRegInA46[25] , \wRegInA46[24] , \wRegInA46[23] , \wRegInA46[22] , 
        \wRegInA46[21] , \wRegInA46[20] , \wRegInA46[19] , \wRegInA46[18] , 
        \wRegInA46[17] , \wRegInA46[16] , \wRegInA46[15] , \wRegInA46[14] , 
        \wRegInA46[13] , \wRegInA46[12] , \wRegInA46[11] , \wRegInA46[10] , 
        \wRegInA46[9] , \wRegInA46[8] , \wRegInA46[7] , \wRegInA46[6] , 
        \wRegInA46[5] , \wRegInA46[4] , \wRegInA46[3] , \wRegInA46[2] , 
        \wRegInA46[1] , \wRegInA46[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_170 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink171[31] , \ScanLink171[30] , \ScanLink171[29] , 
        \ScanLink171[28] , \ScanLink171[27] , \ScanLink171[26] , 
        \ScanLink171[25] , \ScanLink171[24] , \ScanLink171[23] , 
        \ScanLink171[22] , \ScanLink171[21] , \ScanLink171[20] , 
        \ScanLink171[19] , \ScanLink171[18] , \ScanLink171[17] , 
        \ScanLink171[16] , \ScanLink171[15] , \ScanLink171[14] , 
        \ScanLink171[13] , \ScanLink171[12] , \ScanLink171[11] , 
        \ScanLink171[10] , \ScanLink171[9] , \ScanLink171[8] , 
        \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , \ScanLink171[4] , 
        \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , \ScanLink171[0] 
        }), .ScanOut({\ScanLink170[31] , \ScanLink170[30] , \ScanLink170[29] , 
        \ScanLink170[28] , \ScanLink170[27] , \ScanLink170[26] , 
        \ScanLink170[25] , \ScanLink170[24] , \ScanLink170[23] , 
        \ScanLink170[22] , \ScanLink170[21] , \ScanLink170[20] , 
        \ScanLink170[19] , \ScanLink170[18] , \ScanLink170[17] , 
        \ScanLink170[16] , \ScanLink170[15] , \ScanLink170[14] , 
        \ScanLink170[13] , \ScanLink170[12] , \ScanLink170[11] , 
        \ScanLink170[10] , \ScanLink170[9] , \ScanLink170[8] , 
        \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , \ScanLink170[4] , 
        \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , \ScanLink170[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB42[31] , \wRegInB42[30] , \wRegInB42[29] , 
        \wRegInB42[28] , \wRegInB42[27] , \wRegInB42[26] , \wRegInB42[25] , 
        \wRegInB42[24] , \wRegInB42[23] , \wRegInB42[22] , \wRegInB42[21] , 
        \wRegInB42[20] , \wRegInB42[19] , \wRegInB42[18] , \wRegInB42[17] , 
        \wRegInB42[16] , \wRegInB42[15] , \wRegInB42[14] , \wRegInB42[13] , 
        \wRegInB42[12] , \wRegInB42[11] , \wRegInB42[10] , \wRegInB42[9] , 
        \wRegInB42[8] , \wRegInB42[7] , \wRegInB42[6] , \wRegInB42[5] , 
        \wRegInB42[4] , \wRegInB42[3] , \wRegInB42[2] , \wRegInB42[1] , 
        \wRegInB42[0] }), .Out({\wBIn42[31] , \wBIn42[30] , \wBIn42[29] , 
        \wBIn42[28] , \wBIn42[27] , \wBIn42[26] , \wBIn42[25] , \wBIn42[24] , 
        \wBIn42[23] , \wBIn42[22] , \wBIn42[21] , \wBIn42[20] , \wBIn42[19] , 
        \wBIn42[18] , \wBIn42[17] , \wBIn42[16] , \wBIn42[15] , \wBIn42[14] , 
        \wBIn42[13] , \wBIn42[12] , \wBIn42[11] , \wBIn42[10] , \wBIn42[9] , 
        \wBIn42[8] , \wBIn42[7] , \wBIn42[6] , \wBIn42[5] , \wBIn42[4] , 
        \wBIn42[3] , \wBIn42[2] , \wBIn42[1] , \wBIn42[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_20 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink21[31] , \ScanLink21[30] , \ScanLink21[29] , 
        \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , \ScanLink21[25] , 
        \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , \ScanLink21[21] , 
        \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , \ScanLink21[17] , 
        \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , \ScanLink21[13] , 
        \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , \ScanLink21[9] , 
        \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , \ScanLink21[5] , 
        \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , \ScanLink21[1] , 
        \ScanLink21[0] }), .ScanOut({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB117[31] , \wRegInB117[30] , 
        \wRegInB117[29] , \wRegInB117[28] , \wRegInB117[27] , \wRegInB117[26] , 
        \wRegInB117[25] , \wRegInB117[24] , \wRegInB117[23] , \wRegInB117[22] , 
        \wRegInB117[21] , \wRegInB117[20] , \wRegInB117[19] , \wRegInB117[18] , 
        \wRegInB117[17] , \wRegInB117[16] , \wRegInB117[15] , \wRegInB117[14] , 
        \wRegInB117[13] , \wRegInB117[12] , \wRegInB117[11] , \wRegInB117[10] , 
        \wRegInB117[9] , \wRegInB117[8] , \wRegInB117[7] , \wRegInB117[6] , 
        \wRegInB117[5] , \wRegInB117[4] , \wRegInB117[3] , \wRegInB117[2] , 
        \wRegInB117[1] , \wRegInB117[0] }), .Out({\wBIn117[31] , \wBIn117[30] , 
        \wBIn117[29] , \wBIn117[28] , \wBIn117[27] , \wBIn117[26] , 
        \wBIn117[25] , \wBIn117[24] , \wBIn117[23] , \wBIn117[22] , 
        \wBIn117[21] , \wBIn117[20] , \wBIn117[19] , \wBIn117[18] , 
        \wBIn117[17] , \wBIn117[16] , \wBIn117[15] , \wBIn117[14] , 
        \wBIn117[13] , \wBIn117[12] , \wBIn117[11] , \wBIn117[10] , 
        \wBIn117[9] , \wBIn117[8] , \wBIn117[7] , \wBIn117[6] , \wBIn117[5] , 
        \wBIn117[4] , \wBIn117[3] , \wBIn117[2] , \wBIn117[1] , \wBIn117[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn90[31] , \wAIn90[30] , \wAIn90[29] , \wAIn90[28] , \wAIn90[27] , 
        \wAIn90[26] , \wAIn90[25] , \wAIn90[24] , \wAIn90[23] , \wAIn90[22] , 
        \wAIn90[21] , \wAIn90[20] , \wAIn90[19] , \wAIn90[18] , \wAIn90[17] , 
        \wAIn90[16] , \wAIn90[15] , \wAIn90[14] , \wAIn90[13] , \wAIn90[12] , 
        \wAIn90[11] , \wAIn90[10] , \wAIn90[9] , \wAIn90[8] , \wAIn90[7] , 
        \wAIn90[6] , \wAIn90[5] , \wAIn90[4] , \wAIn90[3] , \wAIn90[2] , 
        \wAIn90[1] , \wAIn90[0] }), .BIn({\wBIn90[31] , \wBIn90[30] , 
        \wBIn90[29] , \wBIn90[28] , \wBIn90[27] , \wBIn90[26] , \wBIn90[25] , 
        \wBIn90[24] , \wBIn90[23] , \wBIn90[22] , \wBIn90[21] , \wBIn90[20] , 
        \wBIn90[19] , \wBIn90[18] , \wBIn90[17] , \wBIn90[16] , \wBIn90[15] , 
        \wBIn90[14] , \wBIn90[13] , \wBIn90[12] , \wBIn90[11] , \wBIn90[10] , 
        \wBIn90[9] , \wBIn90[8] , \wBIn90[7] , \wBIn90[6] , \wBIn90[5] , 
        \wBIn90[4] , \wBIn90[3] , \wBIn90[2] , \wBIn90[1] , \wBIn90[0] }), 
        .HiOut({\wBMid89[31] , \wBMid89[30] , \wBMid89[29] , \wBMid89[28] , 
        \wBMid89[27] , \wBMid89[26] , \wBMid89[25] , \wBMid89[24] , 
        \wBMid89[23] , \wBMid89[22] , \wBMid89[21] , \wBMid89[20] , 
        \wBMid89[19] , \wBMid89[18] , \wBMid89[17] , \wBMid89[16] , 
        \wBMid89[15] , \wBMid89[14] , \wBMid89[13] , \wBMid89[12] , 
        \wBMid89[11] , \wBMid89[10] , \wBMid89[9] , \wBMid89[8] , \wBMid89[7] , 
        \wBMid89[6] , \wBMid89[5] , \wBMid89[4] , \wBMid89[3] , \wBMid89[2] , 
        \wBMid89[1] , \wBMid89[0] }), .LoOut({\wAMid90[31] , \wAMid90[30] , 
        \wAMid90[29] , \wAMid90[28] , \wAMid90[27] , \wAMid90[26] , 
        \wAMid90[25] , \wAMid90[24] , \wAMid90[23] , \wAMid90[22] , 
        \wAMid90[21] , \wAMid90[20] , \wAMid90[19] , \wAMid90[18] , 
        \wAMid90[17] , \wAMid90[16] , \wAMid90[15] , \wAMid90[14] , 
        \wAMid90[13] , \wAMid90[12] , \wAMid90[11] , \wAMid90[10] , 
        \wAMid90[9] , \wAMid90[8] , \wAMid90[7] , \wAMid90[6] , \wAMid90[5] , 
        \wAMid90[4] , \wAMid90[3] , \wAMid90[2] , \wAMid90[1] , \wAMid90[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid1[31] , 
        \wAMid1[30] , \wAMid1[29] , \wAMid1[28] , \wAMid1[27] , \wAMid1[26] , 
        \wAMid1[25] , \wAMid1[24] , \wAMid1[23] , \wAMid1[22] , \wAMid1[21] , 
        \wAMid1[20] , \wAMid1[19] , \wAMid1[18] , \wAMid1[17] , \wAMid1[16] , 
        \wAMid1[15] , \wAMid1[14] , \wAMid1[13] , \wAMid1[12] , \wAMid1[11] , 
        \wAMid1[10] , \wAMid1[9] , \wAMid1[8] , \wAMid1[7] , \wAMid1[6] , 
        \wAMid1[5] , \wAMid1[4] , \wAMid1[3] , \wAMid1[2] , \wAMid1[1] , 
        \wAMid1[0] }), .BIn({\wBMid1[31] , \wBMid1[30] , \wBMid1[29] , 
        \wBMid1[28] , \wBMid1[27] , \wBMid1[26] , \wBMid1[25] , \wBMid1[24] , 
        \wBMid1[23] , \wBMid1[22] , \wBMid1[21] , \wBMid1[20] , \wBMid1[19] , 
        \wBMid1[18] , \wBMid1[17] , \wBMid1[16] , \wBMid1[15] , \wBMid1[14] , 
        \wBMid1[13] , \wBMid1[12] , \wBMid1[11] , \wBMid1[10] , \wBMid1[9] , 
        \wBMid1[8] , \wBMid1[7] , \wBMid1[6] , \wBMid1[5] , \wBMid1[4] , 
        \wBMid1[3] , \wBMid1[2] , \wBMid1[1] , \wBMid1[0] }), .HiOut({
        \wRegInB1[31] , \wRegInB1[30] , \wRegInB1[29] , \wRegInB1[28] , 
        \wRegInB1[27] , \wRegInB1[26] , \wRegInB1[25] , \wRegInB1[24] , 
        \wRegInB1[23] , \wRegInB1[22] , \wRegInB1[21] , \wRegInB1[20] , 
        \wRegInB1[19] , \wRegInB1[18] , \wRegInB1[17] , \wRegInB1[16] , 
        \wRegInB1[15] , \wRegInB1[14] , \wRegInB1[13] , \wRegInB1[12] , 
        \wRegInB1[11] , \wRegInB1[10] , \wRegInB1[9] , \wRegInB1[8] , 
        \wRegInB1[7] , \wRegInB1[6] , \wRegInB1[5] , \wRegInB1[4] , 
        \wRegInB1[3] , \wRegInB1[2] , \wRegInB1[1] , \wRegInB1[0] }), .LoOut({
        \wRegInA2[31] , \wRegInA2[30] , \wRegInA2[29] , \wRegInA2[28] , 
        \wRegInA2[27] , \wRegInA2[26] , \wRegInA2[25] , \wRegInA2[24] , 
        \wRegInA2[23] , \wRegInA2[22] , \wRegInA2[21] , \wRegInA2[20] , 
        \wRegInA2[19] , \wRegInA2[18] , \wRegInA2[17] , \wRegInA2[16] , 
        \wRegInA2[15] , \wRegInA2[14] , \wRegInA2[13] , \wRegInA2[12] , 
        \wRegInA2[11] , \wRegInA2[10] , \wRegInA2[9] , \wRegInA2[8] , 
        \wRegInA2[7] , \wRegInA2[6] , \wRegInA2[5] , \wRegInA2[4] , 
        \wRegInA2[3] , \wRegInA2[2] , \wRegInA2[1] , \wRegInA2[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn97[31] , \wAIn97[30] , \wAIn97[29] , \wAIn97[28] , \wAIn97[27] , 
        \wAIn97[26] , \wAIn97[25] , \wAIn97[24] , \wAIn97[23] , \wAIn97[22] , 
        \wAIn97[21] , \wAIn97[20] , \wAIn97[19] , \wAIn97[18] , \wAIn97[17] , 
        \wAIn97[16] , \wAIn97[15] , \wAIn97[14] , \wAIn97[13] , \wAIn97[12] , 
        \wAIn97[11] , \wAIn97[10] , \wAIn97[9] , \wAIn97[8] , \wAIn97[7] , 
        \wAIn97[6] , \wAIn97[5] , \wAIn97[4] , \wAIn97[3] , \wAIn97[2] , 
        \wAIn97[1] , \wAIn97[0] }), .BIn({\wBIn97[31] , \wBIn97[30] , 
        \wBIn97[29] , \wBIn97[28] , \wBIn97[27] , \wBIn97[26] , \wBIn97[25] , 
        \wBIn97[24] , \wBIn97[23] , \wBIn97[22] , \wBIn97[21] , \wBIn97[20] , 
        \wBIn97[19] , \wBIn97[18] , \wBIn97[17] , \wBIn97[16] , \wBIn97[15] , 
        \wBIn97[14] , \wBIn97[13] , \wBIn97[12] , \wBIn97[11] , \wBIn97[10] , 
        \wBIn97[9] , \wBIn97[8] , \wBIn97[7] , \wBIn97[6] , \wBIn97[5] , 
        \wBIn97[4] , \wBIn97[3] , \wBIn97[2] , \wBIn97[1] , \wBIn97[0] }), 
        .HiOut({\wBMid96[31] , \wBMid96[30] , \wBMid96[29] , \wBMid96[28] , 
        \wBMid96[27] , \wBMid96[26] , \wBMid96[25] , \wBMid96[24] , 
        \wBMid96[23] , \wBMid96[22] , \wBMid96[21] , \wBMid96[20] , 
        \wBMid96[19] , \wBMid96[18] , \wBMid96[17] , \wBMid96[16] , 
        \wBMid96[15] , \wBMid96[14] , \wBMid96[13] , \wBMid96[12] , 
        \wBMid96[11] , \wBMid96[10] , \wBMid96[9] , \wBMid96[8] , \wBMid96[7] , 
        \wBMid96[6] , \wBMid96[5] , \wBMid96[4] , \wBMid96[3] , \wBMid96[2] , 
        \wBMid96[1] , \wBMid96[0] }), .LoOut({\wAMid97[31] , \wAMid97[30] , 
        \wAMid97[29] , \wAMid97[28] , \wAMid97[27] , \wAMid97[26] , 
        \wAMid97[25] , \wAMid97[24] , \wAMid97[23] , \wAMid97[22] , 
        \wAMid97[21] , \wAMid97[20] , \wAMid97[19] , \wAMid97[18] , 
        \wAMid97[17] , \wAMid97[16] , \wAMid97[15] , \wAMid97[14] , 
        \wAMid97[13] , \wAMid97[12] , \wAMid97[11] , \wAMid97[10] , 
        \wAMid97[9] , \wAMid97[8] , \wAMid97[7] , \wAMid97[6] , \wAMid97[5] , 
        \wAMid97[4] , \wAMid97[3] , \wAMid97[2] , \wAMid97[1] , \wAMid97[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid80[31] , \wAMid80[30] , \wAMid80[29] , \wAMid80[28] , 
        \wAMid80[27] , \wAMid80[26] , \wAMid80[25] , \wAMid80[24] , 
        \wAMid80[23] , \wAMid80[22] , \wAMid80[21] , \wAMid80[20] , 
        \wAMid80[19] , \wAMid80[18] , \wAMid80[17] , \wAMid80[16] , 
        \wAMid80[15] , \wAMid80[14] , \wAMid80[13] , \wAMid80[12] , 
        \wAMid80[11] , \wAMid80[10] , \wAMid80[9] , \wAMid80[8] , \wAMid80[7] , 
        \wAMid80[6] , \wAMid80[5] , \wAMid80[4] , \wAMid80[3] , \wAMid80[2] , 
        \wAMid80[1] , \wAMid80[0] }), .BIn({\wBMid80[31] , \wBMid80[30] , 
        \wBMid80[29] , \wBMid80[28] , \wBMid80[27] , \wBMid80[26] , 
        \wBMid80[25] , \wBMid80[24] , \wBMid80[23] , \wBMid80[22] , 
        \wBMid80[21] , \wBMid80[20] , \wBMid80[19] , \wBMid80[18] , 
        \wBMid80[17] , \wBMid80[16] , \wBMid80[15] , \wBMid80[14] , 
        \wBMid80[13] , \wBMid80[12] , \wBMid80[11] , \wBMid80[10] , 
        \wBMid80[9] , \wBMid80[8] , \wBMid80[7] , \wBMid80[6] , \wBMid80[5] , 
        \wBMid80[4] , \wBMid80[3] , \wBMid80[2] , \wBMid80[1] , \wBMid80[0] }), 
        .HiOut({\wRegInB80[31] , \wRegInB80[30] , \wRegInB80[29] , 
        \wRegInB80[28] , \wRegInB80[27] , \wRegInB80[26] , \wRegInB80[25] , 
        \wRegInB80[24] , \wRegInB80[23] , \wRegInB80[22] , \wRegInB80[21] , 
        \wRegInB80[20] , \wRegInB80[19] , \wRegInB80[18] , \wRegInB80[17] , 
        \wRegInB80[16] , \wRegInB80[15] , \wRegInB80[14] , \wRegInB80[13] , 
        \wRegInB80[12] , \wRegInB80[11] , \wRegInB80[10] , \wRegInB80[9] , 
        \wRegInB80[8] , \wRegInB80[7] , \wRegInB80[6] , \wRegInB80[5] , 
        \wRegInB80[4] , \wRegInB80[3] , \wRegInB80[2] , \wRegInB80[1] , 
        \wRegInB80[0] }), .LoOut({\wRegInA81[31] , \wRegInA81[30] , 
        \wRegInA81[29] , \wRegInA81[28] , \wRegInA81[27] , \wRegInA81[26] , 
        \wRegInA81[25] , \wRegInA81[24] , \wRegInA81[23] , \wRegInA81[22] , 
        \wRegInA81[21] , \wRegInA81[20] , \wRegInA81[19] , \wRegInA81[18] , 
        \wRegInA81[17] , \wRegInA81[16] , \wRegInA81[15] , \wRegInA81[14] , 
        \wRegInA81[13] , \wRegInA81[12] , \wRegInA81[11] , \wRegInA81[10] , 
        \wRegInA81[9] , \wRegInA81[8] , \wRegInA81[7] , \wRegInA81[6] , 
        \wRegInA81[5] , \wRegInA81[4] , \wRegInA81[3] , \wRegInA81[2] , 
        \wRegInA81[1] , \wRegInA81[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid87[31] , \wAMid87[30] , \wAMid87[29] , \wAMid87[28] , 
        \wAMid87[27] , \wAMid87[26] , \wAMid87[25] , \wAMid87[24] , 
        \wAMid87[23] , \wAMid87[22] , \wAMid87[21] , \wAMid87[20] , 
        \wAMid87[19] , \wAMid87[18] , \wAMid87[17] , \wAMid87[16] , 
        \wAMid87[15] , \wAMid87[14] , \wAMid87[13] , \wAMid87[12] , 
        \wAMid87[11] , \wAMid87[10] , \wAMid87[9] , \wAMid87[8] , \wAMid87[7] , 
        \wAMid87[6] , \wAMid87[5] , \wAMid87[4] , \wAMid87[3] , \wAMid87[2] , 
        \wAMid87[1] , \wAMid87[0] }), .BIn({\wBMid87[31] , \wBMid87[30] , 
        \wBMid87[29] , \wBMid87[28] , \wBMid87[27] , \wBMid87[26] , 
        \wBMid87[25] , \wBMid87[24] , \wBMid87[23] , \wBMid87[22] , 
        \wBMid87[21] , \wBMid87[20] , \wBMid87[19] , \wBMid87[18] , 
        \wBMid87[17] , \wBMid87[16] , \wBMid87[15] , \wBMid87[14] , 
        \wBMid87[13] , \wBMid87[12] , \wBMid87[11] , \wBMid87[10] , 
        \wBMid87[9] , \wBMid87[8] , \wBMid87[7] , \wBMid87[6] , \wBMid87[5] , 
        \wBMid87[4] , \wBMid87[3] , \wBMid87[2] , \wBMid87[1] , \wBMid87[0] }), 
        .HiOut({\wRegInB87[31] , \wRegInB87[30] , \wRegInB87[29] , 
        \wRegInB87[28] , \wRegInB87[27] , \wRegInB87[26] , \wRegInB87[25] , 
        \wRegInB87[24] , \wRegInB87[23] , \wRegInB87[22] , \wRegInB87[21] , 
        \wRegInB87[20] , \wRegInB87[19] , \wRegInB87[18] , \wRegInB87[17] , 
        \wRegInB87[16] , \wRegInB87[15] , \wRegInB87[14] , \wRegInB87[13] , 
        \wRegInB87[12] , \wRegInB87[11] , \wRegInB87[10] , \wRegInB87[9] , 
        \wRegInB87[8] , \wRegInB87[7] , \wRegInB87[6] , \wRegInB87[5] , 
        \wRegInB87[4] , \wRegInB87[3] , \wRegInB87[2] , \wRegInB87[1] , 
        \wRegInB87[0] }), .LoOut({\wRegInA88[31] , \wRegInA88[30] , 
        \wRegInA88[29] , \wRegInA88[28] , \wRegInA88[27] , \wRegInA88[26] , 
        \wRegInA88[25] , \wRegInA88[24] , \wRegInA88[23] , \wRegInA88[22] , 
        \wRegInA88[21] , \wRegInA88[20] , \wRegInA88[19] , \wRegInA88[18] , 
        \wRegInA88[17] , \wRegInA88[16] , \wRegInA88[15] , \wRegInA88[14] , 
        \wRegInA88[13] , \wRegInA88[12] , \wRegInA88[11] , \wRegInA88[10] , 
        \wRegInA88[9] , \wRegInA88[8] , \wRegInA88[7] , \wRegInA88[6] , 
        \wRegInA88[5] , \wRegInA88[4] , \wRegInA88[3] , \wRegInA88[2] , 
        \wRegInA88[1] , \wRegInA88[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_195 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink196[31] , \ScanLink196[30] , \ScanLink196[29] , 
        \ScanLink196[28] , \ScanLink196[27] , \ScanLink196[26] , 
        \ScanLink196[25] , \ScanLink196[24] , \ScanLink196[23] , 
        \ScanLink196[22] , \ScanLink196[21] , \ScanLink196[20] , 
        \ScanLink196[19] , \ScanLink196[18] , \ScanLink196[17] , 
        \ScanLink196[16] , \ScanLink196[15] , \ScanLink196[14] , 
        \ScanLink196[13] , \ScanLink196[12] , \ScanLink196[11] , 
        \ScanLink196[10] , \ScanLink196[9] , \ScanLink196[8] , 
        \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , \ScanLink196[4] , 
        \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , \ScanLink196[0] 
        }), .ScanOut({\ScanLink195[31] , \ScanLink195[30] , \ScanLink195[29] , 
        \ScanLink195[28] , \ScanLink195[27] , \ScanLink195[26] , 
        \ScanLink195[25] , \ScanLink195[24] , \ScanLink195[23] , 
        \ScanLink195[22] , \ScanLink195[21] , \ScanLink195[20] , 
        \ScanLink195[19] , \ScanLink195[18] , \ScanLink195[17] , 
        \ScanLink195[16] , \ScanLink195[15] , \ScanLink195[14] , 
        \ScanLink195[13] , \ScanLink195[12] , \ScanLink195[11] , 
        \ScanLink195[10] , \ScanLink195[9] , \ScanLink195[8] , 
        \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , \ScanLink195[4] , 
        \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , \ScanLink195[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA30[31] , \wRegInA30[30] , \wRegInA30[29] , 
        \wRegInA30[28] , \wRegInA30[27] , \wRegInA30[26] , \wRegInA30[25] , 
        \wRegInA30[24] , \wRegInA30[23] , \wRegInA30[22] , \wRegInA30[21] , 
        \wRegInA30[20] , \wRegInA30[19] , \wRegInA30[18] , \wRegInA30[17] , 
        \wRegInA30[16] , \wRegInA30[15] , \wRegInA30[14] , \wRegInA30[13] , 
        \wRegInA30[12] , \wRegInA30[11] , \wRegInA30[10] , \wRegInA30[9] , 
        \wRegInA30[8] , \wRegInA30[7] , \wRegInA30[6] , \wRegInA30[5] , 
        \wRegInA30[4] , \wRegInA30[3] , \wRegInA30[2] , \wRegInA30[1] , 
        \wRegInA30[0] }), .Out({\wAIn30[31] , \wAIn30[30] , \wAIn30[29] , 
        \wAIn30[28] , \wAIn30[27] , \wAIn30[26] , \wAIn30[25] , \wAIn30[24] , 
        \wAIn30[23] , \wAIn30[22] , \wAIn30[21] , \wAIn30[20] , \wAIn30[19] , 
        \wAIn30[18] , \wAIn30[17] , \wAIn30[16] , \wAIn30[15] , \wAIn30[14] , 
        \wAIn30[13] , \wAIn30[12] , \wAIn30[11] , \wAIn30[10] , \wAIn30[9] , 
        \wAIn30[8] , \wAIn30[7] , \wAIn30[6] , \wAIn30[5] , \wAIn30[4] , 
        \wAIn30[3] , \wAIn30[2] , \wAIn30[1] , \wAIn30[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_209 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink210[31] , \ScanLink210[30] , \ScanLink210[29] , 
        \ScanLink210[28] , \ScanLink210[27] , \ScanLink210[26] , 
        \ScanLink210[25] , \ScanLink210[24] , \ScanLink210[23] , 
        \ScanLink210[22] , \ScanLink210[21] , \ScanLink210[20] , 
        \ScanLink210[19] , \ScanLink210[18] , \ScanLink210[17] , 
        \ScanLink210[16] , \ScanLink210[15] , \ScanLink210[14] , 
        \ScanLink210[13] , \ScanLink210[12] , \ScanLink210[11] , 
        \ScanLink210[10] , \ScanLink210[9] , \ScanLink210[8] , 
        \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , \ScanLink210[4] , 
        \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , \ScanLink210[0] 
        }), .ScanOut({\ScanLink209[31] , \ScanLink209[30] , \ScanLink209[29] , 
        \ScanLink209[28] , \ScanLink209[27] , \ScanLink209[26] , 
        \ScanLink209[25] , \ScanLink209[24] , \ScanLink209[23] , 
        \ScanLink209[22] , \ScanLink209[21] , \ScanLink209[20] , 
        \ScanLink209[19] , \ScanLink209[18] , \ScanLink209[17] , 
        \ScanLink209[16] , \ScanLink209[15] , \ScanLink209[14] , 
        \ScanLink209[13] , \ScanLink209[12] , \ScanLink209[11] , 
        \ScanLink209[10] , \ScanLink209[9] , \ScanLink209[8] , 
        \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , \ScanLink209[4] , 
        \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , \ScanLink209[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA23[31] , \wRegInA23[30] , \wRegInA23[29] , 
        \wRegInA23[28] , \wRegInA23[27] , \wRegInA23[26] , \wRegInA23[25] , 
        \wRegInA23[24] , \wRegInA23[23] , \wRegInA23[22] , \wRegInA23[21] , 
        \wRegInA23[20] , \wRegInA23[19] , \wRegInA23[18] , \wRegInA23[17] , 
        \wRegInA23[16] , \wRegInA23[15] , \wRegInA23[14] , \wRegInA23[13] , 
        \wRegInA23[12] , \wRegInA23[11] , \wRegInA23[10] , \wRegInA23[9] , 
        \wRegInA23[8] , \wRegInA23[7] , \wRegInA23[6] , \wRegInA23[5] , 
        \wRegInA23[4] , \wRegInA23[3] , \wRegInA23[2] , \wRegInA23[1] , 
        \wRegInA23[0] }), .Out({\wAIn23[31] , \wAIn23[30] , \wAIn23[29] , 
        \wAIn23[28] , \wAIn23[27] , \wAIn23[26] , \wAIn23[25] , \wAIn23[24] , 
        \wAIn23[23] , \wAIn23[22] , \wAIn23[21] , \wAIn23[20] , \wAIn23[19] , 
        \wAIn23[18] , \wAIn23[17] , \wAIn23[16] , \wAIn23[15] , \wAIn23[14] , 
        \wAIn23[13] , \wAIn23[12] , \wAIn23[11] , \wAIn23[10] , \wAIn23[9] , 
        \wAIn23[8] , \wAIn23[7] , \wAIn23[6] , \wAIn23[5] , \wAIn23[4] , 
        \wAIn23[3] , \wAIn23[2] , \wAIn23[1] , \wAIn23[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_139 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink140[31] , \ScanLink140[30] , \ScanLink140[29] , 
        \ScanLink140[28] , \ScanLink140[27] , \ScanLink140[26] , 
        \ScanLink140[25] , \ScanLink140[24] , \ScanLink140[23] , 
        \ScanLink140[22] , \ScanLink140[21] , \ScanLink140[20] , 
        \ScanLink140[19] , \ScanLink140[18] , \ScanLink140[17] , 
        \ScanLink140[16] , \ScanLink140[15] , \ScanLink140[14] , 
        \ScanLink140[13] , \ScanLink140[12] , \ScanLink140[11] , 
        \ScanLink140[10] , \ScanLink140[9] , \ScanLink140[8] , 
        \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , \ScanLink140[4] , 
        \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , \ScanLink140[0] 
        }), .ScanOut({\ScanLink139[31] , \ScanLink139[30] , \ScanLink139[29] , 
        \ScanLink139[28] , \ScanLink139[27] , \ScanLink139[26] , 
        \ScanLink139[25] , \ScanLink139[24] , \ScanLink139[23] , 
        \ScanLink139[22] , \ScanLink139[21] , \ScanLink139[20] , 
        \ScanLink139[19] , \ScanLink139[18] , \ScanLink139[17] , 
        \ScanLink139[16] , \ScanLink139[15] , \ScanLink139[14] , 
        \ScanLink139[13] , \ScanLink139[12] , \ScanLink139[11] , 
        \ScanLink139[10] , \ScanLink139[9] , \ScanLink139[8] , 
        \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , \ScanLink139[4] , 
        \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , \ScanLink139[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA58[31] , \wRegInA58[30] , \wRegInA58[29] , 
        \wRegInA58[28] , \wRegInA58[27] , \wRegInA58[26] , \wRegInA58[25] , 
        \wRegInA58[24] , \wRegInA58[23] , \wRegInA58[22] , \wRegInA58[21] , 
        \wRegInA58[20] , \wRegInA58[19] , \wRegInA58[18] , \wRegInA58[17] , 
        \wRegInA58[16] , \wRegInA58[15] , \wRegInA58[14] , \wRegInA58[13] , 
        \wRegInA58[12] , \wRegInA58[11] , \wRegInA58[10] , \wRegInA58[9] , 
        \wRegInA58[8] , \wRegInA58[7] , \wRegInA58[6] , \wRegInA58[5] , 
        \wRegInA58[4] , \wRegInA58[3] , \wRegInA58[2] , \wRegInA58[1] , 
        \wRegInA58[0] }), .Out({\wAIn58[31] , \wAIn58[30] , \wAIn58[29] , 
        \wAIn58[28] , \wAIn58[27] , \wAIn58[26] , \wAIn58[25] , \wAIn58[24] , 
        \wAIn58[23] , \wAIn58[22] , \wAIn58[21] , \wAIn58[20] , \wAIn58[19] , 
        \wAIn58[18] , \wAIn58[17] , \wAIn58[16] , \wAIn58[15] , \wAIn58[14] , 
        \wAIn58[13] , \wAIn58[12] , \wAIn58[11] , \wAIn58[10] , \wAIn58[9] , 
        \wAIn58[8] , \wAIn58[7] , \wAIn58[6] , \wAIn58[5] , \wAIn58[4] , 
        \wAIn58[3] , \wAIn58[2] , \wAIn58[1] , \wAIn58[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_69 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink70[31] , \ScanLink70[30] , \ScanLink70[29] , 
        \ScanLink70[28] , \ScanLink70[27] , \ScanLink70[26] , \ScanLink70[25] , 
        \ScanLink70[24] , \ScanLink70[23] , \ScanLink70[22] , \ScanLink70[21] , 
        \ScanLink70[20] , \ScanLink70[19] , \ScanLink70[18] , \ScanLink70[17] , 
        \ScanLink70[16] , \ScanLink70[15] , \ScanLink70[14] , \ScanLink70[13] , 
        \ScanLink70[12] , \ScanLink70[11] , \ScanLink70[10] , \ScanLink70[9] , 
        \ScanLink70[8] , \ScanLink70[7] , \ScanLink70[6] , \ScanLink70[5] , 
        \ScanLink70[4] , \ScanLink70[3] , \ScanLink70[2] , \ScanLink70[1] , 
        \ScanLink70[0] }), .ScanOut({\ScanLink69[31] , \ScanLink69[30] , 
        \ScanLink69[29] , \ScanLink69[28] , \ScanLink69[27] , \ScanLink69[26] , 
        \ScanLink69[25] , \ScanLink69[24] , \ScanLink69[23] , \ScanLink69[22] , 
        \ScanLink69[21] , \ScanLink69[20] , \ScanLink69[19] , \ScanLink69[18] , 
        \ScanLink69[17] , \ScanLink69[16] , \ScanLink69[15] , \ScanLink69[14] , 
        \ScanLink69[13] , \ScanLink69[12] , \ScanLink69[11] , \ScanLink69[10] , 
        \ScanLink69[9] , \ScanLink69[8] , \ScanLink69[7] , \ScanLink69[6] , 
        \ScanLink69[5] , \ScanLink69[4] , \ScanLink69[3] , \ScanLink69[2] , 
        \ScanLink69[1] , \ScanLink69[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA93[31] , \wRegInA93[30] , 
        \wRegInA93[29] , \wRegInA93[28] , \wRegInA93[27] , \wRegInA93[26] , 
        \wRegInA93[25] , \wRegInA93[24] , \wRegInA93[23] , \wRegInA93[22] , 
        \wRegInA93[21] , \wRegInA93[20] , \wRegInA93[19] , \wRegInA93[18] , 
        \wRegInA93[17] , \wRegInA93[16] , \wRegInA93[15] , \wRegInA93[14] , 
        \wRegInA93[13] , \wRegInA93[12] , \wRegInA93[11] , \wRegInA93[10] , 
        \wRegInA93[9] , \wRegInA93[8] , \wRegInA93[7] , \wRegInA93[6] , 
        \wRegInA93[5] , \wRegInA93[4] , \wRegInA93[3] , \wRegInA93[2] , 
        \wRegInA93[1] , \wRegInA93[0] }), .Out({\wAIn93[31] , \wAIn93[30] , 
        \wAIn93[29] , \wAIn93[28] , \wAIn93[27] , \wAIn93[26] , \wAIn93[25] , 
        \wAIn93[24] , \wAIn93[23] , \wAIn93[22] , \wAIn93[21] , \wAIn93[20] , 
        \wAIn93[19] , \wAIn93[18] , \wAIn93[17] , \wAIn93[16] , \wAIn93[15] , 
        \wAIn93[14] , \wAIn93[13] , \wAIn93[12] , \wAIn93[11] , \wAIn93[10] , 
        \wAIn93[9] , \wAIn93[8] , \wAIn93[7] , \wAIn93[6] , \wAIn93[5] , 
        \wAIn93[4] , \wAIn93[3] , \wAIn93[2] , \wAIn93[1] , \wAIn93[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_192 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink193[31] , \ScanLink193[30] , \ScanLink193[29] , 
        \ScanLink193[28] , \ScanLink193[27] , \ScanLink193[26] , 
        \ScanLink193[25] , \ScanLink193[24] , \ScanLink193[23] , 
        \ScanLink193[22] , \ScanLink193[21] , \ScanLink193[20] , 
        \ScanLink193[19] , \ScanLink193[18] , \ScanLink193[17] , 
        \ScanLink193[16] , \ScanLink193[15] , \ScanLink193[14] , 
        \ScanLink193[13] , \ScanLink193[12] , \ScanLink193[11] , 
        \ScanLink193[10] , \ScanLink193[9] , \ScanLink193[8] , 
        \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , \ScanLink193[4] , 
        \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , \ScanLink193[0] 
        }), .ScanOut({\ScanLink192[31] , \ScanLink192[30] , \ScanLink192[29] , 
        \ScanLink192[28] , \ScanLink192[27] , \ScanLink192[26] , 
        \ScanLink192[25] , \ScanLink192[24] , \ScanLink192[23] , 
        \ScanLink192[22] , \ScanLink192[21] , \ScanLink192[20] , 
        \ScanLink192[19] , \ScanLink192[18] , \ScanLink192[17] , 
        \ScanLink192[16] , \ScanLink192[15] , \ScanLink192[14] , 
        \ScanLink192[13] , \ScanLink192[12] , \ScanLink192[11] , 
        \ScanLink192[10] , \ScanLink192[9] , \ScanLink192[8] , 
        \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , \ScanLink192[4] , 
        \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , \ScanLink192[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB31[31] , \wRegInB31[30] , \wRegInB31[29] , 
        \wRegInB31[28] , \wRegInB31[27] , \wRegInB31[26] , \wRegInB31[25] , 
        \wRegInB31[24] , \wRegInB31[23] , \wRegInB31[22] , \wRegInB31[21] , 
        \wRegInB31[20] , \wRegInB31[19] , \wRegInB31[18] , \wRegInB31[17] , 
        \wRegInB31[16] , \wRegInB31[15] , \wRegInB31[14] , \wRegInB31[13] , 
        \wRegInB31[12] , \wRegInB31[11] , \wRegInB31[10] , \wRegInB31[9] , 
        \wRegInB31[8] , \wRegInB31[7] , \wRegInB31[6] , \wRegInB31[5] , 
        \wRegInB31[4] , \wRegInB31[3] , \wRegInB31[2] , \wRegInB31[1] , 
        \wRegInB31[0] }), .Out({\wBIn31[31] , \wBIn31[30] , \wBIn31[29] , 
        \wBIn31[28] , \wBIn31[27] , \wBIn31[26] , \wBIn31[25] , \wBIn31[24] , 
        \wBIn31[23] , \wBIn31[22] , \wBIn31[21] , \wBIn31[20] , \wBIn31[19] , 
        \wBIn31[18] , \wBIn31[17] , \wBIn31[16] , \wBIn31[15] , \wBIn31[14] , 
        \wBIn31[13] , \wBIn31[12] , \wBIn31[11] , \wBIn31[10] , \wBIn31[9] , 
        \wBIn31[8] , \wBIn31[7] , \wBIn31[6] , \wBIn31[5] , \wBIn31[4] , 
        \wBIn31[3] , \wBIn31[2] , \wBIn31[1] , \wBIn31[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid6[31] , 
        \wAMid6[30] , \wAMid6[29] , \wAMid6[28] , \wAMid6[27] , \wAMid6[26] , 
        \wAMid6[25] , \wAMid6[24] , \wAMid6[23] , \wAMid6[22] , \wAMid6[21] , 
        \wAMid6[20] , \wAMid6[19] , \wAMid6[18] , \wAMid6[17] , \wAMid6[16] , 
        \wAMid6[15] , \wAMid6[14] , \wAMid6[13] , \wAMid6[12] , \wAMid6[11] , 
        \wAMid6[10] , \wAMid6[9] , \wAMid6[8] , \wAMid6[7] , \wAMid6[6] , 
        \wAMid6[5] , \wAMid6[4] , \wAMid6[3] , \wAMid6[2] , \wAMid6[1] , 
        \wAMid6[0] }), .BIn({\wBMid6[31] , \wBMid6[30] , \wBMid6[29] , 
        \wBMid6[28] , \wBMid6[27] , \wBMid6[26] , \wBMid6[25] , \wBMid6[24] , 
        \wBMid6[23] , \wBMid6[22] , \wBMid6[21] , \wBMid6[20] , \wBMid6[19] , 
        \wBMid6[18] , \wBMid6[17] , \wBMid6[16] , \wBMid6[15] , \wBMid6[14] , 
        \wBMid6[13] , \wBMid6[12] , \wBMid6[11] , \wBMid6[10] , \wBMid6[9] , 
        \wBMid6[8] , \wBMid6[7] , \wBMid6[6] , \wBMid6[5] , \wBMid6[4] , 
        \wBMid6[3] , \wBMid6[2] , \wBMid6[1] , \wBMid6[0] }), .HiOut({
        \wRegInB6[31] , \wRegInB6[30] , \wRegInB6[29] , \wRegInB6[28] , 
        \wRegInB6[27] , \wRegInB6[26] , \wRegInB6[25] , \wRegInB6[24] , 
        \wRegInB6[23] , \wRegInB6[22] , \wRegInB6[21] , \wRegInB6[20] , 
        \wRegInB6[19] , \wRegInB6[18] , \wRegInB6[17] , \wRegInB6[16] , 
        \wRegInB6[15] , \wRegInB6[14] , \wRegInB6[13] , \wRegInB6[12] , 
        \wRegInB6[11] , \wRegInB6[10] , \wRegInB6[9] , \wRegInB6[8] , 
        \wRegInB6[7] , \wRegInB6[6] , \wRegInB6[5] , \wRegInB6[4] , 
        \wRegInB6[3] , \wRegInB6[2] , \wRegInB6[1] , \wRegInB6[0] }), .LoOut({
        \wRegInA7[31] , \wRegInA7[30] , \wRegInA7[29] , \wRegInA7[28] , 
        \wRegInA7[27] , \wRegInA7[26] , \wRegInA7[25] , \wRegInA7[24] , 
        \wRegInA7[23] , \wRegInA7[22] , \wRegInA7[21] , \wRegInA7[20] , 
        \wRegInA7[19] , \wRegInA7[18] , \wRegInA7[17] , \wRegInA7[16] , 
        \wRegInA7[15] , \wRegInA7[14] , \wRegInA7[13] , \wRegInA7[12] , 
        \wRegInA7[11] , \wRegInA7[10] , \wRegInA7[9] , \wRegInA7[8] , 
        \wRegInA7[7] , \wRegInA7[6] , \wRegInA7[5] , \wRegInA7[4] , 
        \wRegInA7[3] , \wRegInA7[2] , \wRegInA7[1] , \wRegInA7[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_229 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink230[31] , \ScanLink230[30] , \ScanLink230[29] , 
        \ScanLink230[28] , \ScanLink230[27] , \ScanLink230[26] , 
        \ScanLink230[25] , \ScanLink230[24] , \ScanLink230[23] , 
        \ScanLink230[22] , \ScanLink230[21] , \ScanLink230[20] , 
        \ScanLink230[19] , \ScanLink230[18] , \ScanLink230[17] , 
        \ScanLink230[16] , \ScanLink230[15] , \ScanLink230[14] , 
        \ScanLink230[13] , \ScanLink230[12] , \ScanLink230[11] , 
        \ScanLink230[10] , \ScanLink230[9] , \ScanLink230[8] , 
        \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , \ScanLink230[4] , 
        \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , \ScanLink230[0] 
        }), .ScanOut({\ScanLink229[31] , \ScanLink229[30] , \ScanLink229[29] , 
        \ScanLink229[28] , \ScanLink229[27] , \ScanLink229[26] , 
        \ScanLink229[25] , \ScanLink229[24] , \ScanLink229[23] , 
        \ScanLink229[22] , \ScanLink229[21] , \ScanLink229[20] , 
        \ScanLink229[19] , \ScanLink229[18] , \ScanLink229[17] , 
        \ScanLink229[16] , \ScanLink229[15] , \ScanLink229[14] , 
        \ScanLink229[13] , \ScanLink229[12] , \ScanLink229[11] , 
        \ScanLink229[10] , \ScanLink229[9] , \ScanLink229[8] , 
        \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , \ScanLink229[4] , 
        \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , \ScanLink229[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA13[31] , \wRegInA13[30] , \wRegInA13[29] , 
        \wRegInA13[28] , \wRegInA13[27] , \wRegInA13[26] , \wRegInA13[25] , 
        \wRegInA13[24] , \wRegInA13[23] , \wRegInA13[22] , \wRegInA13[21] , 
        \wRegInA13[20] , \wRegInA13[19] , \wRegInA13[18] , \wRegInA13[17] , 
        \wRegInA13[16] , \wRegInA13[15] , \wRegInA13[14] , \wRegInA13[13] , 
        \wRegInA13[12] , \wRegInA13[11] , \wRegInA13[10] , \wRegInA13[9] , 
        \wRegInA13[8] , \wRegInA13[7] , \wRegInA13[6] , \wRegInA13[5] , 
        \wRegInA13[4] , \wRegInA13[3] , \wRegInA13[2] , \wRegInA13[1] , 
        \wRegInA13[0] }), .Out({\wAIn13[31] , \wAIn13[30] , \wAIn13[29] , 
        \wAIn13[28] , \wAIn13[27] , \wAIn13[26] , \wAIn13[25] , \wAIn13[24] , 
        \wAIn13[23] , \wAIn13[22] , \wAIn13[21] , \wAIn13[20] , \wAIn13[19] , 
        \wAIn13[18] , \wAIn13[17] , \wAIn13[16] , \wAIn13[15] , \wAIn13[14] , 
        \wAIn13[13] , \wAIn13[12] , \wAIn13[11] , \wAIn13[10] , \wAIn13[9] , 
        \wAIn13[8] , \wAIn13[7] , \wAIn13[6] , \wAIn13[5] , \wAIn13[4] , 
        \wAIn13[3] , \wAIn13[2] , \wAIn13[1] , \wAIn13[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_119 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink120[31] , \ScanLink120[30] , \ScanLink120[29] , 
        \ScanLink120[28] , \ScanLink120[27] , \ScanLink120[26] , 
        \ScanLink120[25] , \ScanLink120[24] , \ScanLink120[23] , 
        \ScanLink120[22] , \ScanLink120[21] , \ScanLink120[20] , 
        \ScanLink120[19] , \ScanLink120[18] , \ScanLink120[17] , 
        \ScanLink120[16] , \ScanLink120[15] , \ScanLink120[14] , 
        \ScanLink120[13] , \ScanLink120[12] , \ScanLink120[11] , 
        \ScanLink120[10] , \ScanLink120[9] , \ScanLink120[8] , 
        \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , \ScanLink120[4] , 
        \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , \ScanLink120[0] 
        }), .ScanOut({\ScanLink119[31] , \ScanLink119[30] , \ScanLink119[29] , 
        \ScanLink119[28] , \ScanLink119[27] , \ScanLink119[26] , 
        \ScanLink119[25] , \ScanLink119[24] , \ScanLink119[23] , 
        \ScanLink119[22] , \ScanLink119[21] , \ScanLink119[20] , 
        \ScanLink119[19] , \ScanLink119[18] , \ScanLink119[17] , 
        \ScanLink119[16] , \ScanLink119[15] , \ScanLink119[14] , 
        \ScanLink119[13] , \ScanLink119[12] , \ScanLink119[11] , 
        \ScanLink119[10] , \ScanLink119[9] , \ScanLink119[8] , 
        \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , \ScanLink119[4] , 
        \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , \ScanLink119[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA68[31] , \wRegInA68[30] , \wRegInA68[29] , 
        \wRegInA68[28] , \wRegInA68[27] , \wRegInA68[26] , \wRegInA68[25] , 
        \wRegInA68[24] , \wRegInA68[23] , \wRegInA68[22] , \wRegInA68[21] , 
        \wRegInA68[20] , \wRegInA68[19] , \wRegInA68[18] , \wRegInA68[17] , 
        \wRegInA68[16] , \wRegInA68[15] , \wRegInA68[14] , \wRegInA68[13] , 
        \wRegInA68[12] , \wRegInA68[11] , \wRegInA68[10] , \wRegInA68[9] , 
        \wRegInA68[8] , \wRegInA68[7] , \wRegInA68[6] , \wRegInA68[5] , 
        \wRegInA68[4] , \wRegInA68[3] , \wRegInA68[2] , \wRegInA68[1] , 
        \wRegInA68[0] }), .Out({\wAIn68[31] , \wAIn68[30] , \wAIn68[29] , 
        \wAIn68[28] , \wAIn68[27] , \wAIn68[26] , \wAIn68[25] , \wAIn68[24] , 
        \wAIn68[23] , \wAIn68[22] , \wAIn68[21] , \wAIn68[20] , \wAIn68[19] , 
        \wAIn68[18] , \wAIn68[17] , \wAIn68[16] , \wAIn68[15] , \wAIn68[14] , 
        \wAIn68[13] , \wAIn68[12] , \wAIn68[11] , \wAIn68[10] , \wAIn68[9] , 
        \wAIn68[8] , \wAIn68[7] , \wAIn68[6] , \wAIn68[5] , \wAIn68[4] , 
        \wAIn68[3] , \wAIn68[2] , \wAIn68[1] , \wAIn68[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_49 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink50[31] , \ScanLink50[30] , \ScanLink50[29] , 
        \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , \ScanLink50[25] , 
        \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , \ScanLink50[21] , 
        \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , \ScanLink50[17] , 
        \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , \ScanLink50[13] , 
        \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , \ScanLink50[9] , 
        \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , \ScanLink50[5] , 
        \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , \ScanLink50[1] , 
        \ScanLink50[0] }), .ScanOut({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA103[31] , \wRegInA103[30] , 
        \wRegInA103[29] , \wRegInA103[28] , \wRegInA103[27] , \wRegInA103[26] , 
        \wRegInA103[25] , \wRegInA103[24] , \wRegInA103[23] , \wRegInA103[22] , 
        \wRegInA103[21] , \wRegInA103[20] , \wRegInA103[19] , \wRegInA103[18] , 
        \wRegInA103[17] , \wRegInA103[16] , \wRegInA103[15] , \wRegInA103[14] , 
        \wRegInA103[13] , \wRegInA103[12] , \wRegInA103[11] , \wRegInA103[10] , 
        \wRegInA103[9] , \wRegInA103[8] , \wRegInA103[7] , \wRegInA103[6] , 
        \wRegInA103[5] , \wRegInA103[4] , \wRegInA103[3] , \wRegInA103[2] , 
        \wRegInA103[1] , \wRegInA103[0] }), .Out({\wAIn103[31] , \wAIn103[30] , 
        \wAIn103[29] , \wAIn103[28] , \wAIn103[27] , \wAIn103[26] , 
        \wAIn103[25] , \wAIn103[24] , \wAIn103[23] , \wAIn103[22] , 
        \wAIn103[21] , \wAIn103[20] , \wAIn103[19] , \wAIn103[18] , 
        \wAIn103[17] , \wAIn103[16] , \wAIn103[15] , \wAIn103[14] , 
        \wAIn103[13] , \wAIn103[12] , \wAIn103[11] , \wAIn103[10] , 
        \wAIn103[9] , \wAIn103[8] , \wAIn103[7] , \wAIn103[6] , \wAIn103[5] , 
        \wAIn103[4] , \wAIn103[3] , \wAIn103[2] , \wAIn103[1] , \wAIn103[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn102[31] , \wAIn102[30] , \wAIn102[29] , \wAIn102[28] , 
        \wAIn102[27] , \wAIn102[26] , \wAIn102[25] , \wAIn102[24] , 
        \wAIn102[23] , \wAIn102[22] , \wAIn102[21] , \wAIn102[20] , 
        \wAIn102[19] , \wAIn102[18] , \wAIn102[17] , \wAIn102[16] , 
        \wAIn102[15] , \wAIn102[14] , \wAIn102[13] , \wAIn102[12] , 
        \wAIn102[11] , \wAIn102[10] , \wAIn102[9] , \wAIn102[8] , \wAIn102[7] , 
        \wAIn102[6] , \wAIn102[5] , \wAIn102[4] , \wAIn102[3] , \wAIn102[2] , 
        \wAIn102[1] , \wAIn102[0] }), .BIn({\wBIn102[31] , \wBIn102[30] , 
        \wBIn102[29] , \wBIn102[28] , \wBIn102[27] , \wBIn102[26] , 
        \wBIn102[25] , \wBIn102[24] , \wBIn102[23] , \wBIn102[22] , 
        \wBIn102[21] , \wBIn102[20] , \wBIn102[19] , \wBIn102[18] , 
        \wBIn102[17] , \wBIn102[16] , \wBIn102[15] , \wBIn102[14] , 
        \wBIn102[13] , \wBIn102[12] , \wBIn102[11] , \wBIn102[10] , 
        \wBIn102[9] , \wBIn102[8] , \wBIn102[7] , \wBIn102[6] , \wBIn102[5] , 
        \wBIn102[4] , \wBIn102[3] , \wBIn102[2] , \wBIn102[1] , \wBIn102[0] }), 
        .HiOut({\wBMid101[31] , \wBMid101[30] , \wBMid101[29] , \wBMid101[28] , 
        \wBMid101[27] , \wBMid101[26] , \wBMid101[25] , \wBMid101[24] , 
        \wBMid101[23] , \wBMid101[22] , \wBMid101[21] , \wBMid101[20] , 
        \wBMid101[19] , \wBMid101[18] , \wBMid101[17] , \wBMid101[16] , 
        \wBMid101[15] , \wBMid101[14] , \wBMid101[13] , \wBMid101[12] , 
        \wBMid101[11] , \wBMid101[10] , \wBMid101[9] , \wBMid101[8] , 
        \wBMid101[7] , \wBMid101[6] , \wBMid101[5] , \wBMid101[4] , 
        \wBMid101[3] , \wBMid101[2] , \wBMid101[1] , \wBMid101[0] }), .LoOut({
        \wAMid102[31] , \wAMid102[30] , \wAMid102[29] , \wAMid102[28] , 
        \wAMid102[27] , \wAMid102[26] , \wAMid102[25] , \wAMid102[24] , 
        \wAMid102[23] , \wAMid102[22] , \wAMid102[21] , \wAMid102[20] , 
        \wAMid102[19] , \wAMid102[18] , \wAMid102[17] , \wAMid102[16] , 
        \wAMid102[15] , \wAMid102[14] , \wAMid102[13] , \wAMid102[12] , 
        \wAMid102[11] , \wAMid102[10] , \wAMid102[9] , \wAMid102[8] , 
        \wAMid102[7] , \wAMid102[6] , \wAMid102[5] , \wAMid102[4] , 
        \wAMid102[3] , \wAMid102[2] , \wAMid102[1] , \wAMid102[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid42[31] , \wAMid42[30] , \wAMid42[29] , \wAMid42[28] , 
        \wAMid42[27] , \wAMid42[26] , \wAMid42[25] , \wAMid42[24] , 
        \wAMid42[23] , \wAMid42[22] , \wAMid42[21] , \wAMid42[20] , 
        \wAMid42[19] , \wAMid42[18] , \wAMid42[17] , \wAMid42[16] , 
        \wAMid42[15] , \wAMid42[14] , \wAMid42[13] , \wAMid42[12] , 
        \wAMid42[11] , \wAMid42[10] , \wAMid42[9] , \wAMid42[8] , \wAMid42[7] , 
        \wAMid42[6] , \wAMid42[5] , \wAMid42[4] , \wAMid42[3] , \wAMid42[2] , 
        \wAMid42[1] , \wAMid42[0] }), .BIn({\wBMid42[31] , \wBMid42[30] , 
        \wBMid42[29] , \wBMid42[28] , \wBMid42[27] , \wBMid42[26] , 
        \wBMid42[25] , \wBMid42[24] , \wBMid42[23] , \wBMid42[22] , 
        \wBMid42[21] , \wBMid42[20] , \wBMid42[19] , \wBMid42[18] , 
        \wBMid42[17] , \wBMid42[16] , \wBMid42[15] , \wBMid42[14] , 
        \wBMid42[13] , \wBMid42[12] , \wBMid42[11] , \wBMid42[10] , 
        \wBMid42[9] , \wBMid42[8] , \wBMid42[7] , \wBMid42[6] , \wBMid42[5] , 
        \wBMid42[4] , \wBMid42[3] , \wBMid42[2] , \wBMid42[1] , \wBMid42[0] }), 
        .HiOut({\wRegInB42[31] , \wRegInB42[30] , \wRegInB42[29] , 
        \wRegInB42[28] , \wRegInB42[27] , \wRegInB42[26] , \wRegInB42[25] , 
        \wRegInB42[24] , \wRegInB42[23] , \wRegInB42[22] , \wRegInB42[21] , 
        \wRegInB42[20] , \wRegInB42[19] , \wRegInB42[18] , \wRegInB42[17] , 
        \wRegInB42[16] , \wRegInB42[15] , \wRegInB42[14] , \wRegInB42[13] , 
        \wRegInB42[12] , \wRegInB42[11] , \wRegInB42[10] , \wRegInB42[9] , 
        \wRegInB42[8] , \wRegInB42[7] , \wRegInB42[6] , \wRegInB42[5] , 
        \wRegInB42[4] , \wRegInB42[3] , \wRegInB42[2] , \wRegInB42[1] , 
        \wRegInB42[0] }), .LoOut({\wRegInA43[31] , \wRegInA43[30] , 
        \wRegInA43[29] , \wRegInA43[28] , \wRegInA43[27] , \wRegInA43[26] , 
        \wRegInA43[25] , \wRegInA43[24] , \wRegInA43[23] , \wRegInA43[22] , 
        \wRegInA43[21] , \wRegInA43[20] , \wRegInA43[19] , \wRegInA43[18] , 
        \wRegInA43[17] , \wRegInA43[16] , \wRegInA43[15] , \wRegInA43[14] , 
        \wRegInA43[13] , \wRegInA43[12] , \wRegInA43[11] , \wRegInA43[10] , 
        \wRegInA43[9] , \wRegInA43[8] , \wRegInA43[7] , \wRegInA43[6] , 
        \wRegInA43[5] , \wRegInA43[4] , \wRegInA43[3] , \wRegInA43[2] , 
        \wRegInA43[1] , \wRegInA43[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_177 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink178[31] , \ScanLink178[30] , \ScanLink178[29] , 
        \ScanLink178[28] , \ScanLink178[27] , \ScanLink178[26] , 
        \ScanLink178[25] , \ScanLink178[24] , \ScanLink178[23] , 
        \ScanLink178[22] , \ScanLink178[21] , \ScanLink178[20] , 
        \ScanLink178[19] , \ScanLink178[18] , \ScanLink178[17] , 
        \ScanLink178[16] , \ScanLink178[15] , \ScanLink178[14] , 
        \ScanLink178[13] , \ScanLink178[12] , \ScanLink178[11] , 
        \ScanLink178[10] , \ScanLink178[9] , \ScanLink178[8] , 
        \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , \ScanLink178[4] , 
        \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , \ScanLink178[0] 
        }), .ScanOut({\ScanLink177[31] , \ScanLink177[30] , \ScanLink177[29] , 
        \ScanLink177[28] , \ScanLink177[27] , \ScanLink177[26] , 
        \ScanLink177[25] , \ScanLink177[24] , \ScanLink177[23] , 
        \ScanLink177[22] , \ScanLink177[21] , \ScanLink177[20] , 
        \ScanLink177[19] , \ScanLink177[18] , \ScanLink177[17] , 
        \ScanLink177[16] , \ScanLink177[15] , \ScanLink177[14] , 
        \ScanLink177[13] , \ScanLink177[12] , \ScanLink177[11] , 
        \ScanLink177[10] , \ScanLink177[9] , \ScanLink177[8] , 
        \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , \ScanLink177[4] , 
        \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , \ScanLink177[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA39[31] , \wRegInA39[30] , \wRegInA39[29] , 
        \wRegInA39[28] , \wRegInA39[27] , \wRegInA39[26] , \wRegInA39[25] , 
        \wRegInA39[24] , \wRegInA39[23] , \wRegInA39[22] , \wRegInA39[21] , 
        \wRegInA39[20] , \wRegInA39[19] , \wRegInA39[18] , \wRegInA39[17] , 
        \wRegInA39[16] , \wRegInA39[15] , \wRegInA39[14] , \wRegInA39[13] , 
        \wRegInA39[12] , \wRegInA39[11] , \wRegInA39[10] , \wRegInA39[9] , 
        \wRegInA39[8] , \wRegInA39[7] , \wRegInA39[6] , \wRegInA39[5] , 
        \wRegInA39[4] , \wRegInA39[3] , \wRegInA39[2] , \wRegInA39[1] , 
        \wRegInA39[0] }), .Out({\wAIn39[31] , \wAIn39[30] , \wAIn39[29] , 
        \wAIn39[28] , \wAIn39[27] , \wAIn39[26] , \wAIn39[25] , \wAIn39[24] , 
        \wAIn39[23] , \wAIn39[22] , \wAIn39[21] , \wAIn39[20] , \wAIn39[19] , 
        \wAIn39[18] , \wAIn39[17] , \wAIn39[16] , \wAIn39[15] , \wAIn39[14] , 
        \wAIn39[13] , \wAIn39[12] , \wAIn39[11] , \wAIn39[10] , \wAIn39[9] , 
        \wAIn39[8] , \wAIn39[7] , \wAIn39[6] , \wAIn39[5] , \wAIn39[4] , 
        \wAIn39[3] , \wAIn39[2] , \wAIn39[1] , \wAIn39[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_27 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink28[31] , \ScanLink28[30] , \ScanLink28[29] , 
        \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , \ScanLink28[25] , 
        \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , \ScanLink28[21] , 
        \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , \ScanLink28[17] , 
        \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , \ScanLink28[13] , 
        \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , \ScanLink28[9] , 
        \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , \ScanLink28[5] , 
        \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , \ScanLink28[1] , 
        \ScanLink28[0] }), .ScanOut({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA114[31] , \wRegInA114[30] , 
        \wRegInA114[29] , \wRegInA114[28] , \wRegInA114[27] , \wRegInA114[26] , 
        \wRegInA114[25] , \wRegInA114[24] , \wRegInA114[23] , \wRegInA114[22] , 
        \wRegInA114[21] , \wRegInA114[20] , \wRegInA114[19] , \wRegInA114[18] , 
        \wRegInA114[17] , \wRegInA114[16] , \wRegInA114[15] , \wRegInA114[14] , 
        \wRegInA114[13] , \wRegInA114[12] , \wRegInA114[11] , \wRegInA114[10] , 
        \wRegInA114[9] , \wRegInA114[8] , \wRegInA114[7] , \wRegInA114[6] , 
        \wRegInA114[5] , \wRegInA114[4] , \wRegInA114[3] , \wRegInA114[2] , 
        \wRegInA114[1] , \wRegInA114[0] }), .Out({\wAIn114[31] , \wAIn114[30] , 
        \wAIn114[29] , \wAIn114[28] , \wAIn114[27] , \wAIn114[26] , 
        \wAIn114[25] , \wAIn114[24] , \wAIn114[23] , \wAIn114[22] , 
        \wAIn114[21] , \wAIn114[20] , \wAIn114[19] , \wAIn114[18] , 
        \wAIn114[17] , \wAIn114[16] , \wAIn114[15] , \wAIn114[14] , 
        \wAIn114[13] , \wAIn114[12] , \wAIn114[11] , \wAIn114[10] , 
        \wAIn114[9] , \wAIn114[8] , \wAIn114[7] , \wAIn114[6] , \wAIn114[5] , 
        \wAIn114[4] , \wAIn114[3] , \wAIn114[2] , \wAIn114[1] , \wAIn114[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn125[31] , \wAIn125[30] , \wAIn125[29] , \wAIn125[28] , 
        \wAIn125[27] , \wAIn125[26] , \wAIn125[25] , \wAIn125[24] , 
        \wAIn125[23] , \wAIn125[22] , \wAIn125[21] , \wAIn125[20] , 
        \wAIn125[19] , \wAIn125[18] , \wAIn125[17] , \wAIn125[16] , 
        \wAIn125[15] , \wAIn125[14] , \wAIn125[13] , \wAIn125[12] , 
        \wAIn125[11] , \wAIn125[10] , \wAIn125[9] , \wAIn125[8] , \wAIn125[7] , 
        \wAIn125[6] , \wAIn125[5] , \wAIn125[4] , \wAIn125[3] , \wAIn125[2] , 
        \wAIn125[1] , \wAIn125[0] }), .BIn({\wBIn125[31] , \wBIn125[30] , 
        \wBIn125[29] , \wBIn125[28] , \wBIn125[27] , \wBIn125[26] , 
        \wBIn125[25] , \wBIn125[24] , \wBIn125[23] , \wBIn125[22] , 
        \wBIn125[21] , \wBIn125[20] , \wBIn125[19] , \wBIn125[18] , 
        \wBIn125[17] , \wBIn125[16] , \wBIn125[15] , \wBIn125[14] , 
        \wBIn125[13] , \wBIn125[12] , \wBIn125[11] , \wBIn125[10] , 
        \wBIn125[9] , \wBIn125[8] , \wBIn125[7] , \wBIn125[6] , \wBIn125[5] , 
        \wBIn125[4] , \wBIn125[3] , \wBIn125[2] , \wBIn125[1] , \wBIn125[0] }), 
        .HiOut({\wBMid124[31] , \wBMid124[30] , \wBMid124[29] , \wBMid124[28] , 
        \wBMid124[27] , \wBMid124[26] , \wBMid124[25] , \wBMid124[24] , 
        \wBMid124[23] , \wBMid124[22] , \wBMid124[21] , \wBMid124[20] , 
        \wBMid124[19] , \wBMid124[18] , \wBMid124[17] , \wBMid124[16] , 
        \wBMid124[15] , \wBMid124[14] , \wBMid124[13] , \wBMid124[12] , 
        \wBMid124[11] , \wBMid124[10] , \wBMid124[9] , \wBMid124[8] , 
        \wBMid124[7] , \wBMid124[6] , \wBMid124[5] , \wBMid124[4] , 
        \wBMid124[3] , \wBMid124[2] , \wBMid124[1] , \wBMid124[0] }), .LoOut({
        \wAMid125[31] , \wAMid125[30] , \wAMid125[29] , \wAMid125[28] , 
        \wAMid125[27] , \wAMid125[26] , \wAMid125[25] , \wAMid125[24] , 
        \wAMid125[23] , \wAMid125[22] , \wAMid125[21] , \wAMid125[20] , 
        \wAMid125[19] , \wAMid125[18] , \wAMid125[17] , \wAMid125[16] , 
        \wAMid125[15] , \wAMid125[14] , \wAMid125[13] , \wAMid125[12] , 
        \wAMid125[11] , \wAMid125[10] , \wAMid125[9] , \wAMid125[8] , 
        \wAMid125[7] , \wAMid125[6] , \wAMid125[5] , \wAMid125[4] , 
        \wAMid125[3] , \wAMid125[2] , \wAMid125[1] , \wAMid125[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_247 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink248[31] , \ScanLink248[30] , \ScanLink248[29] , 
        \ScanLink248[28] , \ScanLink248[27] , \ScanLink248[26] , 
        \ScanLink248[25] , \ScanLink248[24] , \ScanLink248[23] , 
        \ScanLink248[22] , \ScanLink248[21] , \ScanLink248[20] , 
        \ScanLink248[19] , \ScanLink248[18] , \ScanLink248[17] , 
        \ScanLink248[16] , \ScanLink248[15] , \ScanLink248[14] , 
        \ScanLink248[13] , \ScanLink248[12] , \ScanLink248[11] , 
        \ScanLink248[10] , \ScanLink248[9] , \ScanLink248[8] , 
        \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , \ScanLink248[4] , 
        \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , \ScanLink248[0] 
        }), .ScanOut({\ScanLink247[31] , \ScanLink247[30] , \ScanLink247[29] , 
        \ScanLink247[28] , \ScanLink247[27] , \ScanLink247[26] , 
        \ScanLink247[25] , \ScanLink247[24] , \ScanLink247[23] , 
        \ScanLink247[22] , \ScanLink247[21] , \ScanLink247[20] , 
        \ScanLink247[19] , \ScanLink247[18] , \ScanLink247[17] , 
        \ScanLink247[16] , \ScanLink247[15] , \ScanLink247[14] , 
        \ScanLink247[13] , \ScanLink247[12] , \ScanLink247[11] , 
        \ScanLink247[10] , \ScanLink247[9] , \ScanLink247[8] , 
        \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , \ScanLink247[4] , 
        \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , \ScanLink247[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA4[31] , \wRegInA4[30] , \wRegInA4[29] , \wRegInA4[28] , 
        \wRegInA4[27] , \wRegInA4[26] , \wRegInA4[25] , \wRegInA4[24] , 
        \wRegInA4[23] , \wRegInA4[22] , \wRegInA4[21] , \wRegInA4[20] , 
        \wRegInA4[19] , \wRegInA4[18] , \wRegInA4[17] , \wRegInA4[16] , 
        \wRegInA4[15] , \wRegInA4[14] , \wRegInA4[13] , \wRegInA4[12] , 
        \wRegInA4[11] , \wRegInA4[10] , \wRegInA4[9] , \wRegInA4[8] , 
        \wRegInA4[7] , \wRegInA4[6] , \wRegInA4[5] , \wRegInA4[4] , 
        \wRegInA4[3] , \wRegInA4[2] , \wRegInA4[1] , \wRegInA4[0] }), .Out({
        \wAIn4[31] , \wAIn4[30] , \wAIn4[29] , \wAIn4[28] , \wAIn4[27] , 
        \wAIn4[26] , \wAIn4[25] , \wAIn4[24] , \wAIn4[23] , \wAIn4[22] , 
        \wAIn4[21] , \wAIn4[20] , \wAIn4[19] , \wAIn4[18] , \wAIn4[17] , 
        \wAIn4[16] , \wAIn4[15] , \wAIn4[14] , \wAIn4[13] , \wAIn4[12] , 
        \wAIn4[11] , \wAIn4[10] , \wAIn4[9] , \wAIn4[8] , \wAIn4[7] , 
        \wAIn4[6] , \wAIn4[5] , \wAIn4[4] , \wAIn4[3] , \wAIn4[2] , \wAIn4[1] , 
        \wAIn4[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn69[31] , \wAIn69[30] , \wAIn69[29] , \wAIn69[28] , \wAIn69[27] , 
        \wAIn69[26] , \wAIn69[25] , \wAIn69[24] , \wAIn69[23] , \wAIn69[22] , 
        \wAIn69[21] , \wAIn69[20] , \wAIn69[19] , \wAIn69[18] , \wAIn69[17] , 
        \wAIn69[16] , \wAIn69[15] , \wAIn69[14] , \wAIn69[13] , \wAIn69[12] , 
        \wAIn69[11] , \wAIn69[10] , \wAIn69[9] , \wAIn69[8] , \wAIn69[7] , 
        \wAIn69[6] , \wAIn69[5] , \wAIn69[4] , \wAIn69[3] , \wAIn69[2] , 
        \wAIn69[1] , \wAIn69[0] }), .BIn({\wBIn69[31] , \wBIn69[30] , 
        \wBIn69[29] , \wBIn69[28] , \wBIn69[27] , \wBIn69[26] , \wBIn69[25] , 
        \wBIn69[24] , \wBIn69[23] , \wBIn69[22] , \wBIn69[21] , \wBIn69[20] , 
        \wBIn69[19] , \wBIn69[18] , \wBIn69[17] , \wBIn69[16] , \wBIn69[15] , 
        \wBIn69[14] , \wBIn69[13] , \wBIn69[12] , \wBIn69[11] , \wBIn69[10] , 
        \wBIn69[9] , \wBIn69[8] , \wBIn69[7] , \wBIn69[6] , \wBIn69[5] , 
        \wBIn69[4] , \wBIn69[3] , \wBIn69[2] , \wBIn69[1] , \wBIn69[0] }), 
        .HiOut({\wBMid68[31] , \wBMid68[30] , \wBMid68[29] , \wBMid68[28] , 
        \wBMid68[27] , \wBMid68[26] , \wBMid68[25] , \wBMid68[24] , 
        \wBMid68[23] , \wBMid68[22] , \wBMid68[21] , \wBMid68[20] , 
        \wBMid68[19] , \wBMid68[18] , \wBMid68[17] , \wBMid68[16] , 
        \wBMid68[15] , \wBMid68[14] , \wBMid68[13] , \wBMid68[12] , 
        \wBMid68[11] , \wBMid68[10] , \wBMid68[9] , \wBMid68[8] , \wBMid68[7] , 
        \wBMid68[6] , \wBMid68[5] , \wBMid68[4] , \wBMid68[3] , \wBMid68[2] , 
        \wBMid68[1] , \wBMid68[0] }), .LoOut({\wAMid69[31] , \wAMid69[30] , 
        \wAMid69[29] , \wAMid69[28] , \wAMid69[27] , \wAMid69[26] , 
        \wAMid69[25] , \wAMid69[24] , \wAMid69[23] , \wAMid69[22] , 
        \wAMid69[21] , \wAMid69[20] , \wAMid69[19] , \wAMid69[18] , 
        \wAMid69[17] , \wAMid69[16] , \wAMid69[15] , \wAMid69[14] , 
        \wAMid69[13] , \wAMid69[12] , \wAMid69[11] , \wAMid69[10] , 
        \wAMid69[9] , \wAMid69[8] , \wAMid69[7] , \wAMid69[6] , \wAMid69[5] , 
        \wAMid69[4] , \wAMid69[3] , \wAMid69[2] , \wAMid69[1] , \wAMid69[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn119[31] , \wAIn119[30] , \wAIn119[29] , \wAIn119[28] , 
        \wAIn119[27] , \wAIn119[26] , \wAIn119[25] , \wAIn119[24] , 
        \wAIn119[23] , \wAIn119[22] , \wAIn119[21] , \wAIn119[20] , 
        \wAIn119[19] , \wAIn119[18] , \wAIn119[17] , \wAIn119[16] , 
        \wAIn119[15] , \wAIn119[14] , \wAIn119[13] , \wAIn119[12] , 
        \wAIn119[11] , \wAIn119[10] , \wAIn119[9] , \wAIn119[8] , \wAIn119[7] , 
        \wAIn119[6] , \wAIn119[5] , \wAIn119[4] , \wAIn119[3] , \wAIn119[2] , 
        \wAIn119[1] , \wAIn119[0] }), .BIn({\wBIn119[31] , \wBIn119[30] , 
        \wBIn119[29] , \wBIn119[28] , \wBIn119[27] , \wBIn119[26] , 
        \wBIn119[25] , \wBIn119[24] , \wBIn119[23] , \wBIn119[22] , 
        \wBIn119[21] , \wBIn119[20] , \wBIn119[19] , \wBIn119[18] , 
        \wBIn119[17] , \wBIn119[16] , \wBIn119[15] , \wBIn119[14] , 
        \wBIn119[13] , \wBIn119[12] , \wBIn119[11] , \wBIn119[10] , 
        \wBIn119[9] , \wBIn119[8] , \wBIn119[7] , \wBIn119[6] , \wBIn119[5] , 
        \wBIn119[4] , \wBIn119[3] , \wBIn119[2] , \wBIn119[1] , \wBIn119[0] }), 
        .HiOut({\wBMid118[31] , \wBMid118[30] , \wBMid118[29] , \wBMid118[28] , 
        \wBMid118[27] , \wBMid118[26] , \wBMid118[25] , \wBMid118[24] , 
        \wBMid118[23] , \wBMid118[22] , \wBMid118[21] , \wBMid118[20] , 
        \wBMid118[19] , \wBMid118[18] , \wBMid118[17] , \wBMid118[16] , 
        \wBMid118[15] , \wBMid118[14] , \wBMid118[13] , \wBMid118[12] , 
        \wBMid118[11] , \wBMid118[10] , \wBMid118[9] , \wBMid118[8] , 
        \wBMid118[7] , \wBMid118[6] , \wBMid118[5] , \wBMid118[4] , 
        \wBMid118[3] , \wBMid118[2] , \wBMid118[1] , \wBMid118[0] }), .LoOut({
        \wAMid119[31] , \wAMid119[30] , \wAMid119[29] , \wAMid119[28] , 
        \wAMid119[27] , \wAMid119[26] , \wAMid119[25] , \wAMid119[24] , 
        \wAMid119[23] , \wAMid119[22] , \wAMid119[21] , \wAMid119[20] , 
        \wAMid119[19] , \wAMid119[18] , \wAMid119[17] , \wAMid119[16] , 
        \wAMid119[15] , \wAMid119[14] , \wAMid119[13] , \wAMid119[12] , 
        \wAMid119[11] , \wAMid119[10] , \wAMid119[9] , \wAMid119[8] , 
        \wAMid119[7] , \wAMid119[6] , \wAMid119[5] , \wAMid119[4] , 
        \wAMid119[3] , \wAMid119[2] , \wAMid119[1] , \wAMid119[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid65[31] , \wAMid65[30] , \wAMid65[29] , \wAMid65[28] , 
        \wAMid65[27] , \wAMid65[26] , \wAMid65[25] , \wAMid65[24] , 
        \wAMid65[23] , \wAMid65[22] , \wAMid65[21] , \wAMid65[20] , 
        \wAMid65[19] , \wAMid65[18] , \wAMid65[17] , \wAMid65[16] , 
        \wAMid65[15] , \wAMid65[14] , \wAMid65[13] , \wAMid65[12] , 
        \wAMid65[11] , \wAMid65[10] , \wAMid65[9] , \wAMid65[8] , \wAMid65[7] , 
        \wAMid65[6] , \wAMid65[5] , \wAMid65[4] , \wAMid65[3] , \wAMid65[2] , 
        \wAMid65[1] , \wAMid65[0] }), .BIn({\wBMid65[31] , \wBMid65[30] , 
        \wBMid65[29] , \wBMid65[28] , \wBMid65[27] , \wBMid65[26] , 
        \wBMid65[25] , \wBMid65[24] , \wBMid65[23] , \wBMid65[22] , 
        \wBMid65[21] , \wBMid65[20] , \wBMid65[19] , \wBMid65[18] , 
        \wBMid65[17] , \wBMid65[16] , \wBMid65[15] , \wBMid65[14] , 
        \wBMid65[13] , \wBMid65[12] , \wBMid65[11] , \wBMid65[10] , 
        \wBMid65[9] , \wBMid65[8] , \wBMid65[7] , \wBMid65[6] , \wBMid65[5] , 
        \wBMid65[4] , \wBMid65[3] , \wBMid65[2] , \wBMid65[1] , \wBMid65[0] }), 
        .HiOut({\wRegInB65[31] , \wRegInB65[30] , \wRegInB65[29] , 
        \wRegInB65[28] , \wRegInB65[27] , \wRegInB65[26] , \wRegInB65[25] , 
        \wRegInB65[24] , \wRegInB65[23] , \wRegInB65[22] , \wRegInB65[21] , 
        \wRegInB65[20] , \wRegInB65[19] , \wRegInB65[18] , \wRegInB65[17] , 
        \wRegInB65[16] , \wRegInB65[15] , \wRegInB65[14] , \wRegInB65[13] , 
        \wRegInB65[12] , \wRegInB65[11] , \wRegInB65[10] , \wRegInB65[9] , 
        \wRegInB65[8] , \wRegInB65[7] , \wRegInB65[6] , \wRegInB65[5] , 
        \wRegInB65[4] , \wRegInB65[3] , \wRegInB65[2] , \wRegInB65[1] , 
        \wRegInB65[0] }), .LoOut({\wRegInA66[31] , \wRegInA66[30] , 
        \wRegInA66[29] , \wRegInA66[28] , \wRegInA66[27] , \wRegInA66[26] , 
        \wRegInA66[25] , \wRegInA66[24] , \wRegInA66[23] , \wRegInA66[22] , 
        \wRegInA66[21] , \wRegInA66[20] , \wRegInA66[19] , \wRegInA66[18] , 
        \wRegInA66[17] , \wRegInA66[16] , \wRegInA66[15] , \wRegInA66[14] , 
        \wRegInA66[13] , \wRegInA66[12] , \wRegInA66[11] , \wRegInA66[10] , 
        \wRegInA66[9] , \wRegInA66[8] , \wRegInA66[7] , \wRegInA66[6] , 
        \wRegInA66[5] , \wRegInA66[4] , \wRegInA66[3] , \wRegInA66[2] , 
        \wRegInA66[1] , \wRegInA66[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_150 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink151[31] , \ScanLink151[30] , \ScanLink151[29] , 
        \ScanLink151[28] , \ScanLink151[27] , \ScanLink151[26] , 
        \ScanLink151[25] , \ScanLink151[24] , \ScanLink151[23] , 
        \ScanLink151[22] , \ScanLink151[21] , \ScanLink151[20] , 
        \ScanLink151[19] , \ScanLink151[18] , \ScanLink151[17] , 
        \ScanLink151[16] , \ScanLink151[15] , \ScanLink151[14] , 
        \ScanLink151[13] , \ScanLink151[12] , \ScanLink151[11] , 
        \ScanLink151[10] , \ScanLink151[9] , \ScanLink151[8] , 
        \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , \ScanLink151[4] , 
        \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , \ScanLink151[0] 
        }), .ScanOut({\ScanLink150[31] , \ScanLink150[30] , \ScanLink150[29] , 
        \ScanLink150[28] , \ScanLink150[27] , \ScanLink150[26] , 
        \ScanLink150[25] , \ScanLink150[24] , \ScanLink150[23] , 
        \ScanLink150[22] , \ScanLink150[21] , \ScanLink150[20] , 
        \ScanLink150[19] , \ScanLink150[18] , \ScanLink150[17] , 
        \ScanLink150[16] , \ScanLink150[15] , \ScanLink150[14] , 
        \ScanLink150[13] , \ScanLink150[12] , \ScanLink150[11] , 
        \ScanLink150[10] , \ScanLink150[9] , \ScanLink150[8] , 
        \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , \ScanLink150[4] , 
        \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , \ScanLink150[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB52[31] , \wRegInB52[30] , \wRegInB52[29] , 
        \wRegInB52[28] , \wRegInB52[27] , \wRegInB52[26] , \wRegInB52[25] , 
        \wRegInB52[24] , \wRegInB52[23] , \wRegInB52[22] , \wRegInB52[21] , 
        \wRegInB52[20] , \wRegInB52[19] , \wRegInB52[18] , \wRegInB52[17] , 
        \wRegInB52[16] , \wRegInB52[15] , \wRegInB52[14] , \wRegInB52[13] , 
        \wRegInB52[12] , \wRegInB52[11] , \wRegInB52[10] , \wRegInB52[9] , 
        \wRegInB52[8] , \wRegInB52[7] , \wRegInB52[6] , \wRegInB52[5] , 
        \wRegInB52[4] , \wRegInB52[3] , \wRegInB52[2] , \wRegInB52[1] , 
        \wRegInB52[0] }), .Out({\wBIn52[31] , \wBIn52[30] , \wBIn52[29] , 
        \wBIn52[28] , \wBIn52[27] , \wBIn52[26] , \wBIn52[25] , \wBIn52[24] , 
        \wBIn52[23] , \wBIn52[22] , \wBIn52[21] , \wBIn52[20] , \wBIn52[19] , 
        \wBIn52[18] , \wBIn52[17] , \wBIn52[16] , \wBIn52[15] , \wBIn52[14] , 
        \wBIn52[13] , \wBIn52[12] , \wBIn52[11] , \wBIn52[10] , \wBIn52[9] , 
        \wBIn52[8] , \wBIn52[7] , \wBIn52[6] , \wBIn52[5] , \wBIn52[4] , 
        \wBIn52[3] , \wBIn52[2] , \wBIn52[1] , \wBIn52[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid108[31] , \wAMid108[30] , \wAMid108[29] , \wAMid108[28] , 
        \wAMid108[27] , \wAMid108[26] , \wAMid108[25] , \wAMid108[24] , 
        \wAMid108[23] , \wAMid108[22] , \wAMid108[21] , \wAMid108[20] , 
        \wAMid108[19] , \wAMid108[18] , \wAMid108[17] , \wAMid108[16] , 
        \wAMid108[15] , \wAMid108[14] , \wAMid108[13] , \wAMid108[12] , 
        \wAMid108[11] , \wAMid108[10] , \wAMid108[9] , \wAMid108[8] , 
        \wAMid108[7] , \wAMid108[6] , \wAMid108[5] , \wAMid108[4] , 
        \wAMid108[3] , \wAMid108[2] , \wAMid108[1] , \wAMid108[0] }), .BIn({
        \wBMid108[31] , \wBMid108[30] , \wBMid108[29] , \wBMid108[28] , 
        \wBMid108[27] , \wBMid108[26] , \wBMid108[25] , \wBMid108[24] , 
        \wBMid108[23] , \wBMid108[22] , \wBMid108[21] , \wBMid108[20] , 
        \wBMid108[19] , \wBMid108[18] , \wBMid108[17] , \wBMid108[16] , 
        \wBMid108[15] , \wBMid108[14] , \wBMid108[13] , \wBMid108[12] , 
        \wBMid108[11] , \wBMid108[10] , \wBMid108[9] , \wBMid108[8] , 
        \wBMid108[7] , \wBMid108[6] , \wBMid108[5] , \wBMid108[4] , 
        \wBMid108[3] , \wBMid108[2] , \wBMid108[1] , \wBMid108[0] }), .HiOut({
        \wRegInB108[31] , \wRegInB108[30] , \wRegInB108[29] , \wRegInB108[28] , 
        \wRegInB108[27] , \wRegInB108[26] , \wRegInB108[25] , \wRegInB108[24] , 
        \wRegInB108[23] , \wRegInB108[22] , \wRegInB108[21] , \wRegInB108[20] , 
        \wRegInB108[19] , \wRegInB108[18] , \wRegInB108[17] , \wRegInB108[16] , 
        \wRegInB108[15] , \wRegInB108[14] , \wRegInB108[13] , \wRegInB108[12] , 
        \wRegInB108[11] , \wRegInB108[10] , \wRegInB108[9] , \wRegInB108[8] , 
        \wRegInB108[7] , \wRegInB108[6] , \wRegInB108[5] , \wRegInB108[4] , 
        \wRegInB108[3] , \wRegInB108[2] , \wRegInB108[1] , \wRegInB108[0] }), 
        .LoOut({\wRegInA109[31] , \wRegInA109[30] , \wRegInA109[29] , 
        \wRegInA109[28] , \wRegInA109[27] , \wRegInA109[26] , \wRegInA109[25] , 
        \wRegInA109[24] , \wRegInA109[23] , \wRegInA109[22] , \wRegInA109[21] , 
        \wRegInA109[20] , \wRegInA109[19] , \wRegInA109[18] , \wRegInA109[17] , 
        \wRegInA109[16] , \wRegInA109[15] , \wRegInA109[14] , \wRegInA109[13] , 
        \wRegInA109[12] , \wRegInA109[11] , \wRegInA109[10] , \wRegInA109[9] , 
        \wRegInA109[8] , \wRegInA109[7] , \wRegInA109[6] , \wRegInA109[5] , 
        \wRegInA109[4] , \wRegInA109[3] , \wRegInA109[2] , \wRegInA109[1] , 
        \wRegInA109[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid113[31] , \wAMid113[30] , \wAMid113[29] , \wAMid113[28] , 
        \wAMid113[27] , \wAMid113[26] , \wAMid113[25] , \wAMid113[24] , 
        \wAMid113[23] , \wAMid113[22] , \wAMid113[21] , \wAMid113[20] , 
        \wAMid113[19] , \wAMid113[18] , \wAMid113[17] , \wAMid113[16] , 
        \wAMid113[15] , \wAMid113[14] , \wAMid113[13] , \wAMid113[12] , 
        \wAMid113[11] , \wAMid113[10] , \wAMid113[9] , \wAMid113[8] , 
        \wAMid113[7] , \wAMid113[6] , \wAMid113[5] , \wAMid113[4] , 
        \wAMid113[3] , \wAMid113[2] , \wAMid113[1] , \wAMid113[0] }), .BIn({
        \wBMid113[31] , \wBMid113[30] , \wBMid113[29] , \wBMid113[28] , 
        \wBMid113[27] , \wBMid113[26] , \wBMid113[25] , \wBMid113[24] , 
        \wBMid113[23] , \wBMid113[22] , \wBMid113[21] , \wBMid113[20] , 
        \wBMid113[19] , \wBMid113[18] , \wBMid113[17] , \wBMid113[16] , 
        \wBMid113[15] , \wBMid113[14] , \wBMid113[13] , \wBMid113[12] , 
        \wBMid113[11] , \wBMid113[10] , \wBMid113[9] , \wBMid113[8] , 
        \wBMid113[7] , \wBMid113[6] , \wBMid113[5] , \wBMid113[4] , 
        \wBMid113[3] , \wBMid113[2] , \wBMid113[1] , \wBMid113[0] }), .HiOut({
        \wRegInB113[31] , \wRegInB113[30] , \wRegInB113[29] , \wRegInB113[28] , 
        \wRegInB113[27] , \wRegInB113[26] , \wRegInB113[25] , \wRegInB113[24] , 
        \wRegInB113[23] , \wRegInB113[22] , \wRegInB113[21] , \wRegInB113[20] , 
        \wRegInB113[19] , \wRegInB113[18] , \wRegInB113[17] , \wRegInB113[16] , 
        \wRegInB113[15] , \wRegInB113[14] , \wRegInB113[13] , \wRegInB113[12] , 
        \wRegInB113[11] , \wRegInB113[10] , \wRegInB113[9] , \wRegInB113[8] , 
        \wRegInB113[7] , \wRegInB113[6] , \wRegInB113[5] , \wRegInB113[4] , 
        \wRegInB113[3] , \wRegInB113[2] , \wRegInB113[1] , \wRegInB113[0] }), 
        .LoOut({\wRegInA114[31] , \wRegInA114[30] , \wRegInA114[29] , 
        \wRegInA114[28] , \wRegInA114[27] , \wRegInA114[26] , \wRegInA114[25] , 
        \wRegInA114[24] , \wRegInA114[23] , \wRegInA114[22] , \wRegInA114[21] , 
        \wRegInA114[20] , \wRegInA114[19] , \wRegInA114[18] , \wRegInA114[17] , 
        \wRegInA114[16] , \wRegInA114[15] , \wRegInA114[14] , \wRegInA114[13] , 
        \wRegInA114[12] , \wRegInA114[11] , \wRegInA114[10] , \wRegInA114[9] , 
        \wRegInA114[8] , \wRegInA114[7] , \wRegInA114[6] , \wRegInA114[5] , 
        \wRegInA114[4] , \wRegInA114[3] , \wRegInA114[2] , \wRegInA114[1] , 
        \wRegInA114[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_90 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink91[31] , \ScanLink91[30] , \ScanLink91[29] , 
        \ScanLink91[28] , \ScanLink91[27] , \ScanLink91[26] , \ScanLink91[25] , 
        \ScanLink91[24] , \ScanLink91[23] , \ScanLink91[22] , \ScanLink91[21] , 
        \ScanLink91[20] , \ScanLink91[19] , \ScanLink91[18] , \ScanLink91[17] , 
        \ScanLink91[16] , \ScanLink91[15] , \ScanLink91[14] , \ScanLink91[13] , 
        \ScanLink91[12] , \ScanLink91[11] , \ScanLink91[10] , \ScanLink91[9] , 
        \ScanLink91[8] , \ScanLink91[7] , \ScanLink91[6] , \ScanLink91[5] , 
        \ScanLink91[4] , \ScanLink91[3] , \ScanLink91[2] , \ScanLink91[1] , 
        \ScanLink91[0] }), .ScanOut({\ScanLink90[31] , \ScanLink90[30] , 
        \ScanLink90[29] , \ScanLink90[28] , \ScanLink90[27] , \ScanLink90[26] , 
        \ScanLink90[25] , \ScanLink90[24] , \ScanLink90[23] , \ScanLink90[22] , 
        \ScanLink90[21] , \ScanLink90[20] , \ScanLink90[19] , \ScanLink90[18] , 
        \ScanLink90[17] , \ScanLink90[16] , \ScanLink90[15] , \ScanLink90[14] , 
        \ScanLink90[13] , \ScanLink90[12] , \ScanLink90[11] , \ScanLink90[10] , 
        \ScanLink90[9] , \ScanLink90[8] , \ScanLink90[7] , \ScanLink90[6] , 
        \ScanLink90[5] , \ScanLink90[4] , \ScanLink90[3] , \ScanLink90[2] , 
        \ScanLink90[1] , \ScanLink90[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB82[31] , \wRegInB82[30] , 
        \wRegInB82[29] , \wRegInB82[28] , \wRegInB82[27] , \wRegInB82[26] , 
        \wRegInB82[25] , \wRegInB82[24] , \wRegInB82[23] , \wRegInB82[22] , 
        \wRegInB82[21] , \wRegInB82[20] , \wRegInB82[19] , \wRegInB82[18] , 
        \wRegInB82[17] , \wRegInB82[16] , \wRegInB82[15] , \wRegInB82[14] , 
        \wRegInB82[13] , \wRegInB82[12] , \wRegInB82[11] , \wRegInB82[10] , 
        \wRegInB82[9] , \wRegInB82[8] , \wRegInB82[7] , \wRegInB82[6] , 
        \wRegInB82[5] , \wRegInB82[4] , \wRegInB82[3] , \wRegInB82[2] , 
        \wRegInB82[1] , \wRegInB82[0] }), .Out({\wBIn82[31] , \wBIn82[30] , 
        \wBIn82[29] , \wBIn82[28] , \wBIn82[27] , \wBIn82[26] , \wBIn82[25] , 
        \wBIn82[24] , \wBIn82[23] , \wBIn82[22] , \wBIn82[21] , \wBIn82[20] , 
        \wBIn82[19] , \wBIn82[18] , \wBIn82[17] , \wBIn82[16] , \wBIn82[15] , 
        \wBIn82[14] , \wBIn82[13] , \wBIn82[12] , \wBIn82[11] , \wBIn82[10] , 
        \wBIn82[9] , \wBIn82[8] , \wBIn82[7] , \wBIn82[6] , \wBIn82[5] , 
        \wBIn82[4] , \wBIn82[3] , \wBIn82[2] , \wBIn82[1] , \wBIn82[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid59[31] , \wAMid59[30] , \wAMid59[29] , \wAMid59[28] , 
        \wAMid59[27] , \wAMid59[26] , \wAMid59[25] , \wAMid59[24] , 
        \wAMid59[23] , \wAMid59[22] , \wAMid59[21] , \wAMid59[20] , 
        \wAMid59[19] , \wAMid59[18] , \wAMid59[17] , \wAMid59[16] , 
        \wAMid59[15] , \wAMid59[14] , \wAMid59[13] , \wAMid59[12] , 
        \wAMid59[11] , \wAMid59[10] , \wAMid59[9] , \wAMid59[8] , \wAMid59[7] , 
        \wAMid59[6] , \wAMid59[5] , \wAMid59[4] , \wAMid59[3] , \wAMid59[2] , 
        \wAMid59[1] , \wAMid59[0] }), .BIn({\wBMid59[31] , \wBMid59[30] , 
        \wBMid59[29] , \wBMid59[28] , \wBMid59[27] , \wBMid59[26] , 
        \wBMid59[25] , \wBMid59[24] , \wBMid59[23] , \wBMid59[22] , 
        \wBMid59[21] , \wBMid59[20] , \wBMid59[19] , \wBMid59[18] , 
        \wBMid59[17] , \wBMid59[16] , \wBMid59[15] , \wBMid59[14] , 
        \wBMid59[13] , \wBMid59[12] , \wBMid59[11] , \wBMid59[10] , 
        \wBMid59[9] , \wBMid59[8] , \wBMid59[7] , \wBMid59[6] , \wBMid59[5] , 
        \wBMid59[4] , \wBMid59[3] , \wBMid59[2] , \wBMid59[1] , \wBMid59[0] }), 
        .HiOut({\wRegInB59[31] , \wRegInB59[30] , \wRegInB59[29] , 
        \wRegInB59[28] , \wRegInB59[27] , \wRegInB59[26] , \wRegInB59[25] , 
        \wRegInB59[24] , \wRegInB59[23] , \wRegInB59[22] , \wRegInB59[21] , 
        \wRegInB59[20] , \wRegInB59[19] , \wRegInB59[18] , \wRegInB59[17] , 
        \wRegInB59[16] , \wRegInB59[15] , \wRegInB59[14] , \wRegInB59[13] , 
        \wRegInB59[12] , \wRegInB59[11] , \wRegInB59[10] , \wRegInB59[9] , 
        \wRegInB59[8] , \wRegInB59[7] , \wRegInB59[6] , \wRegInB59[5] , 
        \wRegInB59[4] , \wRegInB59[3] , \wRegInB59[2] , \wRegInB59[1] , 
        \wRegInB59[0] }), .LoOut({\wRegInA60[31] , \wRegInA60[30] , 
        \wRegInA60[29] , \wRegInA60[28] , \wRegInA60[27] , \wRegInA60[26] , 
        \wRegInA60[25] , \wRegInA60[24] , \wRegInA60[23] , \wRegInA60[22] , 
        \wRegInA60[21] , \wRegInA60[20] , \wRegInA60[19] , \wRegInA60[18] , 
        \wRegInA60[17] , \wRegInA60[16] , \wRegInA60[15] , \wRegInA60[14] , 
        \wRegInA60[13] , \wRegInA60[12] , \wRegInA60[11] , \wRegInA60[10] , 
        \wRegInA60[9] , \wRegInA60[8] , \wRegInA60[7] , \wRegInA60[6] , 
        \wRegInA60[5] , \wRegInA60[4] , \wRegInA60[3] , \wRegInA60[2] , 
        \wRegInA60[1] , \wRegInA60[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid10[31] , \wAMid10[30] , \wAMid10[29] , \wAMid10[28] , 
        \wAMid10[27] , \wAMid10[26] , \wAMid10[25] , \wAMid10[24] , 
        \wAMid10[23] , \wAMid10[22] , \wAMid10[21] , \wAMid10[20] , 
        \wAMid10[19] , \wAMid10[18] , \wAMid10[17] , \wAMid10[16] , 
        \wAMid10[15] , \wAMid10[14] , \wAMid10[13] , \wAMid10[12] , 
        \wAMid10[11] , \wAMid10[10] , \wAMid10[9] , \wAMid10[8] , \wAMid10[7] , 
        \wAMid10[6] , \wAMid10[5] , \wAMid10[4] , \wAMid10[3] , \wAMid10[2] , 
        \wAMid10[1] , \wAMid10[0] }), .BIn({\wBMid10[31] , \wBMid10[30] , 
        \wBMid10[29] , \wBMid10[28] , \wBMid10[27] , \wBMid10[26] , 
        \wBMid10[25] , \wBMid10[24] , \wBMid10[23] , \wBMid10[22] , 
        \wBMid10[21] , \wBMid10[20] , \wBMid10[19] , \wBMid10[18] , 
        \wBMid10[17] , \wBMid10[16] , \wBMid10[15] , \wBMid10[14] , 
        \wBMid10[13] , \wBMid10[12] , \wBMid10[11] , \wBMid10[10] , 
        \wBMid10[9] , \wBMid10[8] , \wBMid10[7] , \wBMid10[6] , \wBMid10[5] , 
        \wBMid10[4] , \wBMid10[3] , \wBMid10[2] , \wBMid10[1] , \wBMid10[0] }), 
        .HiOut({\wRegInB10[31] , \wRegInB10[30] , \wRegInB10[29] , 
        \wRegInB10[28] , \wRegInB10[27] , \wRegInB10[26] , \wRegInB10[25] , 
        \wRegInB10[24] , \wRegInB10[23] , \wRegInB10[22] , \wRegInB10[21] , 
        \wRegInB10[20] , \wRegInB10[19] , \wRegInB10[18] , \wRegInB10[17] , 
        \wRegInB10[16] , \wRegInB10[15] , \wRegInB10[14] , \wRegInB10[13] , 
        \wRegInB10[12] , \wRegInB10[11] , \wRegInB10[10] , \wRegInB10[9] , 
        \wRegInB10[8] , \wRegInB10[7] , \wRegInB10[6] , \wRegInB10[5] , 
        \wRegInB10[4] , \wRegInB10[3] , \wRegInB10[2] , \wRegInB10[1] , 
        \wRegInB10[0] }), .LoOut({\wRegInA11[31] , \wRegInA11[30] , 
        \wRegInA11[29] , \wRegInA11[28] , \wRegInA11[27] , \wRegInA11[26] , 
        \wRegInA11[25] , \wRegInA11[24] , \wRegInA11[23] , \wRegInA11[22] , 
        \wRegInA11[21] , \wRegInA11[20] , \wRegInA11[19] , \wRegInA11[18] , 
        \wRegInA11[17] , \wRegInA11[16] , \wRegInA11[15] , \wRegInA11[14] , 
        \wRegInA11[13] , \wRegInA11[12] , \wRegInA11[11] , \wRegInA11[10] , 
        \wRegInA11[9] , \wRegInA11[8] , \wRegInA11[7] , \wRegInA11[6] , 
        \wRegInA11[5] , \wRegInA11[4] , \wRegInA11[3] , \wRegInA11[2] , 
        \wRegInA11[1] , \wRegInA11[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid37[31] , \wAMid37[30] , \wAMid37[29] , \wAMid37[28] , 
        \wAMid37[27] , \wAMid37[26] , \wAMid37[25] , \wAMid37[24] , 
        \wAMid37[23] , \wAMid37[22] , \wAMid37[21] , \wAMid37[20] , 
        \wAMid37[19] , \wAMid37[18] , \wAMid37[17] , \wAMid37[16] , 
        \wAMid37[15] , \wAMid37[14] , \wAMid37[13] , \wAMid37[12] , 
        \wAMid37[11] , \wAMid37[10] , \wAMid37[9] , \wAMid37[8] , \wAMid37[7] , 
        \wAMid37[6] , \wAMid37[5] , \wAMid37[4] , \wAMid37[3] , \wAMid37[2] , 
        \wAMid37[1] , \wAMid37[0] }), .BIn({\wBMid37[31] , \wBMid37[30] , 
        \wBMid37[29] , \wBMid37[28] , \wBMid37[27] , \wBMid37[26] , 
        \wBMid37[25] , \wBMid37[24] , \wBMid37[23] , \wBMid37[22] , 
        \wBMid37[21] , \wBMid37[20] , \wBMid37[19] , \wBMid37[18] , 
        \wBMid37[17] , \wBMid37[16] , \wBMid37[15] , \wBMid37[14] , 
        \wBMid37[13] , \wBMid37[12] , \wBMid37[11] , \wBMid37[10] , 
        \wBMid37[9] , \wBMid37[8] , \wBMid37[7] , \wBMid37[6] , \wBMid37[5] , 
        \wBMid37[4] , \wBMid37[3] , \wBMid37[2] , \wBMid37[1] , \wBMid37[0] }), 
        .HiOut({\wRegInB37[31] , \wRegInB37[30] , \wRegInB37[29] , 
        \wRegInB37[28] , \wRegInB37[27] , \wRegInB37[26] , \wRegInB37[25] , 
        \wRegInB37[24] , \wRegInB37[23] , \wRegInB37[22] , \wRegInB37[21] , 
        \wRegInB37[20] , \wRegInB37[19] , \wRegInB37[18] , \wRegInB37[17] , 
        \wRegInB37[16] , \wRegInB37[15] , \wRegInB37[14] , \wRegInB37[13] , 
        \wRegInB37[12] , \wRegInB37[11] , \wRegInB37[10] , \wRegInB37[9] , 
        \wRegInB37[8] , \wRegInB37[7] , \wRegInB37[6] , \wRegInB37[5] , 
        \wRegInB37[4] , \wRegInB37[3] , \wRegInB37[2] , \wRegInB37[1] , 
        \wRegInB37[0] }), .LoOut({\wRegInA38[31] , \wRegInA38[30] , 
        \wRegInA38[29] , \wRegInA38[28] , \wRegInA38[27] , \wRegInA38[26] , 
        \wRegInA38[25] , \wRegInA38[24] , \wRegInA38[23] , \wRegInA38[22] , 
        \wRegInA38[21] , \wRegInA38[20] , \wRegInA38[19] , \wRegInA38[18] , 
        \wRegInA38[17] , \wRegInA38[16] , \wRegInA38[15] , \wRegInA38[14] , 
        \wRegInA38[13] , \wRegInA38[12] , \wRegInA38[11] , \wRegInA38[10] , 
        \wRegInA38[9] , \wRegInA38[8] , \wRegInA38[7] , \wRegInA38[6] , 
        \wRegInA38[5] , \wRegInA38[4] , \wRegInA38[3] , \wRegInA38[2] , 
        \wRegInA38[1] , \wRegInA38[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_232 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink233[31] , \ScanLink233[30] , \ScanLink233[29] , 
        \ScanLink233[28] , \ScanLink233[27] , \ScanLink233[26] , 
        \ScanLink233[25] , \ScanLink233[24] , \ScanLink233[23] , 
        \ScanLink233[22] , \ScanLink233[21] , \ScanLink233[20] , 
        \ScanLink233[19] , \ScanLink233[18] , \ScanLink233[17] , 
        \ScanLink233[16] , \ScanLink233[15] , \ScanLink233[14] , 
        \ScanLink233[13] , \ScanLink233[12] , \ScanLink233[11] , 
        \ScanLink233[10] , \ScanLink233[9] , \ScanLink233[8] , 
        \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , \ScanLink233[4] , 
        \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , \ScanLink233[0] 
        }), .ScanOut({\ScanLink232[31] , \ScanLink232[30] , \ScanLink232[29] , 
        \ScanLink232[28] , \ScanLink232[27] , \ScanLink232[26] , 
        \ScanLink232[25] , \ScanLink232[24] , \ScanLink232[23] , 
        \ScanLink232[22] , \ScanLink232[21] , \ScanLink232[20] , 
        \ScanLink232[19] , \ScanLink232[18] , \ScanLink232[17] , 
        \ScanLink232[16] , \ScanLink232[15] , \ScanLink232[14] , 
        \ScanLink232[13] , \ScanLink232[12] , \ScanLink232[11] , 
        \ScanLink232[10] , \ScanLink232[9] , \ScanLink232[8] , 
        \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , \ScanLink232[4] , 
        \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , \ScanLink232[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB11[31] , \wRegInB11[30] , \wRegInB11[29] , 
        \wRegInB11[28] , \wRegInB11[27] , \wRegInB11[26] , \wRegInB11[25] , 
        \wRegInB11[24] , \wRegInB11[23] , \wRegInB11[22] , \wRegInB11[21] , 
        \wRegInB11[20] , \wRegInB11[19] , \wRegInB11[18] , \wRegInB11[17] , 
        \wRegInB11[16] , \wRegInB11[15] , \wRegInB11[14] , \wRegInB11[13] , 
        \wRegInB11[12] , \wRegInB11[11] , \wRegInB11[10] , \wRegInB11[9] , 
        \wRegInB11[8] , \wRegInB11[7] , \wRegInB11[6] , \wRegInB11[5] , 
        \wRegInB11[4] , \wRegInB11[3] , \wRegInB11[2] , \wRegInB11[1] , 
        \wRegInB11[0] }), .Out({\wBIn11[31] , \wBIn11[30] , \wBIn11[29] , 
        \wBIn11[28] , \wBIn11[27] , \wBIn11[26] , \wBIn11[25] , \wBIn11[24] , 
        \wBIn11[23] , \wBIn11[22] , \wBIn11[21] , \wBIn11[20] , \wBIn11[19] , 
        \wBIn11[18] , \wBIn11[17] , \wBIn11[16] , \wBIn11[15] , \wBIn11[14] , 
        \wBIn11[13] , \wBIn11[12] , \wBIn11[11] , \wBIn11[10] , \wBIn11[9] , 
        \wBIn11[8] , \wBIn11[7] , \wBIn11[6] , \wBIn11[5] , \wBIn11[4] , 
        \wBIn11[3] , \wBIn11[2] , \wBIn11[1] , \wBIn11[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_102 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink103[31] , \ScanLink103[30] , \ScanLink103[29] , 
        \ScanLink103[28] , \ScanLink103[27] , \ScanLink103[26] , 
        \ScanLink103[25] , \ScanLink103[24] , \ScanLink103[23] , 
        \ScanLink103[22] , \ScanLink103[21] , \ScanLink103[20] , 
        \ScanLink103[19] , \ScanLink103[18] , \ScanLink103[17] , 
        \ScanLink103[16] , \ScanLink103[15] , \ScanLink103[14] , 
        \ScanLink103[13] , \ScanLink103[12] , \ScanLink103[11] , 
        \ScanLink103[10] , \ScanLink103[9] , \ScanLink103[8] , 
        \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , \ScanLink103[4] , 
        \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , \ScanLink103[0] 
        }), .ScanOut({\ScanLink102[31] , \ScanLink102[30] , \ScanLink102[29] , 
        \ScanLink102[28] , \ScanLink102[27] , \ScanLink102[26] , 
        \ScanLink102[25] , \ScanLink102[24] , \ScanLink102[23] , 
        \ScanLink102[22] , \ScanLink102[21] , \ScanLink102[20] , 
        \ScanLink102[19] , \ScanLink102[18] , \ScanLink102[17] , 
        \ScanLink102[16] , \ScanLink102[15] , \ScanLink102[14] , 
        \ScanLink102[13] , \ScanLink102[12] , \ScanLink102[11] , 
        \ScanLink102[10] , \ScanLink102[9] , \ScanLink102[8] , 
        \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , \ScanLink102[4] , 
        \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , \ScanLink102[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB76[31] , \wRegInB76[30] , \wRegInB76[29] , 
        \wRegInB76[28] , \wRegInB76[27] , \wRegInB76[26] , \wRegInB76[25] , 
        \wRegInB76[24] , \wRegInB76[23] , \wRegInB76[22] , \wRegInB76[21] , 
        \wRegInB76[20] , \wRegInB76[19] , \wRegInB76[18] , \wRegInB76[17] , 
        \wRegInB76[16] , \wRegInB76[15] , \wRegInB76[14] , \wRegInB76[13] , 
        \wRegInB76[12] , \wRegInB76[11] , \wRegInB76[10] , \wRegInB76[9] , 
        \wRegInB76[8] , \wRegInB76[7] , \wRegInB76[6] , \wRegInB76[5] , 
        \wRegInB76[4] , \wRegInB76[3] , \wRegInB76[2] , \wRegInB76[1] , 
        \wRegInB76[0] }), .Out({\wBIn76[31] , \wBIn76[30] , \wBIn76[29] , 
        \wBIn76[28] , \wBIn76[27] , \wBIn76[26] , \wBIn76[25] , \wBIn76[24] , 
        \wBIn76[23] , \wBIn76[22] , \wBIn76[21] , \wBIn76[20] , \wBIn76[19] , 
        \wBIn76[18] , \wBIn76[17] , \wBIn76[16] , \wBIn76[15] , \wBIn76[14] , 
        \wBIn76[13] , \wBIn76[12] , \wBIn76[11] , \wBIn76[10] , \wBIn76[9] , 
        \wBIn76[8] , \wBIn76[7] , \wBIn76[6] , \wBIn76[5] , \wBIn76[4] , 
        \wBIn76[3] , \wBIn76[2] , \wBIn76[1] , \wBIn76[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_125 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink126[31] , \ScanLink126[30] , \ScanLink126[29] , 
        \ScanLink126[28] , \ScanLink126[27] , \ScanLink126[26] , 
        \ScanLink126[25] , \ScanLink126[24] , \ScanLink126[23] , 
        \ScanLink126[22] , \ScanLink126[21] , \ScanLink126[20] , 
        \ScanLink126[19] , \ScanLink126[18] , \ScanLink126[17] , 
        \ScanLink126[16] , \ScanLink126[15] , \ScanLink126[14] , 
        \ScanLink126[13] , \ScanLink126[12] , \ScanLink126[11] , 
        \ScanLink126[10] , \ScanLink126[9] , \ScanLink126[8] , 
        \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , \ScanLink126[4] , 
        \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , \ScanLink126[0] 
        }), .ScanOut({\ScanLink125[31] , \ScanLink125[30] , \ScanLink125[29] , 
        \ScanLink125[28] , \ScanLink125[27] , \ScanLink125[26] , 
        \ScanLink125[25] , \ScanLink125[24] , \ScanLink125[23] , 
        \ScanLink125[22] , \ScanLink125[21] , \ScanLink125[20] , 
        \ScanLink125[19] , \ScanLink125[18] , \ScanLink125[17] , 
        \ScanLink125[16] , \ScanLink125[15] , \ScanLink125[14] , 
        \ScanLink125[13] , \ScanLink125[12] , \ScanLink125[11] , 
        \ScanLink125[10] , \ScanLink125[9] , \ScanLink125[8] , 
        \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , \ScanLink125[4] , 
        \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , \ScanLink125[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA65[31] , \wRegInA65[30] , \wRegInA65[29] , 
        \wRegInA65[28] , \wRegInA65[27] , \wRegInA65[26] , \wRegInA65[25] , 
        \wRegInA65[24] , \wRegInA65[23] , \wRegInA65[22] , \wRegInA65[21] , 
        \wRegInA65[20] , \wRegInA65[19] , \wRegInA65[18] , \wRegInA65[17] , 
        \wRegInA65[16] , \wRegInA65[15] , \wRegInA65[14] , \wRegInA65[13] , 
        \wRegInA65[12] , \wRegInA65[11] , \wRegInA65[10] , \wRegInA65[9] , 
        \wRegInA65[8] , \wRegInA65[7] , \wRegInA65[6] , \wRegInA65[5] , 
        \wRegInA65[4] , \wRegInA65[3] , \wRegInA65[2] , \wRegInA65[1] , 
        \wRegInA65[0] }), .Out({\wAIn65[31] , \wAIn65[30] , \wAIn65[29] , 
        \wAIn65[28] , \wAIn65[27] , \wAIn65[26] , \wAIn65[25] , \wAIn65[24] , 
        \wAIn65[23] , \wAIn65[22] , \wAIn65[21] , \wAIn65[20] , \wAIn65[19] , 
        \wAIn65[18] , \wAIn65[17] , \wAIn65[16] , \wAIn65[15] , \wAIn65[14] , 
        \wAIn65[13] , \wAIn65[12] , \wAIn65[11] , \wAIn65[10] , \wAIn65[9] , 
        \wAIn65[8] , \wAIn65[7] , \wAIn65[6] , \wAIn65[5] , \wAIn65[4] , 
        \wAIn65[3] , \wAIn65[2] , \wAIn65[1] , \wAIn65[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_52 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink53[31] , \ScanLink53[30] , \ScanLink53[29] , 
        \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , \ScanLink53[25] , 
        \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , \ScanLink53[21] , 
        \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , \ScanLink53[17] , 
        \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , \ScanLink53[13] , 
        \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , \ScanLink53[9] , 
        \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , \ScanLink53[5] , 
        \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , \ScanLink53[1] , 
        \ScanLink53[0] }), .ScanOut({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB101[31] , \wRegInB101[30] , 
        \wRegInB101[29] , \wRegInB101[28] , \wRegInB101[27] , \wRegInB101[26] , 
        \wRegInB101[25] , \wRegInB101[24] , \wRegInB101[23] , \wRegInB101[22] , 
        \wRegInB101[21] , \wRegInB101[20] , \wRegInB101[19] , \wRegInB101[18] , 
        \wRegInB101[17] , \wRegInB101[16] , \wRegInB101[15] , \wRegInB101[14] , 
        \wRegInB101[13] , \wRegInB101[12] , \wRegInB101[11] , \wRegInB101[10] , 
        \wRegInB101[9] , \wRegInB101[8] , \wRegInB101[7] , \wRegInB101[6] , 
        \wRegInB101[5] , \wRegInB101[4] , \wRegInB101[3] , \wRegInB101[2] , 
        \wRegInB101[1] , \wRegInB101[0] }), .Out({\wBIn101[31] , \wBIn101[30] , 
        \wBIn101[29] , \wBIn101[28] , \wBIn101[27] , \wBIn101[26] , 
        \wBIn101[25] , \wBIn101[24] , \wBIn101[23] , \wBIn101[22] , 
        \wBIn101[21] , \wBIn101[20] , \wBIn101[19] , \wBIn101[18] , 
        \wBIn101[17] , \wBIn101[16] , \wBIn101[15] , \wBIn101[14] , 
        \wBIn101[13] , \wBIn101[12] , \wBIn101[11] , \wBIn101[10] , 
        \wBIn101[9] , \wBIn101[8] , \wBIn101[7] , \wBIn101[6] , \wBIn101[5] , 
        \wBIn101[4] , \wBIn101[3] , \wBIn101[2] , \wBIn101[1] , \wBIn101[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_75 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink76[31] , \ScanLink76[30] , \ScanLink76[29] , 
        \ScanLink76[28] , \ScanLink76[27] , \ScanLink76[26] , \ScanLink76[25] , 
        \ScanLink76[24] , \ScanLink76[23] , \ScanLink76[22] , \ScanLink76[21] , 
        \ScanLink76[20] , \ScanLink76[19] , \ScanLink76[18] , \ScanLink76[17] , 
        \ScanLink76[16] , \ScanLink76[15] , \ScanLink76[14] , \ScanLink76[13] , 
        \ScanLink76[12] , \ScanLink76[11] , \ScanLink76[10] , \ScanLink76[9] , 
        \ScanLink76[8] , \ScanLink76[7] , \ScanLink76[6] , \ScanLink76[5] , 
        \ScanLink76[4] , \ScanLink76[3] , \ScanLink76[2] , \ScanLink76[1] , 
        \ScanLink76[0] }), .ScanOut({\ScanLink75[31] , \ScanLink75[30] , 
        \ScanLink75[29] , \ScanLink75[28] , \ScanLink75[27] , \ScanLink75[26] , 
        \ScanLink75[25] , \ScanLink75[24] , \ScanLink75[23] , \ScanLink75[22] , 
        \ScanLink75[21] , \ScanLink75[20] , \ScanLink75[19] , \ScanLink75[18] , 
        \ScanLink75[17] , \ScanLink75[16] , \ScanLink75[15] , \ScanLink75[14] , 
        \ScanLink75[13] , \ScanLink75[12] , \ScanLink75[11] , \ScanLink75[10] , 
        \ScanLink75[9] , \ScanLink75[8] , \ScanLink75[7] , \ScanLink75[6] , 
        \ScanLink75[5] , \ScanLink75[4] , \ScanLink75[3] , \ScanLink75[2] , 
        \ScanLink75[1] , \ScanLink75[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA90[31] , \wRegInA90[30] , 
        \wRegInA90[29] , \wRegInA90[28] , \wRegInA90[27] , \wRegInA90[26] , 
        \wRegInA90[25] , \wRegInA90[24] , \wRegInA90[23] , \wRegInA90[22] , 
        \wRegInA90[21] , \wRegInA90[20] , \wRegInA90[19] , \wRegInA90[18] , 
        \wRegInA90[17] , \wRegInA90[16] , \wRegInA90[15] , \wRegInA90[14] , 
        \wRegInA90[13] , \wRegInA90[12] , \wRegInA90[11] , \wRegInA90[10] , 
        \wRegInA90[9] , \wRegInA90[8] , \wRegInA90[7] , \wRegInA90[6] , 
        \wRegInA90[5] , \wRegInA90[4] , \wRegInA90[3] , \wRegInA90[2] , 
        \wRegInA90[1] , \wRegInA90[0] }), .Out({\wAIn90[31] , \wAIn90[30] , 
        \wAIn90[29] , \wAIn90[28] , \wAIn90[27] , \wAIn90[26] , \wAIn90[25] , 
        \wAIn90[24] , \wAIn90[23] , \wAIn90[22] , \wAIn90[21] , \wAIn90[20] , 
        \wAIn90[19] , \wAIn90[18] , \wAIn90[17] , \wAIn90[16] , \wAIn90[15] , 
        \wAIn90[14] , \wAIn90[13] , \wAIn90[12] , \wAIn90[11] , \wAIn90[10] , 
        \wAIn90[9] , \wAIn90[8] , \wAIn90[7] , \wAIn90[6] , \wAIn90[5] , 
        \wAIn90[4] , \wAIn90[3] , \wAIn90[2] , \wAIn90[1] , \wAIn90[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid25[31] , \wAMid25[30] , \wAMid25[29] , \wAMid25[28] , 
        \wAMid25[27] , \wAMid25[26] , \wAMid25[25] , \wAMid25[24] , 
        \wAMid25[23] , \wAMid25[22] , \wAMid25[21] , \wAMid25[20] , 
        \wAMid25[19] , \wAMid25[18] , \wAMid25[17] , \wAMid25[16] , 
        \wAMid25[15] , \wAMid25[14] , \wAMid25[13] , \wAMid25[12] , 
        \wAMid25[11] , \wAMid25[10] , \wAMid25[9] , \wAMid25[8] , \wAMid25[7] , 
        \wAMid25[6] , \wAMid25[5] , \wAMid25[4] , \wAMid25[3] , \wAMid25[2] , 
        \wAMid25[1] , \wAMid25[0] }), .BIn({\wBMid25[31] , \wBMid25[30] , 
        \wBMid25[29] , \wBMid25[28] , \wBMid25[27] , \wBMid25[26] , 
        \wBMid25[25] , \wBMid25[24] , \wBMid25[23] , \wBMid25[22] , 
        \wBMid25[21] , \wBMid25[20] , \wBMid25[19] , \wBMid25[18] , 
        \wBMid25[17] , \wBMid25[16] , \wBMid25[15] , \wBMid25[14] , 
        \wBMid25[13] , \wBMid25[12] , \wBMid25[11] , \wBMid25[10] , 
        \wBMid25[9] , \wBMid25[8] , \wBMid25[7] , \wBMid25[6] , \wBMid25[5] , 
        \wBMid25[4] , \wBMid25[3] , \wBMid25[2] , \wBMid25[1] , \wBMid25[0] }), 
        .HiOut({\wRegInB25[31] , \wRegInB25[30] , \wRegInB25[29] , 
        \wRegInB25[28] , \wRegInB25[27] , \wRegInB25[26] , \wRegInB25[25] , 
        \wRegInB25[24] , \wRegInB25[23] , \wRegInB25[22] , \wRegInB25[21] , 
        \wRegInB25[20] , \wRegInB25[19] , \wRegInB25[18] , \wRegInB25[17] , 
        \wRegInB25[16] , \wRegInB25[15] , \wRegInB25[14] , \wRegInB25[13] , 
        \wRegInB25[12] , \wRegInB25[11] , \wRegInB25[10] , \wRegInB25[9] , 
        \wRegInB25[8] , \wRegInB25[7] , \wRegInB25[6] , \wRegInB25[5] , 
        \wRegInB25[4] , \wRegInB25[3] , \wRegInB25[2] , \wRegInB25[1] , 
        \wRegInB25[0] }), .LoOut({\wRegInA26[31] , \wRegInA26[30] , 
        \wRegInA26[29] , \wRegInA26[28] , \wRegInA26[27] , \wRegInA26[26] , 
        \wRegInA26[25] , \wRegInA26[24] , \wRegInA26[23] , \wRegInA26[22] , 
        \wRegInA26[21] , \wRegInA26[20] , \wRegInA26[19] , \wRegInA26[18] , 
        \wRegInA26[17] , \wRegInA26[16] , \wRegInA26[15] , \wRegInA26[14] , 
        \wRegInA26[13] , \wRegInA26[12] , \wRegInA26[11] , \wRegInA26[10] , 
        \wRegInA26[9] , \wRegInA26[8] , \wRegInA26[7] , \wRegInA26[6] , 
        \wRegInA26[5] , \wRegInA26[4] , \wRegInA26[3] , \wRegInA26[2] , 
        \wRegInA26[1] , \wRegInA26[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid89[31] , \wAMid89[30] , \wAMid89[29] , \wAMid89[28] , 
        \wAMid89[27] , \wAMid89[26] , \wAMid89[25] , \wAMid89[24] , 
        \wAMid89[23] , \wAMid89[22] , \wAMid89[21] , \wAMid89[20] , 
        \wAMid89[19] , \wAMid89[18] , \wAMid89[17] , \wAMid89[16] , 
        \wAMid89[15] , \wAMid89[14] , \wAMid89[13] , \wAMid89[12] , 
        \wAMid89[11] , \wAMid89[10] , \wAMid89[9] , \wAMid89[8] , \wAMid89[7] , 
        \wAMid89[6] , \wAMid89[5] , \wAMid89[4] , \wAMid89[3] , \wAMid89[2] , 
        \wAMid89[1] , \wAMid89[0] }), .BIn({\wBMid89[31] , \wBMid89[30] , 
        \wBMid89[29] , \wBMid89[28] , \wBMid89[27] , \wBMid89[26] , 
        \wBMid89[25] , \wBMid89[24] , \wBMid89[23] , \wBMid89[22] , 
        \wBMid89[21] , \wBMid89[20] , \wBMid89[19] , \wBMid89[18] , 
        \wBMid89[17] , \wBMid89[16] , \wBMid89[15] , \wBMid89[14] , 
        \wBMid89[13] , \wBMid89[12] , \wBMid89[11] , \wBMid89[10] , 
        \wBMid89[9] , \wBMid89[8] , \wBMid89[7] , \wBMid89[6] , \wBMid89[5] , 
        \wBMid89[4] , \wBMid89[3] , \wBMid89[2] , \wBMid89[1] , \wBMid89[0] }), 
        .HiOut({\wRegInB89[31] , \wRegInB89[30] , \wRegInB89[29] , 
        \wRegInB89[28] , \wRegInB89[27] , \wRegInB89[26] , \wRegInB89[25] , 
        \wRegInB89[24] , \wRegInB89[23] , \wRegInB89[22] , \wRegInB89[21] , 
        \wRegInB89[20] , \wRegInB89[19] , \wRegInB89[18] , \wRegInB89[17] , 
        \wRegInB89[16] , \wRegInB89[15] , \wRegInB89[14] , \wRegInB89[13] , 
        \wRegInB89[12] , \wRegInB89[11] , \wRegInB89[10] , \wRegInB89[9] , 
        \wRegInB89[8] , \wRegInB89[7] , \wRegInB89[6] , \wRegInB89[5] , 
        \wRegInB89[4] , \wRegInB89[3] , \wRegInB89[2] , \wRegInB89[1] , 
        \wRegInB89[0] }), .LoOut({\wRegInA90[31] , \wRegInA90[30] , 
        \wRegInA90[29] , \wRegInA90[28] , \wRegInA90[27] , \wRegInA90[26] , 
        \wRegInA90[25] , \wRegInA90[24] , \wRegInA90[23] , \wRegInA90[22] , 
        \wRegInA90[21] , \wRegInA90[20] , \wRegInA90[19] , \wRegInA90[18] , 
        \wRegInA90[17] , \wRegInA90[16] , \wRegInA90[15] , \wRegInA90[14] , 
        \wRegInA90[13] , \wRegInA90[12] , \wRegInA90[11] , \wRegInA90[10] , 
        \wRegInA90[9] , \wRegInA90[8] , \wRegInA90[7] , \wRegInA90[6] , 
        \wRegInA90[5] , \wRegInA90[4] , \wRegInA90[3] , \wRegInA90[2] , 
        \wRegInA90[1] , \wRegInA90[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_215 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink216[31] , \ScanLink216[30] , \ScanLink216[29] , 
        \ScanLink216[28] , \ScanLink216[27] , \ScanLink216[26] , 
        \ScanLink216[25] , \ScanLink216[24] , \ScanLink216[23] , 
        \ScanLink216[22] , \ScanLink216[21] , \ScanLink216[20] , 
        \ScanLink216[19] , \ScanLink216[18] , \ScanLink216[17] , 
        \ScanLink216[16] , \ScanLink216[15] , \ScanLink216[14] , 
        \ScanLink216[13] , \ScanLink216[12] , \ScanLink216[11] , 
        \ScanLink216[10] , \ScanLink216[9] , \ScanLink216[8] , 
        \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , \ScanLink216[4] , 
        \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , \ScanLink216[0] 
        }), .ScanOut({\ScanLink215[31] , \ScanLink215[30] , \ScanLink215[29] , 
        \ScanLink215[28] , \ScanLink215[27] , \ScanLink215[26] , 
        \ScanLink215[25] , \ScanLink215[24] , \ScanLink215[23] , 
        \ScanLink215[22] , \ScanLink215[21] , \ScanLink215[20] , 
        \ScanLink215[19] , \ScanLink215[18] , \ScanLink215[17] , 
        \ScanLink215[16] , \ScanLink215[15] , \ScanLink215[14] , 
        \ScanLink215[13] , \ScanLink215[12] , \ScanLink215[11] , 
        \ScanLink215[10] , \ScanLink215[9] , \ScanLink215[8] , 
        \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , \ScanLink215[4] , 
        \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , \ScanLink215[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA20[31] , \wRegInA20[30] , \wRegInA20[29] , 
        \wRegInA20[28] , \wRegInA20[27] , \wRegInA20[26] , \wRegInA20[25] , 
        \wRegInA20[24] , \wRegInA20[23] , \wRegInA20[22] , \wRegInA20[21] , 
        \wRegInA20[20] , \wRegInA20[19] , \wRegInA20[18] , \wRegInA20[17] , 
        \wRegInA20[16] , \wRegInA20[15] , \wRegInA20[14] , \wRegInA20[13] , 
        \wRegInA20[12] , \wRegInA20[11] , \wRegInA20[10] , \wRegInA20[9] , 
        \wRegInA20[8] , \wRegInA20[7] , \wRegInA20[6] , \wRegInA20[5] , 
        \wRegInA20[4] , \wRegInA20[3] , \wRegInA20[2] , \wRegInA20[1] , 
        \wRegInA20[0] }), .Out({\wAIn20[31] , \wAIn20[30] , \wAIn20[29] , 
        \wAIn20[28] , \wAIn20[27] , \wAIn20[26] , \wAIn20[25] , \wAIn20[24] , 
        \wAIn20[23] , \wAIn20[22] , \wAIn20[21] , \wAIn20[20] , \wAIn20[19] , 
        \wAIn20[18] , \wAIn20[17] , \wAIn20[16] , \wAIn20[15] , \wAIn20[14] , 
        \wAIn20[13] , \wAIn20[12] , \wAIn20[11] , \wAIn20[10] , \wAIn20[9] , 
        \wAIn20[8] , \wAIn20[7] , \wAIn20[6] , \wAIn20[5] , \wAIn20[4] , 
        \wAIn20[3] , \wAIn20[2] , \wAIn20[1] , \wAIn20[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_189 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink190[31] , \ScanLink190[30] , \ScanLink190[29] , 
        \ScanLink190[28] , \ScanLink190[27] , \ScanLink190[26] , 
        \ScanLink190[25] , \ScanLink190[24] , \ScanLink190[23] , 
        \ScanLink190[22] , \ScanLink190[21] , \ScanLink190[20] , 
        \ScanLink190[19] , \ScanLink190[18] , \ScanLink190[17] , 
        \ScanLink190[16] , \ScanLink190[15] , \ScanLink190[14] , 
        \ScanLink190[13] , \ScanLink190[12] , \ScanLink190[11] , 
        \ScanLink190[10] , \ScanLink190[9] , \ScanLink190[8] , 
        \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , \ScanLink190[4] , 
        \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , \ScanLink190[0] 
        }), .ScanOut({\ScanLink189[31] , \ScanLink189[30] , \ScanLink189[29] , 
        \ScanLink189[28] , \ScanLink189[27] , \ScanLink189[26] , 
        \ScanLink189[25] , \ScanLink189[24] , \ScanLink189[23] , 
        \ScanLink189[22] , \ScanLink189[21] , \ScanLink189[20] , 
        \ScanLink189[19] , \ScanLink189[18] , \ScanLink189[17] , 
        \ScanLink189[16] , \ScanLink189[15] , \ScanLink189[14] , 
        \ScanLink189[13] , \ScanLink189[12] , \ScanLink189[11] , 
        \ScanLink189[10] , \ScanLink189[9] , \ScanLink189[8] , 
        \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , \ScanLink189[4] , 
        \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , \ScanLink189[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA33[31] , \wRegInA33[30] , \wRegInA33[29] , 
        \wRegInA33[28] , \wRegInA33[27] , \wRegInA33[26] , \wRegInA33[25] , 
        \wRegInA33[24] , \wRegInA33[23] , \wRegInA33[22] , \wRegInA33[21] , 
        \wRegInA33[20] , \wRegInA33[19] , \wRegInA33[18] , \wRegInA33[17] , 
        \wRegInA33[16] , \wRegInA33[15] , \wRegInA33[14] , \wRegInA33[13] , 
        \wRegInA33[12] , \wRegInA33[11] , \wRegInA33[10] , \wRegInA33[9] , 
        \wRegInA33[8] , \wRegInA33[7] , \wRegInA33[6] , \wRegInA33[5] , 
        \wRegInA33[4] , \wRegInA33[3] , \wRegInA33[2] , \wRegInA33[1] , 
        \wRegInA33[0] }), .Out({\wAIn33[31] , \wAIn33[30] , \wAIn33[29] , 
        \wAIn33[28] , \wAIn33[27] , \wAIn33[26] , \wAIn33[25] , \wAIn33[24] , 
        \wAIn33[23] , \wAIn33[22] , \wAIn33[21] , \wAIn33[20] , \wAIn33[19] , 
        \wAIn33[18] , \wAIn33[17] , \wAIn33[16] , \wAIn33[15] , \wAIn33[14] , 
        \wAIn33[13] , \wAIn33[12] , \wAIn33[11] , \wAIn33[10] , \wAIn33[9] , 
        \wAIn33[8] , \wAIn33[7] , \wAIn33[6] , \wAIn33[5] , \wAIn33[4] , 
        \wAIn33[3] , \wAIn33[2] , \wAIn33[1] , \wAIn33[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_220 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink221[31] , \ScanLink221[30] , \ScanLink221[29] , 
        \ScanLink221[28] , \ScanLink221[27] , \ScanLink221[26] , 
        \ScanLink221[25] , \ScanLink221[24] , \ScanLink221[23] , 
        \ScanLink221[22] , \ScanLink221[21] , \ScanLink221[20] , 
        \ScanLink221[19] , \ScanLink221[18] , \ScanLink221[17] , 
        \ScanLink221[16] , \ScanLink221[15] , \ScanLink221[14] , 
        \ScanLink221[13] , \ScanLink221[12] , \ScanLink221[11] , 
        \ScanLink221[10] , \ScanLink221[9] , \ScanLink221[8] , 
        \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , \ScanLink221[4] , 
        \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , \ScanLink221[0] 
        }), .ScanOut({\ScanLink220[31] , \ScanLink220[30] , \ScanLink220[29] , 
        \ScanLink220[28] , \ScanLink220[27] , \ScanLink220[26] , 
        \ScanLink220[25] , \ScanLink220[24] , \ScanLink220[23] , 
        \ScanLink220[22] , \ScanLink220[21] , \ScanLink220[20] , 
        \ScanLink220[19] , \ScanLink220[18] , \ScanLink220[17] , 
        \ScanLink220[16] , \ScanLink220[15] , \ScanLink220[14] , 
        \ScanLink220[13] , \ScanLink220[12] , \ScanLink220[11] , 
        \ScanLink220[10] , \ScanLink220[9] , \ScanLink220[8] , 
        \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , \ScanLink220[4] , 
        \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , \ScanLink220[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB17[31] , \wRegInB17[30] , \wRegInB17[29] , 
        \wRegInB17[28] , \wRegInB17[27] , \wRegInB17[26] , \wRegInB17[25] , 
        \wRegInB17[24] , \wRegInB17[23] , \wRegInB17[22] , \wRegInB17[21] , 
        \wRegInB17[20] , \wRegInB17[19] , \wRegInB17[18] , \wRegInB17[17] , 
        \wRegInB17[16] , \wRegInB17[15] , \wRegInB17[14] , \wRegInB17[13] , 
        \wRegInB17[12] , \wRegInB17[11] , \wRegInB17[10] , \wRegInB17[9] , 
        \wRegInB17[8] , \wRegInB17[7] , \wRegInB17[6] , \wRegInB17[5] , 
        \wRegInB17[4] , \wRegInB17[3] , \wRegInB17[2] , \wRegInB17[1] , 
        \wRegInB17[0] }), .Out({\wBIn17[31] , \wBIn17[30] , \wBIn17[29] , 
        \wBIn17[28] , \wBIn17[27] , \wBIn17[26] , \wBIn17[25] , \wBIn17[24] , 
        \wBIn17[23] , \wBIn17[22] , \wBIn17[21] , \wBIn17[20] , \wBIn17[19] , 
        \wBIn17[18] , \wBIn17[17] , \wBIn17[16] , \wBIn17[15] , \wBIn17[14] , 
        \wBIn17[13] , \wBIn17[12] , \wBIn17[11] , \wBIn17[10] , \wBIn17[9] , 
        \wBIn17[8] , \wBIn17[7] , \wBIn17[6] , \wBIn17[5] , \wBIn17[4] , 
        \wBIn17[3] , \wBIn17[2] , \wBIn17[1] , \wBIn17[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_110 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink111[31] , \ScanLink111[30] , \ScanLink111[29] , 
        \ScanLink111[28] , \ScanLink111[27] , \ScanLink111[26] , 
        \ScanLink111[25] , \ScanLink111[24] , \ScanLink111[23] , 
        \ScanLink111[22] , \ScanLink111[21] , \ScanLink111[20] , 
        \ScanLink111[19] , \ScanLink111[18] , \ScanLink111[17] , 
        \ScanLink111[16] , \ScanLink111[15] , \ScanLink111[14] , 
        \ScanLink111[13] , \ScanLink111[12] , \ScanLink111[11] , 
        \ScanLink111[10] , \ScanLink111[9] , \ScanLink111[8] , 
        \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , \ScanLink111[4] , 
        \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , \ScanLink111[0] 
        }), .ScanOut({\ScanLink110[31] , \ScanLink110[30] , \ScanLink110[29] , 
        \ScanLink110[28] , \ScanLink110[27] , \ScanLink110[26] , 
        \ScanLink110[25] , \ScanLink110[24] , \ScanLink110[23] , 
        \ScanLink110[22] , \ScanLink110[21] , \ScanLink110[20] , 
        \ScanLink110[19] , \ScanLink110[18] , \ScanLink110[17] , 
        \ScanLink110[16] , \ScanLink110[15] , \ScanLink110[14] , 
        \ScanLink110[13] , \ScanLink110[12] , \ScanLink110[11] , 
        \ScanLink110[10] , \ScanLink110[9] , \ScanLink110[8] , 
        \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , \ScanLink110[4] , 
        \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , \ScanLink110[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB72[31] , \wRegInB72[30] , \wRegInB72[29] , 
        \wRegInB72[28] , \wRegInB72[27] , \wRegInB72[26] , \wRegInB72[25] , 
        \wRegInB72[24] , \wRegInB72[23] , \wRegInB72[22] , \wRegInB72[21] , 
        \wRegInB72[20] , \wRegInB72[19] , \wRegInB72[18] , \wRegInB72[17] , 
        \wRegInB72[16] , \wRegInB72[15] , \wRegInB72[14] , \wRegInB72[13] , 
        \wRegInB72[12] , \wRegInB72[11] , \wRegInB72[10] , \wRegInB72[9] , 
        \wRegInB72[8] , \wRegInB72[7] , \wRegInB72[6] , \wRegInB72[5] , 
        \wRegInB72[4] , \wRegInB72[3] , \wRegInB72[2] , \wRegInB72[1] , 
        \wRegInB72[0] }), .Out({\wBIn72[31] , \wBIn72[30] , \wBIn72[29] , 
        \wBIn72[28] , \wBIn72[27] , \wBIn72[26] , \wBIn72[25] , \wBIn72[24] , 
        \wBIn72[23] , \wBIn72[22] , \wBIn72[21] , \wBIn72[20] , \wBIn72[19] , 
        \wBIn72[18] , \wBIn72[17] , \wBIn72[16] , \wBIn72[15] , \wBIn72[14] , 
        \wBIn72[13] , \wBIn72[12] , \wBIn72[11] , \wBIn72[10] , \wBIn72[9] , 
        \wBIn72[8] , \wBIn72[7] , \wBIn72[6] , \wBIn72[5] , \wBIn72[4] , 
        \wBIn72[3] , \wBIn72[2] , \wBIn72[1] , \wBIn72[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_40 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink41[31] , \ScanLink41[30] , \ScanLink41[29] , 
        \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , \ScanLink41[25] , 
        \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , \ScanLink41[21] , 
        \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , \ScanLink41[17] , 
        \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , \ScanLink41[13] , 
        \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , \ScanLink41[9] , 
        \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , \ScanLink41[5] , 
        \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , \ScanLink41[1] , 
        \ScanLink41[0] }), .ScanOut({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB107[31] , \wRegInB107[30] , 
        \wRegInB107[29] , \wRegInB107[28] , \wRegInB107[27] , \wRegInB107[26] , 
        \wRegInB107[25] , \wRegInB107[24] , \wRegInB107[23] , \wRegInB107[22] , 
        \wRegInB107[21] , \wRegInB107[20] , \wRegInB107[19] , \wRegInB107[18] , 
        \wRegInB107[17] , \wRegInB107[16] , \wRegInB107[15] , \wRegInB107[14] , 
        \wRegInB107[13] , \wRegInB107[12] , \wRegInB107[11] , \wRegInB107[10] , 
        \wRegInB107[9] , \wRegInB107[8] , \wRegInB107[7] , \wRegInB107[6] , 
        \wRegInB107[5] , \wRegInB107[4] , \wRegInB107[3] , \wRegInB107[2] , 
        \wRegInB107[1] , \wRegInB107[0] }), .Out({\wBIn107[31] , \wBIn107[30] , 
        \wBIn107[29] , \wBIn107[28] , \wBIn107[27] , \wBIn107[26] , 
        \wBIn107[25] , \wBIn107[24] , \wBIn107[23] , \wBIn107[22] , 
        \wBIn107[21] , \wBIn107[20] , \wBIn107[19] , \wBIn107[18] , 
        \wBIn107[17] , \wBIn107[16] , \wBIn107[15] , \wBIn107[14] , 
        \wBIn107[13] , \wBIn107[12] , \wBIn107[11] , \wBIn107[10] , 
        \wBIn107[9] , \wBIn107[8] , \wBIn107[7] , \wBIn107[6] , \wBIn107[5] , 
        \wBIn107[4] , \wBIn107[3] , \wBIn107[2] , \wBIn107[1] , \wBIn107[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn29[31] , \wAIn29[30] , \wAIn29[29] , \wAIn29[28] , \wAIn29[27] , 
        \wAIn29[26] , \wAIn29[25] , \wAIn29[24] , \wAIn29[23] , \wAIn29[22] , 
        \wAIn29[21] , \wAIn29[20] , \wAIn29[19] , \wAIn29[18] , \wAIn29[17] , 
        \wAIn29[16] , \wAIn29[15] , \wAIn29[14] , \wAIn29[13] , \wAIn29[12] , 
        \wAIn29[11] , \wAIn29[10] , \wAIn29[9] , \wAIn29[8] , \wAIn29[7] , 
        \wAIn29[6] , \wAIn29[5] , \wAIn29[4] , \wAIn29[3] , \wAIn29[2] , 
        \wAIn29[1] , \wAIn29[0] }), .BIn({\wBIn29[31] , \wBIn29[30] , 
        \wBIn29[29] , \wBIn29[28] , \wBIn29[27] , \wBIn29[26] , \wBIn29[25] , 
        \wBIn29[24] , \wBIn29[23] , \wBIn29[22] , \wBIn29[21] , \wBIn29[20] , 
        \wBIn29[19] , \wBIn29[18] , \wBIn29[17] , \wBIn29[16] , \wBIn29[15] , 
        \wBIn29[14] , \wBIn29[13] , \wBIn29[12] , \wBIn29[11] , \wBIn29[10] , 
        \wBIn29[9] , \wBIn29[8] , \wBIn29[7] , \wBIn29[6] , \wBIn29[5] , 
        \wBIn29[4] , \wBIn29[3] , \wBIn29[2] , \wBIn29[1] , \wBIn29[0] }), 
        .HiOut({\wBMid28[31] , \wBMid28[30] , \wBMid28[29] , \wBMid28[28] , 
        \wBMid28[27] , \wBMid28[26] , \wBMid28[25] , \wBMid28[24] , 
        \wBMid28[23] , \wBMid28[22] , \wBMid28[21] , \wBMid28[20] , 
        \wBMid28[19] , \wBMid28[18] , \wBMid28[17] , \wBMid28[16] , 
        \wBMid28[15] , \wBMid28[14] , \wBMid28[13] , \wBMid28[12] , 
        \wBMid28[11] , \wBMid28[10] , \wBMid28[9] , \wBMid28[8] , \wBMid28[7] , 
        \wBMid28[6] , \wBMid28[5] , \wBMid28[4] , \wBMid28[3] , \wBMid28[2] , 
        \wBMid28[1] , \wBMid28[0] }), .LoOut({\wAMid29[31] , \wAMid29[30] , 
        \wAMid29[29] , \wAMid29[28] , \wAMid29[27] , \wAMid29[26] , 
        \wAMid29[25] , \wAMid29[24] , \wAMid29[23] , \wAMid29[22] , 
        \wAMid29[21] , \wAMid29[20] , \wAMid29[19] , \wAMid29[18] , 
        \wAMid29[17] , \wAMid29[16] , \wAMid29[15] , \wAMid29[14] , 
        \wAMid29[13] , \wAMid29[12] , \wAMid29[11] , \wAMid29[10] , 
        \wAMid29[9] , \wAMid29[8] , \wAMid29[7] , \wAMid29[6] , \wAMid29[5] , 
        \wAMid29[4] , \wAMid29[3] , \wAMid29[2] , \wAMid29[1] , \wAMid29[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn32[31] , \wAIn32[30] , \wAIn32[29] , \wAIn32[28] , \wAIn32[27] , 
        \wAIn32[26] , \wAIn32[25] , \wAIn32[24] , \wAIn32[23] , \wAIn32[22] , 
        \wAIn32[21] , \wAIn32[20] , \wAIn32[19] , \wAIn32[18] , \wAIn32[17] , 
        \wAIn32[16] , \wAIn32[15] , \wAIn32[14] , \wAIn32[13] , \wAIn32[12] , 
        \wAIn32[11] , \wAIn32[10] , \wAIn32[9] , \wAIn32[8] , \wAIn32[7] , 
        \wAIn32[6] , \wAIn32[5] , \wAIn32[4] , \wAIn32[3] , \wAIn32[2] , 
        \wAIn32[1] , \wAIn32[0] }), .BIn({\wBIn32[31] , \wBIn32[30] , 
        \wBIn32[29] , \wBIn32[28] , \wBIn32[27] , \wBIn32[26] , \wBIn32[25] , 
        \wBIn32[24] , \wBIn32[23] , \wBIn32[22] , \wBIn32[21] , \wBIn32[20] , 
        \wBIn32[19] , \wBIn32[18] , \wBIn32[17] , \wBIn32[16] , \wBIn32[15] , 
        \wBIn32[14] , \wBIn32[13] , \wBIn32[12] , \wBIn32[11] , \wBIn32[10] , 
        \wBIn32[9] , \wBIn32[8] , \wBIn32[7] , \wBIn32[6] , \wBIn32[5] , 
        \wBIn32[4] , \wBIn32[3] , \wBIn32[2] , \wBIn32[1] , \wBIn32[0] }), 
        .HiOut({\wBMid31[31] , \wBMid31[30] , \wBMid31[29] , \wBMid31[28] , 
        \wBMid31[27] , \wBMid31[26] , \wBMid31[25] , \wBMid31[24] , 
        \wBMid31[23] , \wBMid31[22] , \wBMid31[21] , \wBMid31[20] , 
        \wBMid31[19] , \wBMid31[18] , \wBMid31[17] , \wBMid31[16] , 
        \wBMid31[15] , \wBMid31[14] , \wBMid31[13] , \wBMid31[12] , 
        \wBMid31[11] , \wBMid31[10] , \wBMid31[9] , \wBMid31[8] , \wBMid31[7] , 
        \wBMid31[6] , \wBMid31[5] , \wBMid31[4] , \wBMid31[3] , \wBMid31[2] , 
        \wBMid31[1] , \wBMid31[0] }), .LoOut({\wAMid32[31] , \wAMid32[30] , 
        \wAMid32[29] , \wAMid32[28] , \wAMid32[27] , \wAMid32[26] , 
        \wAMid32[25] , \wAMid32[24] , \wAMid32[23] , \wAMid32[22] , 
        \wAMid32[21] , \wAMid32[20] , \wAMid32[19] , \wAMid32[18] , 
        \wAMid32[17] , \wAMid32[16] , \wAMid32[15] , \wAMid32[14] , 
        \wAMid32[13] , \wAMid32[12] , \wAMid32[11] , \wAMid32[10] , 
        \wAMid32[9] , \wAMid32[8] , \wAMid32[7] , \wAMid32[6] , \wAMid32[5] , 
        \wAMid32[4] , \wAMid32[3] , \wAMid32[2] , \wAMid32[1] , \wAMid32[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_137 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink138[31] , \ScanLink138[30] , \ScanLink138[29] , 
        \ScanLink138[28] , \ScanLink138[27] , \ScanLink138[26] , 
        \ScanLink138[25] , \ScanLink138[24] , \ScanLink138[23] , 
        \ScanLink138[22] , \ScanLink138[21] , \ScanLink138[20] , 
        \ScanLink138[19] , \ScanLink138[18] , \ScanLink138[17] , 
        \ScanLink138[16] , \ScanLink138[15] , \ScanLink138[14] , 
        \ScanLink138[13] , \ScanLink138[12] , \ScanLink138[11] , 
        \ScanLink138[10] , \ScanLink138[9] , \ScanLink138[8] , 
        \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , \ScanLink138[4] , 
        \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , \ScanLink138[0] 
        }), .ScanOut({\ScanLink137[31] , \ScanLink137[30] , \ScanLink137[29] , 
        \ScanLink137[28] , \ScanLink137[27] , \ScanLink137[26] , 
        \ScanLink137[25] , \ScanLink137[24] , \ScanLink137[23] , 
        \ScanLink137[22] , \ScanLink137[21] , \ScanLink137[20] , 
        \ScanLink137[19] , \ScanLink137[18] , \ScanLink137[17] , 
        \ScanLink137[16] , \ScanLink137[15] , \ScanLink137[14] , 
        \ScanLink137[13] , \ScanLink137[12] , \ScanLink137[11] , 
        \ScanLink137[10] , \ScanLink137[9] , \ScanLink137[8] , 
        \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , \ScanLink137[4] , 
        \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , \ScanLink137[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA59[31] , \wRegInA59[30] , \wRegInA59[29] , 
        \wRegInA59[28] , \wRegInA59[27] , \wRegInA59[26] , \wRegInA59[25] , 
        \wRegInA59[24] , \wRegInA59[23] , \wRegInA59[22] , \wRegInA59[21] , 
        \wRegInA59[20] , \wRegInA59[19] , \wRegInA59[18] , \wRegInA59[17] , 
        \wRegInA59[16] , \wRegInA59[15] , \wRegInA59[14] , \wRegInA59[13] , 
        \wRegInA59[12] , \wRegInA59[11] , \wRegInA59[10] , \wRegInA59[9] , 
        \wRegInA59[8] , \wRegInA59[7] , \wRegInA59[6] , \wRegInA59[5] , 
        \wRegInA59[4] , \wRegInA59[3] , \wRegInA59[2] , \wRegInA59[1] , 
        \wRegInA59[0] }), .Out({\wAIn59[31] , \wAIn59[30] , \wAIn59[29] , 
        \wAIn59[28] , \wAIn59[27] , \wAIn59[26] , \wAIn59[25] , \wAIn59[24] , 
        \wAIn59[23] , \wAIn59[22] , \wAIn59[21] , \wAIn59[20] , \wAIn59[19] , 
        \wAIn59[18] , \wAIn59[17] , \wAIn59[16] , \wAIn59[15] , \wAIn59[14] , 
        \wAIn59[13] , \wAIn59[12] , \wAIn59[11] , \wAIn59[10] , \wAIn59[9] , 
        \wAIn59[8] , \wAIn59[7] , \wAIn59[6] , \wAIn59[5] , \wAIn59[4] , 
        \wAIn59[3] , \wAIn59[2] , \wAIn59[1] , \wAIn59[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_67 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink68[31] , \ScanLink68[30] , \ScanLink68[29] , 
        \ScanLink68[28] , \ScanLink68[27] , \ScanLink68[26] , \ScanLink68[25] , 
        \ScanLink68[24] , \ScanLink68[23] , \ScanLink68[22] , \ScanLink68[21] , 
        \ScanLink68[20] , \ScanLink68[19] , \ScanLink68[18] , \ScanLink68[17] , 
        \ScanLink68[16] , \ScanLink68[15] , \ScanLink68[14] , \ScanLink68[13] , 
        \ScanLink68[12] , \ScanLink68[11] , \ScanLink68[10] , \ScanLink68[9] , 
        \ScanLink68[8] , \ScanLink68[7] , \ScanLink68[6] , \ScanLink68[5] , 
        \ScanLink68[4] , \ScanLink68[3] , \ScanLink68[2] , \ScanLink68[1] , 
        \ScanLink68[0] }), .ScanOut({\ScanLink67[31] , \ScanLink67[30] , 
        \ScanLink67[29] , \ScanLink67[28] , \ScanLink67[27] , \ScanLink67[26] , 
        \ScanLink67[25] , \ScanLink67[24] , \ScanLink67[23] , \ScanLink67[22] , 
        \ScanLink67[21] , \ScanLink67[20] , \ScanLink67[19] , \ScanLink67[18] , 
        \ScanLink67[17] , \ScanLink67[16] , \ScanLink67[15] , \ScanLink67[14] , 
        \ScanLink67[13] , \ScanLink67[12] , \ScanLink67[11] , \ScanLink67[10] , 
        \ScanLink67[9] , \ScanLink67[8] , \ScanLink67[7] , \ScanLink67[6] , 
        \ScanLink67[5] , \ScanLink67[4] , \ScanLink67[3] , \ScanLink67[2] , 
        \ScanLink67[1] , \ScanLink67[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA94[31] , \wRegInA94[30] , 
        \wRegInA94[29] , \wRegInA94[28] , \wRegInA94[27] , \wRegInA94[26] , 
        \wRegInA94[25] , \wRegInA94[24] , \wRegInA94[23] , \wRegInA94[22] , 
        \wRegInA94[21] , \wRegInA94[20] , \wRegInA94[19] , \wRegInA94[18] , 
        \wRegInA94[17] , \wRegInA94[16] , \wRegInA94[15] , \wRegInA94[14] , 
        \wRegInA94[13] , \wRegInA94[12] , \wRegInA94[11] , \wRegInA94[10] , 
        \wRegInA94[9] , \wRegInA94[8] , \wRegInA94[7] , \wRegInA94[6] , 
        \wRegInA94[5] , \wRegInA94[4] , \wRegInA94[3] , \wRegInA94[2] , 
        \wRegInA94[1] , \wRegInA94[0] }), .Out({\wAIn94[31] , \wAIn94[30] , 
        \wAIn94[29] , \wAIn94[28] , \wAIn94[27] , \wAIn94[26] , \wAIn94[25] , 
        \wAIn94[24] , \wAIn94[23] , \wAIn94[22] , \wAIn94[21] , \wAIn94[20] , 
        \wAIn94[19] , \wAIn94[18] , \wAIn94[17] , \wAIn94[16] , \wAIn94[15] , 
        \wAIn94[14] , \wAIn94[13] , \wAIn94[12] , \wAIn94[11] , \wAIn94[10] , 
        \wAIn94[9] , \wAIn94[8] , \wAIn94[7] , \wAIn94[6] , \wAIn94[5] , 
        \wAIn94[4] , \wAIn94[3] , \wAIn94[2] , \wAIn94[1] , \wAIn94[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn47[31] , \wAIn47[30] , \wAIn47[29] , \wAIn47[28] , \wAIn47[27] , 
        \wAIn47[26] , \wAIn47[25] , \wAIn47[24] , \wAIn47[23] , \wAIn47[22] , 
        \wAIn47[21] , \wAIn47[20] , \wAIn47[19] , \wAIn47[18] , \wAIn47[17] , 
        \wAIn47[16] , \wAIn47[15] , \wAIn47[14] , \wAIn47[13] , \wAIn47[12] , 
        \wAIn47[11] , \wAIn47[10] , \wAIn47[9] , \wAIn47[8] , \wAIn47[7] , 
        \wAIn47[6] , \wAIn47[5] , \wAIn47[4] , \wAIn47[3] , \wAIn47[2] , 
        \wAIn47[1] , \wAIn47[0] }), .BIn({\wBIn47[31] , \wBIn47[30] , 
        \wBIn47[29] , \wBIn47[28] , \wBIn47[27] , \wBIn47[26] , \wBIn47[25] , 
        \wBIn47[24] , \wBIn47[23] , \wBIn47[22] , \wBIn47[21] , \wBIn47[20] , 
        \wBIn47[19] , \wBIn47[18] , \wBIn47[17] , \wBIn47[16] , \wBIn47[15] , 
        \wBIn47[14] , \wBIn47[13] , \wBIn47[12] , \wBIn47[11] , \wBIn47[10] , 
        \wBIn47[9] , \wBIn47[8] , \wBIn47[7] , \wBIn47[6] , \wBIn47[5] , 
        \wBIn47[4] , \wBIn47[3] , \wBIn47[2] , \wBIn47[1] , \wBIn47[0] }), 
        .HiOut({\wBMid46[31] , \wBMid46[30] , \wBMid46[29] , \wBMid46[28] , 
        \wBMid46[27] , \wBMid46[26] , \wBMid46[25] , \wBMid46[24] , 
        \wBMid46[23] , \wBMid46[22] , \wBMid46[21] , \wBMid46[20] , 
        \wBMid46[19] , \wBMid46[18] , \wBMid46[17] , \wBMid46[16] , 
        \wBMid46[15] , \wBMid46[14] , \wBMid46[13] , \wBMid46[12] , 
        \wBMid46[11] , \wBMid46[10] , \wBMid46[9] , \wBMid46[8] , \wBMid46[7] , 
        \wBMid46[6] , \wBMid46[5] , \wBMid46[4] , \wBMid46[3] , \wBMid46[2] , 
        \wBMid46[1] , \wBMid46[0] }), .LoOut({\wAMid47[31] , \wAMid47[30] , 
        \wAMid47[29] , \wAMid47[28] , \wAMid47[27] , \wAMid47[26] , 
        \wAMid47[25] , \wAMid47[24] , \wAMid47[23] , \wAMid47[22] , 
        \wAMid47[21] , \wAMid47[20] , \wAMid47[19] , \wAMid47[18] , 
        \wAMid47[17] , \wAMid47[16] , \wAMid47[15] , \wAMid47[14] , 
        \wAMid47[13] , \wAMid47[12] , \wAMid47[11] , \wAMid47[10] , 
        \wAMid47[9] , \wAMid47[8] , \wAMid47[7] , \wAMid47[6] , \wAMid47[5] , 
        \wAMid47[4] , \wAMid47[3] , \wAMid47[2] , \wAMid47[1] , \wAMid47[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn60[31] , \wAIn60[30] , \wAIn60[29] , \wAIn60[28] , \wAIn60[27] , 
        \wAIn60[26] , \wAIn60[25] , \wAIn60[24] , \wAIn60[23] , \wAIn60[22] , 
        \wAIn60[21] , \wAIn60[20] , \wAIn60[19] , \wAIn60[18] , \wAIn60[17] , 
        \wAIn60[16] , \wAIn60[15] , \wAIn60[14] , \wAIn60[13] , \wAIn60[12] , 
        \wAIn60[11] , \wAIn60[10] , \wAIn60[9] , \wAIn60[8] , \wAIn60[7] , 
        \wAIn60[6] , \wAIn60[5] , \wAIn60[4] , \wAIn60[3] , \wAIn60[2] , 
        \wAIn60[1] , \wAIn60[0] }), .BIn({\wBIn60[31] , \wBIn60[30] , 
        \wBIn60[29] , \wBIn60[28] , \wBIn60[27] , \wBIn60[26] , \wBIn60[25] , 
        \wBIn60[24] , \wBIn60[23] , \wBIn60[22] , \wBIn60[21] , \wBIn60[20] , 
        \wBIn60[19] , \wBIn60[18] , \wBIn60[17] , \wBIn60[16] , \wBIn60[15] , 
        \wBIn60[14] , \wBIn60[13] , \wBIn60[12] , \wBIn60[11] , \wBIn60[10] , 
        \wBIn60[9] , \wBIn60[8] , \wBIn60[7] , \wBIn60[6] , \wBIn60[5] , 
        \wBIn60[4] , \wBIn60[3] , \wBIn60[2] , \wBIn60[1] , \wBIn60[0] }), 
        .HiOut({\wBMid59[31] , \wBMid59[30] , \wBMid59[29] , \wBMid59[28] , 
        \wBMid59[27] , \wBMid59[26] , \wBMid59[25] , \wBMid59[24] , 
        \wBMid59[23] , \wBMid59[22] , \wBMid59[21] , \wBMid59[20] , 
        \wBMid59[19] , \wBMid59[18] , \wBMid59[17] , \wBMid59[16] , 
        \wBMid59[15] , \wBMid59[14] , \wBMid59[13] , \wBMid59[12] , 
        \wBMid59[11] , \wBMid59[10] , \wBMid59[9] , \wBMid59[8] , \wBMid59[7] , 
        \wBMid59[6] , \wBMid59[5] , \wBMid59[4] , \wBMid59[3] , \wBMid59[2] , 
        \wBMid59[1] , \wBMid59[0] }), .LoOut({\wAMid60[31] , \wAMid60[30] , 
        \wAMid60[29] , \wAMid60[28] , \wAMid60[27] , \wAMid60[26] , 
        \wAMid60[25] , \wAMid60[24] , \wAMid60[23] , \wAMid60[22] , 
        \wAMid60[21] , \wAMid60[20] , \wAMid60[19] , \wAMid60[18] , 
        \wAMid60[17] , \wAMid60[16] , \wAMid60[15] , \wAMid60[14] , 
        \wAMid60[13] , \wAMid60[12] , \wAMid60[11] , \wAMid60[10] , 
        \wAMid60[9] , \wAMid60[8] , \wAMid60[7] , \wAMid60[6] , \wAMid60[5] , 
        \wAMid60[4] , \wAMid60[3] , \wAMid60[2] , \wAMid60[1] , \wAMid60[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid101[31] , \wAMid101[30] , \wAMid101[29] , \wAMid101[28] , 
        \wAMid101[27] , \wAMid101[26] , \wAMid101[25] , \wAMid101[24] , 
        \wAMid101[23] , \wAMid101[22] , \wAMid101[21] , \wAMid101[20] , 
        \wAMid101[19] , \wAMid101[18] , \wAMid101[17] , \wAMid101[16] , 
        \wAMid101[15] , \wAMid101[14] , \wAMid101[13] , \wAMid101[12] , 
        \wAMid101[11] , \wAMid101[10] , \wAMid101[9] , \wAMid101[8] , 
        \wAMid101[7] , \wAMid101[6] , \wAMid101[5] , \wAMid101[4] , 
        \wAMid101[3] , \wAMid101[2] , \wAMid101[1] , \wAMid101[0] }), .BIn({
        \wBMid101[31] , \wBMid101[30] , \wBMid101[29] , \wBMid101[28] , 
        \wBMid101[27] , \wBMid101[26] , \wBMid101[25] , \wBMid101[24] , 
        \wBMid101[23] , \wBMid101[22] , \wBMid101[21] , \wBMid101[20] , 
        \wBMid101[19] , \wBMid101[18] , \wBMid101[17] , \wBMid101[16] , 
        \wBMid101[15] , \wBMid101[14] , \wBMid101[13] , \wBMid101[12] , 
        \wBMid101[11] , \wBMid101[10] , \wBMid101[9] , \wBMid101[8] , 
        \wBMid101[7] , \wBMid101[6] , \wBMid101[5] , \wBMid101[4] , 
        \wBMid101[3] , \wBMid101[2] , \wBMid101[1] , \wBMid101[0] }), .HiOut({
        \wRegInB101[31] , \wRegInB101[30] , \wRegInB101[29] , \wRegInB101[28] , 
        \wRegInB101[27] , \wRegInB101[26] , \wRegInB101[25] , \wRegInB101[24] , 
        \wRegInB101[23] , \wRegInB101[22] , \wRegInB101[21] , \wRegInB101[20] , 
        \wRegInB101[19] , \wRegInB101[18] , \wRegInB101[17] , \wRegInB101[16] , 
        \wRegInB101[15] , \wRegInB101[14] , \wRegInB101[13] , \wRegInB101[12] , 
        \wRegInB101[11] , \wRegInB101[10] , \wRegInB101[9] , \wRegInB101[8] , 
        \wRegInB101[7] , \wRegInB101[6] , \wRegInB101[5] , \wRegInB101[4] , 
        \wRegInB101[3] , \wRegInB101[2] , \wRegInB101[1] , \wRegInB101[0] }), 
        .LoOut({\wRegInA102[31] , \wRegInA102[30] , \wRegInA102[29] , 
        \wRegInA102[28] , \wRegInA102[27] , \wRegInA102[26] , \wRegInA102[25] , 
        \wRegInA102[24] , \wRegInA102[23] , \wRegInA102[22] , \wRegInA102[21] , 
        \wRegInA102[20] , \wRegInA102[19] , \wRegInA102[18] , \wRegInA102[17] , 
        \wRegInA102[16] , \wRegInA102[15] , \wRegInA102[14] , \wRegInA102[13] , 
        \wRegInA102[12] , \wRegInA102[11] , \wRegInA102[10] , \wRegInA102[9] , 
        \wRegInA102[8] , \wRegInA102[7] , \wRegInA102[6] , \wRegInA102[5] , 
        \wRegInA102[4] , \wRegInA102[3] , \wRegInA102[2] , \wRegInA102[1] , 
        \wRegInA102[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_207 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink208[31] , \ScanLink208[30] , \ScanLink208[29] , 
        \ScanLink208[28] , \ScanLink208[27] , \ScanLink208[26] , 
        \ScanLink208[25] , \ScanLink208[24] , \ScanLink208[23] , 
        \ScanLink208[22] , \ScanLink208[21] , \ScanLink208[20] , 
        \ScanLink208[19] , \ScanLink208[18] , \ScanLink208[17] , 
        \ScanLink208[16] , \ScanLink208[15] , \ScanLink208[14] , 
        \ScanLink208[13] , \ScanLink208[12] , \ScanLink208[11] , 
        \ScanLink208[10] , \ScanLink208[9] , \ScanLink208[8] , 
        \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , \ScanLink208[4] , 
        \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , \ScanLink208[0] 
        }), .ScanOut({\ScanLink207[31] , \ScanLink207[30] , \ScanLink207[29] , 
        \ScanLink207[28] , \ScanLink207[27] , \ScanLink207[26] , 
        \ScanLink207[25] , \ScanLink207[24] , \ScanLink207[23] , 
        \ScanLink207[22] , \ScanLink207[21] , \ScanLink207[20] , 
        \ScanLink207[19] , \ScanLink207[18] , \ScanLink207[17] , 
        \ScanLink207[16] , \ScanLink207[15] , \ScanLink207[14] , 
        \ScanLink207[13] , \ScanLink207[12] , \ScanLink207[11] , 
        \ScanLink207[10] , \ScanLink207[9] , \ScanLink207[8] , 
        \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , \ScanLink207[4] , 
        \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , \ScanLink207[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA24[31] , \wRegInA24[30] , \wRegInA24[29] , 
        \wRegInA24[28] , \wRegInA24[27] , \wRegInA24[26] , \wRegInA24[25] , 
        \wRegInA24[24] , \wRegInA24[23] , \wRegInA24[22] , \wRegInA24[21] , 
        \wRegInA24[20] , \wRegInA24[19] , \wRegInA24[18] , \wRegInA24[17] , 
        \wRegInA24[16] , \wRegInA24[15] , \wRegInA24[14] , \wRegInA24[13] , 
        \wRegInA24[12] , \wRegInA24[11] , \wRegInA24[10] , \wRegInA24[9] , 
        \wRegInA24[8] , \wRegInA24[7] , \wRegInA24[6] , \wRegInA24[5] , 
        \wRegInA24[4] , \wRegInA24[3] , \wRegInA24[2] , \wRegInA24[1] , 
        \wRegInA24[0] }), .Out({\wAIn24[31] , \wAIn24[30] , \wAIn24[29] , 
        \wAIn24[28] , \wAIn24[27] , \wAIn24[26] , \wAIn24[25] , \wAIn24[24] , 
        \wAIn24[23] , \wAIn24[22] , \wAIn24[21] , \wAIn24[20] , \wAIn24[19] , 
        \wAIn24[18] , \wAIn24[17] , \wAIn24[16] , \wAIn24[15] , \wAIn24[14] , 
        \wAIn24[13] , \wAIn24[12] , \wAIn24[11] , \wAIn24[10] , \wAIn24[9] , 
        \wAIn24[8] , \wAIn24[7] , \wAIn24[6] , \wAIn24[5] , \wAIn24[4] , 
        \wAIn24[3] , \wAIn24[2] , \wAIn24[1] , \wAIn24[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_159 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink160[31] , \ScanLink160[30] , \ScanLink160[29] , 
        \ScanLink160[28] , \ScanLink160[27] , \ScanLink160[26] , 
        \ScanLink160[25] , \ScanLink160[24] , \ScanLink160[23] , 
        \ScanLink160[22] , \ScanLink160[21] , \ScanLink160[20] , 
        \ScanLink160[19] , \ScanLink160[18] , \ScanLink160[17] , 
        \ScanLink160[16] , \ScanLink160[15] , \ScanLink160[14] , 
        \ScanLink160[13] , \ScanLink160[12] , \ScanLink160[11] , 
        \ScanLink160[10] , \ScanLink160[9] , \ScanLink160[8] , 
        \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , \ScanLink160[4] , 
        \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , \ScanLink160[0] 
        }), .ScanOut({\ScanLink159[31] , \ScanLink159[30] , \ScanLink159[29] , 
        \ScanLink159[28] , \ScanLink159[27] , \ScanLink159[26] , 
        \ScanLink159[25] , \ScanLink159[24] , \ScanLink159[23] , 
        \ScanLink159[22] , \ScanLink159[21] , \ScanLink159[20] , 
        \ScanLink159[19] , \ScanLink159[18] , \ScanLink159[17] , 
        \ScanLink159[16] , \ScanLink159[15] , \ScanLink159[14] , 
        \ScanLink159[13] , \ScanLink159[12] , \ScanLink159[11] , 
        \ScanLink159[10] , \ScanLink159[9] , \ScanLink159[8] , 
        \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , \ScanLink159[4] , 
        \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , \ScanLink159[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA48[31] , \wRegInA48[30] , \wRegInA48[29] , 
        \wRegInA48[28] , \wRegInA48[27] , \wRegInA48[26] , \wRegInA48[25] , 
        \wRegInA48[24] , \wRegInA48[23] , \wRegInA48[22] , \wRegInA48[21] , 
        \wRegInA48[20] , \wRegInA48[19] , \wRegInA48[18] , \wRegInA48[17] , 
        \wRegInA48[16] , \wRegInA48[15] , \wRegInA48[14] , \wRegInA48[13] , 
        \wRegInA48[12] , \wRegInA48[11] , \wRegInA48[10] , \wRegInA48[9] , 
        \wRegInA48[8] , \wRegInA48[7] , \wRegInA48[6] , \wRegInA48[5] , 
        \wRegInA48[4] , \wRegInA48[3] , \wRegInA48[2] , \wRegInA48[1] , 
        \wRegInA48[0] }), .Out({\wAIn48[31] , \wAIn48[30] , \wAIn48[29] , 
        \wAIn48[28] , \wAIn48[27] , \wAIn48[26] , \wAIn48[25] , \wAIn48[24] , 
        \wAIn48[23] , \wAIn48[22] , \wAIn48[21] , \wAIn48[20] , \wAIn48[19] , 
        \wAIn48[18] , \wAIn48[17] , \wAIn48[16] , \wAIn48[15] , \wAIn48[14] , 
        \wAIn48[13] , \wAIn48[12] , \wAIn48[11] , \wAIn48[10] , \wAIn48[9] , 
        \wAIn48[8] , \wAIn48[7] , \wAIn48[6] , \wAIn48[5] , \wAIn48[4] , 
        \wAIn48[3] , \wAIn48[2] , \wAIn48[1] , \wAIn48[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_3 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[31] , \ScanLink4[30] , \ScanLink4[29] , 
        \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , \ScanLink4[25] , 
        \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , \ScanLink4[21] , 
        \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , \ScanLink4[17] , 
        \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA126[31] , \wRegInA126[30] , 
        \wRegInA126[29] , \wRegInA126[28] , \wRegInA126[27] , \wRegInA126[26] , 
        \wRegInA126[25] , \wRegInA126[24] , \wRegInA126[23] , \wRegInA126[22] , 
        \wRegInA126[21] , \wRegInA126[20] , \wRegInA126[19] , \wRegInA126[18] , 
        \wRegInA126[17] , \wRegInA126[16] , \wRegInA126[15] , \wRegInA126[14] , 
        \wRegInA126[13] , \wRegInA126[12] , \wRegInA126[11] , \wRegInA126[10] , 
        \wRegInA126[9] , \wRegInA126[8] , \wRegInA126[7] , \wRegInA126[6] , 
        \wRegInA126[5] , \wRegInA126[4] , \wRegInA126[3] , \wRegInA126[2] , 
        \wRegInA126[1] , \wRegInA126[0] }), .Out({\wAIn126[31] , \wAIn126[30] , 
        \wAIn126[29] , \wAIn126[28] , \wAIn126[27] , \wAIn126[26] , 
        \wAIn126[25] , \wAIn126[24] , \wAIn126[23] , \wAIn126[22] , 
        \wAIn126[21] , \wAIn126[20] , \wAIn126[19] , \wAIn126[18] , 
        \wAIn126[17] , \wAIn126[16] , \wAIn126[15] , \wAIn126[14] , 
        \wAIn126[13] , \wAIn126[12] , \wAIn126[11] , \wAIn126[10] , 
        \wAIn126[9] , \wAIn126[8] , \wAIn126[7] , \wAIn126[6] , \wAIn126[5] , 
        \wAIn126[4] , \wAIn126[3] , \wAIn126[2] , \wAIn126[1] , \wAIn126[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid126[31] , \wAMid126[30] , \wAMid126[29] , \wAMid126[28] , 
        \wAMid126[27] , \wAMid126[26] , \wAMid126[25] , \wAMid126[24] , 
        \wAMid126[23] , \wAMid126[22] , \wAMid126[21] , \wAMid126[20] , 
        \wAMid126[19] , \wAMid126[18] , \wAMid126[17] , \wAMid126[16] , 
        \wAMid126[15] , \wAMid126[14] , \wAMid126[13] , \wAMid126[12] , 
        \wAMid126[11] , \wAMid126[10] , \wAMid126[9] , \wAMid126[8] , 
        \wAMid126[7] , \wAMid126[6] , \wAMid126[5] , \wAMid126[4] , 
        \wAMid126[3] , \wAMid126[2] , \wAMid126[1] , \wAMid126[0] }), .BIn({
        \wBMid126[31] , \wBMid126[30] , \wBMid126[29] , \wBMid126[28] , 
        \wBMid126[27] , \wBMid126[26] , \wBMid126[25] , \wBMid126[24] , 
        \wBMid126[23] , \wBMid126[22] , \wBMid126[21] , \wBMid126[20] , 
        \wBMid126[19] , \wBMid126[18] , \wBMid126[17] , \wBMid126[16] , 
        \wBMid126[15] , \wBMid126[14] , \wBMid126[13] , \wBMid126[12] , 
        \wBMid126[11] , \wBMid126[10] , \wBMid126[9] , \wBMid126[8] , 
        \wBMid126[7] , \wBMid126[6] , \wBMid126[5] , \wBMid126[4] , 
        \wBMid126[3] , \wBMid126[2] , \wBMid126[1] , \wBMid126[0] }), .HiOut({
        \wRegInB126[31] , \wRegInB126[30] , \wRegInB126[29] , \wRegInB126[28] , 
        \wRegInB126[27] , \wRegInB126[26] , \wRegInB126[25] , \wRegInB126[24] , 
        \wRegInB126[23] , \wRegInB126[22] , \wRegInB126[21] , \wRegInB126[20] , 
        \wRegInB126[19] , \wRegInB126[18] , \wRegInB126[17] , \wRegInB126[16] , 
        \wRegInB126[15] , \wRegInB126[14] , \wRegInB126[13] , \wRegInB126[12] , 
        \wRegInB126[11] , \wRegInB126[10] , \wRegInB126[9] , \wRegInB126[8] , 
        \wRegInB126[7] , \wRegInB126[6] , \wRegInB126[5] , \wRegInB126[4] , 
        \wRegInB126[3] , \wRegInB126[2] , \wRegInB126[1] , \wRegInB126[0] }), 
        .LoOut({\wRegInA127[31] , \wRegInA127[30] , \wRegInA127[29] , 
        \wRegInA127[28] , \wRegInA127[27] , \wRegInA127[26] , \wRegInA127[25] , 
        \wRegInA127[24] , \wRegInA127[23] , \wRegInA127[22] , \wRegInA127[21] , 
        \wRegInA127[20] , \wRegInA127[19] , \wRegInA127[18] , \wRegInA127[17] , 
        \wRegInA127[16] , \wRegInA127[15] , \wRegInA127[14] , \wRegInA127[13] , 
        \wRegInA127[12] , \wRegInA127[11] , \wRegInA127[10] , \wRegInA127[9] , 
        \wRegInA127[8] , \wRegInA127[7] , \wRegInA127[6] , \wRegInA127[5] , 
        \wRegInA127[4] , \wRegInA127[3] , \wRegInA127[2] , \wRegInA127[1] , 
        \wRegInA127[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_82 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink83[31] , \ScanLink83[30] , \ScanLink83[29] , 
        \ScanLink83[28] , \ScanLink83[27] , \ScanLink83[26] , \ScanLink83[25] , 
        \ScanLink83[24] , \ScanLink83[23] , \ScanLink83[22] , \ScanLink83[21] , 
        \ScanLink83[20] , \ScanLink83[19] , \ScanLink83[18] , \ScanLink83[17] , 
        \ScanLink83[16] , \ScanLink83[15] , \ScanLink83[14] , \ScanLink83[13] , 
        \ScanLink83[12] , \ScanLink83[11] , \ScanLink83[10] , \ScanLink83[9] , 
        \ScanLink83[8] , \ScanLink83[7] , \ScanLink83[6] , \ScanLink83[5] , 
        \ScanLink83[4] , \ScanLink83[3] , \ScanLink83[2] , \ScanLink83[1] , 
        \ScanLink83[0] }), .ScanOut({\ScanLink82[31] , \ScanLink82[30] , 
        \ScanLink82[29] , \ScanLink82[28] , \ScanLink82[27] , \ScanLink82[26] , 
        \ScanLink82[25] , \ScanLink82[24] , \ScanLink82[23] , \ScanLink82[22] , 
        \ScanLink82[21] , \ScanLink82[20] , \ScanLink82[19] , \ScanLink82[18] , 
        \ScanLink82[17] , \ScanLink82[16] , \ScanLink82[15] , \ScanLink82[14] , 
        \ScanLink82[13] , \ScanLink82[12] , \ScanLink82[11] , \ScanLink82[10] , 
        \ScanLink82[9] , \ScanLink82[8] , \ScanLink82[7] , \ScanLink82[6] , 
        \ScanLink82[5] , \ScanLink82[4] , \ScanLink82[3] , \ScanLink82[2] , 
        \ScanLink82[1] , \ScanLink82[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB86[31] , \wRegInB86[30] , 
        \wRegInB86[29] , \wRegInB86[28] , \wRegInB86[27] , \wRegInB86[26] , 
        \wRegInB86[25] , \wRegInB86[24] , \wRegInB86[23] , \wRegInB86[22] , 
        \wRegInB86[21] , \wRegInB86[20] , \wRegInB86[19] , \wRegInB86[18] , 
        \wRegInB86[17] , \wRegInB86[16] , \wRegInB86[15] , \wRegInB86[14] , 
        \wRegInB86[13] , \wRegInB86[12] , \wRegInB86[11] , \wRegInB86[10] , 
        \wRegInB86[9] , \wRegInB86[8] , \wRegInB86[7] , \wRegInB86[6] , 
        \wRegInB86[5] , \wRegInB86[4] , \wRegInB86[3] , \wRegInB86[2] , 
        \wRegInB86[1] , \wRegInB86[0] }), .Out({\wBIn86[31] , \wBIn86[30] , 
        \wBIn86[29] , \wBIn86[28] , \wBIn86[27] , \wBIn86[26] , \wBIn86[25] , 
        \wBIn86[24] , \wBIn86[23] , \wBIn86[22] , \wBIn86[21] , \wBIn86[20] , 
        \wBIn86[19] , \wBIn86[18] , \wBIn86[17] , \wBIn86[16] , \wBIn86[15] , 
        \wBIn86[14] , \wBIn86[13] , \wBIn86[12] , \wBIn86[11] , \wBIn86[10] , 
        \wBIn86[9] , \wBIn86[8] , \wBIn86[7] , \wBIn86[6] , \wBIn86[5] , 
        \wBIn86[4] , \wBIn86[3] , \wBIn86[2] , \wBIn86[1] , \wBIn86[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_99 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink100[31] , \ScanLink100[30] , \ScanLink100[29] , 
        \ScanLink100[28] , \ScanLink100[27] , \ScanLink100[26] , 
        \ScanLink100[25] , \ScanLink100[24] , \ScanLink100[23] , 
        \ScanLink100[22] , \ScanLink100[21] , \ScanLink100[20] , 
        \ScanLink100[19] , \ScanLink100[18] , \ScanLink100[17] , 
        \ScanLink100[16] , \ScanLink100[15] , \ScanLink100[14] , 
        \ScanLink100[13] , \ScanLink100[12] , \ScanLink100[11] , 
        \ScanLink100[10] , \ScanLink100[9] , \ScanLink100[8] , 
        \ScanLink100[7] , \ScanLink100[6] , \ScanLink100[5] , \ScanLink100[4] , 
        \ScanLink100[3] , \ScanLink100[2] , \ScanLink100[1] , \ScanLink100[0] 
        }), .ScanOut({\ScanLink99[31] , \ScanLink99[30] , \ScanLink99[29] , 
        \ScanLink99[28] , \ScanLink99[27] , \ScanLink99[26] , \ScanLink99[25] , 
        \ScanLink99[24] , \ScanLink99[23] , \ScanLink99[22] , \ScanLink99[21] , 
        \ScanLink99[20] , \ScanLink99[19] , \ScanLink99[18] , \ScanLink99[17] , 
        \ScanLink99[16] , \ScanLink99[15] , \ScanLink99[14] , \ScanLink99[13] , 
        \ScanLink99[12] , \ScanLink99[11] , \ScanLink99[10] , \ScanLink99[9] , 
        \ScanLink99[8] , \ScanLink99[7] , \ScanLink99[6] , \ScanLink99[5] , 
        \ScanLink99[4] , \ScanLink99[3] , \ScanLink99[2] , \ScanLink99[1] , 
        \ScanLink99[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(
        \wEnable[0] ), .In({\wRegInA78[31] , \wRegInA78[30] , \wRegInA78[29] , 
        \wRegInA78[28] , \wRegInA78[27] , \wRegInA78[26] , \wRegInA78[25] , 
        \wRegInA78[24] , \wRegInA78[23] , \wRegInA78[22] , \wRegInA78[21] , 
        \wRegInA78[20] , \wRegInA78[19] , \wRegInA78[18] , \wRegInA78[17] , 
        \wRegInA78[16] , \wRegInA78[15] , \wRegInA78[14] , \wRegInA78[13] , 
        \wRegInA78[12] , \wRegInA78[11] , \wRegInA78[10] , \wRegInA78[9] , 
        \wRegInA78[8] , \wRegInA78[7] , \wRegInA78[6] , \wRegInA78[5] , 
        \wRegInA78[4] , \wRegInA78[3] , \wRegInA78[2] , \wRegInA78[1] , 
        \wRegInA78[0] }), .Out({\wAIn78[31] , \wAIn78[30] , \wAIn78[29] , 
        \wAIn78[28] , \wAIn78[27] , \wAIn78[26] , \wAIn78[25] , \wAIn78[24] , 
        \wAIn78[23] , \wAIn78[22] , \wAIn78[21] , \wAIn78[20] , \wAIn78[19] , 
        \wAIn78[18] , \wAIn78[17] , \wAIn78[16] , \wAIn78[15] , \wAIn78[14] , 
        \wAIn78[13] , \wAIn78[12] , \wAIn78[11] , \wAIn78[10] , \wAIn78[9] , 
        \wAIn78[8] , \wAIn78[7] , \wAIn78[6] , \wAIn78[5] , \wAIn78[4] , 
        \wAIn78[3] , \wAIn78[2] , \wAIn78[1] , \wAIn78[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn110[31] , \wAIn110[30] , \wAIn110[29] , \wAIn110[28] , 
        \wAIn110[27] , \wAIn110[26] , \wAIn110[25] , \wAIn110[24] , 
        \wAIn110[23] , \wAIn110[22] , \wAIn110[21] , \wAIn110[20] , 
        \wAIn110[19] , \wAIn110[18] , \wAIn110[17] , \wAIn110[16] , 
        \wAIn110[15] , \wAIn110[14] , \wAIn110[13] , \wAIn110[12] , 
        \wAIn110[11] , \wAIn110[10] , \wAIn110[9] , \wAIn110[8] , \wAIn110[7] , 
        \wAIn110[6] , \wAIn110[5] , \wAIn110[4] , \wAIn110[3] , \wAIn110[2] , 
        \wAIn110[1] , \wAIn110[0] }), .BIn({\wBIn110[31] , \wBIn110[30] , 
        \wBIn110[29] , \wBIn110[28] , \wBIn110[27] , \wBIn110[26] , 
        \wBIn110[25] , \wBIn110[24] , \wBIn110[23] , \wBIn110[22] , 
        \wBIn110[21] , \wBIn110[20] , \wBIn110[19] , \wBIn110[18] , 
        \wBIn110[17] , \wBIn110[16] , \wBIn110[15] , \wBIn110[14] , 
        \wBIn110[13] , \wBIn110[12] , \wBIn110[11] , \wBIn110[10] , 
        \wBIn110[9] , \wBIn110[8] , \wBIn110[7] , \wBIn110[6] , \wBIn110[5] , 
        \wBIn110[4] , \wBIn110[3] , \wBIn110[2] , \wBIn110[1] , \wBIn110[0] }), 
        .HiOut({\wBMid109[31] , \wBMid109[30] , \wBMid109[29] , \wBMid109[28] , 
        \wBMid109[27] , \wBMid109[26] , \wBMid109[25] , \wBMid109[24] , 
        \wBMid109[23] , \wBMid109[22] , \wBMid109[21] , \wBMid109[20] , 
        \wBMid109[19] , \wBMid109[18] , \wBMid109[17] , \wBMid109[16] , 
        \wBMid109[15] , \wBMid109[14] , \wBMid109[13] , \wBMid109[12] , 
        \wBMid109[11] , \wBMid109[10] , \wBMid109[9] , \wBMid109[8] , 
        \wBMid109[7] , \wBMid109[6] , \wBMid109[5] , \wBMid109[4] , 
        \wBMid109[3] , \wBMid109[2] , \wBMid109[1] , \wBMid109[0] }), .LoOut({
        \wAMid110[31] , \wAMid110[30] , \wAMid110[29] , \wAMid110[28] , 
        \wAMid110[27] , \wAMid110[26] , \wAMid110[25] , \wAMid110[24] , 
        \wAMid110[23] , \wAMid110[22] , \wAMid110[21] , \wAMid110[20] , 
        \wAMid110[19] , \wAMid110[18] , \wAMid110[17] , \wAMid110[16] , 
        \wAMid110[15] , \wAMid110[14] , \wAMid110[13] , \wAMid110[12] , 
        \wAMid110[11] , \wAMid110[10] , \wAMid110[9] , \wAMid110[8] , 
        \wAMid110[7] , \wAMid110[6] , \wAMid110[5] , \wAMid110[4] , 
        \wAMid110[3] , \wAMid110[2] , \wAMid110[1] , \wAMid110[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid50[31] , \wAMid50[30] , \wAMid50[29] , \wAMid50[28] , 
        \wAMid50[27] , \wAMid50[26] , \wAMid50[25] , \wAMid50[24] , 
        \wAMid50[23] , \wAMid50[22] , \wAMid50[21] , \wAMid50[20] , 
        \wAMid50[19] , \wAMid50[18] , \wAMid50[17] , \wAMid50[16] , 
        \wAMid50[15] , \wAMid50[14] , \wAMid50[13] , \wAMid50[12] , 
        \wAMid50[11] , \wAMid50[10] , \wAMid50[9] , \wAMid50[8] , \wAMid50[7] , 
        \wAMid50[6] , \wAMid50[5] , \wAMid50[4] , \wAMid50[3] , \wAMid50[2] , 
        \wAMid50[1] , \wAMid50[0] }), .BIn({\wBMid50[31] , \wBMid50[30] , 
        \wBMid50[29] , \wBMid50[28] , \wBMid50[27] , \wBMid50[26] , 
        \wBMid50[25] , \wBMid50[24] , \wBMid50[23] , \wBMid50[22] , 
        \wBMid50[21] , \wBMid50[20] , \wBMid50[19] , \wBMid50[18] , 
        \wBMid50[17] , \wBMid50[16] , \wBMid50[15] , \wBMid50[14] , 
        \wBMid50[13] , \wBMid50[12] , \wBMid50[11] , \wBMid50[10] , 
        \wBMid50[9] , \wBMid50[8] , \wBMid50[7] , \wBMid50[6] , \wBMid50[5] , 
        \wBMid50[4] , \wBMid50[3] , \wBMid50[2] , \wBMid50[1] , \wBMid50[0] }), 
        .HiOut({\wRegInB50[31] , \wRegInB50[30] , \wRegInB50[29] , 
        \wRegInB50[28] , \wRegInB50[27] , \wRegInB50[26] , \wRegInB50[25] , 
        \wRegInB50[24] , \wRegInB50[23] , \wRegInB50[22] , \wRegInB50[21] , 
        \wRegInB50[20] , \wRegInB50[19] , \wRegInB50[18] , \wRegInB50[17] , 
        \wRegInB50[16] , \wRegInB50[15] , \wRegInB50[14] , \wRegInB50[13] , 
        \wRegInB50[12] , \wRegInB50[11] , \wRegInB50[10] , \wRegInB50[9] , 
        \wRegInB50[8] , \wRegInB50[7] , \wRegInB50[6] , \wRegInB50[5] , 
        \wRegInB50[4] , \wRegInB50[3] , \wRegInB50[2] , \wRegInB50[1] , 
        \wRegInB50[0] }), .LoOut({\wRegInA51[31] , \wRegInA51[30] , 
        \wRegInA51[29] , \wRegInA51[28] , \wRegInA51[27] , \wRegInA51[26] , 
        \wRegInA51[25] , \wRegInA51[24] , \wRegInA51[23] , \wRegInA51[22] , 
        \wRegInA51[21] , \wRegInA51[20] , \wRegInA51[19] , \wRegInA51[18] , 
        \wRegInA51[17] , \wRegInA51[16] , \wRegInA51[15] , \wRegInA51[14] , 
        \wRegInA51[13] , \wRegInA51[12] , \wRegInA51[11] , \wRegInA51[10] , 
        \wRegInA51[9] , \wRegInA51[8] , \wRegInA51[7] , \wRegInA51[6] , 
        \wRegInA51[5] , \wRegInA51[4] , \wRegInA51[3] , \wRegInA51[2] , 
        \wRegInA51[1] , \wRegInA51[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_165 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink166[31] , \ScanLink166[30] , \ScanLink166[29] , 
        \ScanLink166[28] , \ScanLink166[27] , \ScanLink166[26] , 
        \ScanLink166[25] , \ScanLink166[24] , \ScanLink166[23] , 
        \ScanLink166[22] , \ScanLink166[21] , \ScanLink166[20] , 
        \ScanLink166[19] , \ScanLink166[18] , \ScanLink166[17] , 
        \ScanLink166[16] , \ScanLink166[15] , \ScanLink166[14] , 
        \ScanLink166[13] , \ScanLink166[12] , \ScanLink166[11] , 
        \ScanLink166[10] , \ScanLink166[9] , \ScanLink166[8] , 
        \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , \ScanLink166[4] , 
        \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , \ScanLink166[0] 
        }), .ScanOut({\ScanLink165[31] , \ScanLink165[30] , \ScanLink165[29] , 
        \ScanLink165[28] , \ScanLink165[27] , \ScanLink165[26] , 
        \ScanLink165[25] , \ScanLink165[24] , \ScanLink165[23] , 
        \ScanLink165[22] , \ScanLink165[21] , \ScanLink165[20] , 
        \ScanLink165[19] , \ScanLink165[18] , \ScanLink165[17] , 
        \ScanLink165[16] , \ScanLink165[15] , \ScanLink165[14] , 
        \ScanLink165[13] , \ScanLink165[12] , \ScanLink165[11] , 
        \ScanLink165[10] , \ScanLink165[9] , \ScanLink165[8] , 
        \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , \ScanLink165[4] , 
        \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , \ScanLink165[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA45[31] , \wRegInA45[30] , \wRegInA45[29] , 
        \wRegInA45[28] , \wRegInA45[27] , \wRegInA45[26] , \wRegInA45[25] , 
        \wRegInA45[24] , \wRegInA45[23] , \wRegInA45[22] , \wRegInA45[21] , 
        \wRegInA45[20] , \wRegInA45[19] , \wRegInA45[18] , \wRegInA45[17] , 
        \wRegInA45[16] , \wRegInA45[15] , \wRegInA45[14] , \wRegInA45[13] , 
        \wRegInA45[12] , \wRegInA45[11] , \wRegInA45[10] , \wRegInA45[9] , 
        \wRegInA45[8] , \wRegInA45[7] , \wRegInA45[6] , \wRegInA45[5] , 
        \wRegInA45[4] , \wRegInA45[3] , \wRegInA45[2] , \wRegInA45[1] , 
        \wRegInA45[0] }), .Out({\wAIn45[31] , \wAIn45[30] , \wAIn45[29] , 
        \wAIn45[28] , \wAIn45[27] , \wAIn45[26] , \wAIn45[25] , \wAIn45[24] , 
        \wAIn45[23] , \wAIn45[22] , \wAIn45[21] , \wAIn45[20] , \wAIn45[19] , 
        \wAIn45[18] , \wAIn45[17] , \wAIn45[16] , \wAIn45[15] , \wAIn45[14] , 
        \wAIn45[13] , \wAIn45[12] , \wAIn45[11] , \wAIn45[10] , \wAIn45[9] , 
        \wAIn45[8] , \wAIn45[7] , \wAIn45[6] , \wAIn45[5] , \wAIn45[4] , 
        \wAIn45[3] , \wAIn45[2] , \wAIn45[1] , \wAIn45[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_35 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink36[31] , \ScanLink36[30] , \ScanLink36[29] , 
        \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , \ScanLink36[25] , 
        \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , \ScanLink36[21] , 
        \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , \ScanLink36[17] , 
        \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , \ScanLink36[13] , 
        \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , \ScanLink36[9] , 
        \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , \ScanLink36[5] , 
        \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , \ScanLink36[1] , 
        \ScanLink36[0] }), .ScanOut({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA110[31] , \wRegInA110[30] , 
        \wRegInA110[29] , \wRegInA110[28] , \wRegInA110[27] , \wRegInA110[26] , 
        \wRegInA110[25] , \wRegInA110[24] , \wRegInA110[23] , \wRegInA110[22] , 
        \wRegInA110[21] , \wRegInA110[20] , \wRegInA110[19] , \wRegInA110[18] , 
        \wRegInA110[17] , \wRegInA110[16] , \wRegInA110[15] , \wRegInA110[14] , 
        \wRegInA110[13] , \wRegInA110[12] , \wRegInA110[11] , \wRegInA110[10] , 
        \wRegInA110[9] , \wRegInA110[8] , \wRegInA110[7] , \wRegInA110[6] , 
        \wRegInA110[5] , \wRegInA110[4] , \wRegInA110[3] , \wRegInA110[2] , 
        \wRegInA110[1] , \wRegInA110[0] }), .Out({\wAIn110[31] , \wAIn110[30] , 
        \wAIn110[29] , \wAIn110[28] , \wAIn110[27] , \wAIn110[26] , 
        \wAIn110[25] , \wAIn110[24] , \wAIn110[23] , \wAIn110[22] , 
        \wAIn110[21] , \wAIn110[20] , \wAIn110[19] , \wAIn110[18] , 
        \wAIn110[17] , \wAIn110[16] , \wAIn110[15] , \wAIn110[14] , 
        \wAIn110[13] , \wAIn110[12] , \wAIn110[11] , \wAIn110[10] , 
        \wAIn110[9] , \wAIn110[8] , \wAIn110[7] , \wAIn110[6] , \wAIn110[5] , 
        \wAIn110[4] , \wAIn110[3] , \wAIn110[2] , \wAIn110[1] , \wAIn110[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_255 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink256[31] , \ScanLink256[30] , \ScanLink256[29] , 
        \ScanLink256[28] , \ScanLink256[27] , \ScanLink256[26] , 
        \ScanLink256[25] , \ScanLink256[24] , \ScanLink256[23] , 
        \ScanLink256[22] , \ScanLink256[21] , \ScanLink256[20] , 
        \ScanLink256[19] , \ScanLink256[18] , \ScanLink256[17] , 
        \ScanLink256[16] , \ScanLink256[15] , \ScanLink256[14] , 
        \ScanLink256[13] , \ScanLink256[12] , \ScanLink256[11] , 
        \ScanLink256[10] , \ScanLink256[9] , \ScanLink256[8] , 
        \ScanLink256[7] , \ScanLink256[6] , \ScanLink256[5] , \ScanLink256[4] , 
        \ScanLink256[3] , \ScanLink256[2] , \ScanLink256[1] , \ScanLink256[0] 
        }), .ScanOut({\ScanLink255[31] , \ScanLink255[30] , \ScanLink255[29] , 
        \ScanLink255[28] , \ScanLink255[27] , \ScanLink255[26] , 
        \ScanLink255[25] , \ScanLink255[24] , \ScanLink255[23] , 
        \ScanLink255[22] , \ScanLink255[21] , \ScanLink255[20] , 
        \ScanLink255[19] , \ScanLink255[18] , \ScanLink255[17] , 
        \ScanLink255[16] , \ScanLink255[15] , \ScanLink255[14] , 
        \ScanLink255[13] , \ScanLink255[12] , \ScanLink255[11] , 
        \ScanLink255[10] , \ScanLink255[9] , \ScanLink255[8] , 
        \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , \ScanLink255[4] , 
        \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , \ScanLink255[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA0[31] , \wRegInA0[30] , \wRegInA0[29] , \wRegInA0[28] , 
        \wRegInA0[27] , \wRegInA0[26] , \wRegInA0[25] , \wRegInA0[24] , 
        \wRegInA0[23] , \wRegInA0[22] , \wRegInA0[21] , \wRegInA0[20] , 
        \wRegInA0[19] , \wRegInA0[18] , \wRegInA0[17] , \wRegInA0[16] , 
        \wRegInA0[15] , \wRegInA0[14] , \wRegInA0[13] , \wRegInA0[12] , 
        \wRegInA0[11] , \wRegInA0[10] , \wRegInA0[9] , \wRegInA0[8] , 
        \wRegInA0[7] , \wRegInA0[6] , \wRegInA0[5] , \wRegInA0[4] , 
        \wRegInA0[3] , \wRegInA0[2] , \wRegInA0[1] , \wRegInA0[0] }), .Out({
        \wAIn0[31] , \wAIn0[30] , \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , 
        \wAIn0[26] , \wAIn0[25] , \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , 
        \wAIn0[21] , \wAIn0[20] , \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , 
        \wAIn0[16] , \wAIn0[15] , \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , 
        \wAIn0[11] , \wAIn0[10] , \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , 
        \wAIn0[6] , \wAIn0[5] , \wAIn0[4] , \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , 
        \wAIn0[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid77[31] , \wAMid77[30] , \wAMid77[29] , \wAMid77[28] , 
        \wAMid77[27] , \wAMid77[26] , \wAMid77[25] , \wAMid77[24] , 
        \wAMid77[23] , \wAMid77[22] , \wAMid77[21] , \wAMid77[20] , 
        \wAMid77[19] , \wAMid77[18] , \wAMid77[17] , \wAMid77[16] , 
        \wAMid77[15] , \wAMid77[14] , \wAMid77[13] , \wAMid77[12] , 
        \wAMid77[11] , \wAMid77[10] , \wAMid77[9] , \wAMid77[8] , \wAMid77[7] , 
        \wAMid77[6] , \wAMid77[5] , \wAMid77[4] , \wAMid77[3] , \wAMid77[2] , 
        \wAMid77[1] , \wAMid77[0] }), .BIn({\wBMid77[31] , \wBMid77[30] , 
        \wBMid77[29] , \wBMid77[28] , \wBMid77[27] , \wBMid77[26] , 
        \wBMid77[25] , \wBMid77[24] , \wBMid77[23] , \wBMid77[22] , 
        \wBMid77[21] , \wBMid77[20] , \wBMid77[19] , \wBMid77[18] , 
        \wBMid77[17] , \wBMid77[16] , \wBMid77[15] , \wBMid77[14] , 
        \wBMid77[13] , \wBMid77[12] , \wBMid77[11] , \wBMid77[10] , 
        \wBMid77[9] , \wBMid77[8] , \wBMid77[7] , \wBMid77[6] , \wBMid77[5] , 
        \wBMid77[4] , \wBMid77[3] , \wBMid77[2] , \wBMid77[1] , \wBMid77[0] }), 
        .HiOut({\wRegInB77[31] , \wRegInB77[30] , \wRegInB77[29] , 
        \wRegInB77[28] , \wRegInB77[27] , \wRegInB77[26] , \wRegInB77[25] , 
        \wRegInB77[24] , \wRegInB77[23] , \wRegInB77[22] , \wRegInB77[21] , 
        \wRegInB77[20] , \wRegInB77[19] , \wRegInB77[18] , \wRegInB77[17] , 
        \wRegInB77[16] , \wRegInB77[15] , \wRegInB77[14] , \wRegInB77[13] , 
        \wRegInB77[12] , \wRegInB77[11] , \wRegInB77[10] , \wRegInB77[9] , 
        \wRegInB77[8] , \wRegInB77[7] , \wRegInB77[6] , \wRegInB77[5] , 
        \wRegInB77[4] , \wRegInB77[3] , \wRegInB77[2] , \wRegInB77[1] , 
        \wRegInB77[0] }), .LoOut({\wRegInA78[31] , \wRegInA78[30] , 
        \wRegInA78[29] , \wRegInA78[28] , \wRegInA78[27] , \wRegInA78[26] , 
        \wRegInA78[25] , \wRegInA78[24] , \wRegInA78[23] , \wRegInA78[22] , 
        \wRegInA78[21] , \wRegInA78[20] , \wRegInA78[19] , \wRegInA78[18] , 
        \wRegInA78[17] , \wRegInA78[16] , \wRegInA78[15] , \wRegInA78[14] , 
        \wRegInA78[13] , \wRegInA78[12] , \wRegInA78[11] , \wRegInA78[10] , 
        \wRegInA78[9] , \wRegInA78[8] , \wRegInA78[7] , \wRegInA78[6] , 
        \wRegInA78[5] , \wRegInA78[4] , \wRegInA78[3] , \wRegInA78[2] , 
        \wRegInA78[1] , \wRegInA78[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_12 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[31] , \ScanLink13[30] , \ScanLink13[29] , 
        \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , \ScanLink13[25] , 
        \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , \ScanLink13[21] , 
        \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , \ScanLink13[17] , 
        \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , \ScanLink13[13] , 
        \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , \ScanLink13[9] , 
        \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB121[31] , \wRegInB121[30] , 
        \wRegInB121[29] , \wRegInB121[28] , \wRegInB121[27] , \wRegInB121[26] , 
        \wRegInB121[25] , \wRegInB121[24] , \wRegInB121[23] , \wRegInB121[22] , 
        \wRegInB121[21] , \wRegInB121[20] , \wRegInB121[19] , \wRegInB121[18] , 
        \wRegInB121[17] , \wRegInB121[16] , \wRegInB121[15] , \wRegInB121[14] , 
        \wRegInB121[13] , \wRegInB121[12] , \wRegInB121[11] , \wRegInB121[10] , 
        \wRegInB121[9] , \wRegInB121[8] , \wRegInB121[7] , \wRegInB121[6] , 
        \wRegInB121[5] , \wRegInB121[4] , \wRegInB121[3] , \wRegInB121[2] , 
        \wRegInB121[1] , \wRegInB121[0] }), .Out({\wBIn121[31] , \wBIn121[30] , 
        \wBIn121[29] , \wBIn121[28] , \wBIn121[27] , \wBIn121[26] , 
        \wBIn121[25] , \wBIn121[24] , \wBIn121[23] , \wBIn121[22] , 
        \wBIn121[21] , \wBIn121[20] , \wBIn121[19] , \wBIn121[18] , 
        \wBIn121[17] , \wBIn121[16] , \wBIn121[15] , \wBIn121[14] , 
        \wBIn121[13] , \wBIn121[12] , \wBIn121[11] , \wBIn121[10] , 
        \wBIn121[9] , \wBIn121[8] , \wBIn121[7] , \wBIn121[6] , \wBIn121[5] , 
        \wBIn121[4] , \wBIn121[3] , \wBIn121[2] , \wBIn121[1] , \wBIn121[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_142 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink143[31] , \ScanLink143[30] , \ScanLink143[29] , 
        \ScanLink143[28] , \ScanLink143[27] , \ScanLink143[26] , 
        \ScanLink143[25] , \ScanLink143[24] , \ScanLink143[23] , 
        \ScanLink143[22] , \ScanLink143[21] , \ScanLink143[20] , 
        \ScanLink143[19] , \ScanLink143[18] , \ScanLink143[17] , 
        \ScanLink143[16] , \ScanLink143[15] , \ScanLink143[14] , 
        \ScanLink143[13] , \ScanLink143[12] , \ScanLink143[11] , 
        \ScanLink143[10] , \ScanLink143[9] , \ScanLink143[8] , 
        \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , \ScanLink143[4] , 
        \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , \ScanLink143[0] 
        }), .ScanOut({\ScanLink142[31] , \ScanLink142[30] , \ScanLink142[29] , 
        \ScanLink142[28] , \ScanLink142[27] , \ScanLink142[26] , 
        \ScanLink142[25] , \ScanLink142[24] , \ScanLink142[23] , 
        \ScanLink142[22] , \ScanLink142[21] , \ScanLink142[20] , 
        \ScanLink142[19] , \ScanLink142[18] , \ScanLink142[17] , 
        \ScanLink142[16] , \ScanLink142[15] , \ScanLink142[14] , 
        \ScanLink142[13] , \ScanLink142[12] , \ScanLink142[11] , 
        \ScanLink142[10] , \ScanLink142[9] , \ScanLink142[8] , 
        \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , \ScanLink142[4] , 
        \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , \ScanLink142[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB56[31] , \wRegInB56[30] , \wRegInB56[29] , 
        \wRegInB56[28] , \wRegInB56[27] , \wRegInB56[26] , \wRegInB56[25] , 
        \wRegInB56[24] , \wRegInB56[23] , \wRegInB56[22] , \wRegInB56[21] , 
        \wRegInB56[20] , \wRegInB56[19] , \wRegInB56[18] , \wRegInB56[17] , 
        \wRegInB56[16] , \wRegInB56[15] , \wRegInB56[14] , \wRegInB56[13] , 
        \wRegInB56[12] , \wRegInB56[11] , \wRegInB56[10] , \wRegInB56[9] , 
        \wRegInB56[8] , \wRegInB56[7] , \wRegInB56[6] , \wRegInB56[5] , 
        \wRegInB56[4] , \wRegInB56[3] , \wRegInB56[2] , \wRegInB56[1] , 
        \wRegInB56[0] }), .Out({\wBIn56[31] , \wBIn56[30] , \wBIn56[29] , 
        \wBIn56[28] , \wBIn56[27] , \wBIn56[26] , \wBIn56[25] , \wBIn56[24] , 
        \wBIn56[23] , \wBIn56[22] , \wBIn56[21] , \wBIn56[20] , \wBIn56[19] , 
        \wBIn56[18] , \wBIn56[17] , \wBIn56[16] , \wBIn56[15] , \wBIn56[14] , 
        \wBIn56[13] , \wBIn56[12] , \wBIn56[11] , \wBIn56[10] , \wBIn56[9] , 
        \wBIn56[8] , \wBIn56[7] , \wBIn56[6] , \wBIn56[5] , \wBIn56[4] , 
        \wBIn56[3] , \wBIn56[2] , \wBIn56[1] , \wBIn56[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid19[31] , \wAMid19[30] , \wAMid19[29] , \wAMid19[28] , 
        \wAMid19[27] , \wAMid19[26] , \wAMid19[25] , \wAMid19[24] , 
        \wAMid19[23] , \wAMid19[22] , \wAMid19[21] , \wAMid19[20] , 
        \wAMid19[19] , \wAMid19[18] , \wAMid19[17] , \wAMid19[16] , 
        \wAMid19[15] , \wAMid19[14] , \wAMid19[13] , \wAMid19[12] , 
        \wAMid19[11] , \wAMid19[10] , \wAMid19[9] , \wAMid19[8] , \wAMid19[7] , 
        \wAMid19[6] , \wAMid19[5] , \wAMid19[4] , \wAMid19[3] , \wAMid19[2] , 
        \wAMid19[1] , \wAMid19[0] }), .BIn({\wBMid19[31] , \wBMid19[30] , 
        \wBMid19[29] , \wBMid19[28] , \wBMid19[27] , \wBMid19[26] , 
        \wBMid19[25] , \wBMid19[24] , \wBMid19[23] , \wBMid19[22] , 
        \wBMid19[21] , \wBMid19[20] , \wBMid19[19] , \wBMid19[18] , 
        \wBMid19[17] , \wBMid19[16] , \wBMid19[15] , \wBMid19[14] , 
        \wBMid19[13] , \wBMid19[12] , \wBMid19[11] , \wBMid19[10] , 
        \wBMid19[9] , \wBMid19[8] , \wBMid19[7] , \wBMid19[6] , \wBMid19[5] , 
        \wBMid19[4] , \wBMid19[3] , \wBMid19[2] , \wBMid19[1] , \wBMid19[0] }), 
        .HiOut({\wRegInB19[31] , \wRegInB19[30] , \wRegInB19[29] , 
        \wRegInB19[28] , \wRegInB19[27] , \wRegInB19[26] , \wRegInB19[25] , 
        \wRegInB19[24] , \wRegInB19[23] , \wRegInB19[22] , \wRegInB19[21] , 
        \wRegInB19[20] , \wRegInB19[19] , \wRegInB19[18] , \wRegInB19[17] , 
        \wRegInB19[16] , \wRegInB19[15] , \wRegInB19[14] , \wRegInB19[13] , 
        \wRegInB19[12] , \wRegInB19[11] , \wRegInB19[10] , \wRegInB19[9] , 
        \wRegInB19[8] , \wRegInB19[7] , \wRegInB19[6] , \wRegInB19[5] , 
        \wRegInB19[4] , \wRegInB19[3] , \wRegInB19[2] , \wRegInB19[1] , 
        \wRegInB19[0] }), .LoOut({\wRegInA20[31] , \wRegInA20[30] , 
        \wRegInA20[29] , \wRegInA20[28] , \wRegInA20[27] , \wRegInA20[26] , 
        \wRegInA20[25] , \wRegInA20[24] , \wRegInA20[23] , \wRegInA20[22] , 
        \wRegInA20[21] , \wRegInA20[20] , \wRegInA20[19] , \wRegInA20[18] , 
        \wRegInA20[17] , \wRegInA20[16] , \wRegInA20[15] , \wRegInA20[14] , 
        \wRegInA20[13] , \wRegInA20[12] , \wRegInA20[11] , \wRegInA20[10] , 
        \wRegInA20[9] , \wRegInA20[8] , \wRegInA20[7] , \wRegInA20[6] , 
        \wRegInA20[5] , \wRegInA20[4] , \wRegInA20[3] , \wRegInA20[2] , 
        \wRegInA20[1] , \wRegInA20[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid92[31] , \wAMid92[30] , \wAMid92[29] , \wAMid92[28] , 
        \wAMid92[27] , \wAMid92[26] , \wAMid92[25] , \wAMid92[24] , 
        \wAMid92[23] , \wAMid92[22] , \wAMid92[21] , \wAMid92[20] , 
        \wAMid92[19] , \wAMid92[18] , \wAMid92[17] , \wAMid92[16] , 
        \wAMid92[15] , \wAMid92[14] , \wAMid92[13] , \wAMid92[12] , 
        \wAMid92[11] , \wAMid92[10] , \wAMid92[9] , \wAMid92[8] , \wAMid92[7] , 
        \wAMid92[6] , \wAMid92[5] , \wAMid92[4] , \wAMid92[3] , \wAMid92[2] , 
        \wAMid92[1] , \wAMid92[0] }), .BIn({\wBMid92[31] , \wBMid92[30] , 
        \wBMid92[29] , \wBMid92[28] , \wBMid92[27] , \wBMid92[26] , 
        \wBMid92[25] , \wBMid92[24] , \wBMid92[23] , \wBMid92[22] , 
        \wBMid92[21] , \wBMid92[20] , \wBMid92[19] , \wBMid92[18] , 
        \wBMid92[17] , \wBMid92[16] , \wBMid92[15] , \wBMid92[14] , 
        \wBMid92[13] , \wBMid92[12] , \wBMid92[11] , \wBMid92[10] , 
        \wBMid92[9] , \wBMid92[8] , \wBMid92[7] , \wBMid92[6] , \wBMid92[5] , 
        \wBMid92[4] , \wBMid92[3] , \wBMid92[2] , \wBMid92[1] , \wBMid92[0] }), 
        .HiOut({\wRegInB92[31] , \wRegInB92[30] , \wRegInB92[29] , 
        \wRegInB92[28] , \wRegInB92[27] , \wRegInB92[26] , \wRegInB92[25] , 
        \wRegInB92[24] , \wRegInB92[23] , \wRegInB92[22] , \wRegInB92[21] , 
        \wRegInB92[20] , \wRegInB92[19] , \wRegInB92[18] , \wRegInB92[17] , 
        \wRegInB92[16] , \wRegInB92[15] , \wRegInB92[14] , \wRegInB92[13] , 
        \wRegInB92[12] , \wRegInB92[11] , \wRegInB92[10] , \wRegInB92[9] , 
        \wRegInB92[8] , \wRegInB92[7] , \wRegInB92[6] , \wRegInB92[5] , 
        \wRegInB92[4] , \wRegInB92[3] , \wRegInB92[2] , \wRegInB92[1] , 
        \wRegInB92[0] }), .LoOut({\wRegInA93[31] , \wRegInA93[30] , 
        \wRegInA93[29] , \wRegInA93[28] , \wRegInA93[27] , \wRegInA93[26] , 
        \wRegInA93[25] , \wRegInA93[24] , \wRegInA93[23] , \wRegInA93[22] , 
        \wRegInA93[21] , \wRegInA93[20] , \wRegInA93[19] , \wRegInA93[18] , 
        \wRegInA93[17] , \wRegInA93[16] , \wRegInA93[15] , \wRegInA93[14] , 
        \wRegInA93[13] , \wRegInA93[12] , \wRegInA93[11] , \wRegInA93[10] , 
        \wRegInA93[9] , \wRegInA93[8] , \wRegInA93[7] , \wRegInA93[6] , 
        \wRegInA93[5] , \wRegInA93[4] , \wRegInA93[3] , \wRegInA93[2] , 
        \wRegInA93[1] , \wRegInA93[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn21[31] , \wAIn21[30] , \wAIn21[29] , \wAIn21[28] , \wAIn21[27] , 
        \wAIn21[26] , \wAIn21[25] , \wAIn21[24] , \wAIn21[23] , \wAIn21[22] , 
        \wAIn21[21] , \wAIn21[20] , \wAIn21[19] , \wAIn21[18] , \wAIn21[17] , 
        \wAIn21[16] , \wAIn21[15] , \wAIn21[14] , \wAIn21[13] , \wAIn21[12] , 
        \wAIn21[11] , \wAIn21[10] , \wAIn21[9] , \wAIn21[8] , \wAIn21[7] , 
        \wAIn21[6] , \wAIn21[5] , \wAIn21[4] , \wAIn21[3] , \wAIn21[2] , 
        \wAIn21[1] , \wAIn21[0] }), .BIn({\wBIn21[31] , \wBIn21[30] , 
        \wBIn21[29] , \wBIn21[28] , \wBIn21[27] , \wBIn21[26] , \wBIn21[25] , 
        \wBIn21[24] , \wBIn21[23] , \wBIn21[22] , \wBIn21[21] , \wBIn21[20] , 
        \wBIn21[19] , \wBIn21[18] , \wBIn21[17] , \wBIn21[16] , \wBIn21[15] , 
        \wBIn21[14] , \wBIn21[13] , \wBIn21[12] , \wBIn21[11] , \wBIn21[10] , 
        \wBIn21[9] , \wBIn21[8] , \wBIn21[7] , \wBIn21[6] , \wBIn21[5] , 
        \wBIn21[4] , \wBIn21[3] , \wBIn21[2] , \wBIn21[1] , \wBIn21[0] }), 
        .HiOut({\wBMid20[31] , \wBMid20[30] , \wBMid20[29] , \wBMid20[28] , 
        \wBMid20[27] , \wBMid20[26] , \wBMid20[25] , \wBMid20[24] , 
        \wBMid20[23] , \wBMid20[22] , \wBMid20[21] , \wBMid20[20] , 
        \wBMid20[19] , \wBMid20[18] , \wBMid20[17] , \wBMid20[16] , 
        \wBMid20[15] , \wBMid20[14] , \wBMid20[13] , \wBMid20[12] , 
        \wBMid20[11] , \wBMid20[10] , \wBMid20[9] , \wBMid20[8] , \wBMid20[7] , 
        \wBMid20[6] , \wBMid20[5] , \wBMid20[4] , \wBMid20[3] , \wBMid20[2] , 
        \wBMid20[1] , \wBMid20[0] }), .LoOut({\wAMid21[31] , \wAMid21[30] , 
        \wAMid21[29] , \wAMid21[28] , \wAMid21[27] , \wAMid21[26] , 
        \wAMid21[25] , \wAMid21[24] , \wAMid21[23] , \wAMid21[22] , 
        \wAMid21[21] , \wAMid21[20] , \wAMid21[19] , \wAMid21[18] , 
        \wAMid21[17] , \wAMid21[16] , \wAMid21[15] , \wAMid21[14] , 
        \wAMid21[13] , \wAMid21[12] , \wAMid21[11] , \wAMid21[10] , 
        \wAMid21[9] , \wAMid21[8] , \wAMid21[7] , \wAMid21[6] , \wAMid21[5] , 
        \wAMid21[4] , \wAMid21[3] , \wAMid21[2] , \wAMid21[1] , \wAMid21[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn85[31] , \wAIn85[30] , \wAIn85[29] , \wAIn85[28] , \wAIn85[27] , 
        \wAIn85[26] , \wAIn85[25] , \wAIn85[24] , \wAIn85[23] , \wAIn85[22] , 
        \wAIn85[21] , \wAIn85[20] , \wAIn85[19] , \wAIn85[18] , \wAIn85[17] , 
        \wAIn85[16] , \wAIn85[15] , \wAIn85[14] , \wAIn85[13] , \wAIn85[12] , 
        \wAIn85[11] , \wAIn85[10] , \wAIn85[9] , \wAIn85[8] , \wAIn85[7] , 
        \wAIn85[6] , \wAIn85[5] , \wAIn85[4] , \wAIn85[3] , \wAIn85[2] , 
        \wAIn85[1] , \wAIn85[0] }), .BIn({\wBIn85[31] , \wBIn85[30] , 
        \wBIn85[29] , \wBIn85[28] , \wBIn85[27] , \wBIn85[26] , \wBIn85[25] , 
        \wBIn85[24] , \wBIn85[23] , \wBIn85[22] , \wBIn85[21] , \wBIn85[20] , 
        \wBIn85[19] , \wBIn85[18] , \wBIn85[17] , \wBIn85[16] , \wBIn85[15] , 
        \wBIn85[14] , \wBIn85[13] , \wBIn85[12] , \wBIn85[11] , \wBIn85[10] , 
        \wBIn85[9] , \wBIn85[8] , \wBIn85[7] , \wBIn85[6] , \wBIn85[5] , 
        \wBIn85[4] , \wBIn85[3] , \wBIn85[2] , \wBIn85[1] , \wBIn85[0] }), 
        .HiOut({\wBMid84[31] , \wBMid84[30] , \wBMid84[29] , \wBMid84[28] , 
        \wBMid84[27] , \wBMid84[26] , \wBMid84[25] , \wBMid84[24] , 
        \wBMid84[23] , \wBMid84[22] , \wBMid84[21] , \wBMid84[20] , 
        \wBMid84[19] , \wBMid84[18] , \wBMid84[17] , \wBMid84[16] , 
        \wBMid84[15] , \wBMid84[14] , \wBMid84[13] , \wBMid84[12] , 
        \wBMid84[11] , \wBMid84[10] , \wBMid84[9] , \wBMid84[8] , \wBMid84[7] , 
        \wBMid84[6] , \wBMid84[5] , \wBMid84[4] , \wBMid84[3] , \wBMid84[2] , 
        \wBMid84[1] , \wBMid84[0] }), .LoOut({\wAMid85[31] , \wAMid85[30] , 
        \wAMid85[29] , \wAMid85[28] , \wAMid85[27] , \wAMid85[26] , 
        \wAMid85[25] , \wAMid85[24] , \wAMid85[23] , \wAMid85[22] , 
        \wAMid85[21] , \wAMid85[20] , \wAMid85[19] , \wAMid85[18] , 
        \wAMid85[17] , \wAMid85[16] , \wAMid85[15] , \wAMid85[14] , 
        \wAMid85[13] , \wAMid85[12] , \wAMid85[11] , \wAMid85[10] , 
        \wAMid85[9] , \wAMid85[8] , \wAMid85[7] , \wAMid85[6] , \wAMid85[5] , 
        \wAMid85[4] , \wAMid85[3] , \wAMid85[2] , \wAMid85[1] , \wAMid85[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_180 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink181[31] , \ScanLink181[30] , \ScanLink181[29] , 
        \ScanLink181[28] , \ScanLink181[27] , \ScanLink181[26] , 
        \ScanLink181[25] , \ScanLink181[24] , \ScanLink181[23] , 
        \ScanLink181[22] , \ScanLink181[21] , \ScanLink181[20] , 
        \ScanLink181[19] , \ScanLink181[18] , \ScanLink181[17] , 
        \ScanLink181[16] , \ScanLink181[15] , \ScanLink181[14] , 
        \ScanLink181[13] , \ScanLink181[12] , \ScanLink181[11] , 
        \ScanLink181[10] , \ScanLink181[9] , \ScanLink181[8] , 
        \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , \ScanLink181[4] , 
        \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , \ScanLink181[0] 
        }), .ScanOut({\ScanLink180[31] , \ScanLink180[30] , \ScanLink180[29] , 
        \ScanLink180[28] , \ScanLink180[27] , \ScanLink180[26] , 
        \ScanLink180[25] , \ScanLink180[24] , \ScanLink180[23] , 
        \ScanLink180[22] , \ScanLink180[21] , \ScanLink180[20] , 
        \ScanLink180[19] , \ScanLink180[18] , \ScanLink180[17] , 
        \ScanLink180[16] , \ScanLink180[15] , \ScanLink180[14] , 
        \ScanLink180[13] , \ScanLink180[12] , \ScanLink180[11] , 
        \ScanLink180[10] , \ScanLink180[9] , \ScanLink180[8] , 
        \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , \ScanLink180[4] , 
        \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , \ScanLink180[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB37[31] , \wRegInB37[30] , \wRegInB37[29] , 
        \wRegInB37[28] , \wRegInB37[27] , \wRegInB37[26] , \wRegInB37[25] , 
        \wRegInB37[24] , \wRegInB37[23] , \wRegInB37[22] , \wRegInB37[21] , 
        \wRegInB37[20] , \wRegInB37[19] , \wRegInB37[18] , \wRegInB37[17] , 
        \wRegInB37[16] , \wRegInB37[15] , \wRegInB37[14] , \wRegInB37[13] , 
        \wRegInB37[12] , \wRegInB37[11] , \wRegInB37[10] , \wRegInB37[9] , 
        \wRegInB37[8] , \wRegInB37[7] , \wRegInB37[6] , \wRegInB37[5] , 
        \wRegInB37[4] , \wRegInB37[3] , \wRegInB37[2] , \wRegInB37[1] , 
        \wRegInB37[0] }), .Out({\wBIn37[31] , \wBIn37[30] , \wBIn37[29] , 
        \wBIn37[28] , \wBIn37[27] , \wBIn37[26] , \wBIn37[25] , \wBIn37[24] , 
        \wBIn37[23] , \wBIn37[22] , \wBIn37[21] , \wBIn37[20] , \wBIn37[19] , 
        \wBIn37[18] , \wBIn37[17] , \wBIn37[16] , \wBIn37[15] , \wBIn37[14] , 
        \wBIn37[13] , \wBIn37[12] , \wBIn37[11] , \wBIn37[10] , \wBIn37[9] , 
        \wBIn37[8] , \wBIn37[7] , \wBIn37[6] , \wBIn37[5] , \wBIn37[4] , 
        \wBIn37[3] , \wBIn37[2] , \wBIn37[1] , \wBIn37[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid36[31] , \wAMid36[30] , \wAMid36[29] , \wAMid36[28] , 
        \wAMid36[27] , \wAMid36[26] , \wAMid36[25] , \wAMid36[24] , 
        \wAMid36[23] , \wAMid36[22] , \wAMid36[21] , \wAMid36[20] , 
        \wAMid36[19] , \wAMid36[18] , \wAMid36[17] , \wAMid36[16] , 
        \wAMid36[15] , \wAMid36[14] , \wAMid36[13] , \wAMid36[12] , 
        \wAMid36[11] , \wAMid36[10] , \wAMid36[9] , \wAMid36[8] , \wAMid36[7] , 
        \wAMid36[6] , \wAMid36[5] , \wAMid36[4] , \wAMid36[3] , \wAMid36[2] , 
        \wAMid36[1] , \wAMid36[0] }), .BIn({\wBMid36[31] , \wBMid36[30] , 
        \wBMid36[29] , \wBMid36[28] , \wBMid36[27] , \wBMid36[26] , 
        \wBMid36[25] , \wBMid36[24] , \wBMid36[23] , \wBMid36[22] , 
        \wBMid36[21] , \wBMid36[20] , \wBMid36[19] , \wBMid36[18] , 
        \wBMid36[17] , \wBMid36[16] , \wBMid36[15] , \wBMid36[14] , 
        \wBMid36[13] , \wBMid36[12] , \wBMid36[11] , \wBMid36[10] , 
        \wBMid36[9] , \wBMid36[8] , \wBMid36[7] , \wBMid36[6] , \wBMid36[5] , 
        \wBMid36[4] , \wBMid36[3] , \wBMid36[2] , \wBMid36[1] , \wBMid36[0] }), 
        .HiOut({\wRegInB36[31] , \wRegInB36[30] , \wRegInB36[29] , 
        \wRegInB36[28] , \wRegInB36[27] , \wRegInB36[26] , \wRegInB36[25] , 
        \wRegInB36[24] , \wRegInB36[23] , \wRegInB36[22] , \wRegInB36[21] , 
        \wRegInB36[20] , \wRegInB36[19] , \wRegInB36[18] , \wRegInB36[17] , 
        \wRegInB36[16] , \wRegInB36[15] , \wRegInB36[14] , \wRegInB36[13] , 
        \wRegInB36[12] , \wRegInB36[11] , \wRegInB36[10] , \wRegInB36[9] , 
        \wRegInB36[8] , \wRegInB36[7] , \wRegInB36[6] , \wRegInB36[5] , 
        \wRegInB36[4] , \wRegInB36[3] , \wRegInB36[2] , \wRegInB36[1] , 
        \wRegInB36[0] }), .LoOut({\wRegInA37[31] , \wRegInA37[30] , 
        \wRegInA37[29] , \wRegInA37[28] , \wRegInA37[27] , \wRegInA37[26] , 
        \wRegInA37[25] , \wRegInA37[24] , \wRegInA37[23] , \wRegInA37[22] , 
        \wRegInA37[21] , \wRegInA37[20] , \wRegInA37[19] , \wRegInA37[18] , 
        \wRegInA37[17] , \wRegInA37[16] , \wRegInA37[15] , \wRegInA37[14] , 
        \wRegInA37[13] , \wRegInA37[12] , \wRegInA37[11] , \wRegInA37[10] , 
        \wRegInA37[9] , \wRegInA37[8] , \wRegInA37[7] , \wRegInA37[6] , 
        \wRegInA37[5] , \wRegInA37[4] , \wRegInA37[3] , \wRegInA37[2] , 
        \wRegInA37[1] , \wRegInA37[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_233 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink234[31] , \ScanLink234[30] , \ScanLink234[29] , 
        \ScanLink234[28] , \ScanLink234[27] , \ScanLink234[26] , 
        \ScanLink234[25] , \ScanLink234[24] , \ScanLink234[23] , 
        \ScanLink234[22] , \ScanLink234[21] , \ScanLink234[20] , 
        \ScanLink234[19] , \ScanLink234[18] , \ScanLink234[17] , 
        \ScanLink234[16] , \ScanLink234[15] , \ScanLink234[14] , 
        \ScanLink234[13] , \ScanLink234[12] , \ScanLink234[11] , 
        \ScanLink234[10] , \ScanLink234[9] , \ScanLink234[8] , 
        \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , \ScanLink234[4] , 
        \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , \ScanLink234[0] 
        }), .ScanOut({\ScanLink233[31] , \ScanLink233[30] , \ScanLink233[29] , 
        \ScanLink233[28] , \ScanLink233[27] , \ScanLink233[26] , 
        \ScanLink233[25] , \ScanLink233[24] , \ScanLink233[23] , 
        \ScanLink233[22] , \ScanLink233[21] , \ScanLink233[20] , 
        \ScanLink233[19] , \ScanLink233[18] , \ScanLink233[17] , 
        \ScanLink233[16] , \ScanLink233[15] , \ScanLink233[14] , 
        \ScanLink233[13] , \ScanLink233[12] , \ScanLink233[11] , 
        \ScanLink233[10] , \ScanLink233[9] , \ScanLink233[8] , 
        \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , \ScanLink233[4] , 
        \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , \ScanLink233[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA11[31] , \wRegInA11[30] , \wRegInA11[29] , 
        \wRegInA11[28] , \wRegInA11[27] , \wRegInA11[26] , \wRegInA11[25] , 
        \wRegInA11[24] , \wRegInA11[23] , \wRegInA11[22] , \wRegInA11[21] , 
        \wRegInA11[20] , \wRegInA11[19] , \wRegInA11[18] , \wRegInA11[17] , 
        \wRegInA11[16] , \wRegInA11[15] , \wRegInA11[14] , \wRegInA11[13] , 
        \wRegInA11[12] , \wRegInA11[11] , \wRegInA11[10] , \wRegInA11[9] , 
        \wRegInA11[8] , \wRegInA11[7] , \wRegInA11[6] , \wRegInA11[5] , 
        \wRegInA11[4] , \wRegInA11[3] , \wRegInA11[2] , \wRegInA11[1] , 
        \wRegInA11[0] }), .Out({\wAIn11[31] , \wAIn11[30] , \wAIn11[29] , 
        \wAIn11[28] , \wAIn11[27] , \wAIn11[26] , \wAIn11[25] , \wAIn11[24] , 
        \wAIn11[23] , \wAIn11[22] , \wAIn11[21] , \wAIn11[20] , \wAIn11[19] , 
        \wAIn11[18] , \wAIn11[17] , \wAIn11[16] , \wAIn11[15] , \wAIn11[14] , 
        \wAIn11[13] , \wAIn11[12] , \wAIn11[11] , \wAIn11[10] , \wAIn11[9] , 
        \wAIn11[8] , \wAIn11[7] , \wAIn11[6] , \wAIn11[5] , \wAIn11[4] , 
        \wAIn11[3] , \wAIn11[2] , \wAIn11[1] , \wAIn11[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_103 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink104[31] , \ScanLink104[30] , \ScanLink104[29] , 
        \ScanLink104[28] , \ScanLink104[27] , \ScanLink104[26] , 
        \ScanLink104[25] , \ScanLink104[24] , \ScanLink104[23] , 
        \ScanLink104[22] , \ScanLink104[21] , \ScanLink104[20] , 
        \ScanLink104[19] , \ScanLink104[18] , \ScanLink104[17] , 
        \ScanLink104[16] , \ScanLink104[15] , \ScanLink104[14] , 
        \ScanLink104[13] , \ScanLink104[12] , \ScanLink104[11] , 
        \ScanLink104[10] , \ScanLink104[9] , \ScanLink104[8] , 
        \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , \ScanLink104[4] , 
        \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , \ScanLink104[0] 
        }), .ScanOut({\ScanLink103[31] , \ScanLink103[30] , \ScanLink103[29] , 
        \ScanLink103[28] , \ScanLink103[27] , \ScanLink103[26] , 
        \ScanLink103[25] , \ScanLink103[24] , \ScanLink103[23] , 
        \ScanLink103[22] , \ScanLink103[21] , \ScanLink103[20] , 
        \ScanLink103[19] , \ScanLink103[18] , \ScanLink103[17] , 
        \ScanLink103[16] , \ScanLink103[15] , \ScanLink103[14] , 
        \ScanLink103[13] , \ScanLink103[12] , \ScanLink103[11] , 
        \ScanLink103[10] , \ScanLink103[9] , \ScanLink103[8] , 
        \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , \ScanLink103[4] , 
        \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , \ScanLink103[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA76[31] , \wRegInA76[30] , \wRegInA76[29] , 
        \wRegInA76[28] , \wRegInA76[27] , \wRegInA76[26] , \wRegInA76[25] , 
        \wRegInA76[24] , \wRegInA76[23] , \wRegInA76[22] , \wRegInA76[21] , 
        \wRegInA76[20] , \wRegInA76[19] , \wRegInA76[18] , \wRegInA76[17] , 
        \wRegInA76[16] , \wRegInA76[15] , \wRegInA76[14] , \wRegInA76[13] , 
        \wRegInA76[12] , \wRegInA76[11] , \wRegInA76[10] , \wRegInA76[9] , 
        \wRegInA76[8] , \wRegInA76[7] , \wRegInA76[6] , \wRegInA76[5] , 
        \wRegInA76[4] , \wRegInA76[3] , \wRegInA76[2] , \wRegInA76[1] , 
        \wRegInA76[0] }), .Out({\wAIn76[31] , \wAIn76[30] , \wAIn76[29] , 
        \wAIn76[28] , \wAIn76[27] , \wAIn76[26] , \wAIn76[25] , \wAIn76[24] , 
        \wAIn76[23] , \wAIn76[22] , \wAIn76[21] , \wAIn76[20] , \wAIn76[19] , 
        \wAIn76[18] , \wAIn76[17] , \wAIn76[16] , \wAIn76[15] , \wAIn76[14] , 
        \wAIn76[13] , \wAIn76[12] , \wAIn76[11] , \wAIn76[10] , \wAIn76[9] , 
        \wAIn76[8] , \wAIn76[7] , \wAIn76[6] , \wAIn76[5] , \wAIn76[4] , 
        \wAIn76[3] , \wAIn76[2] , \wAIn76[1] , \wAIn76[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_53 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink54[31] , \ScanLink54[30] , \ScanLink54[29] , 
        \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , \ScanLink54[25] , 
        \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , \ScanLink54[21] , 
        \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , \ScanLink54[17] , 
        \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , \ScanLink54[13] , 
        \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , \ScanLink54[9] , 
        \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , \ScanLink54[5] , 
        \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , \ScanLink54[1] , 
        \ScanLink54[0] }), .ScanOut({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA101[31] , \wRegInA101[30] , 
        \wRegInA101[29] , \wRegInA101[28] , \wRegInA101[27] , \wRegInA101[26] , 
        \wRegInA101[25] , \wRegInA101[24] , \wRegInA101[23] , \wRegInA101[22] , 
        \wRegInA101[21] , \wRegInA101[20] , \wRegInA101[19] , \wRegInA101[18] , 
        \wRegInA101[17] , \wRegInA101[16] , \wRegInA101[15] , \wRegInA101[14] , 
        \wRegInA101[13] , \wRegInA101[12] , \wRegInA101[11] , \wRegInA101[10] , 
        \wRegInA101[9] , \wRegInA101[8] , \wRegInA101[7] , \wRegInA101[6] , 
        \wRegInA101[5] , \wRegInA101[4] , \wRegInA101[3] , \wRegInA101[2] , 
        \wRegInA101[1] , \wRegInA101[0] }), .Out({\wAIn101[31] , \wAIn101[30] , 
        \wAIn101[29] , \wAIn101[28] , \wAIn101[27] , \wAIn101[26] , 
        \wAIn101[25] , \wAIn101[24] , \wAIn101[23] , \wAIn101[22] , 
        \wAIn101[21] , \wAIn101[20] , \wAIn101[19] , \wAIn101[18] , 
        \wAIn101[17] , \wAIn101[16] , \wAIn101[15] , \wAIn101[14] , 
        \wAIn101[13] , \wAIn101[12] , \wAIn101[11] , \wAIn101[10] , 
        \wAIn101[9] , \wAIn101[8] , \wAIn101[7] , \wAIn101[6] , \wAIn101[5] , 
        \wAIn101[4] , \wAIn101[3] , \wAIn101[2] , \wAIn101[1] , \wAIn101[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn28[31] , \wAIn28[30] , \wAIn28[29] , \wAIn28[28] , \wAIn28[27] , 
        \wAIn28[26] , \wAIn28[25] , \wAIn28[24] , \wAIn28[23] , \wAIn28[22] , 
        \wAIn28[21] , \wAIn28[20] , \wAIn28[19] , \wAIn28[18] , \wAIn28[17] , 
        \wAIn28[16] , \wAIn28[15] , \wAIn28[14] , \wAIn28[13] , \wAIn28[12] , 
        \wAIn28[11] , \wAIn28[10] , \wAIn28[9] , \wAIn28[8] , \wAIn28[7] , 
        \wAIn28[6] , \wAIn28[5] , \wAIn28[4] , \wAIn28[3] , \wAIn28[2] , 
        \wAIn28[1] , \wAIn28[0] }), .BIn({\wBIn28[31] , \wBIn28[30] , 
        \wBIn28[29] , \wBIn28[28] , \wBIn28[27] , \wBIn28[26] , \wBIn28[25] , 
        \wBIn28[24] , \wBIn28[23] , \wBIn28[22] , \wBIn28[21] , \wBIn28[20] , 
        \wBIn28[19] , \wBIn28[18] , \wBIn28[17] , \wBIn28[16] , \wBIn28[15] , 
        \wBIn28[14] , \wBIn28[13] , \wBIn28[12] , \wBIn28[11] , \wBIn28[10] , 
        \wBIn28[9] , \wBIn28[8] , \wBIn28[7] , \wBIn28[6] , \wBIn28[5] , 
        \wBIn28[4] , \wBIn28[3] , \wBIn28[2] , \wBIn28[1] , \wBIn28[0] }), 
        .HiOut({\wBMid27[31] , \wBMid27[30] , \wBMid27[29] , \wBMid27[28] , 
        \wBMid27[27] , \wBMid27[26] , \wBMid27[25] , \wBMid27[24] , 
        \wBMid27[23] , \wBMid27[22] , \wBMid27[21] , \wBMid27[20] , 
        \wBMid27[19] , \wBMid27[18] , \wBMid27[17] , \wBMid27[16] , 
        \wBMid27[15] , \wBMid27[14] , \wBMid27[13] , \wBMid27[12] , 
        \wBMid27[11] , \wBMid27[10] , \wBMid27[9] , \wBMid27[8] , \wBMid27[7] , 
        \wBMid27[6] , \wBMid27[5] , \wBMid27[4] , \wBMid27[3] , \wBMid27[2] , 
        \wBMid27[1] , \wBMid27[0] }), .LoOut({\wAMid28[31] , \wAMid28[30] , 
        \wAMid28[29] , \wAMid28[28] , \wAMid28[27] , \wAMid28[26] , 
        \wAMid28[25] , \wAMid28[24] , \wAMid28[23] , \wAMid28[22] , 
        \wAMid28[21] , \wAMid28[20] , \wAMid28[19] , \wAMid28[18] , 
        \wAMid28[17] , \wAMid28[16] , \wAMid28[15] , \wAMid28[14] , 
        \wAMid28[13] , \wAMid28[12] , \wAMid28[11] , \wAMid28[10] , 
        \wAMid28[9] , \wAMid28[8] , \wAMid28[7] , \wAMid28[6] , \wAMid28[5] , 
        \wAMid28[4] , \wAMid28[3] , \wAMid28[2] , \wAMid28[1] , \wAMid28[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn54[31] , \wAIn54[30] , \wAIn54[29] , \wAIn54[28] , \wAIn54[27] , 
        \wAIn54[26] , \wAIn54[25] , \wAIn54[24] , \wAIn54[23] , \wAIn54[22] , 
        \wAIn54[21] , \wAIn54[20] , \wAIn54[19] , \wAIn54[18] , \wAIn54[17] , 
        \wAIn54[16] , \wAIn54[15] , \wAIn54[14] , \wAIn54[13] , \wAIn54[12] , 
        \wAIn54[11] , \wAIn54[10] , \wAIn54[9] , \wAIn54[8] , \wAIn54[7] , 
        \wAIn54[6] , \wAIn54[5] , \wAIn54[4] , \wAIn54[3] , \wAIn54[2] , 
        \wAIn54[1] , \wAIn54[0] }), .BIn({\wBIn54[31] , \wBIn54[30] , 
        \wBIn54[29] , \wBIn54[28] , \wBIn54[27] , \wBIn54[26] , \wBIn54[25] , 
        \wBIn54[24] , \wBIn54[23] , \wBIn54[22] , \wBIn54[21] , \wBIn54[20] , 
        \wBIn54[19] , \wBIn54[18] , \wBIn54[17] , \wBIn54[16] , \wBIn54[15] , 
        \wBIn54[14] , \wBIn54[13] , \wBIn54[12] , \wBIn54[11] , \wBIn54[10] , 
        \wBIn54[9] , \wBIn54[8] , \wBIn54[7] , \wBIn54[6] , \wBIn54[5] , 
        \wBIn54[4] , \wBIn54[3] , \wBIn54[2] , \wBIn54[1] , \wBIn54[0] }), 
        .HiOut({\wBMid53[31] , \wBMid53[30] , \wBMid53[29] , \wBMid53[28] , 
        \wBMid53[27] , \wBMid53[26] , \wBMid53[25] , \wBMid53[24] , 
        \wBMid53[23] , \wBMid53[22] , \wBMid53[21] , \wBMid53[20] , 
        \wBMid53[19] , \wBMid53[18] , \wBMid53[17] , \wBMid53[16] , 
        \wBMid53[15] , \wBMid53[14] , \wBMid53[13] , \wBMid53[12] , 
        \wBMid53[11] , \wBMid53[10] , \wBMid53[9] , \wBMid53[8] , \wBMid53[7] , 
        \wBMid53[6] , \wBMid53[5] , \wBMid53[4] , \wBMid53[3] , \wBMid53[2] , 
        \wBMid53[1] , \wBMid53[0] }), .LoOut({\wAMid54[31] , \wAMid54[30] , 
        \wAMid54[29] , \wAMid54[28] , \wAMid54[27] , \wAMid54[26] , 
        \wAMid54[25] , \wAMid54[24] , \wAMid54[23] , \wAMid54[22] , 
        \wAMid54[21] , \wAMid54[20] , \wAMid54[19] , \wAMid54[18] , 
        \wAMid54[17] , \wAMid54[16] , \wAMid54[15] , \wAMid54[14] , 
        \wAMid54[13] , \wAMid54[12] , \wAMid54[11] , \wAMid54[10] , 
        \wAMid54[9] , \wAMid54[8] , \wAMid54[7] , \wAMid54[6] , \wAMid54[5] , 
        \wAMid54[4] , \wAMid54[3] , \wAMid54[2] , \wAMid54[1] , \wAMid54[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn68[31] , \wAIn68[30] , \wAIn68[29] , \wAIn68[28] , \wAIn68[27] , 
        \wAIn68[26] , \wAIn68[25] , \wAIn68[24] , \wAIn68[23] , \wAIn68[22] , 
        \wAIn68[21] , \wAIn68[20] , \wAIn68[19] , \wAIn68[18] , \wAIn68[17] , 
        \wAIn68[16] , \wAIn68[15] , \wAIn68[14] , \wAIn68[13] , \wAIn68[12] , 
        \wAIn68[11] , \wAIn68[10] , \wAIn68[9] , \wAIn68[8] , \wAIn68[7] , 
        \wAIn68[6] , \wAIn68[5] , \wAIn68[4] , \wAIn68[3] , \wAIn68[2] , 
        \wAIn68[1] , \wAIn68[0] }), .BIn({\wBIn68[31] , \wBIn68[30] , 
        \wBIn68[29] , \wBIn68[28] , \wBIn68[27] , \wBIn68[26] , \wBIn68[25] , 
        \wBIn68[24] , \wBIn68[23] , \wBIn68[22] , \wBIn68[21] , \wBIn68[20] , 
        \wBIn68[19] , \wBIn68[18] , \wBIn68[17] , \wBIn68[16] , \wBIn68[15] , 
        \wBIn68[14] , \wBIn68[13] , \wBIn68[12] , \wBIn68[11] , \wBIn68[10] , 
        \wBIn68[9] , \wBIn68[8] , \wBIn68[7] , \wBIn68[6] , \wBIn68[5] , 
        \wBIn68[4] , \wBIn68[3] , \wBIn68[2] , \wBIn68[1] , \wBIn68[0] }), 
        .HiOut({\wBMid67[31] , \wBMid67[30] , \wBMid67[29] , \wBMid67[28] , 
        \wBMid67[27] , \wBMid67[26] , \wBMid67[25] , \wBMid67[24] , 
        \wBMid67[23] , \wBMid67[22] , \wBMid67[21] , \wBMid67[20] , 
        \wBMid67[19] , \wBMid67[18] , \wBMid67[17] , \wBMid67[16] , 
        \wBMid67[15] , \wBMid67[14] , \wBMid67[13] , \wBMid67[12] , 
        \wBMid67[11] , \wBMid67[10] , \wBMid67[9] , \wBMid67[8] , \wBMid67[7] , 
        \wBMid67[6] , \wBMid67[5] , \wBMid67[4] , \wBMid67[3] , \wBMid67[2] , 
        \wBMid67[1] , \wBMid67[0] }), .LoOut({\wAMid68[31] , \wAMid68[30] , 
        \wAMid68[29] , \wAMid68[28] , \wAMid68[27] , \wAMid68[26] , 
        \wAMid68[25] , \wAMid68[24] , \wAMid68[23] , \wAMid68[22] , 
        \wAMid68[21] , \wAMid68[20] , \wAMid68[19] , \wAMid68[18] , 
        \wAMid68[17] , \wAMid68[16] , \wAMid68[15] , \wAMid68[14] , 
        \wAMid68[13] , \wAMid68[12] , \wAMid68[11] , \wAMid68[10] , 
        \wAMid68[9] , \wAMid68[8] , \wAMid68[7] , \wAMid68[6] , \wAMid68[5] , 
        \wAMid68[4] , \wAMid68[3] , \wAMid68[2] , \wAMid68[1] , \wAMid68[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn118[31] , \wAIn118[30] , \wAIn118[29] , \wAIn118[28] , 
        \wAIn118[27] , \wAIn118[26] , \wAIn118[25] , \wAIn118[24] , 
        \wAIn118[23] , \wAIn118[22] , \wAIn118[21] , \wAIn118[20] , 
        \wAIn118[19] , \wAIn118[18] , \wAIn118[17] , \wAIn118[16] , 
        \wAIn118[15] , \wAIn118[14] , \wAIn118[13] , \wAIn118[12] , 
        \wAIn118[11] , \wAIn118[10] , \wAIn118[9] , \wAIn118[8] , \wAIn118[7] , 
        \wAIn118[6] , \wAIn118[5] , \wAIn118[4] , \wAIn118[3] , \wAIn118[2] , 
        \wAIn118[1] , \wAIn118[0] }), .BIn({\wBIn118[31] , \wBIn118[30] , 
        \wBIn118[29] , \wBIn118[28] , \wBIn118[27] , \wBIn118[26] , 
        \wBIn118[25] , \wBIn118[24] , \wBIn118[23] , \wBIn118[22] , 
        \wBIn118[21] , \wBIn118[20] , \wBIn118[19] , \wBIn118[18] , 
        \wBIn118[17] , \wBIn118[16] , \wBIn118[15] , \wBIn118[14] , 
        \wBIn118[13] , \wBIn118[12] , \wBIn118[11] , \wBIn118[10] , 
        \wBIn118[9] , \wBIn118[8] , \wBIn118[7] , \wBIn118[6] , \wBIn118[5] , 
        \wBIn118[4] , \wBIn118[3] , \wBIn118[2] , \wBIn118[1] , \wBIn118[0] }), 
        .HiOut({\wBMid117[31] , \wBMid117[30] , \wBMid117[29] , \wBMid117[28] , 
        \wBMid117[27] , \wBMid117[26] , \wBMid117[25] , \wBMid117[24] , 
        \wBMid117[23] , \wBMid117[22] , \wBMid117[21] , \wBMid117[20] , 
        \wBMid117[19] , \wBMid117[18] , \wBMid117[17] , \wBMid117[16] , 
        \wBMid117[15] , \wBMid117[14] , \wBMid117[13] , \wBMid117[12] , 
        \wBMid117[11] , \wBMid117[10] , \wBMid117[9] , \wBMid117[8] , 
        \wBMid117[7] , \wBMid117[6] , \wBMid117[5] , \wBMid117[4] , 
        \wBMid117[3] , \wBMid117[2] , \wBMid117[1] , \wBMid117[0] }), .LoOut({
        \wAMid118[31] , \wAMid118[30] , \wAMid118[29] , \wAMid118[28] , 
        \wAMid118[27] , \wAMid118[26] , \wAMid118[25] , \wAMid118[24] , 
        \wAMid118[23] , \wAMid118[22] , \wAMid118[21] , \wAMid118[20] , 
        \wAMid118[19] , \wAMid118[18] , \wAMid118[17] , \wAMid118[16] , 
        \wAMid118[15] , \wAMid118[14] , \wAMid118[13] , \wAMid118[12] , 
        \wAMid118[11] , \wAMid118[10] , \wAMid118[9] , \wAMid118[8] , 
        \wAMid118[7] , \wAMid118[6] , \wAMid118[5] , \wAMid118[4] , 
        \wAMid118[3] , \wAMid118[2] , \wAMid118[1] , \wAMid118[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid11[31] , \wAMid11[30] , \wAMid11[29] , \wAMid11[28] , 
        \wAMid11[27] , \wAMid11[26] , \wAMid11[25] , \wAMid11[24] , 
        \wAMid11[23] , \wAMid11[22] , \wAMid11[21] , \wAMid11[20] , 
        \wAMid11[19] , \wAMid11[18] , \wAMid11[17] , \wAMid11[16] , 
        \wAMid11[15] , \wAMid11[14] , \wAMid11[13] , \wAMid11[12] , 
        \wAMid11[11] , \wAMid11[10] , \wAMid11[9] , \wAMid11[8] , \wAMid11[7] , 
        \wAMid11[6] , \wAMid11[5] , \wAMid11[4] , \wAMid11[3] , \wAMid11[2] , 
        \wAMid11[1] , \wAMid11[0] }), .BIn({\wBMid11[31] , \wBMid11[30] , 
        \wBMid11[29] , \wBMid11[28] , \wBMid11[27] , \wBMid11[26] , 
        \wBMid11[25] , \wBMid11[24] , \wBMid11[23] , \wBMid11[22] , 
        \wBMid11[21] , \wBMid11[20] , \wBMid11[19] , \wBMid11[18] , 
        \wBMid11[17] , \wBMid11[16] , \wBMid11[15] , \wBMid11[14] , 
        \wBMid11[13] , \wBMid11[12] , \wBMid11[11] , \wBMid11[10] , 
        \wBMid11[9] , \wBMid11[8] , \wBMid11[7] , \wBMid11[6] , \wBMid11[5] , 
        \wBMid11[4] , \wBMid11[3] , \wBMid11[2] , \wBMid11[1] , \wBMid11[0] }), 
        .HiOut({\wRegInB11[31] , \wRegInB11[30] , \wRegInB11[29] , 
        \wRegInB11[28] , \wRegInB11[27] , \wRegInB11[26] , \wRegInB11[25] , 
        \wRegInB11[24] , \wRegInB11[23] , \wRegInB11[22] , \wRegInB11[21] , 
        \wRegInB11[20] , \wRegInB11[19] , \wRegInB11[18] , \wRegInB11[17] , 
        \wRegInB11[16] , \wRegInB11[15] , \wRegInB11[14] , \wRegInB11[13] , 
        \wRegInB11[12] , \wRegInB11[11] , \wRegInB11[10] , \wRegInB11[9] , 
        \wRegInB11[8] , \wRegInB11[7] , \wRegInB11[6] , \wRegInB11[5] , 
        \wRegInB11[4] , \wRegInB11[3] , \wRegInB11[2] , \wRegInB11[1] , 
        \wRegInB11[0] }), .LoOut({\wRegInA12[31] , \wRegInA12[30] , 
        \wRegInA12[29] , \wRegInA12[28] , \wRegInA12[27] , \wRegInA12[26] , 
        \wRegInA12[25] , \wRegInA12[24] , \wRegInA12[23] , \wRegInA12[22] , 
        \wRegInA12[21] , \wRegInA12[20] , \wRegInA12[19] , \wRegInA12[18] , 
        \wRegInA12[17] , \wRegInA12[16] , \wRegInA12[15] , \wRegInA12[14] , 
        \wRegInA12[13] , \wRegInA12[12] , \wRegInA12[11] , \wRegInA12[10] , 
        \wRegInA12[9] , \wRegInA12[8] , \wRegInA12[7] , \wRegInA12[6] , 
        \wRegInA12[5] , \wRegInA12[4] , \wRegInA12[3] , \wRegInA12[2] , 
        \wRegInA12[1] , \wRegInA12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_124 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink125[31] , \ScanLink125[30] , \ScanLink125[29] , 
        \ScanLink125[28] , \ScanLink125[27] , \ScanLink125[26] , 
        \ScanLink125[25] , \ScanLink125[24] , \ScanLink125[23] , 
        \ScanLink125[22] , \ScanLink125[21] , \ScanLink125[20] , 
        \ScanLink125[19] , \ScanLink125[18] , \ScanLink125[17] , 
        \ScanLink125[16] , \ScanLink125[15] , \ScanLink125[14] , 
        \ScanLink125[13] , \ScanLink125[12] , \ScanLink125[11] , 
        \ScanLink125[10] , \ScanLink125[9] , \ScanLink125[8] , 
        \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , \ScanLink125[4] , 
        \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , \ScanLink125[0] 
        }), .ScanOut({\ScanLink124[31] , \ScanLink124[30] , \ScanLink124[29] , 
        \ScanLink124[28] , \ScanLink124[27] , \ScanLink124[26] , 
        \ScanLink124[25] , \ScanLink124[24] , \ScanLink124[23] , 
        \ScanLink124[22] , \ScanLink124[21] , \ScanLink124[20] , 
        \ScanLink124[19] , \ScanLink124[18] , \ScanLink124[17] , 
        \ScanLink124[16] , \ScanLink124[15] , \ScanLink124[14] , 
        \ScanLink124[13] , \ScanLink124[12] , \ScanLink124[11] , 
        \ScanLink124[10] , \ScanLink124[9] , \ScanLink124[8] , 
        \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , \ScanLink124[4] , 
        \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , \ScanLink124[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB65[31] , \wRegInB65[30] , \wRegInB65[29] , 
        \wRegInB65[28] , \wRegInB65[27] , \wRegInB65[26] , \wRegInB65[25] , 
        \wRegInB65[24] , \wRegInB65[23] , \wRegInB65[22] , \wRegInB65[21] , 
        \wRegInB65[20] , \wRegInB65[19] , \wRegInB65[18] , \wRegInB65[17] , 
        \wRegInB65[16] , \wRegInB65[15] , \wRegInB65[14] , \wRegInB65[13] , 
        \wRegInB65[12] , \wRegInB65[11] , \wRegInB65[10] , \wRegInB65[9] , 
        \wRegInB65[8] , \wRegInB65[7] , \wRegInB65[6] , \wRegInB65[5] , 
        \wRegInB65[4] , \wRegInB65[3] , \wRegInB65[2] , \wRegInB65[1] , 
        \wRegInB65[0] }), .Out({\wBIn65[31] , \wBIn65[30] , \wBIn65[29] , 
        \wBIn65[28] , \wBIn65[27] , \wBIn65[26] , \wBIn65[25] , \wBIn65[24] , 
        \wBIn65[23] , \wBIn65[22] , \wBIn65[21] , \wBIn65[20] , \wBIn65[19] , 
        \wBIn65[18] , \wBIn65[17] , \wBIn65[16] , \wBIn65[15] , \wBIn65[14] , 
        \wBIn65[13] , \wBIn65[12] , \wBIn65[11] , \wBIn65[10] , \wBIn65[9] , 
        \wBIn65[8] , \wBIn65[7] , \wBIn65[6] , \wBIn65[5] , \wBIn65[4] , 
        \wBIn65[3] , \wBIn65[2] , \wBIn65[1] , \wBIn65[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_74 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink75[31] , \ScanLink75[30] , \ScanLink75[29] , 
        \ScanLink75[28] , \ScanLink75[27] , \ScanLink75[26] , \ScanLink75[25] , 
        \ScanLink75[24] , \ScanLink75[23] , \ScanLink75[22] , \ScanLink75[21] , 
        \ScanLink75[20] , \ScanLink75[19] , \ScanLink75[18] , \ScanLink75[17] , 
        \ScanLink75[16] , \ScanLink75[15] , \ScanLink75[14] , \ScanLink75[13] , 
        \ScanLink75[12] , \ScanLink75[11] , \ScanLink75[10] , \ScanLink75[9] , 
        \ScanLink75[8] , \ScanLink75[7] , \ScanLink75[6] , \ScanLink75[5] , 
        \ScanLink75[4] , \ScanLink75[3] , \ScanLink75[2] , \ScanLink75[1] , 
        \ScanLink75[0] }), .ScanOut({\ScanLink74[31] , \ScanLink74[30] , 
        \ScanLink74[29] , \ScanLink74[28] , \ScanLink74[27] , \ScanLink74[26] , 
        \ScanLink74[25] , \ScanLink74[24] , \ScanLink74[23] , \ScanLink74[22] , 
        \ScanLink74[21] , \ScanLink74[20] , \ScanLink74[19] , \ScanLink74[18] , 
        \ScanLink74[17] , \ScanLink74[16] , \ScanLink74[15] , \ScanLink74[14] , 
        \ScanLink74[13] , \ScanLink74[12] , \ScanLink74[11] , \ScanLink74[10] , 
        \ScanLink74[9] , \ScanLink74[8] , \ScanLink74[7] , \ScanLink74[6] , 
        \ScanLink74[5] , \ScanLink74[4] , \ScanLink74[3] , \ScanLink74[2] , 
        \ScanLink74[1] , \ScanLink74[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB90[31] , \wRegInB90[30] , 
        \wRegInB90[29] , \wRegInB90[28] , \wRegInB90[27] , \wRegInB90[26] , 
        \wRegInB90[25] , \wRegInB90[24] , \wRegInB90[23] , \wRegInB90[22] , 
        \wRegInB90[21] , \wRegInB90[20] , \wRegInB90[19] , \wRegInB90[18] , 
        \wRegInB90[17] , \wRegInB90[16] , \wRegInB90[15] , \wRegInB90[14] , 
        \wRegInB90[13] , \wRegInB90[12] , \wRegInB90[11] , \wRegInB90[10] , 
        \wRegInB90[9] , \wRegInB90[8] , \wRegInB90[7] , \wRegInB90[6] , 
        \wRegInB90[5] , \wRegInB90[4] , \wRegInB90[3] , \wRegInB90[2] , 
        \wRegInB90[1] , \wRegInB90[0] }), .Out({\wBIn90[31] , \wBIn90[30] , 
        \wBIn90[29] , \wBIn90[28] , \wBIn90[27] , \wBIn90[26] , \wBIn90[25] , 
        \wBIn90[24] , \wBIn90[23] , \wBIn90[22] , \wBIn90[21] , \wBIn90[20] , 
        \wBIn90[19] , \wBIn90[18] , \wBIn90[17] , \wBIn90[16] , \wBIn90[15] , 
        \wBIn90[14] , \wBIn90[13] , \wBIn90[12] , \wBIn90[11] , \wBIn90[10] , 
        \wBIn90[9] , \wBIn90[8] , \wBIn90[7] , \wBIn90[6] , \wBIn90[5] , 
        \wBIn90[4] , \wBIn90[3] , \wBIn90[2] , \wBIn90[1] , \wBIn90[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid112[31] , \wAMid112[30] , \wAMid112[29] , \wAMid112[28] , 
        \wAMid112[27] , \wAMid112[26] , \wAMid112[25] , \wAMid112[24] , 
        \wAMid112[23] , \wAMid112[22] , \wAMid112[21] , \wAMid112[20] , 
        \wAMid112[19] , \wAMid112[18] , \wAMid112[17] , \wAMid112[16] , 
        \wAMid112[15] , \wAMid112[14] , \wAMid112[13] , \wAMid112[12] , 
        \wAMid112[11] , \wAMid112[10] , \wAMid112[9] , \wAMid112[8] , 
        \wAMid112[7] , \wAMid112[6] , \wAMid112[5] , \wAMid112[4] , 
        \wAMid112[3] , \wAMid112[2] , \wAMid112[1] , \wAMid112[0] }), .BIn({
        \wBMid112[31] , \wBMid112[30] , \wBMid112[29] , \wBMid112[28] , 
        \wBMid112[27] , \wBMid112[26] , \wBMid112[25] , \wBMid112[24] , 
        \wBMid112[23] , \wBMid112[22] , \wBMid112[21] , \wBMid112[20] , 
        \wBMid112[19] , \wBMid112[18] , \wBMid112[17] , \wBMid112[16] , 
        \wBMid112[15] , \wBMid112[14] , \wBMid112[13] , \wBMid112[12] , 
        \wBMid112[11] , \wBMid112[10] , \wBMid112[9] , \wBMid112[8] , 
        \wBMid112[7] , \wBMid112[6] , \wBMid112[5] , \wBMid112[4] , 
        \wBMid112[3] , \wBMid112[2] , \wBMid112[1] , \wBMid112[0] }), .HiOut({
        \wRegInB112[31] , \wRegInB112[30] , \wRegInB112[29] , \wRegInB112[28] , 
        \wRegInB112[27] , \wRegInB112[26] , \wRegInB112[25] , \wRegInB112[24] , 
        \wRegInB112[23] , \wRegInB112[22] , \wRegInB112[21] , \wRegInB112[20] , 
        \wRegInB112[19] , \wRegInB112[18] , \wRegInB112[17] , \wRegInB112[16] , 
        \wRegInB112[15] , \wRegInB112[14] , \wRegInB112[13] , \wRegInB112[12] , 
        \wRegInB112[11] , \wRegInB112[10] , \wRegInB112[9] , \wRegInB112[8] , 
        \wRegInB112[7] , \wRegInB112[6] , \wRegInB112[5] , \wRegInB112[4] , 
        \wRegInB112[3] , \wRegInB112[2] , \wRegInB112[1] , \wRegInB112[0] }), 
        .LoOut({\wRegInA113[31] , \wRegInA113[30] , \wRegInA113[29] , 
        \wRegInA113[28] , \wRegInA113[27] , \wRegInA113[26] , \wRegInA113[25] , 
        \wRegInA113[24] , \wRegInA113[23] , \wRegInA113[22] , \wRegInA113[21] , 
        \wRegInA113[20] , \wRegInA113[19] , \wRegInA113[18] , \wRegInA113[17] , 
        \wRegInA113[16] , \wRegInA113[15] , \wRegInA113[14] , \wRegInA113[13] , 
        \wRegInA113[12] , \wRegInA113[11] , \wRegInA113[10] , \wRegInA113[9] , 
        \wRegInA113[8] , \wRegInA113[7] , \wRegInA113[6] , \wRegInA113[5] , 
        \wRegInA113[4] , \wRegInA113[3] , \wRegInA113[2] , \wRegInA113[1] , 
        \wRegInA113[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_214 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink215[31] , \ScanLink215[30] , \ScanLink215[29] , 
        \ScanLink215[28] , \ScanLink215[27] , \ScanLink215[26] , 
        \ScanLink215[25] , \ScanLink215[24] , \ScanLink215[23] , 
        \ScanLink215[22] , \ScanLink215[21] , \ScanLink215[20] , 
        \ScanLink215[19] , \ScanLink215[18] , \ScanLink215[17] , 
        \ScanLink215[16] , \ScanLink215[15] , \ScanLink215[14] , 
        \ScanLink215[13] , \ScanLink215[12] , \ScanLink215[11] , 
        \ScanLink215[10] , \ScanLink215[9] , \ScanLink215[8] , 
        \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , \ScanLink215[4] , 
        \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , \ScanLink215[0] 
        }), .ScanOut({\ScanLink214[31] , \ScanLink214[30] , \ScanLink214[29] , 
        \ScanLink214[28] , \ScanLink214[27] , \ScanLink214[26] , 
        \ScanLink214[25] , \ScanLink214[24] , \ScanLink214[23] , 
        \ScanLink214[22] , \ScanLink214[21] , \ScanLink214[20] , 
        \ScanLink214[19] , \ScanLink214[18] , \ScanLink214[17] , 
        \ScanLink214[16] , \ScanLink214[15] , \ScanLink214[14] , 
        \ScanLink214[13] , \ScanLink214[12] , \ScanLink214[11] , 
        \ScanLink214[10] , \ScanLink214[9] , \ScanLink214[8] , 
        \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , \ScanLink214[4] , 
        \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , \ScanLink214[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB20[31] , \wRegInB20[30] , \wRegInB20[29] , 
        \wRegInB20[28] , \wRegInB20[27] , \wRegInB20[26] , \wRegInB20[25] , 
        \wRegInB20[24] , \wRegInB20[23] , \wRegInB20[22] , \wRegInB20[21] , 
        \wRegInB20[20] , \wRegInB20[19] , \wRegInB20[18] , \wRegInB20[17] , 
        \wRegInB20[16] , \wRegInB20[15] , \wRegInB20[14] , \wRegInB20[13] , 
        \wRegInB20[12] , \wRegInB20[11] , \wRegInB20[10] , \wRegInB20[9] , 
        \wRegInB20[8] , \wRegInB20[7] , \wRegInB20[6] , \wRegInB20[5] , 
        \wRegInB20[4] , \wRegInB20[3] , \wRegInB20[2] , \wRegInB20[1] , 
        \wRegInB20[0] }), .Out({\wBIn20[31] , \wBIn20[30] , \wBIn20[29] , 
        \wBIn20[28] , \wBIn20[27] , \wBIn20[26] , \wBIn20[25] , \wBIn20[24] , 
        \wBIn20[23] , \wBIn20[22] , \wBIn20[21] , \wBIn20[20] , \wBIn20[19] , 
        \wBIn20[18] , \wBIn20[17] , \wBIn20[16] , \wBIn20[15] , \wBIn20[14] , 
        \wBIn20[13] , \wBIn20[12] , \wBIn20[11] , \wBIn20[10] , \wBIn20[9] , 
        \wBIn20[8] , \wBIn20[7] , \wBIn20[6] , \wBIn20[5] , \wBIn20[4] , 
        \wBIn20[3] , \wBIn20[2] , \wBIn20[1] , \wBIn20[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_188 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink189[31] , \ScanLink189[30] , \ScanLink189[29] , 
        \ScanLink189[28] , \ScanLink189[27] , \ScanLink189[26] , 
        \ScanLink189[25] , \ScanLink189[24] , \ScanLink189[23] , 
        \ScanLink189[22] , \ScanLink189[21] , \ScanLink189[20] , 
        \ScanLink189[19] , \ScanLink189[18] , \ScanLink189[17] , 
        \ScanLink189[16] , \ScanLink189[15] , \ScanLink189[14] , 
        \ScanLink189[13] , \ScanLink189[12] , \ScanLink189[11] , 
        \ScanLink189[10] , \ScanLink189[9] , \ScanLink189[8] , 
        \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , \ScanLink189[4] , 
        \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , \ScanLink189[0] 
        }), .ScanOut({\ScanLink188[31] , \ScanLink188[30] , \ScanLink188[29] , 
        \ScanLink188[28] , \ScanLink188[27] , \ScanLink188[26] , 
        \ScanLink188[25] , \ScanLink188[24] , \ScanLink188[23] , 
        \ScanLink188[22] , \ScanLink188[21] , \ScanLink188[20] , 
        \ScanLink188[19] , \ScanLink188[18] , \ScanLink188[17] , 
        \ScanLink188[16] , \ScanLink188[15] , \ScanLink188[14] , 
        \ScanLink188[13] , \ScanLink188[12] , \ScanLink188[11] , 
        \ScanLink188[10] , \ScanLink188[9] , \ScanLink188[8] , 
        \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , \ScanLink188[4] , 
        \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , \ScanLink188[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB33[31] , \wRegInB33[30] , \wRegInB33[29] , 
        \wRegInB33[28] , \wRegInB33[27] , \wRegInB33[26] , \wRegInB33[25] , 
        \wRegInB33[24] , \wRegInB33[23] , \wRegInB33[22] , \wRegInB33[21] , 
        \wRegInB33[20] , \wRegInB33[19] , \wRegInB33[18] , \wRegInB33[17] , 
        \wRegInB33[16] , \wRegInB33[15] , \wRegInB33[14] , \wRegInB33[13] , 
        \wRegInB33[12] , \wRegInB33[11] , \wRegInB33[10] , \wRegInB33[9] , 
        \wRegInB33[8] , \wRegInB33[7] , \wRegInB33[6] , \wRegInB33[5] , 
        \wRegInB33[4] , \wRegInB33[3] , \wRegInB33[2] , \wRegInB33[1] , 
        \wRegInB33[0] }), .Out({\wBIn33[31] , \wBIn33[30] , \wBIn33[29] , 
        \wBIn33[28] , \wBIn33[27] , \wBIn33[26] , \wBIn33[25] , \wBIn33[24] , 
        \wBIn33[23] , \wBIn33[22] , \wBIn33[21] , \wBIn33[20] , \wBIn33[19] , 
        \wBIn33[18] , \wBIn33[17] , \wBIn33[16] , \wBIn33[15] , \wBIn33[14] , 
        \wBIn33[13] , \wBIn33[12] , \wBIn33[11] , \wBIn33[10] , \wBIn33[9] , 
        \wBIn33[8] , \wBIn33[7] , \wBIn33[6] , \wBIn33[5] , \wBIn33[4] , 
        \wBIn33[3] , \wBIn33[2] , \wBIn33[1] , \wBIn33[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_91 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink92[31] , \ScanLink92[30] , \ScanLink92[29] , 
        \ScanLink92[28] , \ScanLink92[27] , \ScanLink92[26] , \ScanLink92[25] , 
        \ScanLink92[24] , \ScanLink92[23] , \ScanLink92[22] , \ScanLink92[21] , 
        \ScanLink92[20] , \ScanLink92[19] , \ScanLink92[18] , \ScanLink92[17] , 
        \ScanLink92[16] , \ScanLink92[15] , \ScanLink92[14] , \ScanLink92[13] , 
        \ScanLink92[12] , \ScanLink92[11] , \ScanLink92[10] , \ScanLink92[9] , 
        \ScanLink92[8] , \ScanLink92[7] , \ScanLink92[6] , \ScanLink92[5] , 
        \ScanLink92[4] , \ScanLink92[3] , \ScanLink92[2] , \ScanLink92[1] , 
        \ScanLink92[0] }), .ScanOut({\ScanLink91[31] , \ScanLink91[30] , 
        \ScanLink91[29] , \ScanLink91[28] , \ScanLink91[27] , \ScanLink91[26] , 
        \ScanLink91[25] , \ScanLink91[24] , \ScanLink91[23] , \ScanLink91[22] , 
        \ScanLink91[21] , \ScanLink91[20] , \ScanLink91[19] , \ScanLink91[18] , 
        \ScanLink91[17] , \ScanLink91[16] , \ScanLink91[15] , \ScanLink91[14] , 
        \ScanLink91[13] , \ScanLink91[12] , \ScanLink91[11] , \ScanLink91[10] , 
        \ScanLink91[9] , \ScanLink91[8] , \ScanLink91[7] , \ScanLink91[6] , 
        \ScanLink91[5] , \ScanLink91[4] , \ScanLink91[3] , \ScanLink91[2] , 
        \ScanLink91[1] , \ScanLink91[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA82[31] , \wRegInA82[30] , 
        \wRegInA82[29] , \wRegInA82[28] , \wRegInA82[27] , \wRegInA82[26] , 
        \wRegInA82[25] , \wRegInA82[24] , \wRegInA82[23] , \wRegInA82[22] , 
        \wRegInA82[21] , \wRegInA82[20] , \wRegInA82[19] , \wRegInA82[18] , 
        \wRegInA82[17] , \wRegInA82[16] , \wRegInA82[15] , \wRegInA82[14] , 
        \wRegInA82[13] , \wRegInA82[12] , \wRegInA82[11] , \wRegInA82[10] , 
        \wRegInA82[9] , \wRegInA82[8] , \wRegInA82[7] , \wRegInA82[6] , 
        \wRegInA82[5] , \wRegInA82[4] , \wRegInA82[3] , \wRegInA82[2] , 
        \wRegInA82[1] , \wRegInA82[0] }), .Out({\wAIn82[31] , \wAIn82[30] , 
        \wAIn82[29] , \wAIn82[28] , \wAIn82[27] , \wAIn82[26] , \wAIn82[25] , 
        \wAIn82[24] , \wAIn82[23] , \wAIn82[22] , \wAIn82[21] , \wAIn82[20] , 
        \wAIn82[19] , \wAIn82[18] , \wAIn82[17] , \wAIn82[16] , \wAIn82[15] , 
        \wAIn82[14] , \wAIn82[13] , \wAIn82[12] , \wAIn82[11] , \wAIn82[10] , 
        \wAIn82[9] , \wAIn82[8] , \wAIn82[7] , \wAIn82[6] , \wAIn82[5] , 
        \wAIn82[4] , \wAIn82[3] , \wAIn82[2] , \wAIn82[1] , \wAIn82[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn73[31] , \wAIn73[30] , \wAIn73[29] , \wAIn73[28] , \wAIn73[27] , 
        \wAIn73[26] , \wAIn73[25] , \wAIn73[24] , \wAIn73[23] , \wAIn73[22] , 
        \wAIn73[21] , \wAIn73[20] , \wAIn73[19] , \wAIn73[18] , \wAIn73[17] , 
        \wAIn73[16] , \wAIn73[15] , \wAIn73[14] , \wAIn73[13] , \wAIn73[12] , 
        \wAIn73[11] , \wAIn73[10] , \wAIn73[9] , \wAIn73[8] , \wAIn73[7] , 
        \wAIn73[6] , \wAIn73[5] , \wAIn73[4] , \wAIn73[3] , \wAIn73[2] , 
        \wAIn73[1] , \wAIn73[0] }), .BIn({\wBIn73[31] , \wBIn73[30] , 
        \wBIn73[29] , \wBIn73[28] , \wBIn73[27] , \wBIn73[26] , \wBIn73[25] , 
        \wBIn73[24] , \wBIn73[23] , \wBIn73[22] , \wBIn73[21] , \wBIn73[20] , 
        \wBIn73[19] , \wBIn73[18] , \wBIn73[17] , \wBIn73[16] , \wBIn73[15] , 
        \wBIn73[14] , \wBIn73[13] , \wBIn73[12] , \wBIn73[11] , \wBIn73[10] , 
        \wBIn73[9] , \wBIn73[8] , \wBIn73[7] , \wBIn73[6] , \wBIn73[5] , 
        \wBIn73[4] , \wBIn73[3] , \wBIn73[2] , \wBIn73[1] , \wBIn73[0] }), 
        .HiOut({\wBMid72[31] , \wBMid72[30] , \wBMid72[29] , \wBMid72[28] , 
        \wBMid72[27] , \wBMid72[26] , \wBMid72[25] , \wBMid72[24] , 
        \wBMid72[23] , \wBMid72[22] , \wBMid72[21] , \wBMid72[20] , 
        \wBMid72[19] , \wBMid72[18] , \wBMid72[17] , \wBMid72[16] , 
        \wBMid72[15] , \wBMid72[14] , \wBMid72[13] , \wBMid72[12] , 
        \wBMid72[11] , \wBMid72[10] , \wBMid72[9] , \wBMid72[8] , \wBMid72[7] , 
        \wBMid72[6] , \wBMid72[5] , \wBMid72[4] , \wBMid72[3] , \wBMid72[2] , 
        \wBMid72[1] , \wBMid72[0] }), .LoOut({\wAMid73[31] , \wAMid73[30] , 
        \wAMid73[29] , \wAMid73[28] , \wAMid73[27] , \wAMid73[26] , 
        \wAMid73[25] , \wAMid73[24] , \wAMid73[23] , \wAMid73[22] , 
        \wAMid73[21] , \wAMid73[20] , \wAMid73[19] , \wAMid73[18] , 
        \wAMid73[17] , \wAMid73[16] , \wAMid73[15] , \wAMid73[14] , 
        \wAMid73[13] , \wAMid73[12] , \wAMid73[11] , \wAMid73[10] , 
        \wAMid73[9] , \wAMid73[8] , \wAMid73[7] , \wAMid73[6] , \wAMid73[5] , 
        \wAMid73[4] , \wAMid73[3] , \wAMid73[2] , \wAMid73[1] , \wAMid73[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid43[31] , \wAMid43[30] , \wAMid43[29] , \wAMid43[28] , 
        \wAMid43[27] , \wAMid43[26] , \wAMid43[25] , \wAMid43[24] , 
        \wAMid43[23] , \wAMid43[22] , \wAMid43[21] , \wAMid43[20] , 
        \wAMid43[19] , \wAMid43[18] , \wAMid43[17] , \wAMid43[16] , 
        \wAMid43[15] , \wAMid43[14] , \wAMid43[13] , \wAMid43[12] , 
        \wAMid43[11] , \wAMid43[10] , \wAMid43[9] , \wAMid43[8] , \wAMid43[7] , 
        \wAMid43[6] , \wAMid43[5] , \wAMid43[4] , \wAMid43[3] , \wAMid43[2] , 
        \wAMid43[1] , \wAMid43[0] }), .BIn({\wBMid43[31] , \wBMid43[30] , 
        \wBMid43[29] , \wBMid43[28] , \wBMid43[27] , \wBMid43[26] , 
        \wBMid43[25] , \wBMid43[24] , \wBMid43[23] , \wBMid43[22] , 
        \wBMid43[21] , \wBMid43[20] , \wBMid43[19] , \wBMid43[18] , 
        \wBMid43[17] , \wBMid43[16] , \wBMid43[15] , \wBMid43[14] , 
        \wBMid43[13] , \wBMid43[12] , \wBMid43[11] , \wBMid43[10] , 
        \wBMid43[9] , \wBMid43[8] , \wBMid43[7] , \wBMid43[6] , \wBMid43[5] , 
        \wBMid43[4] , \wBMid43[3] , \wBMid43[2] , \wBMid43[1] , \wBMid43[0] }), 
        .HiOut({\wRegInB43[31] , \wRegInB43[30] , \wRegInB43[29] , 
        \wRegInB43[28] , \wRegInB43[27] , \wRegInB43[26] , \wRegInB43[25] , 
        \wRegInB43[24] , \wRegInB43[23] , \wRegInB43[22] , \wRegInB43[21] , 
        \wRegInB43[20] , \wRegInB43[19] , \wRegInB43[18] , \wRegInB43[17] , 
        \wRegInB43[16] , \wRegInB43[15] , \wRegInB43[14] , \wRegInB43[13] , 
        \wRegInB43[12] , \wRegInB43[11] , \wRegInB43[10] , \wRegInB43[9] , 
        \wRegInB43[8] , \wRegInB43[7] , \wRegInB43[6] , \wRegInB43[5] , 
        \wRegInB43[4] , \wRegInB43[3] , \wRegInB43[2] , \wRegInB43[1] , 
        \wRegInB43[0] }), .LoOut({\wRegInA44[31] , \wRegInA44[30] , 
        \wRegInA44[29] , \wRegInA44[28] , \wRegInA44[27] , \wRegInA44[26] , 
        \wRegInA44[25] , \wRegInA44[24] , \wRegInA44[23] , \wRegInA44[22] , 
        \wRegInA44[21] , \wRegInA44[20] , \wRegInA44[19] , \wRegInA44[18] , 
        \wRegInA44[17] , \wRegInA44[16] , \wRegInA44[15] , \wRegInA44[14] , 
        \wRegInA44[13] , \wRegInA44[12] , \wRegInA44[11] , \wRegInA44[10] , 
        \wRegInA44[9] , \wRegInA44[8] , \wRegInA44[7] , \wRegInA44[6] , 
        \wRegInA44[5] , \wRegInA44[4] , \wRegInA44[3] , \wRegInA44[2] , 
        \wRegInA44[1] , \wRegInA44[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid58[31] , \wAMid58[30] , \wAMid58[29] , \wAMid58[28] , 
        \wAMid58[27] , \wAMid58[26] , \wAMid58[25] , \wAMid58[24] , 
        \wAMid58[23] , \wAMid58[22] , \wAMid58[21] , \wAMid58[20] , 
        \wAMid58[19] , \wAMid58[18] , \wAMid58[17] , \wAMid58[16] , 
        \wAMid58[15] , \wAMid58[14] , \wAMid58[13] , \wAMid58[12] , 
        \wAMid58[11] , \wAMid58[10] , \wAMid58[9] , \wAMid58[8] , \wAMid58[7] , 
        \wAMid58[6] , \wAMid58[5] , \wAMid58[4] , \wAMid58[3] , \wAMid58[2] , 
        \wAMid58[1] , \wAMid58[0] }), .BIn({\wBMid58[31] , \wBMid58[30] , 
        \wBMid58[29] , \wBMid58[28] , \wBMid58[27] , \wBMid58[26] , 
        \wBMid58[25] , \wBMid58[24] , \wBMid58[23] , \wBMid58[22] , 
        \wBMid58[21] , \wBMid58[20] , \wBMid58[19] , \wBMid58[18] , 
        \wBMid58[17] , \wBMid58[16] , \wBMid58[15] , \wBMid58[14] , 
        \wBMid58[13] , \wBMid58[12] , \wBMid58[11] , \wBMid58[10] , 
        \wBMid58[9] , \wBMid58[8] , \wBMid58[7] , \wBMid58[6] , \wBMid58[5] , 
        \wBMid58[4] , \wBMid58[3] , \wBMid58[2] , \wBMid58[1] , \wBMid58[0] }), 
        .HiOut({\wRegInB58[31] , \wRegInB58[30] , \wRegInB58[29] , 
        \wRegInB58[28] , \wRegInB58[27] , \wRegInB58[26] , \wRegInB58[25] , 
        \wRegInB58[24] , \wRegInB58[23] , \wRegInB58[22] , \wRegInB58[21] , 
        \wRegInB58[20] , \wRegInB58[19] , \wRegInB58[18] , \wRegInB58[17] , 
        \wRegInB58[16] , \wRegInB58[15] , \wRegInB58[14] , \wRegInB58[13] , 
        \wRegInB58[12] , \wRegInB58[11] , \wRegInB58[10] , \wRegInB58[9] , 
        \wRegInB58[8] , \wRegInB58[7] , \wRegInB58[6] , \wRegInB58[5] , 
        \wRegInB58[4] , \wRegInB58[3] , \wRegInB58[2] , \wRegInB58[1] , 
        \wRegInB58[0] }), .LoOut({\wRegInA59[31] , \wRegInA59[30] , 
        \wRegInA59[29] , \wRegInA59[28] , \wRegInA59[27] , \wRegInA59[26] , 
        \wRegInA59[25] , \wRegInA59[24] , \wRegInA59[23] , \wRegInA59[22] , 
        \wRegInA59[21] , \wRegInA59[20] , \wRegInA59[19] , \wRegInA59[18] , 
        \wRegInA59[17] , \wRegInA59[16] , \wRegInA59[15] , \wRegInA59[14] , 
        \wRegInA59[13] , \wRegInA59[12] , \wRegInA59[11] , \wRegInA59[10] , 
        \wRegInA59[9] , \wRegInA59[8] , \wRegInA59[7] , \wRegInA59[6] , 
        \wRegInA59[5] , \wRegInA59[4] , \wRegInA59[3] , \wRegInA59[2] , 
        \wRegInA59[1] , \wRegInA59[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_176 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink177[31] , \ScanLink177[30] , \ScanLink177[29] , 
        \ScanLink177[28] , \ScanLink177[27] , \ScanLink177[26] , 
        \ScanLink177[25] , \ScanLink177[24] , \ScanLink177[23] , 
        \ScanLink177[22] , \ScanLink177[21] , \ScanLink177[20] , 
        \ScanLink177[19] , \ScanLink177[18] , \ScanLink177[17] , 
        \ScanLink177[16] , \ScanLink177[15] , \ScanLink177[14] , 
        \ScanLink177[13] , \ScanLink177[12] , \ScanLink177[11] , 
        \ScanLink177[10] , \ScanLink177[9] , \ScanLink177[8] , 
        \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , \ScanLink177[4] , 
        \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , \ScanLink177[0] 
        }), .ScanOut({\ScanLink176[31] , \ScanLink176[30] , \ScanLink176[29] , 
        \ScanLink176[28] , \ScanLink176[27] , \ScanLink176[26] , 
        \ScanLink176[25] , \ScanLink176[24] , \ScanLink176[23] , 
        \ScanLink176[22] , \ScanLink176[21] , \ScanLink176[20] , 
        \ScanLink176[19] , \ScanLink176[18] , \ScanLink176[17] , 
        \ScanLink176[16] , \ScanLink176[15] , \ScanLink176[14] , 
        \ScanLink176[13] , \ScanLink176[12] , \ScanLink176[11] , 
        \ScanLink176[10] , \ScanLink176[9] , \ScanLink176[8] , 
        \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , \ScanLink176[4] , 
        \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , \ScanLink176[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB39[31] , \wRegInB39[30] , \wRegInB39[29] , 
        \wRegInB39[28] , \wRegInB39[27] , \wRegInB39[26] , \wRegInB39[25] , 
        \wRegInB39[24] , \wRegInB39[23] , \wRegInB39[22] , \wRegInB39[21] , 
        \wRegInB39[20] , \wRegInB39[19] , \wRegInB39[18] , \wRegInB39[17] , 
        \wRegInB39[16] , \wRegInB39[15] , \wRegInB39[14] , \wRegInB39[13] , 
        \wRegInB39[12] , \wRegInB39[11] , \wRegInB39[10] , \wRegInB39[9] , 
        \wRegInB39[8] , \wRegInB39[7] , \wRegInB39[6] , \wRegInB39[5] , 
        \wRegInB39[4] , \wRegInB39[3] , \wRegInB39[2] , \wRegInB39[1] , 
        \wRegInB39[0] }), .Out({\wBIn39[31] , \wBIn39[30] , \wBIn39[29] , 
        \wBIn39[28] , \wBIn39[27] , \wBIn39[26] , \wBIn39[25] , \wBIn39[24] , 
        \wBIn39[23] , \wBIn39[22] , \wBIn39[21] , \wBIn39[20] , \wBIn39[19] , 
        \wBIn39[18] , \wBIn39[17] , \wBIn39[16] , \wBIn39[15] , \wBIn39[14] , 
        \wBIn39[13] , \wBIn39[12] , \wBIn39[11] , \wBIn39[10] , \wBIn39[9] , 
        \wBIn39[8] , \wBIn39[7] , \wBIn39[6] , \wBIn39[5] , \wBIn39[4] , 
        \wBIn39[3] , \wBIn39[2] , \wBIn39[1] , \wBIn39[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_26 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink27[31] , \ScanLink27[30] , \ScanLink27[29] , 
        \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , \ScanLink27[25] , 
        \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , \ScanLink27[21] , 
        \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , \ScanLink27[17] , 
        \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , \ScanLink27[13] , 
        \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , \ScanLink27[9] , 
        \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , \ScanLink27[5] , 
        \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , \ScanLink27[1] , 
        \ScanLink27[0] }), .ScanOut({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB114[31] , \wRegInB114[30] , 
        \wRegInB114[29] , \wRegInB114[28] , \wRegInB114[27] , \wRegInB114[26] , 
        \wRegInB114[25] , \wRegInB114[24] , \wRegInB114[23] , \wRegInB114[22] , 
        \wRegInB114[21] , \wRegInB114[20] , \wRegInB114[19] , \wRegInB114[18] , 
        \wRegInB114[17] , \wRegInB114[16] , \wRegInB114[15] , \wRegInB114[14] , 
        \wRegInB114[13] , \wRegInB114[12] , \wRegInB114[11] , \wRegInB114[10] , 
        \wRegInB114[9] , \wRegInB114[8] , \wRegInB114[7] , \wRegInB114[6] , 
        \wRegInB114[5] , \wRegInB114[4] , \wRegInB114[3] , \wRegInB114[2] , 
        \wRegInB114[1] , \wRegInB114[0] }), .Out({\wBIn114[31] , \wBIn114[30] , 
        \wBIn114[29] , \wBIn114[28] , \wBIn114[27] , \wBIn114[26] , 
        \wBIn114[25] , \wBIn114[24] , \wBIn114[23] , \wBIn114[22] , 
        \wBIn114[21] , \wBIn114[20] , \wBIn114[19] , \wBIn114[18] , 
        \wBIn114[17] , \wBIn114[16] , \wBIn114[15] , \wBIn114[14] , 
        \wBIn114[13] , \wBIn114[12] , \wBIn114[11] , \wBIn114[10] , 
        \wBIn114[9] , \wBIn114[8] , \wBIn114[7] , \wBIn114[6] , \wBIn114[5] , 
        \wBIn114[4] , \wBIn114[3] , \wBIn114[2] , \wBIn114[1] , \wBIn114[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn103[31] , \wAIn103[30] , \wAIn103[29] , \wAIn103[28] , 
        \wAIn103[27] , \wAIn103[26] , \wAIn103[25] , \wAIn103[24] , 
        \wAIn103[23] , \wAIn103[22] , \wAIn103[21] , \wAIn103[20] , 
        \wAIn103[19] , \wAIn103[18] , \wAIn103[17] , \wAIn103[16] , 
        \wAIn103[15] , \wAIn103[14] , \wAIn103[13] , \wAIn103[12] , 
        \wAIn103[11] , \wAIn103[10] , \wAIn103[9] , \wAIn103[8] , \wAIn103[7] , 
        \wAIn103[6] , \wAIn103[5] , \wAIn103[4] , \wAIn103[3] , \wAIn103[2] , 
        \wAIn103[1] , \wAIn103[0] }), .BIn({\wBIn103[31] , \wBIn103[30] , 
        \wBIn103[29] , \wBIn103[28] , \wBIn103[27] , \wBIn103[26] , 
        \wBIn103[25] , \wBIn103[24] , \wBIn103[23] , \wBIn103[22] , 
        \wBIn103[21] , \wBIn103[20] , \wBIn103[19] , \wBIn103[18] , 
        \wBIn103[17] , \wBIn103[16] , \wBIn103[15] , \wBIn103[14] , 
        \wBIn103[13] , \wBIn103[12] , \wBIn103[11] , \wBIn103[10] , 
        \wBIn103[9] , \wBIn103[8] , \wBIn103[7] , \wBIn103[6] , \wBIn103[5] , 
        \wBIn103[4] , \wBIn103[3] , \wBIn103[2] , \wBIn103[1] , \wBIn103[0] }), 
        .HiOut({\wBMid102[31] , \wBMid102[30] , \wBMid102[29] , \wBMid102[28] , 
        \wBMid102[27] , \wBMid102[26] , \wBMid102[25] , \wBMid102[24] , 
        \wBMid102[23] , \wBMid102[22] , \wBMid102[21] , \wBMid102[20] , 
        \wBMid102[19] , \wBMid102[18] , \wBMid102[17] , \wBMid102[16] , 
        \wBMid102[15] , \wBMid102[14] , \wBMid102[13] , \wBMid102[12] , 
        \wBMid102[11] , \wBMid102[10] , \wBMid102[9] , \wBMid102[8] , 
        \wBMid102[7] , \wBMid102[6] , \wBMid102[5] , \wBMid102[4] , 
        \wBMid102[3] , \wBMid102[2] , \wBMid102[1] , \wBMid102[0] }), .LoOut({
        \wAMid103[31] , \wAMid103[30] , \wAMid103[29] , \wAMid103[28] , 
        \wAMid103[27] , \wAMid103[26] , \wAMid103[25] , \wAMid103[24] , 
        \wAMid103[23] , \wAMid103[22] , \wAMid103[21] , \wAMid103[20] , 
        \wAMid103[19] , \wAMid103[18] , \wAMid103[17] , \wAMid103[16] , 
        \wAMid103[15] , \wAMid103[14] , \wAMid103[13] , \wAMid103[12] , 
        \wAMid103[11] , \wAMid103[10] , \wAMid103[9] , \wAMid103[8] , 
        \wAMid103[7] , \wAMid103[6] , \wAMid103[5] , \wAMid103[4] , 
        \wAMid103[3] , \wAMid103[2] , \wAMid103[1] , \wAMid103[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_246 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink247[31] , \ScanLink247[30] , \ScanLink247[29] , 
        \ScanLink247[28] , \ScanLink247[27] , \ScanLink247[26] , 
        \ScanLink247[25] , \ScanLink247[24] , \ScanLink247[23] , 
        \ScanLink247[22] , \ScanLink247[21] , \ScanLink247[20] , 
        \ScanLink247[19] , \ScanLink247[18] , \ScanLink247[17] , 
        \ScanLink247[16] , \ScanLink247[15] , \ScanLink247[14] , 
        \ScanLink247[13] , \ScanLink247[12] , \ScanLink247[11] , 
        \ScanLink247[10] , \ScanLink247[9] , \ScanLink247[8] , 
        \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , \ScanLink247[4] , 
        \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , \ScanLink247[0] 
        }), .ScanOut({\ScanLink246[31] , \ScanLink246[30] , \ScanLink246[29] , 
        \ScanLink246[28] , \ScanLink246[27] , \ScanLink246[26] , 
        \ScanLink246[25] , \ScanLink246[24] , \ScanLink246[23] , 
        \ScanLink246[22] , \ScanLink246[21] , \ScanLink246[20] , 
        \ScanLink246[19] , \ScanLink246[18] , \ScanLink246[17] , 
        \ScanLink246[16] , \ScanLink246[15] , \ScanLink246[14] , 
        \ScanLink246[13] , \ScanLink246[12] , \ScanLink246[11] , 
        \ScanLink246[10] , \ScanLink246[9] , \ScanLink246[8] , 
        \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , \ScanLink246[4] , 
        \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , \ScanLink246[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB4[31] , \wRegInB4[30] , \wRegInB4[29] , \wRegInB4[28] , 
        \wRegInB4[27] , \wRegInB4[26] , \wRegInB4[25] , \wRegInB4[24] , 
        \wRegInB4[23] , \wRegInB4[22] , \wRegInB4[21] , \wRegInB4[20] , 
        \wRegInB4[19] , \wRegInB4[18] , \wRegInB4[17] , \wRegInB4[16] , 
        \wRegInB4[15] , \wRegInB4[14] , \wRegInB4[13] , \wRegInB4[12] , 
        \wRegInB4[11] , \wRegInB4[10] , \wRegInB4[9] , \wRegInB4[8] , 
        \wRegInB4[7] , \wRegInB4[6] , \wRegInB4[5] , \wRegInB4[4] , 
        \wRegInB4[3] , \wRegInB4[2] , \wRegInB4[1] , \wRegInB4[0] }), .Out({
        \wBIn4[31] , \wBIn4[30] , \wBIn4[29] , \wBIn4[28] , \wBIn4[27] , 
        \wBIn4[26] , \wBIn4[25] , \wBIn4[24] , \wBIn4[23] , \wBIn4[22] , 
        \wBIn4[21] , \wBIn4[20] , \wBIn4[19] , \wBIn4[18] , \wBIn4[17] , 
        \wBIn4[16] , \wBIn4[15] , \wBIn4[14] , \wBIn4[13] , \wBIn4[12] , 
        \wBIn4[11] , \wBIn4[10] , \wBIn4[9] , \wBIn4[8] , \wBIn4[7] , 
        \wBIn4[6] , \wBIn4[5] , \wBIn4[4] , \wBIn4[3] , \wBIn4[2] , \wBIn4[1] , 
        \wBIn4[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn124[31] , \wAIn124[30] , \wAIn124[29] , \wAIn124[28] , 
        \wAIn124[27] , \wAIn124[26] , \wAIn124[25] , \wAIn124[24] , 
        \wAIn124[23] , \wAIn124[22] , \wAIn124[21] , \wAIn124[20] , 
        \wAIn124[19] , \wAIn124[18] , \wAIn124[17] , \wAIn124[16] , 
        \wAIn124[15] , \wAIn124[14] , \wAIn124[13] , \wAIn124[12] , 
        \wAIn124[11] , \wAIn124[10] , \wAIn124[9] , \wAIn124[8] , \wAIn124[7] , 
        \wAIn124[6] , \wAIn124[5] , \wAIn124[4] , \wAIn124[3] , \wAIn124[2] , 
        \wAIn124[1] , \wAIn124[0] }), .BIn({\wBIn124[31] , \wBIn124[30] , 
        \wBIn124[29] , \wBIn124[28] , \wBIn124[27] , \wBIn124[26] , 
        \wBIn124[25] , \wBIn124[24] , \wBIn124[23] , \wBIn124[22] , 
        \wBIn124[21] , \wBIn124[20] , \wBIn124[19] , \wBIn124[18] , 
        \wBIn124[17] , \wBIn124[16] , \wBIn124[15] , \wBIn124[14] , 
        \wBIn124[13] , \wBIn124[12] , \wBIn124[11] , \wBIn124[10] , 
        \wBIn124[9] , \wBIn124[8] , \wBIn124[7] , \wBIn124[6] , \wBIn124[5] , 
        \wBIn124[4] , \wBIn124[3] , \wBIn124[2] , \wBIn124[1] , \wBIn124[0] }), 
        .HiOut({\wBMid123[31] , \wBMid123[30] , \wBMid123[29] , \wBMid123[28] , 
        \wBMid123[27] , \wBMid123[26] , \wBMid123[25] , \wBMid123[24] , 
        \wBMid123[23] , \wBMid123[22] , \wBMid123[21] , \wBMid123[20] , 
        \wBMid123[19] , \wBMid123[18] , \wBMid123[17] , \wBMid123[16] , 
        \wBMid123[15] , \wBMid123[14] , \wBMid123[13] , \wBMid123[12] , 
        \wBMid123[11] , \wBMid123[10] , \wBMid123[9] , \wBMid123[8] , 
        \wBMid123[7] , \wBMid123[6] , \wBMid123[5] , \wBMid123[4] , 
        \wBMid123[3] , \wBMid123[2] , \wBMid123[1] , \wBMid123[0] }), .LoOut({
        \wAMid124[31] , \wAMid124[30] , \wAMid124[29] , \wAMid124[28] , 
        \wAMid124[27] , \wAMid124[26] , \wAMid124[25] , \wAMid124[24] , 
        \wAMid124[23] , \wAMid124[22] , \wAMid124[21] , \wAMid124[20] , 
        \wAMid124[19] , \wAMid124[18] , \wAMid124[17] , \wAMid124[16] , 
        \wAMid124[15] , \wAMid124[14] , \wAMid124[13] , \wAMid124[12] , 
        \wAMid124[11] , \wAMid124[10] , \wAMid124[9] , \wAMid124[8] , 
        \wAMid124[7] , \wAMid124[6] , \wAMid124[5] , \wAMid124[4] , 
        \wAMid124[3] , \wAMid124[2] , \wAMid124[1] , \wAMid124[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid64[31] , \wAMid64[30] , \wAMid64[29] , \wAMid64[28] , 
        \wAMid64[27] , \wAMid64[26] , \wAMid64[25] , \wAMid64[24] , 
        \wAMid64[23] , \wAMid64[22] , \wAMid64[21] , \wAMid64[20] , 
        \wAMid64[19] , \wAMid64[18] , \wAMid64[17] , \wAMid64[16] , 
        \wAMid64[15] , \wAMid64[14] , \wAMid64[13] , \wAMid64[12] , 
        \wAMid64[11] , \wAMid64[10] , \wAMid64[9] , \wAMid64[8] , \wAMid64[7] , 
        \wAMid64[6] , \wAMid64[5] , \wAMid64[4] , \wAMid64[3] , \wAMid64[2] , 
        \wAMid64[1] , \wAMid64[0] }), .BIn({\wBMid64[31] , \wBMid64[30] , 
        \wBMid64[29] , \wBMid64[28] , \wBMid64[27] , \wBMid64[26] , 
        \wBMid64[25] , \wBMid64[24] , \wBMid64[23] , \wBMid64[22] , 
        \wBMid64[21] , \wBMid64[20] , \wBMid64[19] , \wBMid64[18] , 
        \wBMid64[17] , \wBMid64[16] , \wBMid64[15] , \wBMid64[14] , 
        \wBMid64[13] , \wBMid64[12] , \wBMid64[11] , \wBMid64[10] , 
        \wBMid64[9] , \wBMid64[8] , \wBMid64[7] , \wBMid64[6] , \wBMid64[5] , 
        \wBMid64[4] , \wBMid64[3] , \wBMid64[2] , \wBMid64[1] , \wBMid64[0] }), 
        .HiOut({\wRegInB64[31] , \wRegInB64[30] , \wRegInB64[29] , 
        \wRegInB64[28] , \wRegInB64[27] , \wRegInB64[26] , \wRegInB64[25] , 
        \wRegInB64[24] , \wRegInB64[23] , \wRegInB64[22] , \wRegInB64[21] , 
        \wRegInB64[20] , \wRegInB64[19] , \wRegInB64[18] , \wRegInB64[17] , 
        \wRegInB64[16] , \wRegInB64[15] , \wRegInB64[14] , \wRegInB64[13] , 
        \wRegInB64[12] , \wRegInB64[11] , \wRegInB64[10] , \wRegInB64[9] , 
        \wRegInB64[8] , \wRegInB64[7] , \wRegInB64[6] , \wRegInB64[5] , 
        \wRegInB64[4] , \wRegInB64[3] , \wRegInB64[2] , \wRegInB64[1] , 
        \wRegInB64[0] }), .LoOut({\wRegInA65[31] , \wRegInA65[30] , 
        \wRegInA65[29] , \wRegInA65[28] , \wRegInA65[27] , \wRegInA65[26] , 
        \wRegInA65[25] , \wRegInA65[24] , \wRegInA65[23] , \wRegInA65[22] , 
        \wRegInA65[21] , \wRegInA65[20] , \wRegInA65[19] , \wRegInA65[18] , 
        \wRegInA65[17] , \wRegInA65[16] , \wRegInA65[15] , \wRegInA65[14] , 
        \wRegInA65[13] , \wRegInA65[12] , \wRegInA65[11] , \wRegInA65[10] , 
        \wRegInA65[9] , \wRegInA65[8] , \wRegInA65[7] , \wRegInA65[6] , 
        \wRegInA65[5] , \wRegInA65[4] , \wRegInA65[3] , \wRegInA65[2] , 
        \wRegInA65[1] , \wRegInA65[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_151 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink152[31] , \ScanLink152[30] , \ScanLink152[29] , 
        \ScanLink152[28] , \ScanLink152[27] , \ScanLink152[26] , 
        \ScanLink152[25] , \ScanLink152[24] , \ScanLink152[23] , 
        \ScanLink152[22] , \ScanLink152[21] , \ScanLink152[20] , 
        \ScanLink152[19] , \ScanLink152[18] , \ScanLink152[17] , 
        \ScanLink152[16] , \ScanLink152[15] , \ScanLink152[14] , 
        \ScanLink152[13] , \ScanLink152[12] , \ScanLink152[11] , 
        \ScanLink152[10] , \ScanLink152[9] , \ScanLink152[8] , 
        \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , \ScanLink152[4] , 
        \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , \ScanLink152[0] 
        }), .ScanOut({\ScanLink151[31] , \ScanLink151[30] , \ScanLink151[29] , 
        \ScanLink151[28] , \ScanLink151[27] , \ScanLink151[26] , 
        \ScanLink151[25] , \ScanLink151[24] , \ScanLink151[23] , 
        \ScanLink151[22] , \ScanLink151[21] , \ScanLink151[20] , 
        \ScanLink151[19] , \ScanLink151[18] , \ScanLink151[17] , 
        \ScanLink151[16] , \ScanLink151[15] , \ScanLink151[14] , 
        \ScanLink151[13] , \ScanLink151[12] , \ScanLink151[11] , 
        \ScanLink151[10] , \ScanLink151[9] , \ScanLink151[8] , 
        \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , \ScanLink151[4] , 
        \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , \ScanLink151[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA52[31] , \wRegInA52[30] , \wRegInA52[29] , 
        \wRegInA52[28] , \wRegInA52[27] , \wRegInA52[26] , \wRegInA52[25] , 
        \wRegInA52[24] , \wRegInA52[23] , \wRegInA52[22] , \wRegInA52[21] , 
        \wRegInA52[20] , \wRegInA52[19] , \wRegInA52[18] , \wRegInA52[17] , 
        \wRegInA52[16] , \wRegInA52[15] , \wRegInA52[14] , \wRegInA52[13] , 
        \wRegInA52[12] , \wRegInA52[11] , \wRegInA52[10] , \wRegInA52[9] , 
        \wRegInA52[8] , \wRegInA52[7] , \wRegInA52[6] , \wRegInA52[5] , 
        \wRegInA52[4] , \wRegInA52[3] , \wRegInA52[2] , \wRegInA52[1] , 
        \wRegInA52[0] }), .Out({\wAIn52[31] , \wAIn52[30] , \wAIn52[29] , 
        \wAIn52[28] , \wAIn52[27] , \wAIn52[26] , \wAIn52[25] , \wAIn52[24] , 
        \wAIn52[23] , \wAIn52[22] , \wAIn52[21] , \wAIn52[20] , \wAIn52[19] , 
        \wAIn52[18] , \wAIn52[17] , \wAIn52[16] , \wAIn52[15] , \wAIn52[14] , 
        \wAIn52[13] , \wAIn52[12] , \wAIn52[11] , \wAIn52[10] , \wAIn52[9] , 
        \wAIn52[8] , \wAIn52[7] , \wAIn52[6] , \wAIn52[5] , \wAIn52[4] , 
        \wAIn52[3] , \wAIn52[2] , \wAIn52[1] , \wAIn52[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn96[31] , \wAIn96[30] , \wAIn96[29] , \wAIn96[28] , \wAIn96[27] , 
        \wAIn96[26] , \wAIn96[25] , \wAIn96[24] , \wAIn96[23] , \wAIn96[22] , 
        \wAIn96[21] , \wAIn96[20] , \wAIn96[19] , \wAIn96[18] , \wAIn96[17] , 
        \wAIn96[16] , \wAIn96[15] , \wAIn96[14] , \wAIn96[13] , \wAIn96[12] , 
        \wAIn96[11] , \wAIn96[10] , \wAIn96[9] , \wAIn96[8] , \wAIn96[7] , 
        \wAIn96[6] , \wAIn96[5] , \wAIn96[4] , \wAIn96[3] , \wAIn96[2] , 
        \wAIn96[1] , \wAIn96[0] }), .BIn({\wBIn96[31] , \wBIn96[30] , 
        \wBIn96[29] , \wBIn96[28] , \wBIn96[27] , \wBIn96[26] , \wBIn96[25] , 
        \wBIn96[24] , \wBIn96[23] , \wBIn96[22] , \wBIn96[21] , \wBIn96[20] , 
        \wBIn96[19] , \wBIn96[18] , \wBIn96[17] , \wBIn96[16] , \wBIn96[15] , 
        \wBIn96[14] , \wBIn96[13] , \wBIn96[12] , \wBIn96[11] , \wBIn96[10] , 
        \wBIn96[9] , \wBIn96[8] , \wBIn96[7] , \wBIn96[6] , \wBIn96[5] , 
        \wBIn96[4] , \wBIn96[3] , \wBIn96[2] , \wBIn96[1] , \wBIn96[0] }), 
        .HiOut({\wBMid95[31] , \wBMid95[30] , \wBMid95[29] , \wBMid95[28] , 
        \wBMid95[27] , \wBMid95[26] , \wBMid95[25] , \wBMid95[24] , 
        \wBMid95[23] , \wBMid95[22] , \wBMid95[21] , \wBMid95[20] , 
        \wBMid95[19] , \wBMid95[18] , \wBMid95[17] , \wBMid95[16] , 
        \wBMid95[15] , \wBMid95[14] , \wBMid95[13] , \wBMid95[12] , 
        \wBMid95[11] , \wBMid95[10] , \wBMid95[9] , \wBMid95[8] , \wBMid95[7] , 
        \wBMid95[6] , \wBMid95[5] , \wBMid95[4] , \wBMid95[3] , \wBMid95[2] , 
        \wBMid95[1] , \wBMid95[0] }), .LoOut({\wAMid96[31] , \wAMid96[30] , 
        \wAMid96[29] , \wAMid96[28] , \wAMid96[27] , \wAMid96[26] , 
        \wAMid96[25] , \wAMid96[24] , \wAMid96[23] , \wAMid96[22] , 
        \wAMid96[21] , \wAMid96[20] , \wAMid96[19] , \wAMid96[18] , 
        \wAMid96[17] , \wAMid96[16] , \wAMid96[15] , \wAMid96[14] , 
        \wAMid96[13] , \wAMid96[12] , \wAMid96[11] , \wAMid96[10] , 
        \wAMid96[9] , \wAMid96[8] , \wAMid96[7] , \wAMid96[6] , \wAMid96[5] , 
        \wAMid96[4] , \wAMid96[3] , \wAMid96[2] , \wAMid96[1] , \wAMid96[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid81[31] , \wAMid81[30] , \wAMid81[29] , \wAMid81[28] , 
        \wAMid81[27] , \wAMid81[26] , \wAMid81[25] , \wAMid81[24] , 
        \wAMid81[23] , \wAMid81[22] , \wAMid81[21] , \wAMid81[20] , 
        \wAMid81[19] , \wAMid81[18] , \wAMid81[17] , \wAMid81[16] , 
        \wAMid81[15] , \wAMid81[14] , \wAMid81[13] , \wAMid81[12] , 
        \wAMid81[11] , \wAMid81[10] , \wAMid81[9] , \wAMid81[8] , \wAMid81[7] , 
        \wAMid81[6] , \wAMid81[5] , \wAMid81[4] , \wAMid81[3] , \wAMid81[2] , 
        \wAMid81[1] , \wAMid81[0] }), .BIn({\wBMid81[31] , \wBMid81[30] , 
        \wBMid81[29] , \wBMid81[28] , \wBMid81[27] , \wBMid81[26] , 
        \wBMid81[25] , \wBMid81[24] , \wBMid81[23] , \wBMid81[22] , 
        \wBMid81[21] , \wBMid81[20] , \wBMid81[19] , \wBMid81[18] , 
        \wBMid81[17] , \wBMid81[16] , \wBMid81[15] , \wBMid81[14] , 
        \wBMid81[13] , \wBMid81[12] , \wBMid81[11] , \wBMid81[10] , 
        \wBMid81[9] , \wBMid81[8] , \wBMid81[7] , \wBMid81[6] , \wBMid81[5] , 
        \wBMid81[4] , \wBMid81[3] , \wBMid81[2] , \wBMid81[1] , \wBMid81[0] }), 
        .HiOut({\wRegInB81[31] , \wRegInB81[30] , \wRegInB81[29] , 
        \wRegInB81[28] , \wRegInB81[27] , \wRegInB81[26] , \wRegInB81[25] , 
        \wRegInB81[24] , \wRegInB81[23] , \wRegInB81[22] , \wRegInB81[21] , 
        \wRegInB81[20] , \wRegInB81[19] , \wRegInB81[18] , \wRegInB81[17] , 
        \wRegInB81[16] , \wRegInB81[15] , \wRegInB81[14] , \wRegInB81[13] , 
        \wRegInB81[12] , \wRegInB81[11] , \wRegInB81[10] , \wRegInB81[9] , 
        \wRegInB81[8] , \wRegInB81[7] , \wRegInB81[6] , \wRegInB81[5] , 
        \wRegInB81[4] , \wRegInB81[3] , \wRegInB81[2] , \wRegInB81[1] , 
        \wRegInB81[0] }), .LoOut({\wRegInA82[31] , \wRegInA82[30] , 
        \wRegInA82[29] , \wRegInA82[28] , \wRegInA82[27] , \wRegInA82[26] , 
        \wRegInA82[25] , \wRegInA82[24] , \wRegInA82[23] , \wRegInA82[22] , 
        \wRegInA82[21] , \wRegInA82[20] , \wRegInA82[19] , \wRegInA82[18] , 
        \wRegInA82[17] , \wRegInA82[16] , \wRegInA82[15] , \wRegInA82[14] , 
        \wRegInA82[13] , \wRegInA82[12] , \wRegInA82[11] , \wRegInA82[10] , 
        \wRegInA82[9] , \wRegInA82[8] , \wRegInA82[7] , \wRegInA82[6] , 
        \wRegInA82[5] , \wRegInA82[4] , \wRegInA82[3] , \wRegInA82[2] , 
        \wRegInA82[1] , \wRegInA82[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid109[31] , \wAMid109[30] , \wAMid109[29] , \wAMid109[28] , 
        \wAMid109[27] , \wAMid109[26] , \wAMid109[25] , \wAMid109[24] , 
        \wAMid109[23] , \wAMid109[22] , \wAMid109[21] , \wAMid109[20] , 
        \wAMid109[19] , \wAMid109[18] , \wAMid109[17] , \wAMid109[16] , 
        \wAMid109[15] , \wAMid109[14] , \wAMid109[13] , \wAMid109[12] , 
        \wAMid109[11] , \wAMid109[10] , \wAMid109[9] , \wAMid109[8] , 
        \wAMid109[7] , \wAMid109[6] , \wAMid109[5] , \wAMid109[4] , 
        \wAMid109[3] , \wAMid109[2] , \wAMid109[1] , \wAMid109[0] }), .BIn({
        \wBMid109[31] , \wBMid109[30] , \wBMid109[29] , \wBMid109[28] , 
        \wBMid109[27] , \wBMid109[26] , \wBMid109[25] , \wBMid109[24] , 
        \wBMid109[23] , \wBMid109[22] , \wBMid109[21] , \wBMid109[20] , 
        \wBMid109[19] , \wBMid109[18] , \wBMid109[17] , \wBMid109[16] , 
        \wBMid109[15] , \wBMid109[14] , \wBMid109[13] , \wBMid109[12] , 
        \wBMid109[11] , \wBMid109[10] , \wBMid109[9] , \wBMid109[8] , 
        \wBMid109[7] , \wBMid109[6] , \wBMid109[5] , \wBMid109[4] , 
        \wBMid109[3] , \wBMid109[2] , \wBMid109[1] , \wBMid109[0] }), .HiOut({
        \wRegInB109[31] , \wRegInB109[30] , \wRegInB109[29] , \wRegInB109[28] , 
        \wRegInB109[27] , \wRegInB109[26] , \wRegInB109[25] , \wRegInB109[24] , 
        \wRegInB109[23] , \wRegInB109[22] , \wRegInB109[21] , \wRegInB109[20] , 
        \wRegInB109[19] , \wRegInB109[18] , \wRegInB109[17] , \wRegInB109[16] , 
        \wRegInB109[15] , \wRegInB109[14] , \wRegInB109[13] , \wRegInB109[12] , 
        \wRegInB109[11] , \wRegInB109[10] , \wRegInB109[9] , \wRegInB109[8] , 
        \wRegInB109[7] , \wRegInB109[6] , \wRegInB109[5] , \wRegInB109[4] , 
        \wRegInB109[3] , \wRegInB109[2] , \wRegInB109[1] , \wRegInB109[0] }), 
        .LoOut({\wRegInA110[31] , \wRegInA110[30] , \wRegInA110[29] , 
        \wRegInA110[28] , \wRegInA110[27] , \wRegInA110[26] , \wRegInA110[25] , 
        \wRegInA110[24] , \wRegInA110[23] , \wRegInA110[22] , \wRegInA110[21] , 
        \wRegInA110[20] , \wRegInA110[19] , \wRegInA110[18] , \wRegInA110[17] , 
        \wRegInA110[16] , \wRegInA110[15] , \wRegInA110[14] , \wRegInA110[13] , 
        \wRegInA110[12] , \wRegInA110[11] , \wRegInA110[10] , \wRegInA110[9] , 
        \wRegInA110[8] , \wRegInA110[7] , \wRegInA110[6] , \wRegInA110[5] , 
        \wRegInA110[4] , \wRegInA110[3] , \wRegInA110[2] , \wRegInA110[1] , 
        \wRegInA110[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid7[31] , 
        \wAMid7[30] , \wAMid7[29] , \wAMid7[28] , \wAMid7[27] , \wAMid7[26] , 
        \wAMid7[25] , \wAMid7[24] , \wAMid7[23] , \wAMid7[22] , \wAMid7[21] , 
        \wAMid7[20] , \wAMid7[19] , \wAMid7[18] , \wAMid7[17] , \wAMid7[16] , 
        \wAMid7[15] , \wAMid7[14] , \wAMid7[13] , \wAMid7[12] , \wAMid7[11] , 
        \wAMid7[10] , \wAMid7[9] , \wAMid7[8] , \wAMid7[7] , \wAMid7[6] , 
        \wAMid7[5] , \wAMid7[4] , \wAMid7[3] , \wAMid7[2] , \wAMid7[1] , 
        \wAMid7[0] }), .BIn({\wBMid7[31] , \wBMid7[30] , \wBMid7[29] , 
        \wBMid7[28] , \wBMid7[27] , \wBMid7[26] , \wBMid7[25] , \wBMid7[24] , 
        \wBMid7[23] , \wBMid7[22] , \wBMid7[21] , \wBMid7[20] , \wBMid7[19] , 
        \wBMid7[18] , \wBMid7[17] , \wBMid7[16] , \wBMid7[15] , \wBMid7[14] , 
        \wBMid7[13] , \wBMid7[12] , \wBMid7[11] , \wBMid7[10] , \wBMid7[9] , 
        \wBMid7[8] , \wBMid7[7] , \wBMid7[6] , \wBMid7[5] , \wBMid7[4] , 
        \wBMid7[3] , \wBMid7[2] , \wBMid7[1] , \wBMid7[0] }), .HiOut({
        \wRegInB7[31] , \wRegInB7[30] , \wRegInB7[29] , \wRegInB7[28] , 
        \wRegInB7[27] , \wRegInB7[26] , \wRegInB7[25] , \wRegInB7[24] , 
        \wRegInB7[23] , \wRegInB7[22] , \wRegInB7[21] , \wRegInB7[20] , 
        \wRegInB7[19] , \wRegInB7[18] , \wRegInB7[17] , \wRegInB7[16] , 
        \wRegInB7[15] , \wRegInB7[14] , \wRegInB7[13] , \wRegInB7[12] , 
        \wRegInB7[11] , \wRegInB7[10] , \wRegInB7[9] , \wRegInB7[8] , 
        \wRegInB7[7] , \wRegInB7[6] , \wRegInB7[5] , \wRegInB7[4] , 
        \wRegInB7[3] , \wRegInB7[2] , \wRegInB7[1] , \wRegInB7[0] }), .LoOut({
        \wRegInA8[31] , \wRegInA8[30] , \wRegInA8[29] , \wRegInA8[28] , 
        \wRegInA8[27] , \wRegInA8[26] , \wRegInA8[25] , \wRegInA8[24] , 
        \wRegInA8[23] , \wRegInA8[22] , \wRegInA8[21] , \wRegInA8[20] , 
        \wRegInA8[19] , \wRegInA8[18] , \wRegInA8[17] , \wRegInA8[16] , 
        \wRegInA8[15] , \wRegInA8[14] , \wRegInA8[13] , \wRegInA8[12] , 
        \wRegInA8[11] , \wRegInA8[10] , \wRegInA8[9] , \wRegInA8[8] , 
        \wRegInA8[7] , \wRegInA8[6] , \wRegInA8[5] , \wRegInA8[4] , 
        \wRegInA8[3] , \wRegInA8[2] , \wRegInA8[1] , \wRegInA8[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_193 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink194[31] , \ScanLink194[30] , \ScanLink194[29] , 
        \ScanLink194[28] , \ScanLink194[27] , \ScanLink194[26] , 
        \ScanLink194[25] , \ScanLink194[24] , \ScanLink194[23] , 
        \ScanLink194[22] , \ScanLink194[21] , \ScanLink194[20] , 
        \ScanLink194[19] , \ScanLink194[18] , \ScanLink194[17] , 
        \ScanLink194[16] , \ScanLink194[15] , \ScanLink194[14] , 
        \ScanLink194[13] , \ScanLink194[12] , \ScanLink194[11] , 
        \ScanLink194[10] , \ScanLink194[9] , \ScanLink194[8] , 
        \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , \ScanLink194[4] , 
        \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , \ScanLink194[0] 
        }), .ScanOut({\ScanLink193[31] , \ScanLink193[30] , \ScanLink193[29] , 
        \ScanLink193[28] , \ScanLink193[27] , \ScanLink193[26] , 
        \ScanLink193[25] , \ScanLink193[24] , \ScanLink193[23] , 
        \ScanLink193[22] , \ScanLink193[21] , \ScanLink193[20] , 
        \ScanLink193[19] , \ScanLink193[18] , \ScanLink193[17] , 
        \ScanLink193[16] , \ScanLink193[15] , \ScanLink193[14] , 
        \ScanLink193[13] , \ScanLink193[12] , \ScanLink193[11] , 
        \ScanLink193[10] , \ScanLink193[9] , \ScanLink193[8] , 
        \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , \ScanLink193[4] , 
        \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , \ScanLink193[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA31[31] , \wRegInA31[30] , \wRegInA31[29] , 
        \wRegInA31[28] , \wRegInA31[27] , \wRegInA31[26] , \wRegInA31[25] , 
        \wRegInA31[24] , \wRegInA31[23] , \wRegInA31[22] , \wRegInA31[21] , 
        \wRegInA31[20] , \wRegInA31[19] , \wRegInA31[18] , \wRegInA31[17] , 
        \wRegInA31[16] , \wRegInA31[15] , \wRegInA31[14] , \wRegInA31[13] , 
        \wRegInA31[12] , \wRegInA31[11] , \wRegInA31[10] , \wRegInA31[9] , 
        \wRegInA31[8] , \wRegInA31[7] , \wRegInA31[6] , \wRegInA31[5] , 
        \wRegInA31[4] , \wRegInA31[3] , \wRegInA31[2] , \wRegInA31[1] , 
        \wRegInA31[0] }), .Out({\wAIn31[31] , \wAIn31[30] , \wAIn31[29] , 
        \wAIn31[28] , \wAIn31[27] , \wAIn31[26] , \wAIn31[25] , \wAIn31[24] , 
        \wAIn31[23] , \wAIn31[22] , \wAIn31[21] , \wAIn31[20] , \wAIn31[19] , 
        \wAIn31[18] , \wAIn31[17] , \wAIn31[16] , \wAIn31[15] , \wAIn31[14] , 
        \wAIn31[13] , \wAIn31[12] , \wAIn31[11] , \wAIn31[10] , \wAIn31[9] , 
        \wAIn31[8] , \wAIn31[7] , \wAIn31[6] , \wAIn31[5] , \wAIn31[4] , 
        \wAIn31[3] , \wAIn31[2] , \wAIn31[1] , \wAIn31[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid18[31] , \wAMid18[30] , \wAMid18[29] , \wAMid18[28] , 
        \wAMid18[27] , \wAMid18[26] , \wAMid18[25] , \wAMid18[24] , 
        \wAMid18[23] , \wAMid18[22] , \wAMid18[21] , \wAMid18[20] , 
        \wAMid18[19] , \wAMid18[18] , \wAMid18[17] , \wAMid18[16] , 
        \wAMid18[15] , \wAMid18[14] , \wAMid18[13] , \wAMid18[12] , 
        \wAMid18[11] , \wAMid18[10] , \wAMid18[9] , \wAMid18[8] , \wAMid18[7] , 
        \wAMid18[6] , \wAMid18[5] , \wAMid18[4] , \wAMid18[3] , \wAMid18[2] , 
        \wAMid18[1] , \wAMid18[0] }), .BIn({\wBMid18[31] , \wBMid18[30] , 
        \wBMid18[29] , \wBMid18[28] , \wBMid18[27] , \wBMid18[26] , 
        \wBMid18[25] , \wBMid18[24] , \wBMid18[23] , \wBMid18[22] , 
        \wBMid18[21] , \wBMid18[20] , \wBMid18[19] , \wBMid18[18] , 
        \wBMid18[17] , \wBMid18[16] , \wBMid18[15] , \wBMid18[14] , 
        \wBMid18[13] , \wBMid18[12] , \wBMid18[11] , \wBMid18[10] , 
        \wBMid18[9] , \wBMid18[8] , \wBMid18[7] , \wBMid18[6] , \wBMid18[5] , 
        \wBMid18[4] , \wBMid18[3] , \wBMid18[2] , \wBMid18[1] , \wBMid18[0] }), 
        .HiOut({\wRegInB18[31] , \wRegInB18[30] , \wRegInB18[29] , 
        \wRegInB18[28] , \wRegInB18[27] , \wRegInB18[26] , \wRegInB18[25] , 
        \wRegInB18[24] , \wRegInB18[23] , \wRegInB18[22] , \wRegInB18[21] , 
        \wRegInB18[20] , \wRegInB18[19] , \wRegInB18[18] , \wRegInB18[17] , 
        \wRegInB18[16] , \wRegInB18[15] , \wRegInB18[14] , \wRegInB18[13] , 
        \wRegInB18[12] , \wRegInB18[11] , \wRegInB18[10] , \wRegInB18[9] , 
        \wRegInB18[8] , \wRegInB18[7] , \wRegInB18[6] , \wRegInB18[5] , 
        \wRegInB18[4] , \wRegInB18[3] , \wRegInB18[2] , \wRegInB18[1] , 
        \wRegInB18[0] }), .LoOut({\wRegInA19[31] , \wRegInA19[30] , 
        \wRegInA19[29] , \wRegInA19[28] , \wRegInA19[27] , \wRegInA19[26] , 
        \wRegInA19[25] , \wRegInA19[24] , \wRegInA19[23] , \wRegInA19[22] , 
        \wRegInA19[21] , \wRegInA19[20] , \wRegInA19[19] , \wRegInA19[18] , 
        \wRegInA19[17] , \wRegInA19[16] , \wRegInA19[15] , \wRegInA19[14] , 
        \wRegInA19[13] , \wRegInA19[12] , \wRegInA19[11] , \wRegInA19[10] , 
        \wRegInA19[9] , \wRegInA19[8] , \wRegInA19[7] , \wRegInA19[6] , 
        \wRegInA19[5] , \wRegInA19[4] , \wRegInA19[3] , \wRegInA19[2] , 
        \wRegInA19[1] , \wRegInA19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_228 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink229[31] , \ScanLink229[30] , \ScanLink229[29] , 
        \ScanLink229[28] , \ScanLink229[27] , \ScanLink229[26] , 
        \ScanLink229[25] , \ScanLink229[24] , \ScanLink229[23] , 
        \ScanLink229[22] , \ScanLink229[21] , \ScanLink229[20] , 
        \ScanLink229[19] , \ScanLink229[18] , \ScanLink229[17] , 
        \ScanLink229[16] , \ScanLink229[15] , \ScanLink229[14] , 
        \ScanLink229[13] , \ScanLink229[12] , \ScanLink229[11] , 
        \ScanLink229[10] , \ScanLink229[9] , \ScanLink229[8] , 
        \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , \ScanLink229[4] , 
        \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , \ScanLink229[0] 
        }), .ScanOut({\ScanLink228[31] , \ScanLink228[30] , \ScanLink228[29] , 
        \ScanLink228[28] , \ScanLink228[27] , \ScanLink228[26] , 
        \ScanLink228[25] , \ScanLink228[24] , \ScanLink228[23] , 
        \ScanLink228[22] , \ScanLink228[21] , \ScanLink228[20] , 
        \ScanLink228[19] , \ScanLink228[18] , \ScanLink228[17] , 
        \ScanLink228[16] , \ScanLink228[15] , \ScanLink228[14] , 
        \ScanLink228[13] , \ScanLink228[12] , \ScanLink228[11] , 
        \ScanLink228[10] , \ScanLink228[9] , \ScanLink228[8] , 
        \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , \ScanLink228[4] , 
        \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , \ScanLink228[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB13[31] , \wRegInB13[30] , \wRegInB13[29] , 
        \wRegInB13[28] , \wRegInB13[27] , \wRegInB13[26] , \wRegInB13[25] , 
        \wRegInB13[24] , \wRegInB13[23] , \wRegInB13[22] , \wRegInB13[21] , 
        \wRegInB13[20] , \wRegInB13[19] , \wRegInB13[18] , \wRegInB13[17] , 
        \wRegInB13[16] , \wRegInB13[15] , \wRegInB13[14] , \wRegInB13[13] , 
        \wRegInB13[12] , \wRegInB13[11] , \wRegInB13[10] , \wRegInB13[9] , 
        \wRegInB13[8] , \wRegInB13[7] , \wRegInB13[6] , \wRegInB13[5] , 
        \wRegInB13[4] , \wRegInB13[3] , \wRegInB13[2] , \wRegInB13[1] , 
        \wRegInB13[0] }), .Out({\wBIn13[31] , \wBIn13[30] , \wBIn13[29] , 
        \wBIn13[28] , \wBIn13[27] , \wBIn13[26] , \wBIn13[25] , \wBIn13[24] , 
        \wBIn13[23] , \wBIn13[22] , \wBIn13[21] , \wBIn13[20] , \wBIn13[19] , 
        \wBIn13[18] , \wBIn13[17] , \wBIn13[16] , \wBIn13[15] , \wBIn13[14] , 
        \wBIn13[13] , \wBIn13[12] , \wBIn13[11] , \wBIn13[10] , \wBIn13[9] , 
        \wBIn13[8] , \wBIn13[7] , \wBIn13[6] , \wBIn13[5] , \wBIn13[4] , 
        \wBIn13[3] , \wBIn13[2] , \wBIn13[1] , \wBIn13[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_118 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink119[31] , \ScanLink119[30] , \ScanLink119[29] , 
        \ScanLink119[28] , \ScanLink119[27] , \ScanLink119[26] , 
        \ScanLink119[25] , \ScanLink119[24] , \ScanLink119[23] , 
        \ScanLink119[22] , \ScanLink119[21] , \ScanLink119[20] , 
        \ScanLink119[19] , \ScanLink119[18] , \ScanLink119[17] , 
        \ScanLink119[16] , \ScanLink119[15] , \ScanLink119[14] , 
        \ScanLink119[13] , \ScanLink119[12] , \ScanLink119[11] , 
        \ScanLink119[10] , \ScanLink119[9] , \ScanLink119[8] , 
        \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , \ScanLink119[4] , 
        \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , \ScanLink119[0] 
        }), .ScanOut({\ScanLink118[31] , \ScanLink118[30] , \ScanLink118[29] , 
        \ScanLink118[28] , \ScanLink118[27] , \ScanLink118[26] , 
        \ScanLink118[25] , \ScanLink118[24] , \ScanLink118[23] , 
        \ScanLink118[22] , \ScanLink118[21] , \ScanLink118[20] , 
        \ScanLink118[19] , \ScanLink118[18] , \ScanLink118[17] , 
        \ScanLink118[16] , \ScanLink118[15] , \ScanLink118[14] , 
        \ScanLink118[13] , \ScanLink118[12] , \ScanLink118[11] , 
        \ScanLink118[10] , \ScanLink118[9] , \ScanLink118[8] , 
        \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , \ScanLink118[4] , 
        \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , \ScanLink118[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB68[31] , \wRegInB68[30] , \wRegInB68[29] , 
        \wRegInB68[28] , \wRegInB68[27] , \wRegInB68[26] , \wRegInB68[25] , 
        \wRegInB68[24] , \wRegInB68[23] , \wRegInB68[22] , \wRegInB68[21] , 
        \wRegInB68[20] , \wRegInB68[19] , \wRegInB68[18] , \wRegInB68[17] , 
        \wRegInB68[16] , \wRegInB68[15] , \wRegInB68[14] , \wRegInB68[13] , 
        \wRegInB68[12] , \wRegInB68[11] , \wRegInB68[10] , \wRegInB68[9] , 
        \wRegInB68[8] , \wRegInB68[7] , \wRegInB68[6] , \wRegInB68[5] , 
        \wRegInB68[4] , \wRegInB68[3] , \wRegInB68[2] , \wRegInB68[1] , 
        \wRegInB68[0] }), .Out({\wBIn68[31] , \wBIn68[30] , \wBIn68[29] , 
        \wBIn68[28] , \wBIn68[27] , \wBIn68[26] , \wBIn68[25] , \wBIn68[24] , 
        \wBIn68[23] , \wBIn68[22] , \wBIn68[21] , \wBIn68[20] , \wBIn68[19] , 
        \wBIn68[18] , \wBIn68[17] , \wBIn68[16] , \wBIn68[15] , \wBIn68[14] , 
        \wBIn68[13] , \wBIn68[12] , \wBIn68[11] , \wBIn68[10] , \wBIn68[9] , 
        \wBIn68[8] , \wBIn68[7] , \wBIn68[6] , \wBIn68[5] , \wBIn68[4] , 
        \wBIn68[3] , \wBIn68[2] , \wBIn68[1] , \wBIn68[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_48 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink49[31] , \ScanLink49[30] , \ScanLink49[29] , 
        \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , \ScanLink49[25] , 
        \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , \ScanLink49[21] , 
        \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , \ScanLink49[17] , 
        \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , \ScanLink49[13] , 
        \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , \ScanLink49[9] , 
        \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , \ScanLink49[5] , 
        \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , \ScanLink49[1] , 
        \ScanLink49[0] }), .ScanOut({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB103[31] , \wRegInB103[30] , 
        \wRegInB103[29] , \wRegInB103[28] , \wRegInB103[27] , \wRegInB103[26] , 
        \wRegInB103[25] , \wRegInB103[24] , \wRegInB103[23] , \wRegInB103[22] , 
        \wRegInB103[21] , \wRegInB103[20] , \wRegInB103[19] , \wRegInB103[18] , 
        \wRegInB103[17] , \wRegInB103[16] , \wRegInB103[15] , \wRegInB103[14] , 
        \wRegInB103[13] , \wRegInB103[12] , \wRegInB103[11] , \wRegInB103[10] , 
        \wRegInB103[9] , \wRegInB103[8] , \wRegInB103[7] , \wRegInB103[6] , 
        \wRegInB103[5] , \wRegInB103[4] , \wRegInB103[3] , \wRegInB103[2] , 
        \wRegInB103[1] , \wRegInB103[0] }), .Out({\wBIn103[31] , \wBIn103[30] , 
        \wBIn103[29] , \wBIn103[28] , \wBIn103[27] , \wBIn103[26] , 
        \wBIn103[25] , \wBIn103[24] , \wBIn103[23] , \wBIn103[22] , 
        \wBIn103[21] , \wBIn103[20] , \wBIn103[19] , \wBIn103[18] , 
        \wBIn103[17] , \wBIn103[16] , \wBIn103[15] , \wBIn103[14] , 
        \wBIn103[13] , \wBIn103[12] , \wBIn103[11] , \wBIn103[10] , 
        \wBIn103[9] , \wBIn103[8] , \wBIn103[7] , \wBIn103[6] , \wBIn103[5] , 
        \wBIn103[4] , \wBIn103[3] , \wBIn103[2] , \wBIn103[1] , \wBIn103[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn5[31] , 
        \wAIn5[30] , \wAIn5[29] , \wAIn5[28] , \wAIn5[27] , \wAIn5[26] , 
        \wAIn5[25] , \wAIn5[24] , \wAIn5[23] , \wAIn5[22] , \wAIn5[21] , 
        \wAIn5[20] , \wAIn5[19] , \wAIn5[18] , \wAIn5[17] , \wAIn5[16] , 
        \wAIn5[15] , \wAIn5[14] , \wAIn5[13] , \wAIn5[12] , \wAIn5[11] , 
        \wAIn5[10] , \wAIn5[9] , \wAIn5[8] , \wAIn5[7] , \wAIn5[6] , 
        \wAIn5[5] , \wAIn5[4] , \wAIn5[3] , \wAIn5[2] , \wAIn5[1] , \wAIn5[0] 
        }), .BIn({\wBIn5[31] , \wBIn5[30] , \wBIn5[29] , \wBIn5[28] , 
        \wBIn5[27] , \wBIn5[26] , \wBIn5[25] , \wBIn5[24] , \wBIn5[23] , 
        \wBIn5[22] , \wBIn5[21] , \wBIn5[20] , \wBIn5[19] , \wBIn5[18] , 
        \wBIn5[17] , \wBIn5[16] , \wBIn5[15] , \wBIn5[14] , \wBIn5[13] , 
        \wBIn5[12] , \wBIn5[11] , \wBIn5[10] , \wBIn5[9] , \wBIn5[8] , 
        \wBIn5[7] , \wBIn5[6] , \wBIn5[5] , \wBIn5[4] , \wBIn5[3] , \wBIn5[2] , 
        \wBIn5[1] , \wBIn5[0] }), .HiOut({\wBMid4[31] , \wBMid4[30] , 
        \wBMid4[29] , \wBMid4[28] , \wBMid4[27] , \wBMid4[26] , \wBMid4[25] , 
        \wBMid4[24] , \wBMid4[23] , \wBMid4[22] , \wBMid4[21] , \wBMid4[20] , 
        \wBMid4[19] , \wBMid4[18] , \wBMid4[17] , \wBMid4[16] , \wBMid4[15] , 
        \wBMid4[14] , \wBMid4[13] , \wBMid4[12] , \wBMid4[11] , \wBMid4[10] , 
        \wBMid4[9] , \wBMid4[8] , \wBMid4[7] , \wBMid4[6] , \wBMid4[5] , 
        \wBMid4[4] , \wBMid4[3] , \wBMid4[2] , \wBMid4[1] , \wBMid4[0] }), 
        .LoOut({\wAMid5[31] , \wAMid5[30] , \wAMid5[29] , \wAMid5[28] , 
        \wAMid5[27] , \wAMid5[26] , \wAMid5[25] , \wAMid5[24] , \wAMid5[23] , 
        \wAMid5[22] , \wAMid5[21] , \wAMid5[20] , \wAMid5[19] , \wAMid5[18] , 
        \wAMid5[17] , \wAMid5[16] , \wAMid5[15] , \wAMid5[14] , \wAMid5[13] , 
        \wAMid5[12] , \wAMid5[11] , \wAMid5[10] , \wAMid5[9] , \wAMid5[8] , 
        \wAMid5[7] , \wAMid5[6] , \wAMid5[5] , \wAMid5[4] , \wAMid5[3] , 
        \wAMid5[2] , \wAMid5[1] , \wAMid5[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn13[31] , \wAIn13[30] , \wAIn13[29] , \wAIn13[28] , \wAIn13[27] , 
        \wAIn13[26] , \wAIn13[25] , \wAIn13[24] , \wAIn13[23] , \wAIn13[22] , 
        \wAIn13[21] , \wAIn13[20] , \wAIn13[19] , \wAIn13[18] , \wAIn13[17] , 
        \wAIn13[16] , \wAIn13[15] , \wAIn13[14] , \wAIn13[13] , \wAIn13[12] , 
        \wAIn13[11] , \wAIn13[10] , \wAIn13[9] , \wAIn13[8] , \wAIn13[7] , 
        \wAIn13[6] , \wAIn13[5] , \wAIn13[4] , \wAIn13[3] , \wAIn13[2] , 
        \wAIn13[1] , \wAIn13[0] }), .BIn({\wBIn13[31] , \wBIn13[30] , 
        \wBIn13[29] , \wBIn13[28] , \wBIn13[27] , \wBIn13[26] , \wBIn13[25] , 
        \wBIn13[24] , \wBIn13[23] , \wBIn13[22] , \wBIn13[21] , \wBIn13[20] , 
        \wBIn13[19] , \wBIn13[18] , \wBIn13[17] , \wBIn13[16] , \wBIn13[15] , 
        \wBIn13[14] , \wBIn13[13] , \wBIn13[12] , \wBIn13[11] , \wBIn13[10] , 
        \wBIn13[9] , \wBIn13[8] , \wBIn13[7] , \wBIn13[6] , \wBIn13[5] , 
        \wBIn13[4] , \wBIn13[3] , \wBIn13[2] , \wBIn13[1] , \wBIn13[0] }), 
        .HiOut({\wBMid12[31] , \wBMid12[30] , \wBMid12[29] , \wBMid12[28] , 
        \wBMid12[27] , \wBMid12[26] , \wBMid12[25] , \wBMid12[24] , 
        \wBMid12[23] , \wBMid12[22] , \wBMid12[21] , \wBMid12[20] , 
        \wBMid12[19] , \wBMid12[18] , \wBMid12[17] , \wBMid12[16] , 
        \wBMid12[15] , \wBMid12[14] , \wBMid12[13] , \wBMid12[12] , 
        \wBMid12[11] , \wBMid12[10] , \wBMid12[9] , \wBMid12[8] , \wBMid12[7] , 
        \wBMid12[6] , \wBMid12[5] , \wBMid12[4] , \wBMid12[3] , \wBMid12[2] , 
        \wBMid12[1] , \wBMid12[0] }), .LoOut({\wAMid13[31] , \wAMid13[30] , 
        \wAMid13[29] , \wAMid13[28] , \wAMid13[27] , \wAMid13[26] , 
        \wAMid13[25] , \wAMid13[24] , \wAMid13[23] , \wAMid13[22] , 
        \wAMid13[21] , \wAMid13[20] , \wAMid13[19] , \wAMid13[18] , 
        \wAMid13[17] , \wAMid13[16] , \wAMid13[15] , \wAMid13[14] , 
        \wAMid13[13] , \wAMid13[12] , \wAMid13[11] , \wAMid13[10] , 
        \wAMid13[9] , \wAMid13[8] , \wAMid13[7] , \wAMid13[6] , \wAMid13[5] , 
        \wAMid13[4] , \wAMid13[3] , \wAMid13[2] , \wAMid13[1] , \wAMid13[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn14[31] , \wAIn14[30] , \wAIn14[29] , \wAIn14[28] , \wAIn14[27] , 
        \wAIn14[26] , \wAIn14[25] , \wAIn14[24] , \wAIn14[23] , \wAIn14[22] , 
        \wAIn14[21] , \wAIn14[20] , \wAIn14[19] , \wAIn14[18] , \wAIn14[17] , 
        \wAIn14[16] , \wAIn14[15] , \wAIn14[14] , \wAIn14[13] , \wAIn14[12] , 
        \wAIn14[11] , \wAIn14[10] , \wAIn14[9] , \wAIn14[8] , \wAIn14[7] , 
        \wAIn14[6] , \wAIn14[5] , \wAIn14[4] , \wAIn14[3] , \wAIn14[2] , 
        \wAIn14[1] , \wAIn14[0] }), .BIn({\wBIn14[31] , \wBIn14[30] , 
        \wBIn14[29] , \wBIn14[28] , \wBIn14[27] , \wBIn14[26] , \wBIn14[25] , 
        \wBIn14[24] , \wBIn14[23] , \wBIn14[22] , \wBIn14[21] , \wBIn14[20] , 
        \wBIn14[19] , \wBIn14[18] , \wBIn14[17] , \wBIn14[16] , \wBIn14[15] , 
        \wBIn14[14] , \wBIn14[13] , \wBIn14[12] , \wBIn14[11] , \wBIn14[10] , 
        \wBIn14[9] , \wBIn14[8] , \wBIn14[7] , \wBIn14[6] , \wBIn14[5] , 
        \wBIn14[4] , \wBIn14[3] , \wBIn14[2] , \wBIn14[1] , \wBIn14[0] }), 
        .HiOut({\wBMid13[31] , \wBMid13[30] , \wBMid13[29] , \wBMid13[28] , 
        \wBMid13[27] , \wBMid13[26] , \wBMid13[25] , \wBMid13[24] , 
        \wBMid13[23] , \wBMid13[22] , \wBMid13[21] , \wBMid13[20] , 
        \wBMid13[19] , \wBMid13[18] , \wBMid13[17] , \wBMid13[16] , 
        \wBMid13[15] , \wBMid13[14] , \wBMid13[13] , \wBMid13[12] , 
        \wBMid13[11] , \wBMid13[10] , \wBMid13[9] , \wBMid13[8] , \wBMid13[7] , 
        \wBMid13[6] , \wBMid13[5] , \wBMid13[4] , \wBMid13[3] , \wBMid13[2] , 
        \wBMid13[1] , \wBMid13[0] }), .LoOut({\wAMid14[31] , \wAMid14[30] , 
        \wAMid14[29] , \wAMid14[28] , \wAMid14[27] , \wAMid14[26] , 
        \wAMid14[25] , \wAMid14[24] , \wAMid14[23] , \wAMid14[22] , 
        \wAMid14[21] , \wAMid14[20] , \wAMid14[19] , \wAMid14[18] , 
        \wAMid14[17] , \wAMid14[16] , \wAMid14[15] , \wAMid14[14] , 
        \wAMid14[13] , \wAMid14[12] , \wAMid14[11] , \wAMid14[10] , 
        \wAMid14[9] , \wAMid14[8] , \wAMid14[7] , \wAMid14[6] , \wAMid14[5] , 
        \wAMid14[4] , \wAMid14[3] , \wAMid14[2] , \wAMid14[1] , \wAMid14[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn46[31] , \wAIn46[30] , \wAIn46[29] , \wAIn46[28] , \wAIn46[27] , 
        \wAIn46[26] , \wAIn46[25] , \wAIn46[24] , \wAIn46[23] , \wAIn46[22] , 
        \wAIn46[21] , \wAIn46[20] , \wAIn46[19] , \wAIn46[18] , \wAIn46[17] , 
        \wAIn46[16] , \wAIn46[15] , \wAIn46[14] , \wAIn46[13] , \wAIn46[12] , 
        \wAIn46[11] , \wAIn46[10] , \wAIn46[9] , \wAIn46[8] , \wAIn46[7] , 
        \wAIn46[6] , \wAIn46[5] , \wAIn46[4] , \wAIn46[3] , \wAIn46[2] , 
        \wAIn46[1] , \wAIn46[0] }), .BIn({\wBIn46[31] , \wBIn46[30] , 
        \wBIn46[29] , \wBIn46[28] , \wBIn46[27] , \wBIn46[26] , \wBIn46[25] , 
        \wBIn46[24] , \wBIn46[23] , \wBIn46[22] , \wBIn46[21] , \wBIn46[20] , 
        \wBIn46[19] , \wBIn46[18] , \wBIn46[17] , \wBIn46[16] , \wBIn46[15] , 
        \wBIn46[14] , \wBIn46[13] , \wBIn46[12] , \wBIn46[11] , \wBIn46[10] , 
        \wBIn46[9] , \wBIn46[8] , \wBIn46[7] , \wBIn46[6] , \wBIn46[5] , 
        \wBIn46[4] , \wBIn46[3] , \wBIn46[2] , \wBIn46[1] , \wBIn46[0] }), 
        .HiOut({\wBMid45[31] , \wBMid45[30] , \wBMid45[29] , \wBMid45[28] , 
        \wBMid45[27] , \wBMid45[26] , \wBMid45[25] , \wBMid45[24] , 
        \wBMid45[23] , \wBMid45[22] , \wBMid45[21] , \wBMid45[20] , 
        \wBMid45[19] , \wBMid45[18] , \wBMid45[17] , \wBMid45[16] , 
        \wBMid45[15] , \wBMid45[14] , \wBMid45[13] , \wBMid45[12] , 
        \wBMid45[11] , \wBMid45[10] , \wBMid45[9] , \wBMid45[8] , \wBMid45[7] , 
        \wBMid45[6] , \wBMid45[5] , \wBMid45[4] , \wBMid45[3] , \wBMid45[2] , 
        \wBMid45[1] , \wBMid45[0] }), .LoOut({\wAMid46[31] , \wAMid46[30] , 
        \wAMid46[29] , \wAMid46[28] , \wAMid46[27] , \wAMid46[26] , 
        \wAMid46[25] , \wAMid46[24] , \wAMid46[23] , \wAMid46[22] , 
        \wAMid46[21] , \wAMid46[20] , \wAMid46[19] , \wAMid46[18] , 
        \wAMid46[17] , \wAMid46[16] , \wAMid46[15] , \wAMid46[14] , 
        \wAMid46[13] , \wAMid46[12] , \wAMid46[11] , \wAMid46[10] , 
        \wAMid46[9] , \wAMid46[8] , \wAMid46[7] , \wAMid46[6] , \wAMid46[5] , 
        \wAMid46[4] , \wAMid46[3] , \wAMid46[2] , \wAMid46[1] , \wAMid46[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn61[31] , \wAIn61[30] , \wAIn61[29] , \wAIn61[28] , \wAIn61[27] , 
        \wAIn61[26] , \wAIn61[25] , \wAIn61[24] , \wAIn61[23] , \wAIn61[22] , 
        \wAIn61[21] , \wAIn61[20] , \wAIn61[19] , \wAIn61[18] , \wAIn61[17] , 
        \wAIn61[16] , \wAIn61[15] , \wAIn61[14] , \wAIn61[13] , \wAIn61[12] , 
        \wAIn61[11] , \wAIn61[10] , \wAIn61[9] , \wAIn61[8] , \wAIn61[7] , 
        \wAIn61[6] , \wAIn61[5] , \wAIn61[4] , \wAIn61[3] , \wAIn61[2] , 
        \wAIn61[1] , \wAIn61[0] }), .BIn({\wBIn61[31] , \wBIn61[30] , 
        \wBIn61[29] , \wBIn61[28] , \wBIn61[27] , \wBIn61[26] , \wBIn61[25] , 
        \wBIn61[24] , \wBIn61[23] , \wBIn61[22] , \wBIn61[21] , \wBIn61[20] , 
        \wBIn61[19] , \wBIn61[18] , \wBIn61[17] , \wBIn61[16] , \wBIn61[15] , 
        \wBIn61[14] , \wBIn61[13] , \wBIn61[12] , \wBIn61[11] , \wBIn61[10] , 
        \wBIn61[9] , \wBIn61[8] , \wBIn61[7] , \wBIn61[6] , \wBIn61[5] , 
        \wBIn61[4] , \wBIn61[3] , \wBIn61[2] , \wBIn61[1] , \wBIn61[0] }), 
        .HiOut({\wBMid60[31] , \wBMid60[30] , \wBMid60[29] , \wBMid60[28] , 
        \wBMid60[27] , \wBMid60[26] , \wBMid60[25] , \wBMid60[24] , 
        \wBMid60[23] , \wBMid60[22] , \wBMid60[21] , \wBMid60[20] , 
        \wBMid60[19] , \wBMid60[18] , \wBMid60[17] , \wBMid60[16] , 
        \wBMid60[15] , \wBMid60[14] , \wBMid60[13] , \wBMid60[12] , 
        \wBMid60[11] , \wBMid60[10] , \wBMid60[9] , \wBMid60[8] , \wBMid60[7] , 
        \wBMid60[6] , \wBMid60[5] , \wBMid60[4] , \wBMid60[3] , \wBMid60[2] , 
        \wBMid60[1] , \wBMid60[0] }), .LoOut({\wAMid61[31] , \wAMid61[30] , 
        \wAMid61[29] , \wAMid61[28] , \wAMid61[27] , \wAMid61[26] , 
        \wAMid61[25] , \wAMid61[24] , \wAMid61[23] , \wAMid61[22] , 
        \wAMid61[21] , \wAMid61[20] , \wAMid61[19] , \wAMid61[18] , 
        \wAMid61[17] , \wAMid61[16] , \wAMid61[15] , \wAMid61[14] , 
        \wAMid61[13] , \wAMid61[12] , \wAMid61[11] , \wAMid61[10] , 
        \wAMid61[9] , \wAMid61[8] , \wAMid61[7] , \wAMid61[6] , \wAMid61[5] , 
        \wAMid61[4] , \wAMid61[3] , \wAMid61[2] , \wAMid61[1] , \wAMid61[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn84[31] , \wAIn84[30] , \wAIn84[29] , \wAIn84[28] , \wAIn84[27] , 
        \wAIn84[26] , \wAIn84[25] , \wAIn84[24] , \wAIn84[23] , \wAIn84[22] , 
        \wAIn84[21] , \wAIn84[20] , \wAIn84[19] , \wAIn84[18] , \wAIn84[17] , 
        \wAIn84[16] , \wAIn84[15] , \wAIn84[14] , \wAIn84[13] , \wAIn84[12] , 
        \wAIn84[11] , \wAIn84[10] , \wAIn84[9] , \wAIn84[8] , \wAIn84[7] , 
        \wAIn84[6] , \wAIn84[5] , \wAIn84[4] , \wAIn84[3] , \wAIn84[2] , 
        \wAIn84[1] , \wAIn84[0] }), .BIn({\wBIn84[31] , \wBIn84[30] , 
        \wBIn84[29] , \wBIn84[28] , \wBIn84[27] , \wBIn84[26] , \wBIn84[25] , 
        \wBIn84[24] , \wBIn84[23] , \wBIn84[22] , \wBIn84[21] , \wBIn84[20] , 
        \wBIn84[19] , \wBIn84[18] , \wBIn84[17] , \wBIn84[16] , \wBIn84[15] , 
        \wBIn84[14] , \wBIn84[13] , \wBIn84[12] , \wBIn84[11] , \wBIn84[10] , 
        \wBIn84[9] , \wBIn84[8] , \wBIn84[7] , \wBIn84[6] , \wBIn84[5] , 
        \wBIn84[4] , \wBIn84[3] , \wBIn84[2] , \wBIn84[1] , \wBIn84[0] }), 
        .HiOut({\wBMid83[31] , \wBMid83[30] , \wBMid83[29] , \wBMid83[28] , 
        \wBMid83[27] , \wBMid83[26] , \wBMid83[25] , \wBMid83[24] , 
        \wBMid83[23] , \wBMid83[22] , \wBMid83[21] , \wBMid83[20] , 
        \wBMid83[19] , \wBMid83[18] , \wBMid83[17] , \wBMid83[16] , 
        \wBMid83[15] , \wBMid83[14] , \wBMid83[13] , \wBMid83[12] , 
        \wBMid83[11] , \wBMid83[10] , \wBMid83[9] , \wBMid83[8] , \wBMid83[7] , 
        \wBMid83[6] , \wBMid83[5] , \wBMid83[4] , \wBMid83[3] , \wBMid83[2] , 
        \wBMid83[1] , \wBMid83[0] }), .LoOut({\wAMid84[31] , \wAMid84[30] , 
        \wAMid84[29] , \wAMid84[28] , \wAMid84[27] , \wAMid84[26] , 
        \wAMid84[25] , \wAMid84[24] , \wAMid84[23] , \wAMid84[22] , 
        \wAMid84[21] , \wAMid84[20] , \wAMid84[19] , \wAMid84[18] , 
        \wAMid84[17] , \wAMid84[16] , \wAMid84[15] , \wAMid84[14] , 
        \wAMid84[13] , \wAMid84[12] , \wAMid84[11] , \wAMid84[10] , 
        \wAMid84[9] , \wAMid84[8] , \wAMid84[7] , \wAMid84[6] , \wAMid84[5] , 
        \wAMid84[4] , \wAMid84[3] , \wAMid84[2] , \wAMid84[1] , \wAMid84[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid93[31] , \wAMid93[30] , \wAMid93[29] , \wAMid93[28] , 
        \wAMid93[27] , \wAMid93[26] , \wAMid93[25] , \wAMid93[24] , 
        \wAMid93[23] , \wAMid93[22] , \wAMid93[21] , \wAMid93[20] , 
        \wAMid93[19] , \wAMid93[18] , \wAMid93[17] , \wAMid93[16] , 
        \wAMid93[15] , \wAMid93[14] , \wAMid93[13] , \wAMid93[12] , 
        \wAMid93[11] , \wAMid93[10] , \wAMid93[9] , \wAMid93[8] , \wAMid93[7] , 
        \wAMid93[6] , \wAMid93[5] , \wAMid93[4] , \wAMid93[3] , \wAMid93[2] , 
        \wAMid93[1] , \wAMid93[0] }), .BIn({\wBMid93[31] , \wBMid93[30] , 
        \wBMid93[29] , \wBMid93[28] , \wBMid93[27] , \wBMid93[26] , 
        \wBMid93[25] , \wBMid93[24] , \wBMid93[23] , \wBMid93[22] , 
        \wBMid93[21] , \wBMid93[20] , \wBMid93[19] , \wBMid93[18] , 
        \wBMid93[17] , \wBMid93[16] , \wBMid93[15] , \wBMid93[14] , 
        \wBMid93[13] , \wBMid93[12] , \wBMid93[11] , \wBMid93[10] , 
        \wBMid93[9] , \wBMid93[8] , \wBMid93[7] , \wBMid93[6] , \wBMid93[5] , 
        \wBMid93[4] , \wBMid93[3] , \wBMid93[2] , \wBMid93[1] , \wBMid93[0] }), 
        .HiOut({\wRegInB93[31] , \wRegInB93[30] , \wRegInB93[29] , 
        \wRegInB93[28] , \wRegInB93[27] , \wRegInB93[26] , \wRegInB93[25] , 
        \wRegInB93[24] , \wRegInB93[23] , \wRegInB93[22] , \wRegInB93[21] , 
        \wRegInB93[20] , \wRegInB93[19] , \wRegInB93[18] , \wRegInB93[17] , 
        \wRegInB93[16] , \wRegInB93[15] , \wRegInB93[14] , \wRegInB93[13] , 
        \wRegInB93[12] , \wRegInB93[11] , \wRegInB93[10] , \wRegInB93[9] , 
        \wRegInB93[8] , \wRegInB93[7] , \wRegInB93[6] , \wRegInB93[5] , 
        \wRegInB93[4] , \wRegInB93[3] , \wRegInB93[2] , \wRegInB93[1] , 
        \wRegInB93[0] }), .LoOut({\wRegInA94[31] , \wRegInA94[30] , 
        \wRegInA94[29] , \wRegInA94[28] , \wRegInA94[27] , \wRegInA94[26] , 
        \wRegInA94[25] , \wRegInA94[24] , \wRegInA94[23] , \wRegInA94[22] , 
        \wRegInA94[21] , \wRegInA94[20] , \wRegInA94[19] , \wRegInA94[18] , 
        \wRegInA94[17] , \wRegInA94[16] , \wRegInA94[15] , \wRegInA94[14] , 
        \wRegInA94[13] , \wRegInA94[12] , \wRegInA94[11] , \wRegInA94[10] , 
        \wRegInA94[9] , \wRegInA94[8] , \wRegInA94[7] , \wRegInA94[6] , 
        \wRegInA94[5] , \wRegInA94[4] , \wRegInA94[3] , \wRegInA94[2] , 
        \wRegInA94[1] , \wRegInA94[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid51[31] , \wAMid51[30] , \wAMid51[29] , \wAMid51[28] , 
        \wAMid51[27] , \wAMid51[26] , \wAMid51[25] , \wAMid51[24] , 
        \wAMid51[23] , \wAMid51[22] , \wAMid51[21] , \wAMid51[20] , 
        \wAMid51[19] , \wAMid51[18] , \wAMid51[17] , \wAMid51[16] , 
        \wAMid51[15] , \wAMid51[14] , \wAMid51[13] , \wAMid51[12] , 
        \wAMid51[11] , \wAMid51[10] , \wAMid51[9] , \wAMid51[8] , \wAMid51[7] , 
        \wAMid51[6] , \wAMid51[5] , \wAMid51[4] , \wAMid51[3] , \wAMid51[2] , 
        \wAMid51[1] , \wAMid51[0] }), .BIn({\wBMid51[31] , \wBMid51[30] , 
        \wBMid51[29] , \wBMid51[28] , \wBMid51[27] , \wBMid51[26] , 
        \wBMid51[25] , \wBMid51[24] , \wBMid51[23] , \wBMid51[22] , 
        \wBMid51[21] , \wBMid51[20] , \wBMid51[19] , \wBMid51[18] , 
        \wBMid51[17] , \wBMid51[16] , \wBMid51[15] , \wBMid51[14] , 
        \wBMid51[13] , \wBMid51[12] , \wBMid51[11] , \wBMid51[10] , 
        \wBMid51[9] , \wBMid51[8] , \wBMid51[7] , \wBMid51[6] , \wBMid51[5] , 
        \wBMid51[4] , \wBMid51[3] , \wBMid51[2] , \wBMid51[1] , \wBMid51[0] }), 
        .HiOut({\wRegInB51[31] , \wRegInB51[30] , \wRegInB51[29] , 
        \wRegInB51[28] , \wRegInB51[27] , \wRegInB51[26] , \wRegInB51[25] , 
        \wRegInB51[24] , \wRegInB51[23] , \wRegInB51[22] , \wRegInB51[21] , 
        \wRegInB51[20] , \wRegInB51[19] , \wRegInB51[18] , \wRegInB51[17] , 
        \wRegInB51[16] , \wRegInB51[15] , \wRegInB51[14] , \wRegInB51[13] , 
        \wRegInB51[12] , \wRegInB51[11] , \wRegInB51[10] , \wRegInB51[9] , 
        \wRegInB51[8] , \wRegInB51[7] , \wRegInB51[6] , \wRegInB51[5] , 
        \wRegInB51[4] , \wRegInB51[3] , \wRegInB51[2] , \wRegInB51[1] , 
        \wRegInB51[0] }), .LoOut({\wRegInA52[31] , \wRegInA52[30] , 
        \wRegInA52[29] , \wRegInA52[28] , \wRegInA52[27] , \wRegInA52[26] , 
        \wRegInA52[25] , \wRegInA52[24] , \wRegInA52[23] , \wRegInA52[22] , 
        \wRegInA52[21] , \wRegInA52[20] , \wRegInA52[19] , \wRegInA52[18] , 
        \wRegInA52[17] , \wRegInA52[16] , \wRegInA52[15] , \wRegInA52[14] , 
        \wRegInA52[13] , \wRegInA52[12] , \wRegInA52[11] , \wRegInA52[10] , 
        \wRegInA52[9] , \wRegInA52[8] , \wRegInA52[7] , \wRegInA52[6] , 
        \wRegInA52[5] , \wRegInA52[4] , \wRegInA52[3] , \wRegInA52[2] , 
        \wRegInA52[1] , \wRegInA52[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_181 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink182[31] , \ScanLink182[30] , \ScanLink182[29] , 
        \ScanLink182[28] , \ScanLink182[27] , \ScanLink182[26] , 
        \ScanLink182[25] , \ScanLink182[24] , \ScanLink182[23] , 
        \ScanLink182[22] , \ScanLink182[21] , \ScanLink182[20] , 
        \ScanLink182[19] , \ScanLink182[18] , \ScanLink182[17] , 
        \ScanLink182[16] , \ScanLink182[15] , \ScanLink182[14] , 
        \ScanLink182[13] , \ScanLink182[12] , \ScanLink182[11] , 
        \ScanLink182[10] , \ScanLink182[9] , \ScanLink182[8] , 
        \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , \ScanLink182[4] , 
        \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , \ScanLink182[0] 
        }), .ScanOut({\ScanLink181[31] , \ScanLink181[30] , \ScanLink181[29] , 
        \ScanLink181[28] , \ScanLink181[27] , \ScanLink181[26] , 
        \ScanLink181[25] , \ScanLink181[24] , \ScanLink181[23] , 
        \ScanLink181[22] , \ScanLink181[21] , \ScanLink181[20] , 
        \ScanLink181[19] , \ScanLink181[18] , \ScanLink181[17] , 
        \ScanLink181[16] , \ScanLink181[15] , \ScanLink181[14] , 
        \ScanLink181[13] , \ScanLink181[12] , \ScanLink181[11] , 
        \ScanLink181[10] , \ScanLink181[9] , \ScanLink181[8] , 
        \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , \ScanLink181[4] , 
        \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , \ScanLink181[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA37[31] , \wRegInA37[30] , \wRegInA37[29] , 
        \wRegInA37[28] , \wRegInA37[27] , \wRegInA37[26] , \wRegInA37[25] , 
        \wRegInA37[24] , \wRegInA37[23] , \wRegInA37[22] , \wRegInA37[21] , 
        \wRegInA37[20] , \wRegInA37[19] , \wRegInA37[18] , \wRegInA37[17] , 
        \wRegInA37[16] , \wRegInA37[15] , \wRegInA37[14] , \wRegInA37[13] , 
        \wRegInA37[12] , \wRegInA37[11] , \wRegInA37[10] , \wRegInA37[9] , 
        \wRegInA37[8] , \wRegInA37[7] , \wRegInA37[6] , \wRegInA37[5] , 
        \wRegInA37[4] , \wRegInA37[3] , \wRegInA37[2] , \wRegInA37[1] , 
        \wRegInA37[0] }), .Out({\wAIn37[31] , \wAIn37[30] , \wAIn37[29] , 
        \wAIn37[28] , \wAIn37[27] , \wAIn37[26] , \wAIn37[25] , \wAIn37[24] , 
        \wAIn37[23] , \wAIn37[22] , \wAIn37[21] , \wAIn37[20] , \wAIn37[19] , 
        \wAIn37[18] , \wAIn37[17] , \wAIn37[16] , \wAIn37[15] , \wAIn37[14] , 
        \wAIn37[13] , \wAIn37[12] , \wAIn37[11] , \wAIn37[10] , \wAIn37[9] , 
        \wAIn37[8] , \wAIn37[7] , \wAIn37[6] , \wAIn37[5] , \wAIn37[4] , 
        \wAIn37[3] , \wAIn37[2] , \wAIn37[1] , \wAIn37[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_98 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink99[31] , \ScanLink99[30] , \ScanLink99[29] , 
        \ScanLink99[28] , \ScanLink99[27] , \ScanLink99[26] , \ScanLink99[25] , 
        \ScanLink99[24] , \ScanLink99[23] , \ScanLink99[22] , \ScanLink99[21] , 
        \ScanLink99[20] , \ScanLink99[19] , \ScanLink99[18] , \ScanLink99[17] , 
        \ScanLink99[16] , \ScanLink99[15] , \ScanLink99[14] , \ScanLink99[13] , 
        \ScanLink99[12] , \ScanLink99[11] , \ScanLink99[10] , \ScanLink99[9] , 
        \ScanLink99[8] , \ScanLink99[7] , \ScanLink99[6] , \ScanLink99[5] , 
        \ScanLink99[4] , \ScanLink99[3] , \ScanLink99[2] , \ScanLink99[1] , 
        \ScanLink99[0] }), .ScanOut({\ScanLink98[31] , \ScanLink98[30] , 
        \ScanLink98[29] , \ScanLink98[28] , \ScanLink98[27] , \ScanLink98[26] , 
        \ScanLink98[25] , \ScanLink98[24] , \ScanLink98[23] , \ScanLink98[22] , 
        \ScanLink98[21] , \ScanLink98[20] , \ScanLink98[19] , \ScanLink98[18] , 
        \ScanLink98[17] , \ScanLink98[16] , \ScanLink98[15] , \ScanLink98[14] , 
        \ScanLink98[13] , \ScanLink98[12] , \ScanLink98[11] , \ScanLink98[10] , 
        \ScanLink98[9] , \ScanLink98[8] , \ScanLink98[7] , \ScanLink98[6] , 
        \ScanLink98[5] , \ScanLink98[4] , \ScanLink98[3] , \ScanLink98[2] , 
        \ScanLink98[1] , \ScanLink98[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB78[31] , \wRegInB78[30] , 
        \wRegInB78[29] , \wRegInB78[28] , \wRegInB78[27] , \wRegInB78[26] , 
        \wRegInB78[25] , \wRegInB78[24] , \wRegInB78[23] , \wRegInB78[22] , 
        \wRegInB78[21] , \wRegInB78[20] , \wRegInB78[19] , \wRegInB78[18] , 
        \wRegInB78[17] , \wRegInB78[16] , \wRegInB78[15] , \wRegInB78[14] , 
        \wRegInB78[13] , \wRegInB78[12] , \wRegInB78[11] , \wRegInB78[10] , 
        \wRegInB78[9] , \wRegInB78[8] , \wRegInB78[7] , \wRegInB78[6] , 
        \wRegInB78[5] , \wRegInB78[4] , \wRegInB78[3] , \wRegInB78[2] , 
        \wRegInB78[1] , \wRegInB78[0] }), .Out({\wBIn78[31] , \wBIn78[30] , 
        \wBIn78[29] , \wBIn78[28] , \wBIn78[27] , \wBIn78[26] , \wBIn78[25] , 
        \wBIn78[24] , \wBIn78[23] , \wBIn78[22] , \wBIn78[21] , \wBIn78[20] , 
        \wBIn78[19] , \wBIn78[18] , \wBIn78[17] , \wBIn78[16] , \wBIn78[15] , 
        \wBIn78[14] , \wBIn78[13] , \wBIn78[12] , \wBIn78[11] , \wBIn78[10] , 
        \wBIn78[9] , \wBIn78[8] , \wBIn78[7] , \wBIn78[6] , \wBIn78[5] , 
        \wBIn78[4] , \wBIn78[3] , \wBIn78[2] , \wBIn78[1] , \wBIn78[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_164 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink165[31] , \ScanLink165[30] , \ScanLink165[29] , 
        \ScanLink165[28] , \ScanLink165[27] , \ScanLink165[26] , 
        \ScanLink165[25] , \ScanLink165[24] , \ScanLink165[23] , 
        \ScanLink165[22] , \ScanLink165[21] , \ScanLink165[20] , 
        \ScanLink165[19] , \ScanLink165[18] , \ScanLink165[17] , 
        \ScanLink165[16] , \ScanLink165[15] , \ScanLink165[14] , 
        \ScanLink165[13] , \ScanLink165[12] , \ScanLink165[11] , 
        \ScanLink165[10] , \ScanLink165[9] , \ScanLink165[8] , 
        \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , \ScanLink165[4] , 
        \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , \ScanLink165[0] 
        }), .ScanOut({\ScanLink164[31] , \ScanLink164[30] , \ScanLink164[29] , 
        \ScanLink164[28] , \ScanLink164[27] , \ScanLink164[26] , 
        \ScanLink164[25] , \ScanLink164[24] , \ScanLink164[23] , 
        \ScanLink164[22] , \ScanLink164[21] , \ScanLink164[20] , 
        \ScanLink164[19] , \ScanLink164[18] , \ScanLink164[17] , 
        \ScanLink164[16] , \ScanLink164[15] , \ScanLink164[14] , 
        \ScanLink164[13] , \ScanLink164[12] , \ScanLink164[11] , 
        \ScanLink164[10] , \ScanLink164[9] , \ScanLink164[8] , 
        \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , \ScanLink164[4] , 
        \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , \ScanLink164[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB45[31] , \wRegInB45[30] , \wRegInB45[29] , 
        \wRegInB45[28] , \wRegInB45[27] , \wRegInB45[26] , \wRegInB45[25] , 
        \wRegInB45[24] , \wRegInB45[23] , \wRegInB45[22] , \wRegInB45[21] , 
        \wRegInB45[20] , \wRegInB45[19] , \wRegInB45[18] , \wRegInB45[17] , 
        \wRegInB45[16] , \wRegInB45[15] , \wRegInB45[14] , \wRegInB45[13] , 
        \wRegInB45[12] , \wRegInB45[11] , \wRegInB45[10] , \wRegInB45[9] , 
        \wRegInB45[8] , \wRegInB45[7] , \wRegInB45[6] , \wRegInB45[5] , 
        \wRegInB45[4] , \wRegInB45[3] , \wRegInB45[2] , \wRegInB45[1] , 
        \wRegInB45[0] }), .Out({\wBIn45[31] , \wBIn45[30] , \wBIn45[29] , 
        \wBIn45[28] , \wBIn45[27] , \wBIn45[26] , \wBIn45[25] , \wBIn45[24] , 
        \wBIn45[23] , \wBIn45[22] , \wBIn45[21] , \wBIn45[20] , \wBIn45[19] , 
        \wBIn45[18] , \wBIn45[17] , \wBIn45[16] , \wBIn45[15] , \wBIn45[14] , 
        \wBIn45[13] , \wBIn45[12] , \wBIn45[11] , \wBIn45[10] , \wBIn45[9] , 
        \wBIn45[8] , \wBIn45[7] , \wBIn45[6] , \wBIn45[5] , \wBIn45[4] , 
        \wBIn45[3] , \wBIn45[2] , \wBIn45[1] , \wBIn45[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_34 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink35[31] , \ScanLink35[30] , \ScanLink35[29] , 
        \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , \ScanLink35[25] , 
        \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , \ScanLink35[21] , 
        \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , \ScanLink35[17] , 
        \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , \ScanLink35[13] , 
        \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , \ScanLink35[9] , 
        \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , \ScanLink35[5] , 
        \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , \ScanLink35[1] , 
        \ScanLink35[0] }), .ScanOut({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB110[31] , \wRegInB110[30] , 
        \wRegInB110[29] , \wRegInB110[28] , \wRegInB110[27] , \wRegInB110[26] , 
        \wRegInB110[25] , \wRegInB110[24] , \wRegInB110[23] , \wRegInB110[22] , 
        \wRegInB110[21] , \wRegInB110[20] , \wRegInB110[19] , \wRegInB110[18] , 
        \wRegInB110[17] , \wRegInB110[16] , \wRegInB110[15] , \wRegInB110[14] , 
        \wRegInB110[13] , \wRegInB110[12] , \wRegInB110[11] , \wRegInB110[10] , 
        \wRegInB110[9] , \wRegInB110[8] , \wRegInB110[7] , \wRegInB110[6] , 
        \wRegInB110[5] , \wRegInB110[4] , \wRegInB110[3] , \wRegInB110[2] , 
        \wRegInB110[1] , \wRegInB110[0] }), .Out({\wBIn110[31] , \wBIn110[30] , 
        \wBIn110[29] , \wBIn110[28] , \wBIn110[27] , \wBIn110[26] , 
        \wBIn110[25] , \wBIn110[24] , \wBIn110[23] , \wBIn110[22] , 
        \wBIn110[21] , \wBIn110[20] , \wBIn110[19] , \wBIn110[18] , 
        \wBIn110[17] , \wBIn110[16] , \wBIn110[15] , \wBIn110[14] , 
        \wBIn110[13] , \wBIn110[12] , \wBIn110[11] , \wBIn110[10] , 
        \wBIn110[9] , \wBIn110[8] , \wBIn110[7] , \wBIn110[6] , \wBIn110[5] , 
        \wBIn110[4] , \wBIn110[3] , \wBIn110[2] , \wBIn110[1] , \wBIn110[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn111[31] , \wAIn111[30] , \wAIn111[29] , \wAIn111[28] , 
        \wAIn111[27] , \wAIn111[26] , \wAIn111[25] , \wAIn111[24] , 
        \wAIn111[23] , \wAIn111[22] , \wAIn111[21] , \wAIn111[20] , 
        \wAIn111[19] , \wAIn111[18] , \wAIn111[17] , \wAIn111[16] , 
        \wAIn111[15] , \wAIn111[14] , \wAIn111[13] , \wAIn111[12] , 
        \wAIn111[11] , \wAIn111[10] , \wAIn111[9] , \wAIn111[8] , \wAIn111[7] , 
        \wAIn111[6] , \wAIn111[5] , \wAIn111[4] , \wAIn111[3] , \wAIn111[2] , 
        \wAIn111[1] , \wAIn111[0] }), .BIn({\wBIn111[31] , \wBIn111[30] , 
        \wBIn111[29] , \wBIn111[28] , \wBIn111[27] , \wBIn111[26] , 
        \wBIn111[25] , \wBIn111[24] , \wBIn111[23] , \wBIn111[22] , 
        \wBIn111[21] , \wBIn111[20] , \wBIn111[19] , \wBIn111[18] , 
        \wBIn111[17] , \wBIn111[16] , \wBIn111[15] , \wBIn111[14] , 
        \wBIn111[13] , \wBIn111[12] , \wBIn111[11] , \wBIn111[10] , 
        \wBIn111[9] , \wBIn111[8] , \wBIn111[7] , \wBIn111[6] , \wBIn111[5] , 
        \wBIn111[4] , \wBIn111[3] , \wBIn111[2] , \wBIn111[1] , \wBIn111[0] }), 
        .HiOut({\wBMid110[31] , \wBMid110[30] , \wBMid110[29] , \wBMid110[28] , 
        \wBMid110[27] , \wBMid110[26] , \wBMid110[25] , \wBMid110[24] , 
        \wBMid110[23] , \wBMid110[22] , \wBMid110[21] , \wBMid110[20] , 
        \wBMid110[19] , \wBMid110[18] , \wBMid110[17] , \wBMid110[16] , 
        \wBMid110[15] , \wBMid110[14] , \wBMid110[13] , \wBMid110[12] , 
        \wBMid110[11] , \wBMid110[10] , \wBMid110[9] , \wBMid110[8] , 
        \wBMid110[7] , \wBMid110[6] , \wBMid110[5] , \wBMid110[4] , 
        \wBMid110[3] , \wBMid110[2] , \wBMid110[1] , \wBMid110[0] }), .LoOut({
        \wAMid111[31] , \wAMid111[30] , \wAMid111[29] , \wAMid111[28] , 
        \wAMid111[27] , \wAMid111[26] , \wAMid111[25] , \wAMid111[24] , 
        \wAMid111[23] , \wAMid111[22] , \wAMid111[21] , \wAMid111[20] , 
        \wAMid111[19] , \wAMid111[18] , \wAMid111[17] , \wAMid111[16] , 
        \wAMid111[15] , \wAMid111[14] , \wAMid111[13] , \wAMid111[12] , 
        \wAMid111[11] , \wAMid111[10] , \wAMid111[9] , \wAMid111[8] , 
        \wAMid111[7] , \wAMid111[6] , \wAMid111[5] , \wAMid111[4] , 
        \wAMid111[3] , \wAMid111[2] , \wAMid111[1] , \wAMid111[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_254 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink255[31] , \ScanLink255[30] , \ScanLink255[29] , 
        \ScanLink255[28] , \ScanLink255[27] , \ScanLink255[26] , 
        \ScanLink255[25] , \ScanLink255[24] , \ScanLink255[23] , 
        \ScanLink255[22] , \ScanLink255[21] , \ScanLink255[20] , 
        \ScanLink255[19] , \ScanLink255[18] , \ScanLink255[17] , 
        \ScanLink255[16] , \ScanLink255[15] , \ScanLink255[14] , 
        \ScanLink255[13] , \ScanLink255[12] , \ScanLink255[11] , 
        \ScanLink255[10] , \ScanLink255[9] , \ScanLink255[8] , 
        \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , \ScanLink255[4] , 
        \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , \ScanLink255[0] 
        }), .ScanOut({\ScanLink254[31] , \ScanLink254[30] , \ScanLink254[29] , 
        \ScanLink254[28] , \ScanLink254[27] , \ScanLink254[26] , 
        \ScanLink254[25] , \ScanLink254[24] , \ScanLink254[23] , 
        \ScanLink254[22] , \ScanLink254[21] , \ScanLink254[20] , 
        \ScanLink254[19] , \ScanLink254[18] , \ScanLink254[17] , 
        \ScanLink254[16] , \ScanLink254[15] , \ScanLink254[14] , 
        \ScanLink254[13] , \ScanLink254[12] , \ScanLink254[11] , 
        \ScanLink254[10] , \ScanLink254[9] , \ScanLink254[8] , 
        \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , \ScanLink254[4] , 
        \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , \ScanLink254[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB0[31] , \wRegInB0[30] , \wRegInB0[29] , \wRegInB0[28] , 
        \wRegInB0[27] , \wRegInB0[26] , \wRegInB0[25] , \wRegInB0[24] , 
        \wRegInB0[23] , \wRegInB0[22] , \wRegInB0[21] , \wRegInB0[20] , 
        \wRegInB0[19] , \wRegInB0[18] , \wRegInB0[17] , \wRegInB0[16] , 
        \wRegInB0[15] , \wRegInB0[14] , \wRegInB0[13] , \wRegInB0[12] , 
        \wRegInB0[11] , \wRegInB0[10] , \wRegInB0[9] , \wRegInB0[8] , 
        \wRegInB0[7] , \wRegInB0[6] , \wRegInB0[5] , \wRegInB0[4] , 
        \wRegInB0[3] , \wRegInB0[2] , \wRegInB0[1] , \wRegInB0[0] }), .Out({
        \wBIn0[31] , \wBIn0[30] , \wBIn0[29] , \wBIn0[28] , \wBIn0[27] , 
        \wBIn0[26] , \wBIn0[25] , \wBIn0[24] , \wBIn0[23] , \wBIn0[22] , 
        \wBIn0[21] , \wBIn0[20] , \wBIn0[19] , \wBIn0[18] , \wBIn0[17] , 
        \wBIn0[16] , \wBIn0[15] , \wBIn0[14] , \wBIn0[13] , \wBIn0[12] , 
        \wBIn0[11] , \wBIn0[10] , \wBIn0[9] , \wBIn0[8] , \wBIn0[7] , 
        \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , \wBIn0[3] , \wBIn0[2] , \wBIn0[1] , 
        \wBIn0[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid76[31] , \wAMid76[30] , \wAMid76[29] , \wAMid76[28] , 
        \wAMid76[27] , \wAMid76[26] , \wAMid76[25] , \wAMid76[24] , 
        \wAMid76[23] , \wAMid76[22] , \wAMid76[21] , \wAMid76[20] , 
        \wAMid76[19] , \wAMid76[18] , \wAMid76[17] , \wAMid76[16] , 
        \wAMid76[15] , \wAMid76[14] , \wAMid76[13] , \wAMid76[12] , 
        \wAMid76[11] , \wAMid76[10] , \wAMid76[9] , \wAMid76[8] , \wAMid76[7] , 
        \wAMid76[6] , \wAMid76[5] , \wAMid76[4] , \wAMid76[3] , \wAMid76[2] , 
        \wAMid76[1] , \wAMid76[0] }), .BIn({\wBMid76[31] , \wBMid76[30] , 
        \wBMid76[29] , \wBMid76[28] , \wBMid76[27] , \wBMid76[26] , 
        \wBMid76[25] , \wBMid76[24] , \wBMid76[23] , \wBMid76[22] , 
        \wBMid76[21] , \wBMid76[20] , \wBMid76[19] , \wBMid76[18] , 
        \wBMid76[17] , \wBMid76[16] , \wBMid76[15] , \wBMid76[14] , 
        \wBMid76[13] , \wBMid76[12] , \wBMid76[11] , \wBMid76[10] , 
        \wBMid76[9] , \wBMid76[8] , \wBMid76[7] , \wBMid76[6] , \wBMid76[5] , 
        \wBMid76[4] , \wBMid76[3] , \wBMid76[2] , \wBMid76[1] , \wBMid76[0] }), 
        .HiOut({\wRegInB76[31] , \wRegInB76[30] , \wRegInB76[29] , 
        \wRegInB76[28] , \wRegInB76[27] , \wRegInB76[26] , \wRegInB76[25] , 
        \wRegInB76[24] , \wRegInB76[23] , \wRegInB76[22] , \wRegInB76[21] , 
        \wRegInB76[20] , \wRegInB76[19] , \wRegInB76[18] , \wRegInB76[17] , 
        \wRegInB76[16] , \wRegInB76[15] , \wRegInB76[14] , \wRegInB76[13] , 
        \wRegInB76[12] , \wRegInB76[11] , \wRegInB76[10] , \wRegInB76[9] , 
        \wRegInB76[8] , \wRegInB76[7] , \wRegInB76[6] , \wRegInB76[5] , 
        \wRegInB76[4] , \wRegInB76[3] , \wRegInB76[2] , \wRegInB76[1] , 
        \wRegInB76[0] }), .LoOut({\wRegInA77[31] , \wRegInA77[30] , 
        \wRegInA77[29] , \wRegInA77[28] , \wRegInA77[27] , \wRegInA77[26] , 
        \wRegInA77[25] , \wRegInA77[24] , \wRegInA77[23] , \wRegInA77[22] , 
        \wRegInA77[21] , \wRegInA77[20] , \wRegInA77[19] , \wRegInA77[18] , 
        \wRegInA77[17] , \wRegInA77[16] , \wRegInA77[15] , \wRegInA77[14] , 
        \wRegInA77[13] , \wRegInA77[12] , \wRegInA77[11] , \wRegInA77[10] , 
        \wRegInA77[9] , \wRegInA77[8] , \wRegInA77[7] , \wRegInA77[6] , 
        \wRegInA77[5] , \wRegInA77[4] , \wRegInA77[3] , \wRegInA77[2] , 
        \wRegInA77[1] , \wRegInA77[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_13 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[31] , \ScanLink14[30] , \ScanLink14[29] , 
        \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , \ScanLink14[25] , 
        \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , \ScanLink14[21] , 
        \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , \ScanLink14[17] , 
        \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , \ScanLink14[13] , 
        \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , \ScanLink14[9] , 
        \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA121[31] , \wRegInA121[30] , 
        \wRegInA121[29] , \wRegInA121[28] , \wRegInA121[27] , \wRegInA121[26] , 
        \wRegInA121[25] , \wRegInA121[24] , \wRegInA121[23] , \wRegInA121[22] , 
        \wRegInA121[21] , \wRegInA121[20] , \wRegInA121[19] , \wRegInA121[18] , 
        \wRegInA121[17] , \wRegInA121[16] , \wRegInA121[15] , \wRegInA121[14] , 
        \wRegInA121[13] , \wRegInA121[12] , \wRegInA121[11] , \wRegInA121[10] , 
        \wRegInA121[9] , \wRegInA121[8] , \wRegInA121[7] , \wRegInA121[6] , 
        \wRegInA121[5] , \wRegInA121[4] , \wRegInA121[3] , \wRegInA121[2] , 
        \wRegInA121[1] , \wRegInA121[0] }), .Out({\wAIn121[31] , \wAIn121[30] , 
        \wAIn121[29] , \wAIn121[28] , \wAIn121[27] , \wAIn121[26] , 
        \wAIn121[25] , \wAIn121[24] , \wAIn121[23] , \wAIn121[22] , 
        \wAIn121[21] , \wAIn121[20] , \wAIn121[19] , \wAIn121[18] , 
        \wAIn121[17] , \wAIn121[16] , \wAIn121[15] , \wAIn121[14] , 
        \wAIn121[13] , \wAIn121[12] , \wAIn121[11] , \wAIn121[10] , 
        \wAIn121[9] , \wAIn121[8] , \wAIn121[7] , \wAIn121[6] , \wAIn121[5] , 
        \wAIn121[4] , \wAIn121[3] , \wAIn121[2] , \wAIn121[1] , \wAIn121[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_143 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink144[31] , \ScanLink144[30] , \ScanLink144[29] , 
        \ScanLink144[28] , \ScanLink144[27] , \ScanLink144[26] , 
        \ScanLink144[25] , \ScanLink144[24] , \ScanLink144[23] , 
        \ScanLink144[22] , \ScanLink144[21] , \ScanLink144[20] , 
        \ScanLink144[19] , \ScanLink144[18] , \ScanLink144[17] , 
        \ScanLink144[16] , \ScanLink144[15] , \ScanLink144[14] , 
        \ScanLink144[13] , \ScanLink144[12] , \ScanLink144[11] , 
        \ScanLink144[10] , \ScanLink144[9] , \ScanLink144[8] , 
        \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , \ScanLink144[4] , 
        \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , \ScanLink144[0] 
        }), .ScanOut({\ScanLink143[31] , \ScanLink143[30] , \ScanLink143[29] , 
        \ScanLink143[28] , \ScanLink143[27] , \ScanLink143[26] , 
        \ScanLink143[25] , \ScanLink143[24] , \ScanLink143[23] , 
        \ScanLink143[22] , \ScanLink143[21] , \ScanLink143[20] , 
        \ScanLink143[19] , \ScanLink143[18] , \ScanLink143[17] , 
        \ScanLink143[16] , \ScanLink143[15] , \ScanLink143[14] , 
        \ScanLink143[13] , \ScanLink143[12] , \ScanLink143[11] , 
        \ScanLink143[10] , \ScanLink143[9] , \ScanLink143[8] , 
        \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , \ScanLink143[4] , 
        \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , \ScanLink143[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA56[31] , \wRegInA56[30] , \wRegInA56[29] , 
        \wRegInA56[28] , \wRegInA56[27] , \wRegInA56[26] , \wRegInA56[25] , 
        \wRegInA56[24] , \wRegInA56[23] , \wRegInA56[22] , \wRegInA56[21] , 
        \wRegInA56[20] , \wRegInA56[19] , \wRegInA56[18] , \wRegInA56[17] , 
        \wRegInA56[16] , \wRegInA56[15] , \wRegInA56[14] , \wRegInA56[13] , 
        \wRegInA56[12] , \wRegInA56[11] , \wRegInA56[10] , \wRegInA56[9] , 
        \wRegInA56[8] , \wRegInA56[7] , \wRegInA56[6] , \wRegInA56[5] , 
        \wRegInA56[4] , \wRegInA56[3] , \wRegInA56[2] , \wRegInA56[1] , 
        \wRegInA56[0] }), .Out({\wAIn56[31] , \wAIn56[30] , \wAIn56[29] , 
        \wAIn56[28] , \wAIn56[27] , \wAIn56[26] , \wAIn56[25] , \wAIn56[24] , 
        \wAIn56[23] , \wAIn56[22] , \wAIn56[21] , \wAIn56[20] , \wAIn56[19] , 
        \wAIn56[18] , \wAIn56[17] , \wAIn56[16] , \wAIn56[15] , \wAIn56[14] , 
        \wAIn56[13] , \wAIn56[12] , \wAIn56[11] , \wAIn56[10] , \wAIn56[9] , 
        \wAIn56[8] , \wAIn56[7] , \wAIn56[6] , \wAIn56[5] , \wAIn56[4] , 
        \wAIn56[3] , \wAIn56[2] , \wAIn56[1] , \wAIn56[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid88[31] , \wAMid88[30] , \wAMid88[29] , \wAMid88[28] , 
        \wAMid88[27] , \wAMid88[26] , \wAMid88[25] , \wAMid88[24] , 
        \wAMid88[23] , \wAMid88[22] , \wAMid88[21] , \wAMid88[20] , 
        \wAMid88[19] , \wAMid88[18] , \wAMid88[17] , \wAMid88[16] , 
        \wAMid88[15] , \wAMid88[14] , \wAMid88[13] , \wAMid88[12] , 
        \wAMid88[11] , \wAMid88[10] , \wAMid88[9] , \wAMid88[8] , \wAMid88[7] , 
        \wAMid88[6] , \wAMid88[5] , \wAMid88[4] , \wAMid88[3] , \wAMid88[2] , 
        \wAMid88[1] , \wAMid88[0] }), .BIn({\wBMid88[31] , \wBMid88[30] , 
        \wBMid88[29] , \wBMid88[28] , \wBMid88[27] , \wBMid88[26] , 
        \wBMid88[25] , \wBMid88[24] , \wBMid88[23] , \wBMid88[22] , 
        \wBMid88[21] , \wBMid88[20] , \wBMid88[19] , \wBMid88[18] , 
        \wBMid88[17] , \wBMid88[16] , \wBMid88[15] , \wBMid88[14] , 
        \wBMid88[13] , \wBMid88[12] , \wBMid88[11] , \wBMid88[10] , 
        \wBMid88[9] , \wBMid88[8] , \wBMid88[7] , \wBMid88[6] , \wBMid88[5] , 
        \wBMid88[4] , \wBMid88[3] , \wBMid88[2] , \wBMid88[1] , \wBMid88[0] }), 
        .HiOut({\wRegInB88[31] , \wRegInB88[30] , \wRegInB88[29] , 
        \wRegInB88[28] , \wRegInB88[27] , \wRegInB88[26] , \wRegInB88[25] , 
        \wRegInB88[24] , \wRegInB88[23] , \wRegInB88[22] , \wRegInB88[21] , 
        \wRegInB88[20] , \wRegInB88[19] , \wRegInB88[18] , \wRegInB88[17] , 
        \wRegInB88[16] , \wRegInB88[15] , \wRegInB88[14] , \wRegInB88[13] , 
        \wRegInB88[12] , \wRegInB88[11] , \wRegInB88[10] , \wRegInB88[9] , 
        \wRegInB88[8] , \wRegInB88[7] , \wRegInB88[6] , \wRegInB88[5] , 
        \wRegInB88[4] , \wRegInB88[3] , \wRegInB88[2] , \wRegInB88[1] , 
        \wRegInB88[0] }), .LoOut({\wRegInA89[31] , \wRegInA89[30] , 
        \wRegInA89[29] , \wRegInA89[28] , \wRegInA89[27] , \wRegInA89[26] , 
        \wRegInA89[25] , \wRegInA89[24] , \wRegInA89[23] , \wRegInA89[22] , 
        \wRegInA89[21] , \wRegInA89[20] , \wRegInA89[19] , \wRegInA89[18] , 
        \wRegInA89[17] , \wRegInA89[16] , \wRegInA89[15] , \wRegInA89[14] , 
        \wRegInA89[13] , \wRegInA89[12] , \wRegInA89[11] , \wRegInA89[10] , 
        \wRegInA89[9] , \wRegInA89[8] , \wRegInA89[7] , \wRegInA89[6] , 
        \wRegInA89[5] , \wRegInA89[4] , \wRegInA89[3] , \wRegInA89[2] , 
        \wRegInA89[1] , \wRegInA89[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid100[31] , \wAMid100[30] , \wAMid100[29] , \wAMid100[28] , 
        \wAMid100[27] , \wAMid100[26] , \wAMid100[25] , \wAMid100[24] , 
        \wAMid100[23] , \wAMid100[22] , \wAMid100[21] , \wAMid100[20] , 
        \wAMid100[19] , \wAMid100[18] , \wAMid100[17] , \wAMid100[16] , 
        \wAMid100[15] , \wAMid100[14] , \wAMid100[13] , \wAMid100[12] , 
        \wAMid100[11] , \wAMid100[10] , \wAMid100[9] , \wAMid100[8] , 
        \wAMid100[7] , \wAMid100[6] , \wAMid100[5] , \wAMid100[4] , 
        \wAMid100[3] , \wAMid100[2] , \wAMid100[1] , \wAMid100[0] }), .BIn({
        \wBMid100[31] , \wBMid100[30] , \wBMid100[29] , \wBMid100[28] , 
        \wBMid100[27] , \wBMid100[26] , \wBMid100[25] , \wBMid100[24] , 
        \wBMid100[23] , \wBMid100[22] , \wBMid100[21] , \wBMid100[20] , 
        \wBMid100[19] , \wBMid100[18] , \wBMid100[17] , \wBMid100[16] , 
        \wBMid100[15] , \wBMid100[14] , \wBMid100[13] , \wBMid100[12] , 
        \wBMid100[11] , \wBMid100[10] , \wBMid100[9] , \wBMid100[8] , 
        \wBMid100[7] , \wBMid100[6] , \wBMid100[5] , \wBMid100[4] , 
        \wBMid100[3] , \wBMid100[2] , \wBMid100[1] , \wBMid100[0] }), .HiOut({
        \wRegInB100[31] , \wRegInB100[30] , \wRegInB100[29] , \wRegInB100[28] , 
        \wRegInB100[27] , \wRegInB100[26] , \wRegInB100[25] , \wRegInB100[24] , 
        \wRegInB100[23] , \wRegInB100[22] , \wRegInB100[21] , \wRegInB100[20] , 
        \wRegInB100[19] , \wRegInB100[18] , \wRegInB100[17] , \wRegInB100[16] , 
        \wRegInB100[15] , \wRegInB100[14] , \wRegInB100[13] , \wRegInB100[12] , 
        \wRegInB100[11] , \wRegInB100[10] , \wRegInB100[9] , \wRegInB100[8] , 
        \wRegInB100[7] , \wRegInB100[6] , \wRegInB100[5] , \wRegInB100[4] , 
        \wRegInB100[3] , \wRegInB100[2] , \wRegInB100[1] , \wRegInB100[0] }), 
        .LoOut({\wRegInA101[31] , \wRegInA101[30] , \wRegInA101[29] , 
        \wRegInA101[28] , \wRegInA101[27] , \wRegInA101[26] , \wRegInA101[25] , 
        \wRegInA101[24] , \wRegInA101[23] , \wRegInA101[22] , \wRegInA101[21] , 
        \wRegInA101[20] , \wRegInA101[19] , \wRegInA101[18] , \wRegInA101[17] , 
        \wRegInA101[16] , \wRegInA101[15] , \wRegInA101[14] , \wRegInA101[13] , 
        \wRegInA101[12] , \wRegInA101[11] , \wRegInA101[10] , \wRegInA101[9] , 
        \wRegInA101[8] , \wRegInA101[7] , \wRegInA101[6] , \wRegInA101[5] , 
        \wRegInA101[4] , \wRegInA101[3] , \wRegInA101[2] , \wRegInA101[1] , 
        \wRegInA101[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_158 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink159[31] , \ScanLink159[30] , \ScanLink159[29] , 
        \ScanLink159[28] , \ScanLink159[27] , \ScanLink159[26] , 
        \ScanLink159[25] , \ScanLink159[24] , \ScanLink159[23] , 
        \ScanLink159[22] , \ScanLink159[21] , \ScanLink159[20] , 
        \ScanLink159[19] , \ScanLink159[18] , \ScanLink159[17] , 
        \ScanLink159[16] , \ScanLink159[15] , \ScanLink159[14] , 
        \ScanLink159[13] , \ScanLink159[12] , \ScanLink159[11] , 
        \ScanLink159[10] , \ScanLink159[9] , \ScanLink159[8] , 
        \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , \ScanLink159[4] , 
        \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , \ScanLink159[0] 
        }), .ScanOut({\ScanLink158[31] , \ScanLink158[30] , \ScanLink158[29] , 
        \ScanLink158[28] , \ScanLink158[27] , \ScanLink158[26] , 
        \ScanLink158[25] , \ScanLink158[24] , \ScanLink158[23] , 
        \ScanLink158[22] , \ScanLink158[21] , \ScanLink158[20] , 
        \ScanLink158[19] , \ScanLink158[18] , \ScanLink158[17] , 
        \ScanLink158[16] , \ScanLink158[15] , \ScanLink158[14] , 
        \ScanLink158[13] , \ScanLink158[12] , \ScanLink158[11] , 
        \ScanLink158[10] , \ScanLink158[9] , \ScanLink158[8] , 
        \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , \ScanLink158[4] , 
        \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , \ScanLink158[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB48[31] , \wRegInB48[30] , \wRegInB48[29] , 
        \wRegInB48[28] , \wRegInB48[27] , \wRegInB48[26] , \wRegInB48[25] , 
        \wRegInB48[24] , \wRegInB48[23] , \wRegInB48[22] , \wRegInB48[21] , 
        \wRegInB48[20] , \wRegInB48[19] , \wRegInB48[18] , \wRegInB48[17] , 
        \wRegInB48[16] , \wRegInB48[15] , \wRegInB48[14] , \wRegInB48[13] , 
        \wRegInB48[12] , \wRegInB48[11] , \wRegInB48[10] , \wRegInB48[9] , 
        \wRegInB48[8] , \wRegInB48[7] , \wRegInB48[6] , \wRegInB48[5] , 
        \wRegInB48[4] , \wRegInB48[3] , \wRegInB48[2] , \wRegInB48[1] , 
        \wRegInB48[0] }), .Out({\wBIn48[31] , \wBIn48[30] , \wBIn48[29] , 
        \wBIn48[28] , \wBIn48[27] , \wBIn48[26] , \wBIn48[25] , \wBIn48[24] , 
        \wBIn48[23] , \wBIn48[22] , \wBIn48[21] , \wBIn48[20] , \wBIn48[19] , 
        \wBIn48[18] , \wBIn48[17] , \wBIn48[16] , \wBIn48[15] , \wBIn48[14] , 
        \wBIn48[13] , \wBIn48[12] , \wBIn48[11] , \wBIn48[10] , \wBIn48[9] , 
        \wBIn48[8] , \wBIn48[7] , \wBIn48[6] , \wBIn48[5] , \wBIn48[4] , 
        \wBIn48[3] , \wBIn48[2] , \wBIn48[1] , \wBIn48[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_83 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink84[31] , \ScanLink84[30] , \ScanLink84[29] , 
        \ScanLink84[28] , \ScanLink84[27] , \ScanLink84[26] , \ScanLink84[25] , 
        \ScanLink84[24] , \ScanLink84[23] , \ScanLink84[22] , \ScanLink84[21] , 
        \ScanLink84[20] , \ScanLink84[19] , \ScanLink84[18] , \ScanLink84[17] , 
        \ScanLink84[16] , \ScanLink84[15] , \ScanLink84[14] , \ScanLink84[13] , 
        \ScanLink84[12] , \ScanLink84[11] , \ScanLink84[10] , \ScanLink84[9] , 
        \ScanLink84[8] , \ScanLink84[7] , \ScanLink84[6] , \ScanLink84[5] , 
        \ScanLink84[4] , \ScanLink84[3] , \ScanLink84[2] , \ScanLink84[1] , 
        \ScanLink84[0] }), .ScanOut({\ScanLink83[31] , \ScanLink83[30] , 
        \ScanLink83[29] , \ScanLink83[28] , \ScanLink83[27] , \ScanLink83[26] , 
        \ScanLink83[25] , \ScanLink83[24] , \ScanLink83[23] , \ScanLink83[22] , 
        \ScanLink83[21] , \ScanLink83[20] , \ScanLink83[19] , \ScanLink83[18] , 
        \ScanLink83[17] , \ScanLink83[16] , \ScanLink83[15] , \ScanLink83[14] , 
        \ScanLink83[13] , \ScanLink83[12] , \ScanLink83[11] , \ScanLink83[10] , 
        \ScanLink83[9] , \ScanLink83[8] , \ScanLink83[7] , \ScanLink83[6] , 
        \ScanLink83[5] , \ScanLink83[4] , \ScanLink83[3] , \ScanLink83[2] , 
        \ScanLink83[1] , \ScanLink83[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA86[31] , \wRegInA86[30] , 
        \wRegInA86[29] , \wRegInA86[28] , \wRegInA86[27] , \wRegInA86[26] , 
        \wRegInA86[25] , \wRegInA86[24] , \wRegInA86[23] , \wRegInA86[22] , 
        \wRegInA86[21] , \wRegInA86[20] , \wRegInA86[19] , \wRegInA86[18] , 
        \wRegInA86[17] , \wRegInA86[16] , \wRegInA86[15] , \wRegInA86[14] , 
        \wRegInA86[13] , \wRegInA86[12] , \wRegInA86[11] , \wRegInA86[10] , 
        \wRegInA86[9] , \wRegInA86[8] , \wRegInA86[7] , \wRegInA86[6] , 
        \wRegInA86[5] , \wRegInA86[4] , \wRegInA86[3] , \wRegInA86[2] , 
        \wRegInA86[1] , \wRegInA86[0] }), .Out({\wAIn86[31] , \wAIn86[30] , 
        \wAIn86[29] , \wAIn86[28] , \wAIn86[27] , \wAIn86[26] , \wAIn86[25] , 
        \wAIn86[24] , \wAIn86[23] , \wAIn86[22] , \wAIn86[21] , \wAIn86[20] , 
        \wAIn86[19] , \wAIn86[18] , \wAIn86[17] , \wAIn86[16] , \wAIn86[15] , 
        \wAIn86[14] , \wAIn86[13] , \wAIn86[12] , \wAIn86[11] , \wAIn86[10] , 
        \wAIn86[9] , \wAIn86[8] , \wAIn86[7] , \wAIn86[6] , \wAIn86[5] , 
        \wAIn86[4] , \wAIn86[3] , \wAIn86[2] , \wAIn86[1] , \wAIn86[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_221 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink222[31] , \ScanLink222[30] , \ScanLink222[29] , 
        \ScanLink222[28] , \ScanLink222[27] , \ScanLink222[26] , 
        \ScanLink222[25] , \ScanLink222[24] , \ScanLink222[23] , 
        \ScanLink222[22] , \ScanLink222[21] , \ScanLink222[20] , 
        \ScanLink222[19] , \ScanLink222[18] , \ScanLink222[17] , 
        \ScanLink222[16] , \ScanLink222[15] , \ScanLink222[14] , 
        \ScanLink222[13] , \ScanLink222[12] , \ScanLink222[11] , 
        \ScanLink222[10] , \ScanLink222[9] , \ScanLink222[8] , 
        \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , \ScanLink222[4] , 
        \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , \ScanLink222[0] 
        }), .ScanOut({\ScanLink221[31] , \ScanLink221[30] , \ScanLink221[29] , 
        \ScanLink221[28] , \ScanLink221[27] , \ScanLink221[26] , 
        \ScanLink221[25] , \ScanLink221[24] , \ScanLink221[23] , 
        \ScanLink221[22] , \ScanLink221[21] , \ScanLink221[20] , 
        \ScanLink221[19] , \ScanLink221[18] , \ScanLink221[17] , 
        \ScanLink221[16] , \ScanLink221[15] , \ScanLink221[14] , 
        \ScanLink221[13] , \ScanLink221[12] , \ScanLink221[11] , 
        \ScanLink221[10] , \ScanLink221[9] , \ScanLink221[8] , 
        \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , \ScanLink221[4] , 
        \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , \ScanLink221[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA17[31] , \wRegInA17[30] , \wRegInA17[29] , 
        \wRegInA17[28] , \wRegInA17[27] , \wRegInA17[26] , \wRegInA17[25] , 
        \wRegInA17[24] , \wRegInA17[23] , \wRegInA17[22] , \wRegInA17[21] , 
        \wRegInA17[20] , \wRegInA17[19] , \wRegInA17[18] , \wRegInA17[17] , 
        \wRegInA17[16] , \wRegInA17[15] , \wRegInA17[14] , \wRegInA17[13] , 
        \wRegInA17[12] , \wRegInA17[11] , \wRegInA17[10] , \wRegInA17[9] , 
        \wRegInA17[8] , \wRegInA17[7] , \wRegInA17[6] , \wRegInA17[5] , 
        \wRegInA17[4] , \wRegInA17[3] , \wRegInA17[2] , \wRegInA17[1] , 
        \wRegInA17[0] }), .Out({\wAIn17[31] , \wAIn17[30] , \wAIn17[29] , 
        \wAIn17[28] , \wAIn17[27] , \wAIn17[26] , \wAIn17[25] , \wAIn17[24] , 
        \wAIn17[23] , \wAIn17[22] , \wAIn17[21] , \wAIn17[20] , \wAIn17[19] , 
        \wAIn17[18] , \wAIn17[17] , \wAIn17[16] , \wAIn17[15] , \wAIn17[14] , 
        \wAIn17[13] , \wAIn17[12] , \wAIn17[11] , \wAIn17[10] , \wAIn17[9] , 
        \wAIn17[8] , \wAIn17[7] , \wAIn17[6] , \wAIn17[5] , \wAIn17[4] , 
        \wAIn17[3] , \wAIn17[2] , \wAIn17[1] , \wAIn17[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn33[31] , \wAIn33[30] , \wAIn33[29] , \wAIn33[28] , \wAIn33[27] , 
        \wAIn33[26] , \wAIn33[25] , \wAIn33[24] , \wAIn33[23] , \wAIn33[22] , 
        \wAIn33[21] , \wAIn33[20] , \wAIn33[19] , \wAIn33[18] , \wAIn33[17] , 
        \wAIn33[16] , \wAIn33[15] , \wAIn33[14] , \wAIn33[13] , \wAIn33[12] , 
        \wAIn33[11] , \wAIn33[10] , \wAIn33[9] , \wAIn33[8] , \wAIn33[7] , 
        \wAIn33[6] , \wAIn33[5] , \wAIn33[4] , \wAIn33[3] , \wAIn33[2] , 
        \wAIn33[1] , \wAIn33[0] }), .BIn({\wBIn33[31] , \wBIn33[30] , 
        \wBIn33[29] , \wBIn33[28] , \wBIn33[27] , \wBIn33[26] , \wBIn33[25] , 
        \wBIn33[24] , \wBIn33[23] , \wBIn33[22] , \wBIn33[21] , \wBIn33[20] , 
        \wBIn33[19] , \wBIn33[18] , \wBIn33[17] , \wBIn33[16] , \wBIn33[15] , 
        \wBIn33[14] , \wBIn33[13] , \wBIn33[12] , \wBIn33[11] , \wBIn33[10] , 
        \wBIn33[9] , \wBIn33[8] , \wBIn33[7] , \wBIn33[6] , \wBIn33[5] , 
        \wBIn33[4] , \wBIn33[3] , \wBIn33[2] , \wBIn33[1] , \wBIn33[0] }), 
        .HiOut({\wBMid32[31] , \wBMid32[30] , \wBMid32[29] , \wBMid32[28] , 
        \wBMid32[27] , \wBMid32[26] , \wBMid32[25] , \wBMid32[24] , 
        \wBMid32[23] , \wBMid32[22] , \wBMid32[21] , \wBMid32[20] , 
        \wBMid32[19] , \wBMid32[18] , \wBMid32[17] , \wBMid32[16] , 
        \wBMid32[15] , \wBMid32[14] , \wBMid32[13] , \wBMid32[12] , 
        \wBMid32[11] , \wBMid32[10] , \wBMid32[9] , \wBMid32[8] , \wBMid32[7] , 
        \wBMid32[6] , \wBMid32[5] , \wBMid32[4] , \wBMid32[3] , \wBMid32[2] , 
        \wBMid32[1] , \wBMid32[0] }), .LoOut({\wAMid33[31] , \wAMid33[30] , 
        \wAMid33[29] , \wAMid33[28] , \wAMid33[27] , \wAMid33[26] , 
        \wAMid33[25] , \wAMid33[24] , \wAMid33[23] , \wAMid33[22] , 
        \wAMid33[21] , \wAMid33[20] , \wAMid33[19] , \wAMid33[18] , 
        \wAMid33[17] , \wAMid33[16] , \wAMid33[15] , \wAMid33[14] , 
        \wAMid33[13] , \wAMid33[12] , \wAMid33[11] , \wAMid33[10] , 
        \wAMid33[9] , \wAMid33[8] , \wAMid33[7] , \wAMid33[6] , \wAMid33[5] , 
        \wAMid33[4] , \wAMid33[3] , \wAMid33[2] , \wAMid33[1] , \wAMid33[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid24[31] , \wAMid24[30] , \wAMid24[29] , \wAMid24[28] , 
        \wAMid24[27] , \wAMid24[26] , \wAMid24[25] , \wAMid24[24] , 
        \wAMid24[23] , \wAMid24[22] , \wAMid24[21] , \wAMid24[20] , 
        \wAMid24[19] , \wAMid24[18] , \wAMid24[17] , \wAMid24[16] , 
        \wAMid24[15] , \wAMid24[14] , \wAMid24[13] , \wAMid24[12] , 
        \wAMid24[11] , \wAMid24[10] , \wAMid24[9] , \wAMid24[8] , \wAMid24[7] , 
        \wAMid24[6] , \wAMid24[5] , \wAMid24[4] , \wAMid24[3] , \wAMid24[2] , 
        \wAMid24[1] , \wAMid24[0] }), .BIn({\wBMid24[31] , \wBMid24[30] , 
        \wBMid24[29] , \wBMid24[28] , \wBMid24[27] , \wBMid24[26] , 
        \wBMid24[25] , \wBMid24[24] , \wBMid24[23] , \wBMid24[22] , 
        \wBMid24[21] , \wBMid24[20] , \wBMid24[19] , \wBMid24[18] , 
        \wBMid24[17] , \wBMid24[16] , \wBMid24[15] , \wBMid24[14] , 
        \wBMid24[13] , \wBMid24[12] , \wBMid24[11] , \wBMid24[10] , 
        \wBMid24[9] , \wBMid24[8] , \wBMid24[7] , \wBMid24[6] , \wBMid24[5] , 
        \wBMid24[4] , \wBMid24[3] , \wBMid24[2] , \wBMid24[1] , \wBMid24[0] }), 
        .HiOut({\wRegInB24[31] , \wRegInB24[30] , \wRegInB24[29] , 
        \wRegInB24[28] , \wRegInB24[27] , \wRegInB24[26] , \wRegInB24[25] , 
        \wRegInB24[24] , \wRegInB24[23] , \wRegInB24[22] , \wRegInB24[21] , 
        \wRegInB24[20] , \wRegInB24[19] , \wRegInB24[18] , \wRegInB24[17] , 
        \wRegInB24[16] , \wRegInB24[15] , \wRegInB24[14] , \wRegInB24[13] , 
        \wRegInB24[12] , \wRegInB24[11] , \wRegInB24[10] , \wRegInB24[9] , 
        \wRegInB24[8] , \wRegInB24[7] , \wRegInB24[6] , \wRegInB24[5] , 
        \wRegInB24[4] , \wRegInB24[3] , \wRegInB24[2] , \wRegInB24[1] , 
        \wRegInB24[0] }), .LoOut({\wRegInA25[31] , \wRegInA25[30] , 
        \wRegInA25[29] , \wRegInA25[28] , \wRegInA25[27] , \wRegInA25[26] , 
        \wRegInA25[25] , \wRegInA25[24] , \wRegInA25[23] , \wRegInA25[22] , 
        \wRegInA25[21] , \wRegInA25[20] , \wRegInA25[19] , \wRegInA25[18] , 
        \wRegInA25[17] , \wRegInA25[16] , \wRegInA25[15] , \wRegInA25[14] , 
        \wRegInA25[13] , \wRegInA25[12] , \wRegInA25[11] , \wRegInA25[10] , 
        \wRegInA25[9] , \wRegInA25[8] , \wRegInA25[7] , \wRegInA25[6] , 
        \wRegInA25[5] , \wRegInA25[4] , \wRegInA25[3] , \wRegInA25[2] , 
        \wRegInA25[1] , \wRegInA25[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_111 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink112[31] , \ScanLink112[30] , \ScanLink112[29] , 
        \ScanLink112[28] , \ScanLink112[27] , \ScanLink112[26] , 
        \ScanLink112[25] , \ScanLink112[24] , \ScanLink112[23] , 
        \ScanLink112[22] , \ScanLink112[21] , \ScanLink112[20] , 
        \ScanLink112[19] , \ScanLink112[18] , \ScanLink112[17] , 
        \ScanLink112[16] , \ScanLink112[15] , \ScanLink112[14] , 
        \ScanLink112[13] , \ScanLink112[12] , \ScanLink112[11] , 
        \ScanLink112[10] , \ScanLink112[9] , \ScanLink112[8] , 
        \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , \ScanLink112[4] , 
        \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , \ScanLink112[0] 
        }), .ScanOut({\ScanLink111[31] , \ScanLink111[30] , \ScanLink111[29] , 
        \ScanLink111[28] , \ScanLink111[27] , \ScanLink111[26] , 
        \ScanLink111[25] , \ScanLink111[24] , \ScanLink111[23] , 
        \ScanLink111[22] , \ScanLink111[21] , \ScanLink111[20] , 
        \ScanLink111[19] , \ScanLink111[18] , \ScanLink111[17] , 
        \ScanLink111[16] , \ScanLink111[15] , \ScanLink111[14] , 
        \ScanLink111[13] , \ScanLink111[12] , \ScanLink111[11] , 
        \ScanLink111[10] , \ScanLink111[9] , \ScanLink111[8] , 
        \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , \ScanLink111[4] , 
        \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , \ScanLink111[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA72[31] , \wRegInA72[30] , \wRegInA72[29] , 
        \wRegInA72[28] , \wRegInA72[27] , \wRegInA72[26] , \wRegInA72[25] , 
        \wRegInA72[24] , \wRegInA72[23] , \wRegInA72[22] , \wRegInA72[21] , 
        \wRegInA72[20] , \wRegInA72[19] , \wRegInA72[18] , \wRegInA72[17] , 
        \wRegInA72[16] , \wRegInA72[15] , \wRegInA72[14] , \wRegInA72[13] , 
        \wRegInA72[12] , \wRegInA72[11] , \wRegInA72[10] , \wRegInA72[9] , 
        \wRegInA72[8] , \wRegInA72[7] , \wRegInA72[6] , \wRegInA72[5] , 
        \wRegInA72[4] , \wRegInA72[3] , \wRegInA72[2] , \wRegInA72[1] , 
        \wRegInA72[0] }), .Out({\wAIn72[31] , \wAIn72[30] , \wAIn72[29] , 
        \wAIn72[28] , \wAIn72[27] , \wAIn72[26] , \wAIn72[25] , \wAIn72[24] , 
        \wAIn72[23] , \wAIn72[22] , \wAIn72[21] , \wAIn72[20] , \wAIn72[19] , 
        \wAIn72[18] , \wAIn72[17] , \wAIn72[16] , \wAIn72[15] , \wAIn72[14] , 
        \wAIn72[13] , \wAIn72[12] , \wAIn72[11] , \wAIn72[10] , \wAIn72[9] , 
        \wAIn72[8] , \wAIn72[7] , \wAIn72[6] , \wAIn72[5] , \wAIn72[4] , 
        \wAIn72[3] , \wAIn72[2] , \wAIn72[1] , \wAIn72[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_41 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink42[31] , \ScanLink42[30] , \ScanLink42[29] , 
        \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , \ScanLink42[25] , 
        \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , \ScanLink42[21] , 
        \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , \ScanLink42[17] , 
        \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , \ScanLink42[13] , 
        \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , \ScanLink42[9] , 
        \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , \ScanLink42[5] , 
        \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , \ScanLink42[1] , 
        \ScanLink42[0] }), .ScanOut({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA107[31] , \wRegInA107[30] , 
        \wRegInA107[29] , \wRegInA107[28] , \wRegInA107[27] , \wRegInA107[26] , 
        \wRegInA107[25] , \wRegInA107[24] , \wRegInA107[23] , \wRegInA107[22] , 
        \wRegInA107[21] , \wRegInA107[20] , \wRegInA107[19] , \wRegInA107[18] , 
        \wRegInA107[17] , \wRegInA107[16] , \wRegInA107[15] , \wRegInA107[14] , 
        \wRegInA107[13] , \wRegInA107[12] , \wRegInA107[11] , \wRegInA107[10] , 
        \wRegInA107[9] , \wRegInA107[8] , \wRegInA107[7] , \wRegInA107[6] , 
        \wRegInA107[5] , \wRegInA107[4] , \wRegInA107[3] , \wRegInA107[2] , 
        \wRegInA107[1] , \wRegInA107[0] }), .Out({\wAIn107[31] , \wAIn107[30] , 
        \wAIn107[29] , \wAIn107[28] , \wAIn107[27] , \wAIn107[26] , 
        \wAIn107[25] , \wAIn107[24] , \wAIn107[23] , \wAIn107[22] , 
        \wAIn107[21] , \wAIn107[20] , \wAIn107[19] , \wAIn107[18] , 
        \wAIn107[17] , \wAIn107[16] , \wAIn107[15] , \wAIn107[14] , 
        \wAIn107[13] , \wAIn107[12] , \wAIn107[11] , \wAIn107[10] , 
        \wAIn107[9] , \wAIn107[8] , \wAIn107[7] , \wAIn107[6] , \wAIn107[5] , 
        \wAIn107[4] , \wAIn107[3] , \wAIn107[2] , \wAIn107[1] , \wAIn107[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn34[31] , \wAIn34[30] , \wAIn34[29] , \wAIn34[28] , \wAIn34[27] , 
        \wAIn34[26] , \wAIn34[25] , \wAIn34[24] , \wAIn34[23] , \wAIn34[22] , 
        \wAIn34[21] , \wAIn34[20] , \wAIn34[19] , \wAIn34[18] , \wAIn34[17] , 
        \wAIn34[16] , \wAIn34[15] , \wAIn34[14] , \wAIn34[13] , \wAIn34[12] , 
        \wAIn34[11] , \wAIn34[10] , \wAIn34[9] , \wAIn34[8] , \wAIn34[7] , 
        \wAIn34[6] , \wAIn34[5] , \wAIn34[4] , \wAIn34[3] , \wAIn34[2] , 
        \wAIn34[1] , \wAIn34[0] }), .BIn({\wBIn34[31] , \wBIn34[30] , 
        \wBIn34[29] , \wBIn34[28] , \wBIn34[27] , \wBIn34[26] , \wBIn34[25] , 
        \wBIn34[24] , \wBIn34[23] , \wBIn34[22] , \wBIn34[21] , \wBIn34[20] , 
        \wBIn34[19] , \wBIn34[18] , \wBIn34[17] , \wBIn34[16] , \wBIn34[15] , 
        \wBIn34[14] , \wBIn34[13] , \wBIn34[12] , \wBIn34[11] , \wBIn34[10] , 
        \wBIn34[9] , \wBIn34[8] , \wBIn34[7] , \wBIn34[6] , \wBIn34[5] , 
        \wBIn34[4] , \wBIn34[3] , \wBIn34[2] , \wBIn34[1] , \wBIn34[0] }), 
        .HiOut({\wBMid33[31] , \wBMid33[30] , \wBMid33[29] , \wBMid33[28] , 
        \wBMid33[27] , \wBMid33[26] , \wBMid33[25] , \wBMid33[24] , 
        \wBMid33[23] , \wBMid33[22] , \wBMid33[21] , \wBMid33[20] , 
        \wBMid33[19] , \wBMid33[18] , \wBMid33[17] , \wBMid33[16] , 
        \wBMid33[15] , \wBMid33[14] , \wBMid33[13] , \wBMid33[12] , 
        \wBMid33[11] , \wBMid33[10] , \wBMid33[9] , \wBMid33[8] , \wBMid33[7] , 
        \wBMid33[6] , \wBMid33[5] , \wBMid33[4] , \wBMid33[3] , \wBMid33[2] , 
        \wBMid33[1] , \wBMid33[0] }), .LoOut({\wAMid34[31] , \wAMid34[30] , 
        \wAMid34[29] , \wAMid34[28] , \wAMid34[27] , \wAMid34[26] , 
        \wAMid34[25] , \wAMid34[24] , \wAMid34[23] , \wAMid34[22] , 
        \wAMid34[21] , \wAMid34[20] , \wAMid34[19] , \wAMid34[18] , 
        \wAMid34[17] , \wAMid34[16] , \wAMid34[15] , \wAMid34[14] , 
        \wAMid34[13] , \wAMid34[12] , \wAMid34[11] , \wAMid34[10] , 
        \wAMid34[9] , \wAMid34[8] , \wAMid34[7] , \wAMid34[6] , \wAMid34[5] , 
        \wAMid34[4] , \wAMid34[3] , \wAMid34[2] , \wAMid34[1] , \wAMid34[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn98[31] , \wAIn98[30] , \wAIn98[29] , \wAIn98[28] , \wAIn98[27] , 
        \wAIn98[26] , \wAIn98[25] , \wAIn98[24] , \wAIn98[23] , \wAIn98[22] , 
        \wAIn98[21] , \wAIn98[20] , \wAIn98[19] , \wAIn98[18] , \wAIn98[17] , 
        \wAIn98[16] , \wAIn98[15] , \wAIn98[14] , \wAIn98[13] , \wAIn98[12] , 
        \wAIn98[11] , \wAIn98[10] , \wAIn98[9] , \wAIn98[8] , \wAIn98[7] , 
        \wAIn98[6] , \wAIn98[5] , \wAIn98[4] , \wAIn98[3] , \wAIn98[2] , 
        \wAIn98[1] , \wAIn98[0] }), .BIn({\wBIn98[31] , \wBIn98[30] , 
        \wBIn98[29] , \wBIn98[28] , \wBIn98[27] , \wBIn98[26] , \wBIn98[25] , 
        \wBIn98[24] , \wBIn98[23] , \wBIn98[22] , \wBIn98[21] , \wBIn98[20] , 
        \wBIn98[19] , \wBIn98[18] , \wBIn98[17] , \wBIn98[16] , \wBIn98[15] , 
        \wBIn98[14] , \wBIn98[13] , \wBIn98[12] , \wBIn98[11] , \wBIn98[10] , 
        \wBIn98[9] , \wBIn98[8] , \wBIn98[7] , \wBIn98[6] , \wBIn98[5] , 
        \wBIn98[4] , \wBIn98[3] , \wBIn98[2] , \wBIn98[1] , \wBIn98[0] }), 
        .HiOut({\wBMid97[31] , \wBMid97[30] , \wBMid97[29] , \wBMid97[28] , 
        \wBMid97[27] , \wBMid97[26] , \wBMid97[25] , \wBMid97[24] , 
        \wBMid97[23] , \wBMid97[22] , \wBMid97[21] , \wBMid97[20] , 
        \wBMid97[19] , \wBMid97[18] , \wBMid97[17] , \wBMid97[16] , 
        \wBMid97[15] , \wBMid97[14] , \wBMid97[13] , \wBMid97[12] , 
        \wBMid97[11] , \wBMid97[10] , \wBMid97[9] , \wBMid97[8] , \wBMid97[7] , 
        \wBMid97[6] , \wBMid97[5] , \wBMid97[4] , \wBMid97[3] , \wBMid97[2] , 
        \wBMid97[1] , \wBMid97[0] }), .LoOut({\wAMid98[31] , \wAMid98[30] , 
        \wAMid98[29] , \wAMid98[28] , \wAMid98[27] , \wAMid98[26] , 
        \wAMid98[25] , \wAMid98[24] , \wAMid98[23] , \wAMid98[22] , 
        \wAMid98[21] , \wAMid98[20] , \wAMid98[19] , \wAMid98[18] , 
        \wAMid98[17] , \wAMid98[16] , \wAMid98[15] , \wAMid98[14] , 
        \wAMid98[13] , \wAMid98[12] , \wAMid98[11] , \wAMid98[10] , 
        \wAMid98[9] , \wAMid98[8] , \wAMid98[7] , \wAMid98[6] , \wAMid98[5] , 
        \wAMid98[4] , \wAMid98[3] , \wAMid98[2] , \wAMid98[1] , \wAMid98[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_206 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink207[31] , \ScanLink207[30] , \ScanLink207[29] , 
        \ScanLink207[28] , \ScanLink207[27] , \ScanLink207[26] , 
        \ScanLink207[25] , \ScanLink207[24] , \ScanLink207[23] , 
        \ScanLink207[22] , \ScanLink207[21] , \ScanLink207[20] , 
        \ScanLink207[19] , \ScanLink207[18] , \ScanLink207[17] , 
        \ScanLink207[16] , \ScanLink207[15] , \ScanLink207[14] , 
        \ScanLink207[13] , \ScanLink207[12] , \ScanLink207[11] , 
        \ScanLink207[10] , \ScanLink207[9] , \ScanLink207[8] , 
        \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , \ScanLink207[4] , 
        \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , \ScanLink207[0] 
        }), .ScanOut({\ScanLink206[31] , \ScanLink206[30] , \ScanLink206[29] , 
        \ScanLink206[28] , \ScanLink206[27] , \ScanLink206[26] , 
        \ScanLink206[25] , \ScanLink206[24] , \ScanLink206[23] , 
        \ScanLink206[22] , \ScanLink206[21] , \ScanLink206[20] , 
        \ScanLink206[19] , \ScanLink206[18] , \ScanLink206[17] , 
        \ScanLink206[16] , \ScanLink206[15] , \ScanLink206[14] , 
        \ScanLink206[13] , \ScanLink206[12] , \ScanLink206[11] , 
        \ScanLink206[10] , \ScanLink206[9] , \ScanLink206[8] , 
        \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , \ScanLink206[4] , 
        \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , \ScanLink206[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB24[31] , \wRegInB24[30] , \wRegInB24[29] , 
        \wRegInB24[28] , \wRegInB24[27] , \wRegInB24[26] , \wRegInB24[25] , 
        \wRegInB24[24] , \wRegInB24[23] , \wRegInB24[22] , \wRegInB24[21] , 
        \wRegInB24[20] , \wRegInB24[19] , \wRegInB24[18] , \wRegInB24[17] , 
        \wRegInB24[16] , \wRegInB24[15] , \wRegInB24[14] , \wRegInB24[13] , 
        \wRegInB24[12] , \wRegInB24[11] , \wRegInB24[10] , \wRegInB24[9] , 
        \wRegInB24[8] , \wRegInB24[7] , \wRegInB24[6] , \wRegInB24[5] , 
        \wRegInB24[4] , \wRegInB24[3] , \wRegInB24[2] , \wRegInB24[1] , 
        \wRegInB24[0] }), .Out({\wBIn24[31] , \wBIn24[30] , \wBIn24[29] , 
        \wBIn24[28] , \wBIn24[27] , \wBIn24[26] , \wBIn24[25] , \wBIn24[24] , 
        \wBIn24[23] , \wBIn24[22] , \wBIn24[21] , \wBIn24[20] , \wBIn24[19] , 
        \wBIn24[18] , \wBIn24[17] , \wBIn24[16] , \wBIn24[15] , \wBIn24[14] , 
        \wBIn24[13] , \wBIn24[12] , \wBIn24[11] , \wBIn24[10] , \wBIn24[9] , 
        \wBIn24[8] , \wBIn24[7] , \wBIn24[6] , \wBIn24[5] , \wBIn24[4] , 
        \wBIn24[3] , \wBIn24[2] , \wBIn24[1] , \wBIn24[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_136 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink137[31] , \ScanLink137[30] , \ScanLink137[29] , 
        \ScanLink137[28] , \ScanLink137[27] , \ScanLink137[26] , 
        \ScanLink137[25] , \ScanLink137[24] , \ScanLink137[23] , 
        \ScanLink137[22] , \ScanLink137[21] , \ScanLink137[20] , 
        \ScanLink137[19] , \ScanLink137[18] , \ScanLink137[17] , 
        \ScanLink137[16] , \ScanLink137[15] , \ScanLink137[14] , 
        \ScanLink137[13] , \ScanLink137[12] , \ScanLink137[11] , 
        \ScanLink137[10] , \ScanLink137[9] , \ScanLink137[8] , 
        \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , \ScanLink137[4] , 
        \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , \ScanLink137[0] 
        }), .ScanOut({\ScanLink136[31] , \ScanLink136[30] , \ScanLink136[29] , 
        \ScanLink136[28] , \ScanLink136[27] , \ScanLink136[26] , 
        \ScanLink136[25] , \ScanLink136[24] , \ScanLink136[23] , 
        \ScanLink136[22] , \ScanLink136[21] , \ScanLink136[20] , 
        \ScanLink136[19] , \ScanLink136[18] , \ScanLink136[17] , 
        \ScanLink136[16] , \ScanLink136[15] , \ScanLink136[14] , 
        \ScanLink136[13] , \ScanLink136[12] , \ScanLink136[11] , 
        \ScanLink136[10] , \ScanLink136[9] , \ScanLink136[8] , 
        \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , \ScanLink136[4] , 
        \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , \ScanLink136[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB59[31] , \wRegInB59[30] , \wRegInB59[29] , 
        \wRegInB59[28] , \wRegInB59[27] , \wRegInB59[26] , \wRegInB59[25] , 
        \wRegInB59[24] , \wRegInB59[23] , \wRegInB59[22] , \wRegInB59[21] , 
        \wRegInB59[20] , \wRegInB59[19] , \wRegInB59[18] , \wRegInB59[17] , 
        \wRegInB59[16] , \wRegInB59[15] , \wRegInB59[14] , \wRegInB59[13] , 
        \wRegInB59[12] , \wRegInB59[11] , \wRegInB59[10] , \wRegInB59[9] , 
        \wRegInB59[8] , \wRegInB59[7] , \wRegInB59[6] , \wRegInB59[5] , 
        \wRegInB59[4] , \wRegInB59[3] , \wRegInB59[2] , \wRegInB59[1] , 
        \wRegInB59[0] }), .Out({\wBIn59[31] , \wBIn59[30] , \wBIn59[29] , 
        \wBIn59[28] , \wBIn59[27] , \wBIn59[26] , \wBIn59[25] , \wBIn59[24] , 
        \wBIn59[23] , \wBIn59[22] , \wBIn59[21] , \wBIn59[20] , \wBIn59[19] , 
        \wBIn59[18] , \wBIn59[17] , \wBIn59[16] , \wBIn59[15] , \wBIn59[14] , 
        \wBIn59[13] , \wBIn59[12] , \wBIn59[11] , \wBIn59[10] , \wBIn59[9] , 
        \wBIn59[8] , \wBIn59[7] , \wBIn59[6] , \wBIn59[5] , \wBIn59[4] , 
        \wBIn59[3] , \wBIn59[2] , \wBIn59[1] , \wBIn59[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_66 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink67[31] , \ScanLink67[30] , \ScanLink67[29] , 
        \ScanLink67[28] , \ScanLink67[27] , \ScanLink67[26] , \ScanLink67[25] , 
        \ScanLink67[24] , \ScanLink67[23] , \ScanLink67[22] , \ScanLink67[21] , 
        \ScanLink67[20] , \ScanLink67[19] , \ScanLink67[18] , \ScanLink67[17] , 
        \ScanLink67[16] , \ScanLink67[15] , \ScanLink67[14] , \ScanLink67[13] , 
        \ScanLink67[12] , \ScanLink67[11] , \ScanLink67[10] , \ScanLink67[9] , 
        \ScanLink67[8] , \ScanLink67[7] , \ScanLink67[6] , \ScanLink67[5] , 
        \ScanLink67[4] , \ScanLink67[3] , \ScanLink67[2] , \ScanLink67[1] , 
        \ScanLink67[0] }), .ScanOut({\ScanLink66[31] , \ScanLink66[30] , 
        \ScanLink66[29] , \ScanLink66[28] , \ScanLink66[27] , \ScanLink66[26] , 
        \ScanLink66[25] , \ScanLink66[24] , \ScanLink66[23] , \ScanLink66[22] , 
        \ScanLink66[21] , \ScanLink66[20] , \ScanLink66[19] , \ScanLink66[18] , 
        \ScanLink66[17] , \ScanLink66[16] , \ScanLink66[15] , \ScanLink66[14] , 
        \ScanLink66[13] , \ScanLink66[12] , \ScanLink66[11] , \ScanLink66[10] , 
        \ScanLink66[9] , \ScanLink66[8] , \ScanLink66[7] , \ScanLink66[6] , 
        \ScanLink66[5] , \ScanLink66[4] , \ScanLink66[3] , \ScanLink66[2] , 
        \ScanLink66[1] , \ScanLink66[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB94[31] , \wRegInB94[30] , 
        \wRegInB94[29] , \wRegInB94[28] , \wRegInB94[27] , \wRegInB94[26] , 
        \wRegInB94[25] , \wRegInB94[24] , \wRegInB94[23] , \wRegInB94[22] , 
        \wRegInB94[21] , \wRegInB94[20] , \wRegInB94[19] , \wRegInB94[18] , 
        \wRegInB94[17] , \wRegInB94[16] , \wRegInB94[15] , \wRegInB94[14] , 
        \wRegInB94[13] , \wRegInB94[12] , \wRegInB94[11] , \wRegInB94[10] , 
        \wRegInB94[9] , \wRegInB94[8] , \wRegInB94[7] , \wRegInB94[6] , 
        \wRegInB94[5] , \wRegInB94[4] , \wRegInB94[3] , \wRegInB94[2] , 
        \wRegInB94[1] , \wRegInB94[0] }), .Out({\wBIn94[31] , \wBIn94[30] , 
        \wBIn94[29] , \wBIn94[28] , \wBIn94[27] , \wBIn94[26] , \wBIn94[25] , 
        \wBIn94[24] , \wBIn94[23] , \wBIn94[22] , \wBIn94[21] , \wBIn94[20] , 
        \wBIn94[19] , \wBIn94[18] , \wBIn94[17] , \wBIn94[16] , \wBIn94[15] , 
        \wBIn94[14] , \wBIn94[13] , \wBIn94[12] , \wBIn94[11] , \wBIn94[10] , 
        \wBIn94[9] , \wBIn94[8] , \wBIn94[7] , \wBIn94[6] , \wBIn94[5] , 
        \wBIn94[4] , \wBIn94[3] , \wBIn94[2] , \wBIn94[1] , \wBIn94[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_2 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB126[31] , \wRegInB126[30] , 
        \wRegInB126[29] , \wRegInB126[28] , \wRegInB126[27] , \wRegInB126[26] , 
        \wRegInB126[25] , \wRegInB126[24] , \wRegInB126[23] , \wRegInB126[22] , 
        \wRegInB126[21] , \wRegInB126[20] , \wRegInB126[19] , \wRegInB126[18] , 
        \wRegInB126[17] , \wRegInB126[16] , \wRegInB126[15] , \wRegInB126[14] , 
        \wRegInB126[13] , \wRegInB126[12] , \wRegInB126[11] , \wRegInB126[10] , 
        \wRegInB126[9] , \wRegInB126[8] , \wRegInB126[7] , \wRegInB126[6] , 
        \wRegInB126[5] , \wRegInB126[4] , \wRegInB126[3] , \wRegInB126[2] , 
        \wRegInB126[1] , \wRegInB126[0] }), .Out({\wBIn126[31] , \wBIn126[30] , 
        \wBIn126[29] , \wBIn126[28] , \wBIn126[27] , \wBIn126[26] , 
        \wBIn126[25] , \wBIn126[24] , \wBIn126[23] , \wBIn126[22] , 
        \wBIn126[21] , \wBIn126[20] , \wBIn126[19] , \wBIn126[18] , 
        \wBIn126[17] , \wBIn126[16] , \wBIn126[15] , \wBIn126[14] , 
        \wBIn126[13] , \wBIn126[12] , \wBIn126[11] , \wBIn126[10] , 
        \wBIn126[9] , \wBIn126[8] , \wBIn126[7] , \wBIn126[6] , \wBIn126[5] , 
        \wBIn126[4] , \wBIn126[3] , \wBIn126[2] , \wBIn126[1] , \wBIn126[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid9[31] , 
        \wAMid9[30] , \wAMid9[29] , \wAMid9[28] , \wAMid9[27] , \wAMid9[26] , 
        \wAMid9[25] , \wAMid9[24] , \wAMid9[23] , \wAMid9[22] , \wAMid9[21] , 
        \wAMid9[20] , \wAMid9[19] , \wAMid9[18] , \wAMid9[17] , \wAMid9[16] , 
        \wAMid9[15] , \wAMid9[14] , \wAMid9[13] , \wAMid9[12] , \wAMid9[11] , 
        \wAMid9[10] , \wAMid9[9] , \wAMid9[8] , \wAMid9[7] , \wAMid9[6] , 
        \wAMid9[5] , \wAMid9[4] , \wAMid9[3] , \wAMid9[2] , \wAMid9[1] , 
        \wAMid9[0] }), .BIn({\wBMid9[31] , \wBMid9[30] , \wBMid9[29] , 
        \wBMid9[28] , \wBMid9[27] , \wBMid9[26] , \wBMid9[25] , \wBMid9[24] , 
        \wBMid9[23] , \wBMid9[22] , \wBMid9[21] , \wBMid9[20] , \wBMid9[19] , 
        \wBMid9[18] , \wBMid9[17] , \wBMid9[16] , \wBMid9[15] , \wBMid9[14] , 
        \wBMid9[13] , \wBMid9[12] , \wBMid9[11] , \wBMid9[10] , \wBMid9[9] , 
        \wBMid9[8] , \wBMid9[7] , \wBMid9[6] , \wBMid9[5] , \wBMid9[4] , 
        \wBMid9[3] , \wBMid9[2] , \wBMid9[1] , \wBMid9[0] }), .HiOut({
        \wRegInB9[31] , \wRegInB9[30] , \wRegInB9[29] , \wRegInB9[28] , 
        \wRegInB9[27] , \wRegInB9[26] , \wRegInB9[25] , \wRegInB9[24] , 
        \wRegInB9[23] , \wRegInB9[22] , \wRegInB9[21] , \wRegInB9[20] , 
        \wRegInB9[19] , \wRegInB9[18] , \wRegInB9[17] , \wRegInB9[16] , 
        \wRegInB9[15] , \wRegInB9[14] , \wRegInB9[13] , \wRegInB9[12] , 
        \wRegInB9[11] , \wRegInB9[10] , \wRegInB9[9] , \wRegInB9[8] , 
        \wRegInB9[7] , \wRegInB9[6] , \wRegInB9[5] , \wRegInB9[4] , 
        \wRegInB9[3] , \wRegInB9[2] , \wRegInB9[1] , \wRegInB9[0] }), .LoOut({
        \wRegInA10[31] , \wRegInA10[30] , \wRegInA10[29] , \wRegInA10[28] , 
        \wRegInA10[27] , \wRegInA10[26] , \wRegInA10[25] , \wRegInA10[24] , 
        \wRegInA10[23] , \wRegInA10[22] , \wRegInA10[21] , \wRegInA10[20] , 
        \wRegInA10[19] , \wRegInA10[18] , \wRegInA10[17] , \wRegInA10[16] , 
        \wRegInA10[15] , \wRegInA10[14] , \wRegInA10[13] , \wRegInA10[12] , 
        \wRegInA10[11] , \wRegInA10[10] , \wRegInA10[9] , \wRegInA10[8] , 
        \wRegInA10[7] , \wRegInA10[6] , \wRegInA10[5] , \wRegInA10[4] , 
        \wRegInA10[3] , \wRegInA10[2] , \wRegInA10[1] , \wRegInA10[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_201 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink202[31] , \ScanLink202[30] , \ScanLink202[29] , 
        \ScanLink202[28] , \ScanLink202[27] , \ScanLink202[26] , 
        \ScanLink202[25] , \ScanLink202[24] , \ScanLink202[23] , 
        \ScanLink202[22] , \ScanLink202[21] , \ScanLink202[20] , 
        \ScanLink202[19] , \ScanLink202[18] , \ScanLink202[17] , 
        \ScanLink202[16] , \ScanLink202[15] , \ScanLink202[14] , 
        \ScanLink202[13] , \ScanLink202[12] , \ScanLink202[11] , 
        \ScanLink202[10] , \ScanLink202[9] , \ScanLink202[8] , 
        \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , \ScanLink202[4] , 
        \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , \ScanLink202[0] 
        }), .ScanOut({\ScanLink201[31] , \ScanLink201[30] , \ScanLink201[29] , 
        \ScanLink201[28] , \ScanLink201[27] , \ScanLink201[26] , 
        \ScanLink201[25] , \ScanLink201[24] , \ScanLink201[23] , 
        \ScanLink201[22] , \ScanLink201[21] , \ScanLink201[20] , 
        \ScanLink201[19] , \ScanLink201[18] , \ScanLink201[17] , 
        \ScanLink201[16] , \ScanLink201[15] , \ScanLink201[14] , 
        \ScanLink201[13] , \ScanLink201[12] , \ScanLink201[11] , 
        \ScanLink201[10] , \ScanLink201[9] , \ScanLink201[8] , 
        \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , \ScanLink201[4] , 
        \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , \ScanLink201[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA27[31] , \wRegInA27[30] , \wRegInA27[29] , 
        \wRegInA27[28] , \wRegInA27[27] , \wRegInA27[26] , \wRegInA27[25] , 
        \wRegInA27[24] , \wRegInA27[23] , \wRegInA27[22] , \wRegInA27[21] , 
        \wRegInA27[20] , \wRegInA27[19] , \wRegInA27[18] , \wRegInA27[17] , 
        \wRegInA27[16] , \wRegInA27[15] , \wRegInA27[14] , \wRegInA27[13] , 
        \wRegInA27[12] , \wRegInA27[11] , \wRegInA27[10] , \wRegInA27[9] , 
        \wRegInA27[8] , \wRegInA27[7] , \wRegInA27[6] , \wRegInA27[5] , 
        \wRegInA27[4] , \wRegInA27[3] , \wRegInA27[2] , \wRegInA27[1] , 
        \wRegInA27[0] }), .Out({\wAIn27[31] , \wAIn27[30] , \wAIn27[29] , 
        \wAIn27[28] , \wAIn27[27] , \wAIn27[26] , \wAIn27[25] , \wAIn27[24] , 
        \wAIn27[23] , \wAIn27[22] , \wAIn27[21] , \wAIn27[20] , \wAIn27[19] , 
        \wAIn27[18] , \wAIn27[17] , \wAIn27[16] , \wAIn27[15] , \wAIn27[14] , 
        \wAIn27[13] , \wAIn27[12] , \wAIn27[11] , \wAIn27[10] , \wAIn27[9] , 
        \wAIn27[8] , \wAIn27[7] , \wAIn27[6] , \wAIn27[5] , \wAIn27[4] , 
        \wAIn27[3] , \wAIn27[2] , \wAIn27[1] , \wAIn27[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_5 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[31] , \ScanLink6[30] , \ScanLink6[29] , 
        \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , \ScanLink6[25] , 
        \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , \ScanLink6[21] , 
        \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , \ScanLink6[17] , 
        \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , \ScanLink6[13] , 
        \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , \ScanLink6[9] , 
        \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA125[31] , \wRegInA125[30] , 
        \wRegInA125[29] , \wRegInA125[28] , \wRegInA125[27] , \wRegInA125[26] , 
        \wRegInA125[25] , \wRegInA125[24] , \wRegInA125[23] , \wRegInA125[22] , 
        \wRegInA125[21] , \wRegInA125[20] , \wRegInA125[19] , \wRegInA125[18] , 
        \wRegInA125[17] , \wRegInA125[16] , \wRegInA125[15] , \wRegInA125[14] , 
        \wRegInA125[13] , \wRegInA125[12] , \wRegInA125[11] , \wRegInA125[10] , 
        \wRegInA125[9] , \wRegInA125[8] , \wRegInA125[7] , \wRegInA125[6] , 
        \wRegInA125[5] , \wRegInA125[4] , \wRegInA125[3] , \wRegInA125[2] , 
        \wRegInA125[1] , \wRegInA125[0] }), .Out({\wAIn125[31] , \wAIn125[30] , 
        \wAIn125[29] , \wAIn125[28] , \wAIn125[27] , \wAIn125[26] , 
        \wAIn125[25] , \wAIn125[24] , \wAIn125[23] , \wAIn125[22] , 
        \wAIn125[21] , \wAIn125[20] , \wAIn125[19] , \wAIn125[18] , 
        \wAIn125[17] , \wAIn125[16] , \wAIn125[15] , \wAIn125[14] , 
        \wAIn125[13] , \wAIn125[12] , \wAIn125[11] , \wAIn125[10] , 
        \wAIn125[9] , \wAIn125[8] , \wAIn125[7] , \wAIn125[6] , \wAIn125[5] , 
        \wAIn125[4] , \wAIn125[3] , \wAIn125[2] , \wAIn125[1] , \wAIn125[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_131 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink132[31] , \ScanLink132[30] , \ScanLink132[29] , 
        \ScanLink132[28] , \ScanLink132[27] , \ScanLink132[26] , 
        \ScanLink132[25] , \ScanLink132[24] , \ScanLink132[23] , 
        \ScanLink132[22] , \ScanLink132[21] , \ScanLink132[20] , 
        \ScanLink132[19] , \ScanLink132[18] , \ScanLink132[17] , 
        \ScanLink132[16] , \ScanLink132[15] , \ScanLink132[14] , 
        \ScanLink132[13] , \ScanLink132[12] , \ScanLink132[11] , 
        \ScanLink132[10] , \ScanLink132[9] , \ScanLink132[8] , 
        \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , \ScanLink132[4] , 
        \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , \ScanLink132[0] 
        }), .ScanOut({\ScanLink131[31] , \ScanLink131[30] , \ScanLink131[29] , 
        \ScanLink131[28] , \ScanLink131[27] , \ScanLink131[26] , 
        \ScanLink131[25] , \ScanLink131[24] , \ScanLink131[23] , 
        \ScanLink131[22] , \ScanLink131[21] , \ScanLink131[20] , 
        \ScanLink131[19] , \ScanLink131[18] , \ScanLink131[17] , 
        \ScanLink131[16] , \ScanLink131[15] , \ScanLink131[14] , 
        \ScanLink131[13] , \ScanLink131[12] , \ScanLink131[11] , 
        \ScanLink131[10] , \ScanLink131[9] , \ScanLink131[8] , 
        \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , \ScanLink131[4] , 
        \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , \ScanLink131[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA62[31] , \wRegInA62[30] , \wRegInA62[29] , 
        \wRegInA62[28] , \wRegInA62[27] , \wRegInA62[26] , \wRegInA62[25] , 
        \wRegInA62[24] , \wRegInA62[23] , \wRegInA62[22] , \wRegInA62[21] , 
        \wRegInA62[20] , \wRegInA62[19] , \wRegInA62[18] , \wRegInA62[17] , 
        \wRegInA62[16] , \wRegInA62[15] , \wRegInA62[14] , \wRegInA62[13] , 
        \wRegInA62[12] , \wRegInA62[11] , \wRegInA62[10] , \wRegInA62[9] , 
        \wRegInA62[8] , \wRegInA62[7] , \wRegInA62[6] , \wRegInA62[5] , 
        \wRegInA62[4] , \wRegInA62[3] , \wRegInA62[2] , \wRegInA62[1] , 
        \wRegInA62[0] }), .Out({\wAIn62[31] , \wAIn62[30] , \wAIn62[29] , 
        \wAIn62[28] , \wAIn62[27] , \wAIn62[26] , \wAIn62[25] , \wAIn62[24] , 
        \wAIn62[23] , \wAIn62[22] , \wAIn62[21] , \wAIn62[20] , \wAIn62[19] , 
        \wAIn62[18] , \wAIn62[17] , \wAIn62[16] , \wAIn62[15] , \wAIn62[14] , 
        \wAIn62[13] , \wAIn62[12] , \wAIn62[11] , \wAIn62[10] , \wAIn62[9] , 
        \wAIn62[8] , \wAIn62[7] , \wAIn62[6] , \wAIn62[5] , \wAIn62[4] , 
        \wAIn62[3] , \wAIn62[2] , \wAIn62[1] , \wAIn62[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_61 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink62[31] , \ScanLink62[30] , \ScanLink62[29] , 
        \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , \ScanLink62[25] , 
        \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , \ScanLink62[21] , 
        \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , \ScanLink62[17] , 
        \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , \ScanLink62[13] , 
        \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , \ScanLink62[9] , 
        \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , \ScanLink62[5] , 
        \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , \ScanLink62[1] , 
        \ScanLink62[0] }), .ScanOut({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA97[31] , \wRegInA97[30] , 
        \wRegInA97[29] , \wRegInA97[28] , \wRegInA97[27] , \wRegInA97[26] , 
        \wRegInA97[25] , \wRegInA97[24] , \wRegInA97[23] , \wRegInA97[22] , 
        \wRegInA97[21] , \wRegInA97[20] , \wRegInA97[19] , \wRegInA97[18] , 
        \wRegInA97[17] , \wRegInA97[16] , \wRegInA97[15] , \wRegInA97[14] , 
        \wRegInA97[13] , \wRegInA97[12] , \wRegInA97[11] , \wRegInA97[10] , 
        \wRegInA97[9] , \wRegInA97[8] , \wRegInA97[7] , \wRegInA97[6] , 
        \wRegInA97[5] , \wRegInA97[4] , \wRegInA97[3] , \wRegInA97[2] , 
        \wRegInA97[1] , \wRegInA97[0] }), .Out({\wAIn97[31] , \wAIn97[30] , 
        \wAIn97[29] , \wAIn97[28] , \wAIn97[27] , \wAIn97[26] , \wAIn97[25] , 
        \wAIn97[24] , \wAIn97[23] , \wAIn97[22] , \wAIn97[21] , \wAIn97[20] , 
        \wAIn97[19] , \wAIn97[18] , \wAIn97[17] , \wAIn97[16] , \wAIn97[15] , 
        \wAIn97[14] , \wAIn97[13] , \wAIn97[12] , \wAIn97[11] , \wAIn97[10] , 
        \wAIn97[9] , \wAIn97[8] , \wAIn97[7] , \wAIn97[6] , \wAIn97[5] , 
        \wAIn97[4] , \wAIn97[3] , \wAIn97[2] , \wAIn97[1] , \wAIn97[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid23[31] , \wAMid23[30] , \wAMid23[29] , \wAMid23[28] , 
        \wAMid23[27] , \wAMid23[26] , \wAMid23[25] , \wAMid23[24] , 
        \wAMid23[23] , \wAMid23[22] , \wAMid23[21] , \wAMid23[20] , 
        \wAMid23[19] , \wAMid23[18] , \wAMid23[17] , \wAMid23[16] , 
        \wAMid23[15] , \wAMid23[14] , \wAMid23[13] , \wAMid23[12] , 
        \wAMid23[11] , \wAMid23[10] , \wAMid23[9] , \wAMid23[8] , \wAMid23[7] , 
        \wAMid23[6] , \wAMid23[5] , \wAMid23[4] , \wAMid23[3] , \wAMid23[2] , 
        \wAMid23[1] , \wAMid23[0] }), .BIn({\wBMid23[31] , \wBMid23[30] , 
        \wBMid23[29] , \wBMid23[28] , \wBMid23[27] , \wBMid23[26] , 
        \wBMid23[25] , \wBMid23[24] , \wBMid23[23] , \wBMid23[22] , 
        \wBMid23[21] , \wBMid23[20] , \wBMid23[19] , \wBMid23[18] , 
        \wBMid23[17] , \wBMid23[16] , \wBMid23[15] , \wBMid23[14] , 
        \wBMid23[13] , \wBMid23[12] , \wBMid23[11] , \wBMid23[10] , 
        \wBMid23[9] , \wBMid23[8] , \wBMid23[7] , \wBMid23[6] , \wBMid23[5] , 
        \wBMid23[4] , \wBMid23[3] , \wBMid23[2] , \wBMid23[1] , \wBMid23[0] }), 
        .HiOut({\wRegInB23[31] , \wRegInB23[30] , \wRegInB23[29] , 
        \wRegInB23[28] , \wRegInB23[27] , \wRegInB23[26] , \wRegInB23[25] , 
        \wRegInB23[24] , \wRegInB23[23] , \wRegInB23[22] , \wRegInB23[21] , 
        \wRegInB23[20] , \wRegInB23[19] , \wRegInB23[18] , \wRegInB23[17] , 
        \wRegInB23[16] , \wRegInB23[15] , \wRegInB23[14] , \wRegInB23[13] , 
        \wRegInB23[12] , \wRegInB23[11] , \wRegInB23[10] , \wRegInB23[9] , 
        \wRegInB23[8] , \wRegInB23[7] , \wRegInB23[6] , \wRegInB23[5] , 
        \wRegInB23[4] , \wRegInB23[3] , \wRegInB23[2] , \wRegInB23[1] , 
        \wRegInB23[0] }), .LoOut({\wRegInA24[31] , \wRegInA24[30] , 
        \wRegInA24[29] , \wRegInA24[28] , \wRegInA24[27] , \wRegInA24[26] , 
        \wRegInA24[25] , \wRegInA24[24] , \wRegInA24[23] , \wRegInA24[22] , 
        \wRegInA24[21] , \wRegInA24[20] , \wRegInA24[19] , \wRegInA24[18] , 
        \wRegInA24[17] , \wRegInA24[16] , \wRegInA24[15] , \wRegInA24[14] , 
        \wRegInA24[13] , \wRegInA24[12] , \wRegInA24[11] , \wRegInA24[10] , 
        \wRegInA24[9] , \wRegInA24[8] , \wRegInA24[7] , \wRegInA24[6] , 
        \wRegInA24[5] , \wRegInA24[4] , \wRegInA24[3] , \wRegInA24[2] , 
        \wRegInA24[1] , \wRegInA24[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_116 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink117[31] , \ScanLink117[30] , \ScanLink117[29] , 
        \ScanLink117[28] , \ScanLink117[27] , \ScanLink117[26] , 
        \ScanLink117[25] , \ScanLink117[24] , \ScanLink117[23] , 
        \ScanLink117[22] , \ScanLink117[21] , \ScanLink117[20] , 
        \ScanLink117[19] , \ScanLink117[18] , \ScanLink117[17] , 
        \ScanLink117[16] , \ScanLink117[15] , \ScanLink117[14] , 
        \ScanLink117[13] , \ScanLink117[12] , \ScanLink117[11] , 
        \ScanLink117[10] , \ScanLink117[9] , \ScanLink117[8] , 
        \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , \ScanLink117[4] , 
        \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , \ScanLink117[0] 
        }), .ScanOut({\ScanLink116[31] , \ScanLink116[30] , \ScanLink116[29] , 
        \ScanLink116[28] , \ScanLink116[27] , \ScanLink116[26] , 
        \ScanLink116[25] , \ScanLink116[24] , \ScanLink116[23] , 
        \ScanLink116[22] , \ScanLink116[21] , \ScanLink116[20] , 
        \ScanLink116[19] , \ScanLink116[18] , \ScanLink116[17] , 
        \ScanLink116[16] , \ScanLink116[15] , \ScanLink116[14] , 
        \ScanLink116[13] , \ScanLink116[12] , \ScanLink116[11] , 
        \ScanLink116[10] , \ScanLink116[9] , \ScanLink116[8] , 
        \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , \ScanLink116[4] , 
        \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , \ScanLink116[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB69[31] , \wRegInB69[30] , \wRegInB69[29] , 
        \wRegInB69[28] , \wRegInB69[27] , \wRegInB69[26] , \wRegInB69[25] , 
        \wRegInB69[24] , \wRegInB69[23] , \wRegInB69[22] , \wRegInB69[21] , 
        \wRegInB69[20] , \wRegInB69[19] , \wRegInB69[18] , \wRegInB69[17] , 
        \wRegInB69[16] , \wRegInB69[15] , \wRegInB69[14] , \wRegInB69[13] , 
        \wRegInB69[12] , \wRegInB69[11] , \wRegInB69[10] , \wRegInB69[9] , 
        \wRegInB69[8] , \wRegInB69[7] , \wRegInB69[6] , \wRegInB69[5] , 
        \wRegInB69[4] , \wRegInB69[3] , \wRegInB69[2] , \wRegInB69[1] , 
        \wRegInB69[0] }), .Out({\wBIn69[31] , \wBIn69[30] , \wBIn69[29] , 
        \wBIn69[28] , \wBIn69[27] , \wBIn69[26] , \wBIn69[25] , \wBIn69[24] , 
        \wBIn69[23] , \wBIn69[22] , \wBIn69[21] , \wBIn69[20] , \wBIn69[19] , 
        \wBIn69[18] , \wBIn69[17] , \wBIn69[16] , \wBIn69[15] , \wBIn69[14] , 
        \wBIn69[13] , \wBIn69[12] , \wBIn69[11] , \wBIn69[10] , \wBIn69[9] , 
        \wBIn69[8] , \wBIn69[7] , \wBIn69[6] , \wBIn69[5] , \wBIn69[4] , 
        \wBIn69[3] , \wBIn69[2] , \wBIn69[1] , \wBIn69[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_46 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink47[31] , \ScanLink47[30] , \ScanLink47[29] , 
        \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , \ScanLink47[25] , 
        \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , \ScanLink47[21] , 
        \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , \ScanLink47[17] , 
        \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , \ScanLink47[13] , 
        \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , \ScanLink47[9] , 
        \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , \ScanLink47[5] , 
        \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , \ScanLink47[1] , 
        \ScanLink47[0] }), .ScanOut({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB104[31] , \wRegInB104[30] , 
        \wRegInB104[29] , \wRegInB104[28] , \wRegInB104[27] , \wRegInB104[26] , 
        \wRegInB104[25] , \wRegInB104[24] , \wRegInB104[23] , \wRegInB104[22] , 
        \wRegInB104[21] , \wRegInB104[20] , \wRegInB104[19] , \wRegInB104[18] , 
        \wRegInB104[17] , \wRegInB104[16] , \wRegInB104[15] , \wRegInB104[14] , 
        \wRegInB104[13] , \wRegInB104[12] , \wRegInB104[11] , \wRegInB104[10] , 
        \wRegInB104[9] , \wRegInB104[8] , \wRegInB104[7] , \wRegInB104[6] , 
        \wRegInB104[5] , \wRegInB104[4] , \wRegInB104[3] , \wRegInB104[2] , 
        \wRegInB104[1] , \wRegInB104[0] }), .Out({\wBIn104[31] , \wBIn104[30] , 
        \wBIn104[29] , \wBIn104[28] , \wBIn104[27] , \wBIn104[26] , 
        \wBIn104[25] , \wBIn104[24] , \wBIn104[23] , \wBIn104[22] , 
        \wBIn104[21] , \wBIn104[20] , \wBIn104[19] , \wBIn104[18] , 
        \wBIn104[17] , \wBIn104[16] , \wBIn104[15] , \wBIn104[14] , 
        \wBIn104[13] , \wBIn104[12] , \wBIn104[11] , \wBIn104[10] , 
        \wBIn104[9] , \wBIn104[8] , \wBIn104[7] , \wBIn104[6] , \wBIn104[5] , 
        \wBIn104[4] , \wBIn104[3] , \wBIn104[2] , \wBIn104[1] , \wBIn104[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn41[31] , \wAIn41[30] , \wAIn41[29] , \wAIn41[28] , \wAIn41[27] , 
        \wAIn41[26] , \wAIn41[25] , \wAIn41[24] , \wAIn41[23] , \wAIn41[22] , 
        \wAIn41[21] , \wAIn41[20] , \wAIn41[19] , \wAIn41[18] , \wAIn41[17] , 
        \wAIn41[16] , \wAIn41[15] , \wAIn41[14] , \wAIn41[13] , \wAIn41[12] , 
        \wAIn41[11] , \wAIn41[10] , \wAIn41[9] , \wAIn41[8] , \wAIn41[7] , 
        \wAIn41[6] , \wAIn41[5] , \wAIn41[4] , \wAIn41[3] , \wAIn41[2] , 
        \wAIn41[1] , \wAIn41[0] }), .BIn({\wBIn41[31] , \wBIn41[30] , 
        \wBIn41[29] , \wBIn41[28] , \wBIn41[27] , \wBIn41[26] , \wBIn41[25] , 
        \wBIn41[24] , \wBIn41[23] , \wBIn41[22] , \wBIn41[21] , \wBIn41[20] , 
        \wBIn41[19] , \wBIn41[18] , \wBIn41[17] , \wBIn41[16] , \wBIn41[15] , 
        \wBIn41[14] , \wBIn41[13] , \wBIn41[12] , \wBIn41[11] , \wBIn41[10] , 
        \wBIn41[9] , \wBIn41[8] , \wBIn41[7] , \wBIn41[6] , \wBIn41[5] , 
        \wBIn41[4] , \wBIn41[3] , \wBIn41[2] , \wBIn41[1] , \wBIn41[0] }), 
        .HiOut({\wBMid40[31] , \wBMid40[30] , \wBMid40[29] , \wBMid40[28] , 
        \wBMid40[27] , \wBMid40[26] , \wBMid40[25] , \wBMid40[24] , 
        \wBMid40[23] , \wBMid40[22] , \wBMid40[21] , \wBMid40[20] , 
        \wBMid40[19] , \wBMid40[18] , \wBMid40[17] , \wBMid40[16] , 
        \wBMid40[15] , \wBMid40[14] , \wBMid40[13] , \wBMid40[12] , 
        \wBMid40[11] , \wBMid40[10] , \wBMid40[9] , \wBMid40[8] , \wBMid40[7] , 
        \wBMid40[6] , \wBMid40[5] , \wBMid40[4] , \wBMid40[3] , \wBMid40[2] , 
        \wBMid40[1] , \wBMid40[0] }), .LoOut({\wAMid41[31] , \wAMid41[30] , 
        \wAMid41[29] , \wAMid41[28] , \wAMid41[27] , \wAMid41[26] , 
        \wAMid41[25] , \wAMid41[24] , \wAMid41[23] , \wAMid41[22] , 
        \wAMid41[21] , \wAMid41[20] , \wAMid41[19] , \wAMid41[18] , 
        \wAMid41[17] , \wAMid41[16] , \wAMid41[15] , \wAMid41[14] , 
        \wAMid41[13] , \wAMid41[12] , \wAMid41[11] , \wAMid41[10] , 
        \wAMid41[9] , \wAMid41[8] , \wAMid41[7] , \wAMid41[6] , \wAMid41[5] , 
        \wAMid41[4] , \wAMid41[3] , \wAMid41[2] , \wAMid41[1] , \wAMid41[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid107[31] , \wAMid107[30] , \wAMid107[29] , \wAMid107[28] , 
        \wAMid107[27] , \wAMid107[26] , \wAMid107[25] , \wAMid107[24] , 
        \wAMid107[23] , \wAMid107[22] , \wAMid107[21] , \wAMid107[20] , 
        \wAMid107[19] , \wAMid107[18] , \wAMid107[17] , \wAMid107[16] , 
        \wAMid107[15] , \wAMid107[14] , \wAMid107[13] , \wAMid107[12] , 
        \wAMid107[11] , \wAMid107[10] , \wAMid107[9] , \wAMid107[8] , 
        \wAMid107[7] , \wAMid107[6] , \wAMid107[5] , \wAMid107[4] , 
        \wAMid107[3] , \wAMid107[2] , \wAMid107[1] , \wAMid107[0] }), .BIn({
        \wBMid107[31] , \wBMid107[30] , \wBMid107[29] , \wBMid107[28] , 
        \wBMid107[27] , \wBMid107[26] , \wBMid107[25] , \wBMid107[24] , 
        \wBMid107[23] , \wBMid107[22] , \wBMid107[21] , \wBMid107[20] , 
        \wBMid107[19] , \wBMid107[18] , \wBMid107[17] , \wBMid107[16] , 
        \wBMid107[15] , \wBMid107[14] , \wBMid107[13] , \wBMid107[12] , 
        \wBMid107[11] , \wBMid107[10] , \wBMid107[9] , \wBMid107[8] , 
        \wBMid107[7] , \wBMid107[6] , \wBMid107[5] , \wBMid107[4] , 
        \wBMid107[3] , \wBMid107[2] , \wBMid107[1] , \wBMid107[0] }), .HiOut({
        \wRegInB107[31] , \wRegInB107[30] , \wRegInB107[29] , \wRegInB107[28] , 
        \wRegInB107[27] , \wRegInB107[26] , \wRegInB107[25] , \wRegInB107[24] , 
        \wRegInB107[23] , \wRegInB107[22] , \wRegInB107[21] , \wRegInB107[20] , 
        \wRegInB107[19] , \wRegInB107[18] , \wRegInB107[17] , \wRegInB107[16] , 
        \wRegInB107[15] , \wRegInB107[14] , \wRegInB107[13] , \wRegInB107[12] , 
        \wRegInB107[11] , \wRegInB107[10] , \wRegInB107[9] , \wRegInB107[8] , 
        \wRegInB107[7] , \wRegInB107[6] , \wRegInB107[5] , \wRegInB107[4] , 
        \wRegInB107[3] , \wRegInB107[2] , \wRegInB107[1] , \wRegInB107[0] }), 
        .LoOut({\wRegInA108[31] , \wRegInA108[30] , \wRegInA108[29] , 
        \wRegInA108[28] , \wRegInA108[27] , \wRegInA108[26] , \wRegInA108[25] , 
        \wRegInA108[24] , \wRegInA108[23] , \wRegInA108[22] , \wRegInA108[21] , 
        \wRegInA108[20] , \wRegInA108[19] , \wRegInA108[18] , \wRegInA108[17] , 
        \wRegInA108[16] , \wRegInA108[15] , \wRegInA108[14] , \wRegInA108[13] , 
        \wRegInA108[12] , \wRegInA108[11] , \wRegInA108[10] , \wRegInA108[9] , 
        \wRegInA108[8] , \wRegInA108[7] , \wRegInA108[6] , \wRegInA108[5] , 
        \wRegInA108[4] , \wRegInA108[3] , \wRegInA108[2] , \wRegInA108[1] , 
        \wRegInA108[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid120[31] , \wAMid120[30] , \wAMid120[29] , \wAMid120[28] , 
        \wAMid120[27] , \wAMid120[26] , \wAMid120[25] , \wAMid120[24] , 
        \wAMid120[23] , \wAMid120[22] , \wAMid120[21] , \wAMid120[20] , 
        \wAMid120[19] , \wAMid120[18] , \wAMid120[17] , \wAMid120[16] , 
        \wAMid120[15] , \wAMid120[14] , \wAMid120[13] , \wAMid120[12] , 
        \wAMid120[11] , \wAMid120[10] , \wAMid120[9] , \wAMid120[8] , 
        \wAMid120[7] , \wAMid120[6] , \wAMid120[5] , \wAMid120[4] , 
        \wAMid120[3] , \wAMid120[2] , \wAMid120[1] , \wAMid120[0] }), .BIn({
        \wBMid120[31] , \wBMid120[30] , \wBMid120[29] , \wBMid120[28] , 
        \wBMid120[27] , \wBMid120[26] , \wBMid120[25] , \wBMid120[24] , 
        \wBMid120[23] , \wBMid120[22] , \wBMid120[21] , \wBMid120[20] , 
        \wBMid120[19] , \wBMid120[18] , \wBMid120[17] , \wBMid120[16] , 
        \wBMid120[15] , \wBMid120[14] , \wBMid120[13] , \wBMid120[12] , 
        \wBMid120[11] , \wBMid120[10] , \wBMid120[9] , \wBMid120[8] , 
        \wBMid120[7] , \wBMid120[6] , \wBMid120[5] , \wBMid120[4] , 
        \wBMid120[3] , \wBMid120[2] , \wBMid120[1] , \wBMid120[0] }), .HiOut({
        \wRegInB120[31] , \wRegInB120[30] , \wRegInB120[29] , \wRegInB120[28] , 
        \wRegInB120[27] , \wRegInB120[26] , \wRegInB120[25] , \wRegInB120[24] , 
        \wRegInB120[23] , \wRegInB120[22] , \wRegInB120[21] , \wRegInB120[20] , 
        \wRegInB120[19] , \wRegInB120[18] , \wRegInB120[17] , \wRegInB120[16] , 
        \wRegInB120[15] , \wRegInB120[14] , \wRegInB120[13] , \wRegInB120[12] , 
        \wRegInB120[11] , \wRegInB120[10] , \wRegInB120[9] , \wRegInB120[8] , 
        \wRegInB120[7] , \wRegInB120[6] , \wRegInB120[5] , \wRegInB120[4] , 
        \wRegInB120[3] , \wRegInB120[2] , \wRegInB120[1] , \wRegInB120[0] }), 
        .LoOut({\wRegInA121[31] , \wRegInA121[30] , \wRegInA121[29] , 
        \wRegInA121[28] , \wRegInA121[27] , \wRegInA121[26] , \wRegInA121[25] , 
        \wRegInA121[24] , \wRegInA121[23] , \wRegInA121[22] , \wRegInA121[21] , 
        \wRegInA121[20] , \wRegInA121[19] , \wRegInA121[18] , \wRegInA121[17] , 
        \wRegInA121[16] , \wRegInA121[15] , \wRegInA121[14] , \wRegInA121[13] , 
        \wRegInA121[12] , \wRegInA121[11] , \wRegInA121[10] , \wRegInA121[9] , 
        \wRegInA121[8] , \wRegInA121[7] , \wRegInA121[6] , \wRegInA121[5] , 
        \wRegInA121[4] , \wRegInA121[3] , \wRegInA121[2] , \wRegInA121[1] , 
        \wRegInA121[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_248 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink249[31] , \ScanLink249[30] , \ScanLink249[29] , 
        \ScanLink249[28] , \ScanLink249[27] , \ScanLink249[26] , 
        \ScanLink249[25] , \ScanLink249[24] , \ScanLink249[23] , 
        \ScanLink249[22] , \ScanLink249[21] , \ScanLink249[20] , 
        \ScanLink249[19] , \ScanLink249[18] , \ScanLink249[17] , 
        \ScanLink249[16] , \ScanLink249[15] , \ScanLink249[14] , 
        \ScanLink249[13] , \ScanLink249[12] , \ScanLink249[11] , 
        \ScanLink249[10] , \ScanLink249[9] , \ScanLink249[8] , 
        \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , \ScanLink249[4] , 
        \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , \ScanLink249[0] 
        }), .ScanOut({\ScanLink248[31] , \ScanLink248[30] , \ScanLink248[29] , 
        \ScanLink248[28] , \ScanLink248[27] , \ScanLink248[26] , 
        \ScanLink248[25] , \ScanLink248[24] , \ScanLink248[23] , 
        \ScanLink248[22] , \ScanLink248[21] , \ScanLink248[20] , 
        \ScanLink248[19] , \ScanLink248[18] , \ScanLink248[17] , 
        \ScanLink248[16] , \ScanLink248[15] , \ScanLink248[14] , 
        \ScanLink248[13] , \ScanLink248[12] , \ScanLink248[11] , 
        \ScanLink248[10] , \ScanLink248[9] , \ScanLink248[8] , 
        \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , \ScanLink248[4] , 
        \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , \ScanLink248[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB3[31] , \wRegInB3[30] , \wRegInB3[29] , \wRegInB3[28] , 
        \wRegInB3[27] , \wRegInB3[26] , \wRegInB3[25] , \wRegInB3[24] , 
        \wRegInB3[23] , \wRegInB3[22] , \wRegInB3[21] , \wRegInB3[20] , 
        \wRegInB3[19] , \wRegInB3[18] , \wRegInB3[17] , \wRegInB3[16] , 
        \wRegInB3[15] , \wRegInB3[14] , \wRegInB3[13] , \wRegInB3[12] , 
        \wRegInB3[11] , \wRegInB3[10] , \wRegInB3[9] , \wRegInB3[8] , 
        \wRegInB3[7] , \wRegInB3[6] , \wRegInB3[5] , \wRegInB3[4] , 
        \wRegInB3[3] , \wRegInB3[2] , \wRegInB3[1] , \wRegInB3[0] }), .Out({
        \wBIn3[31] , \wBIn3[30] , \wBIn3[29] , \wBIn3[28] , \wBIn3[27] , 
        \wBIn3[26] , \wBIn3[25] , \wBIn3[24] , \wBIn3[23] , \wBIn3[22] , 
        \wBIn3[21] , \wBIn3[20] , \wBIn3[19] , \wBIn3[18] , \wBIn3[17] , 
        \wBIn3[16] , \wBIn3[15] , \wBIn3[14] , \wBIn3[13] , \wBIn3[12] , 
        \wBIn3[11] , \wBIn3[10] , \wBIn3[9] , \wBIn3[8] , \wBIn3[7] , 
        \wBIn3[6] , \wBIn3[5] , \wBIn3[4] , \wBIn3[3] , \wBIn3[2] , \wBIn3[1] , 
        \wBIn3[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_226 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink227[31] , \ScanLink227[30] , \ScanLink227[29] , 
        \ScanLink227[28] , \ScanLink227[27] , \ScanLink227[26] , 
        \ScanLink227[25] , \ScanLink227[24] , \ScanLink227[23] , 
        \ScanLink227[22] , \ScanLink227[21] , \ScanLink227[20] , 
        \ScanLink227[19] , \ScanLink227[18] , \ScanLink227[17] , 
        \ScanLink227[16] , \ScanLink227[15] , \ScanLink227[14] , 
        \ScanLink227[13] , \ScanLink227[12] , \ScanLink227[11] , 
        \ScanLink227[10] , \ScanLink227[9] , \ScanLink227[8] , 
        \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , \ScanLink227[4] , 
        \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , \ScanLink227[0] 
        }), .ScanOut({\ScanLink226[31] , \ScanLink226[30] , \ScanLink226[29] , 
        \ScanLink226[28] , \ScanLink226[27] , \ScanLink226[26] , 
        \ScanLink226[25] , \ScanLink226[24] , \ScanLink226[23] , 
        \ScanLink226[22] , \ScanLink226[21] , \ScanLink226[20] , 
        \ScanLink226[19] , \ScanLink226[18] , \ScanLink226[17] , 
        \ScanLink226[16] , \ScanLink226[15] , \ScanLink226[14] , 
        \ScanLink226[13] , \ScanLink226[12] , \ScanLink226[11] , 
        \ScanLink226[10] , \ScanLink226[9] , \ScanLink226[8] , 
        \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , \ScanLink226[4] , 
        \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , \ScanLink226[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB14[31] , \wRegInB14[30] , \wRegInB14[29] , 
        \wRegInB14[28] , \wRegInB14[27] , \wRegInB14[26] , \wRegInB14[25] , 
        \wRegInB14[24] , \wRegInB14[23] , \wRegInB14[22] , \wRegInB14[21] , 
        \wRegInB14[20] , \wRegInB14[19] , \wRegInB14[18] , \wRegInB14[17] , 
        \wRegInB14[16] , \wRegInB14[15] , \wRegInB14[14] , \wRegInB14[13] , 
        \wRegInB14[12] , \wRegInB14[11] , \wRegInB14[10] , \wRegInB14[9] , 
        \wRegInB14[8] , \wRegInB14[7] , \wRegInB14[6] , \wRegInB14[5] , 
        \wRegInB14[4] , \wRegInB14[3] , \wRegInB14[2] , \wRegInB14[1] , 
        \wRegInB14[0] }), .Out({\wBIn14[31] , \wBIn14[30] , \wBIn14[29] , 
        \wBIn14[28] , \wBIn14[27] , \wBIn14[26] , \wBIn14[25] , \wBIn14[24] , 
        \wBIn14[23] , \wBIn14[22] , \wBIn14[21] , \wBIn14[20] , \wBIn14[19] , 
        \wBIn14[18] , \wBIn14[17] , \wBIn14[16] , \wBIn14[15] , \wBIn14[14] , 
        \wBIn14[13] , \wBIn14[12] , \wBIn14[11] , \wBIn14[10] , \wBIn14[9] , 
        \wBIn14[8] , \wBIn14[7] , \wBIn14[6] , \wBIn14[5] , \wBIn14[4] , 
        \wBIn14[3] , \wBIn14[2] , \wBIn14[1] , \wBIn14[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_178 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink179[31] , \ScanLink179[30] , \ScanLink179[29] , 
        \ScanLink179[28] , \ScanLink179[27] , \ScanLink179[26] , 
        \ScanLink179[25] , \ScanLink179[24] , \ScanLink179[23] , 
        \ScanLink179[22] , \ScanLink179[21] , \ScanLink179[20] , 
        \ScanLink179[19] , \ScanLink179[18] , \ScanLink179[17] , 
        \ScanLink179[16] , \ScanLink179[15] , \ScanLink179[14] , 
        \ScanLink179[13] , \ScanLink179[12] , \ScanLink179[11] , 
        \ScanLink179[10] , \ScanLink179[9] , \ScanLink179[8] , 
        \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , \ScanLink179[4] , 
        \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , \ScanLink179[0] 
        }), .ScanOut({\ScanLink178[31] , \ScanLink178[30] , \ScanLink178[29] , 
        \ScanLink178[28] , \ScanLink178[27] , \ScanLink178[26] , 
        \ScanLink178[25] , \ScanLink178[24] , \ScanLink178[23] , 
        \ScanLink178[22] , \ScanLink178[21] , \ScanLink178[20] , 
        \ScanLink178[19] , \ScanLink178[18] , \ScanLink178[17] , 
        \ScanLink178[16] , \ScanLink178[15] , \ScanLink178[14] , 
        \ScanLink178[13] , \ScanLink178[12] , \ScanLink178[11] , 
        \ScanLink178[10] , \ScanLink178[9] , \ScanLink178[8] , 
        \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , \ScanLink178[4] , 
        \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , \ScanLink178[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB38[31] , \wRegInB38[30] , \wRegInB38[29] , 
        \wRegInB38[28] , \wRegInB38[27] , \wRegInB38[26] , \wRegInB38[25] , 
        \wRegInB38[24] , \wRegInB38[23] , \wRegInB38[22] , \wRegInB38[21] , 
        \wRegInB38[20] , \wRegInB38[19] , \wRegInB38[18] , \wRegInB38[17] , 
        \wRegInB38[16] , \wRegInB38[15] , \wRegInB38[14] , \wRegInB38[13] , 
        \wRegInB38[12] , \wRegInB38[11] , \wRegInB38[10] , \wRegInB38[9] , 
        \wRegInB38[8] , \wRegInB38[7] , \wRegInB38[6] , \wRegInB38[5] , 
        \wRegInB38[4] , \wRegInB38[3] , \wRegInB38[2] , \wRegInB38[1] , 
        \wRegInB38[0] }), .Out({\wBIn38[31] , \wBIn38[30] , \wBIn38[29] , 
        \wBIn38[28] , \wBIn38[27] , \wBIn38[26] , \wBIn38[25] , \wBIn38[24] , 
        \wBIn38[23] , \wBIn38[22] , \wBIn38[21] , \wBIn38[20] , \wBIn38[19] , 
        \wBIn38[18] , \wBIn38[17] , \wBIn38[16] , \wBIn38[15] , \wBIn38[14] , 
        \wBIn38[13] , \wBIn38[12] , \wBIn38[11] , \wBIn38[10] , \wBIn38[9] , 
        \wBIn38[8] , \wBIn38[7] , \wBIn38[6] , \wBIn38[5] , \wBIn38[4] , 
        \wBIn38[3] , \wBIn38[2] , \wBIn38[1] , \wBIn38[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_28 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink29[31] , \ScanLink29[30] , \ScanLink29[29] , 
        \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , \ScanLink29[25] , 
        \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , \ScanLink29[21] , 
        \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , \ScanLink29[17] , 
        \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , \ScanLink29[13] , 
        \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , \ScanLink29[9] , 
        \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , \ScanLink29[5] , 
        \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , \ScanLink29[1] , 
        \ScanLink29[0] }), .ScanOut({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB113[31] , \wRegInB113[30] , 
        \wRegInB113[29] , \wRegInB113[28] , \wRegInB113[27] , \wRegInB113[26] , 
        \wRegInB113[25] , \wRegInB113[24] , \wRegInB113[23] , \wRegInB113[22] , 
        \wRegInB113[21] , \wRegInB113[20] , \wRegInB113[19] , \wRegInB113[18] , 
        \wRegInB113[17] , \wRegInB113[16] , \wRegInB113[15] , \wRegInB113[14] , 
        \wRegInB113[13] , \wRegInB113[12] , \wRegInB113[11] , \wRegInB113[10] , 
        \wRegInB113[9] , \wRegInB113[8] , \wRegInB113[7] , \wRegInB113[6] , 
        \wRegInB113[5] , \wRegInB113[4] , \wRegInB113[3] , \wRegInB113[2] , 
        \wRegInB113[1] , \wRegInB113[0] }), .Out({\wBIn113[31] , \wBIn113[30] , 
        \wBIn113[29] , \wBIn113[28] , \wBIn113[27] , \wBIn113[26] , 
        \wBIn113[25] , \wBIn113[24] , \wBIn113[23] , \wBIn113[22] , 
        \wBIn113[21] , \wBIn113[20] , \wBIn113[19] , \wBIn113[18] , 
        \wBIn113[17] , \wBIn113[16] , \wBIn113[15] , \wBIn113[14] , 
        \wBIn113[13] , \wBIn113[12] , \wBIn113[11] , \wBIn113[10] , 
        \wBIn113[9] , \wBIn113[8] , \wBIn113[7] , \wBIn113[6] , \wBIn113[5] , 
        \wBIn113[4] , \wBIn113[3] , \wBIn113[2] , \wBIn113[1] , \wBIn113[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_84 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink85[31] , \ScanLink85[30] , \ScanLink85[29] , 
        \ScanLink85[28] , \ScanLink85[27] , \ScanLink85[26] , \ScanLink85[25] , 
        \ScanLink85[24] , \ScanLink85[23] , \ScanLink85[22] , \ScanLink85[21] , 
        \ScanLink85[20] , \ScanLink85[19] , \ScanLink85[18] , \ScanLink85[17] , 
        \ScanLink85[16] , \ScanLink85[15] , \ScanLink85[14] , \ScanLink85[13] , 
        \ScanLink85[12] , \ScanLink85[11] , \ScanLink85[10] , \ScanLink85[9] , 
        \ScanLink85[8] , \ScanLink85[7] , \ScanLink85[6] , \ScanLink85[5] , 
        \ScanLink85[4] , \ScanLink85[3] , \ScanLink85[2] , \ScanLink85[1] , 
        \ScanLink85[0] }), .ScanOut({\ScanLink84[31] , \ScanLink84[30] , 
        \ScanLink84[29] , \ScanLink84[28] , \ScanLink84[27] , \ScanLink84[26] , 
        \ScanLink84[25] , \ScanLink84[24] , \ScanLink84[23] , \ScanLink84[22] , 
        \ScanLink84[21] , \ScanLink84[20] , \ScanLink84[19] , \ScanLink84[18] , 
        \ScanLink84[17] , \ScanLink84[16] , \ScanLink84[15] , \ScanLink84[14] , 
        \ScanLink84[13] , \ScanLink84[12] , \ScanLink84[11] , \ScanLink84[10] , 
        \ScanLink84[9] , \ScanLink84[8] , \ScanLink84[7] , \ScanLink84[6] , 
        \ScanLink84[5] , \ScanLink84[4] , \ScanLink84[3] , \ScanLink84[2] , 
        \ScanLink84[1] , \ScanLink84[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB85[31] , \wRegInB85[30] , 
        \wRegInB85[29] , \wRegInB85[28] , \wRegInB85[27] , \wRegInB85[26] , 
        \wRegInB85[25] , \wRegInB85[24] , \wRegInB85[23] , \wRegInB85[22] , 
        \wRegInB85[21] , \wRegInB85[20] , \wRegInB85[19] , \wRegInB85[18] , 
        \wRegInB85[17] , \wRegInB85[16] , \wRegInB85[15] , \wRegInB85[14] , 
        \wRegInB85[13] , \wRegInB85[12] , \wRegInB85[11] , \wRegInB85[10] , 
        \wRegInB85[9] , \wRegInB85[8] , \wRegInB85[7] , \wRegInB85[6] , 
        \wRegInB85[5] , \wRegInB85[4] , \wRegInB85[3] , \wRegInB85[2] , 
        \wRegInB85[1] , \wRegInB85[0] }), .Out({\wBIn85[31] , \wBIn85[30] , 
        \wBIn85[29] , \wBIn85[28] , \wBIn85[27] , \wBIn85[26] , \wBIn85[25] , 
        \wBIn85[24] , \wBIn85[23] , \wBIn85[22] , \wBIn85[21] , \wBIn85[20] , 
        \wBIn85[19] , \wBIn85[18] , \wBIn85[17] , \wBIn85[16] , \wBIn85[15] , 
        \wBIn85[14] , \wBIn85[13] , \wBIn85[12] , \wBIn85[11] , \wBIn85[10] , 
        \wBIn85[9] , \wBIn85[8] , \wBIn85[7] , \wBIn85[6] , \wBIn85[5] , 
        \wBIn85[4] , \wBIn85[3] , \wBIn85[2] , \wBIn85[1] , \wBIn85[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn66[31] , \wAIn66[30] , \wAIn66[29] , \wAIn66[28] , \wAIn66[27] , 
        \wAIn66[26] , \wAIn66[25] , \wAIn66[24] , \wAIn66[23] , \wAIn66[22] , 
        \wAIn66[21] , \wAIn66[20] , \wAIn66[19] , \wAIn66[18] , \wAIn66[17] , 
        \wAIn66[16] , \wAIn66[15] , \wAIn66[14] , \wAIn66[13] , \wAIn66[12] , 
        \wAIn66[11] , \wAIn66[10] , \wAIn66[9] , \wAIn66[8] , \wAIn66[7] , 
        \wAIn66[6] , \wAIn66[5] , \wAIn66[4] , \wAIn66[3] , \wAIn66[2] , 
        \wAIn66[1] , \wAIn66[0] }), .BIn({\wBIn66[31] , \wBIn66[30] , 
        \wBIn66[29] , \wBIn66[28] , \wBIn66[27] , \wBIn66[26] , \wBIn66[25] , 
        \wBIn66[24] , \wBIn66[23] , \wBIn66[22] , \wBIn66[21] , \wBIn66[20] , 
        \wBIn66[19] , \wBIn66[18] , \wBIn66[17] , \wBIn66[16] , \wBIn66[15] , 
        \wBIn66[14] , \wBIn66[13] , \wBIn66[12] , \wBIn66[11] , \wBIn66[10] , 
        \wBIn66[9] , \wBIn66[8] , \wBIn66[7] , \wBIn66[6] , \wBIn66[5] , 
        \wBIn66[4] , \wBIn66[3] , \wBIn66[2] , \wBIn66[1] , \wBIn66[0] }), 
        .HiOut({\wBMid65[31] , \wBMid65[30] , \wBMid65[29] , \wBMid65[28] , 
        \wBMid65[27] , \wBMid65[26] , \wBMid65[25] , \wBMid65[24] , 
        \wBMid65[23] , \wBMid65[22] , \wBMid65[21] , \wBMid65[20] , 
        \wBMid65[19] , \wBMid65[18] , \wBMid65[17] , \wBMid65[16] , 
        \wBMid65[15] , \wBMid65[14] , \wBMid65[13] , \wBMid65[12] , 
        \wBMid65[11] , \wBMid65[10] , \wBMid65[9] , \wBMid65[8] , \wBMid65[7] , 
        \wBMid65[6] , \wBMid65[5] , \wBMid65[4] , \wBMid65[3] , \wBMid65[2] , 
        \wBMid65[1] , \wBMid65[0] }), .LoOut({\wAMid66[31] , \wAMid66[30] , 
        \wAMid66[29] , \wAMid66[28] , \wAMid66[27] , \wAMid66[26] , 
        \wAMid66[25] , \wAMid66[24] , \wAMid66[23] , \wAMid66[22] , 
        \wAMid66[21] , \wAMid66[20] , \wAMid66[19] , \wAMid66[18] , 
        \wAMid66[17] , \wAMid66[16] , \wAMid66[15] , \wAMid66[14] , 
        \wAMid66[13] , \wAMid66[12] , \wAMid66[11] , \wAMid66[10] , 
        \wAMid66[9] , \wAMid66[8] , \wAMid66[7] , \wAMid66[6] , \wAMid66[5] , 
        \wAMid66[4] , \wAMid66[3] , \wAMid66[2] , \wAMid66[1] , \wAMid66[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn116[31] , \wAIn116[30] , \wAIn116[29] , \wAIn116[28] , 
        \wAIn116[27] , \wAIn116[26] , \wAIn116[25] , \wAIn116[24] , 
        \wAIn116[23] , \wAIn116[22] , \wAIn116[21] , \wAIn116[20] , 
        \wAIn116[19] , \wAIn116[18] , \wAIn116[17] , \wAIn116[16] , 
        \wAIn116[15] , \wAIn116[14] , \wAIn116[13] , \wAIn116[12] , 
        \wAIn116[11] , \wAIn116[10] , \wAIn116[9] , \wAIn116[8] , \wAIn116[7] , 
        \wAIn116[6] , \wAIn116[5] , \wAIn116[4] , \wAIn116[3] , \wAIn116[2] , 
        \wAIn116[1] , \wAIn116[0] }), .BIn({\wBIn116[31] , \wBIn116[30] , 
        \wBIn116[29] , \wBIn116[28] , \wBIn116[27] , \wBIn116[26] , 
        \wBIn116[25] , \wBIn116[24] , \wBIn116[23] , \wBIn116[22] , 
        \wBIn116[21] , \wBIn116[20] , \wBIn116[19] , \wBIn116[18] , 
        \wBIn116[17] , \wBIn116[16] , \wBIn116[15] , \wBIn116[14] , 
        \wBIn116[13] , \wBIn116[12] , \wBIn116[11] , \wBIn116[10] , 
        \wBIn116[9] , \wBIn116[8] , \wBIn116[7] , \wBIn116[6] , \wBIn116[5] , 
        \wBIn116[4] , \wBIn116[3] , \wBIn116[2] , \wBIn116[1] , \wBIn116[0] }), 
        .HiOut({\wBMid115[31] , \wBMid115[30] , \wBMid115[29] , \wBMid115[28] , 
        \wBMid115[27] , \wBMid115[26] , \wBMid115[25] , \wBMid115[24] , 
        \wBMid115[23] , \wBMid115[22] , \wBMid115[21] , \wBMid115[20] , 
        \wBMid115[19] , \wBMid115[18] , \wBMid115[17] , \wBMid115[16] , 
        \wBMid115[15] , \wBMid115[14] , \wBMid115[13] , \wBMid115[12] , 
        \wBMid115[11] , \wBMid115[10] , \wBMid115[9] , \wBMid115[8] , 
        \wBMid115[7] , \wBMid115[6] , \wBMid115[5] , \wBMid115[4] , 
        \wBMid115[3] , \wBMid115[2] , \wBMid115[1] , \wBMid115[0] }), .LoOut({
        \wAMid116[31] , \wAMid116[30] , \wAMid116[29] , \wAMid116[28] , 
        \wAMid116[27] , \wAMid116[26] , \wAMid116[25] , \wAMid116[24] , 
        \wAMid116[23] , \wAMid116[22] , \wAMid116[21] , \wAMid116[20] , 
        \wAMid116[19] , \wAMid116[18] , \wAMid116[17] , \wAMid116[16] , 
        \wAMid116[15] , \wAMid116[14] , \wAMid116[13] , \wAMid116[12] , 
        \wAMid116[11] , \wAMid116[10] , \wAMid116[9] , \wAMid116[8] , 
        \wAMid116[7] , \wAMid116[6] , \wAMid116[5] , \wAMid116[4] , 
        \wAMid116[3] , \wAMid116[2] , \wAMid116[1] , \wAMid116[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid71[31] , \wAMid71[30] , \wAMid71[29] , \wAMid71[28] , 
        \wAMid71[27] , \wAMid71[26] , \wAMid71[25] , \wAMid71[24] , 
        \wAMid71[23] , \wAMid71[22] , \wAMid71[21] , \wAMid71[20] , 
        \wAMid71[19] , \wAMid71[18] , \wAMid71[17] , \wAMid71[16] , 
        \wAMid71[15] , \wAMid71[14] , \wAMid71[13] , \wAMid71[12] , 
        \wAMid71[11] , \wAMid71[10] , \wAMid71[9] , \wAMid71[8] , \wAMid71[7] , 
        \wAMid71[6] , \wAMid71[5] , \wAMid71[4] , \wAMid71[3] , \wAMid71[2] , 
        \wAMid71[1] , \wAMid71[0] }), .BIn({\wBMid71[31] , \wBMid71[30] , 
        \wBMid71[29] , \wBMid71[28] , \wBMid71[27] , \wBMid71[26] , 
        \wBMid71[25] , \wBMid71[24] , \wBMid71[23] , \wBMid71[22] , 
        \wBMid71[21] , \wBMid71[20] , \wBMid71[19] , \wBMid71[18] , 
        \wBMid71[17] , \wBMid71[16] , \wBMid71[15] , \wBMid71[14] , 
        \wBMid71[13] , \wBMid71[12] , \wBMid71[11] , \wBMid71[10] , 
        \wBMid71[9] , \wBMid71[8] , \wBMid71[7] , \wBMid71[6] , \wBMid71[5] , 
        \wBMid71[4] , \wBMid71[3] , \wBMid71[2] , \wBMid71[1] , \wBMid71[0] }), 
        .HiOut({\wRegInB71[31] , \wRegInB71[30] , \wRegInB71[29] , 
        \wRegInB71[28] , \wRegInB71[27] , \wRegInB71[26] , \wRegInB71[25] , 
        \wRegInB71[24] , \wRegInB71[23] , \wRegInB71[22] , \wRegInB71[21] , 
        \wRegInB71[20] , \wRegInB71[19] , \wRegInB71[18] , \wRegInB71[17] , 
        \wRegInB71[16] , \wRegInB71[15] , \wRegInB71[14] , \wRegInB71[13] , 
        \wRegInB71[12] , \wRegInB71[11] , \wRegInB71[10] , \wRegInB71[9] , 
        \wRegInB71[8] , \wRegInB71[7] , \wRegInB71[6] , \wRegInB71[5] , 
        \wRegInB71[4] , \wRegInB71[3] , \wRegInB71[2] , \wRegInB71[1] , 
        \wRegInB71[0] }), .LoOut({\wRegInA72[31] , \wRegInA72[30] , 
        \wRegInA72[29] , \wRegInA72[28] , \wRegInA72[27] , \wRegInA72[26] , 
        \wRegInA72[25] , \wRegInA72[24] , \wRegInA72[23] , \wRegInA72[22] , 
        \wRegInA72[21] , \wRegInA72[20] , \wRegInA72[19] , \wRegInA72[18] , 
        \wRegInA72[17] , \wRegInA72[16] , \wRegInA72[15] , \wRegInA72[14] , 
        \wRegInA72[13] , \wRegInA72[12] , \wRegInA72[11] , \wRegInA72[10] , 
        \wRegInA72[9] , \wRegInA72[8] , \wRegInA72[7] , \wRegInA72[6] , 
        \wRegInA72[5] , \wRegInA72[4] , \wRegInA72[3] , \wRegInA72[2] , 
        \wRegInA72[1] , \wRegInA72[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_144 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink145[31] , \ScanLink145[30] , \ScanLink145[29] , 
        \ScanLink145[28] , \ScanLink145[27] , \ScanLink145[26] , 
        \ScanLink145[25] , \ScanLink145[24] , \ScanLink145[23] , 
        \ScanLink145[22] , \ScanLink145[21] , \ScanLink145[20] , 
        \ScanLink145[19] , \ScanLink145[18] , \ScanLink145[17] , 
        \ScanLink145[16] , \ScanLink145[15] , \ScanLink145[14] , 
        \ScanLink145[13] , \ScanLink145[12] , \ScanLink145[11] , 
        \ScanLink145[10] , \ScanLink145[9] , \ScanLink145[8] , 
        \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , \ScanLink145[4] , 
        \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , \ScanLink145[0] 
        }), .ScanOut({\ScanLink144[31] , \ScanLink144[30] , \ScanLink144[29] , 
        \ScanLink144[28] , \ScanLink144[27] , \ScanLink144[26] , 
        \ScanLink144[25] , \ScanLink144[24] , \ScanLink144[23] , 
        \ScanLink144[22] , \ScanLink144[21] , \ScanLink144[20] , 
        \ScanLink144[19] , \ScanLink144[18] , \ScanLink144[17] , 
        \ScanLink144[16] , \ScanLink144[15] , \ScanLink144[14] , 
        \ScanLink144[13] , \ScanLink144[12] , \ScanLink144[11] , 
        \ScanLink144[10] , \ScanLink144[9] , \ScanLink144[8] , 
        \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , \ScanLink144[4] , 
        \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , \ScanLink144[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB55[31] , \wRegInB55[30] , \wRegInB55[29] , 
        \wRegInB55[28] , \wRegInB55[27] , \wRegInB55[26] , \wRegInB55[25] , 
        \wRegInB55[24] , \wRegInB55[23] , \wRegInB55[22] , \wRegInB55[21] , 
        \wRegInB55[20] , \wRegInB55[19] , \wRegInB55[18] , \wRegInB55[17] , 
        \wRegInB55[16] , \wRegInB55[15] , \wRegInB55[14] , \wRegInB55[13] , 
        \wRegInB55[12] , \wRegInB55[11] , \wRegInB55[10] , \wRegInB55[9] , 
        \wRegInB55[8] , \wRegInB55[7] , \wRegInB55[6] , \wRegInB55[5] , 
        \wRegInB55[4] , \wRegInB55[3] , \wRegInB55[2] , \wRegInB55[1] , 
        \wRegInB55[0] }), .Out({\wBIn55[31] , \wBIn55[30] , \wBIn55[29] , 
        \wBIn55[28] , \wBIn55[27] , \wBIn55[26] , \wBIn55[25] , \wBIn55[24] , 
        \wBIn55[23] , \wBIn55[22] , \wBIn55[21] , \wBIn55[20] , \wBIn55[19] , 
        \wBIn55[18] , \wBIn55[17] , \wBIn55[16] , \wBIn55[15] , \wBIn55[14] , 
        \wBIn55[13] , \wBIn55[12] , \wBIn55[11] , \wBIn55[10] , \wBIn55[9] , 
        \wBIn55[8] , \wBIn55[7] , \wBIn55[6] , \wBIn55[5] , \wBIn55[4] , 
        \wBIn55[3] , \wBIn55[2] , \wBIn55[1] , \wBIn55[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_14 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[31] , \ScanLink15[30] , \ScanLink15[29] , 
        \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , \ScanLink15[25] , 
        \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , \ScanLink15[21] , 
        \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , \ScanLink15[17] , 
        \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , \ScanLink15[13] , 
        \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , \ScanLink15[9] , 
        \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB120[31] , \wRegInB120[30] , 
        \wRegInB120[29] , \wRegInB120[28] , \wRegInB120[27] , \wRegInB120[26] , 
        \wRegInB120[25] , \wRegInB120[24] , \wRegInB120[23] , \wRegInB120[22] , 
        \wRegInB120[21] , \wRegInB120[20] , \wRegInB120[19] , \wRegInB120[18] , 
        \wRegInB120[17] , \wRegInB120[16] , \wRegInB120[15] , \wRegInB120[14] , 
        \wRegInB120[13] , \wRegInB120[12] , \wRegInB120[11] , \wRegInB120[10] , 
        \wRegInB120[9] , \wRegInB120[8] , \wRegInB120[7] , \wRegInB120[6] , 
        \wRegInB120[5] , \wRegInB120[4] , \wRegInB120[3] , \wRegInB120[2] , 
        \wRegInB120[1] , \wRegInB120[0] }), .Out({\wBIn120[31] , \wBIn120[30] , 
        \wBIn120[29] , \wBIn120[28] , \wBIn120[27] , \wBIn120[26] , 
        \wBIn120[25] , \wBIn120[24] , \wBIn120[23] , \wBIn120[22] , 
        \wBIn120[21] , \wBIn120[20] , \wBIn120[19] , \wBIn120[18] , 
        \wBIn120[17] , \wBIn120[16] , \wBIn120[15] , \wBIn120[14] , 
        \wBIn120[13] , \wBIn120[12] , \wBIn120[11] , \wBIn120[10] , 
        \wBIn120[9] , \wBIn120[8] , \wBIn120[7] , \wBIn120[6] , \wBIn120[5] , 
        \wBIn120[4] , \wBIn120[3] , \wBIn120[2] , \wBIn120[1] , \wBIn120[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_253 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink254[31] , \ScanLink254[30] , \ScanLink254[29] , 
        \ScanLink254[28] , \ScanLink254[27] , \ScanLink254[26] , 
        \ScanLink254[25] , \ScanLink254[24] , \ScanLink254[23] , 
        \ScanLink254[22] , \ScanLink254[21] , \ScanLink254[20] , 
        \ScanLink254[19] , \ScanLink254[18] , \ScanLink254[17] , 
        \ScanLink254[16] , \ScanLink254[15] , \ScanLink254[14] , 
        \ScanLink254[13] , \ScanLink254[12] , \ScanLink254[11] , 
        \ScanLink254[10] , \ScanLink254[9] , \ScanLink254[8] , 
        \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , \ScanLink254[4] , 
        \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , \ScanLink254[0] 
        }), .ScanOut({\ScanLink253[31] , \ScanLink253[30] , \ScanLink253[29] , 
        \ScanLink253[28] , \ScanLink253[27] , \ScanLink253[26] , 
        \ScanLink253[25] , \ScanLink253[24] , \ScanLink253[23] , 
        \ScanLink253[22] , \ScanLink253[21] , \ScanLink253[20] , 
        \ScanLink253[19] , \ScanLink253[18] , \ScanLink253[17] , 
        \ScanLink253[16] , \ScanLink253[15] , \ScanLink253[14] , 
        \ScanLink253[13] , \ScanLink253[12] , \ScanLink253[11] , 
        \ScanLink253[10] , \ScanLink253[9] , \ScanLink253[8] , 
        \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , \ScanLink253[4] , 
        \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , \ScanLink253[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA1[31] , \wRegInA1[30] , \wRegInA1[29] , \wRegInA1[28] , 
        \wRegInA1[27] , \wRegInA1[26] , \wRegInA1[25] , \wRegInA1[24] , 
        \wRegInA1[23] , \wRegInA1[22] , \wRegInA1[21] , \wRegInA1[20] , 
        \wRegInA1[19] , \wRegInA1[18] , \wRegInA1[17] , \wRegInA1[16] , 
        \wRegInA1[15] , \wRegInA1[14] , \wRegInA1[13] , \wRegInA1[12] , 
        \wRegInA1[11] , \wRegInA1[10] , \wRegInA1[9] , \wRegInA1[8] , 
        \wRegInA1[7] , \wRegInA1[6] , \wRegInA1[5] , \wRegInA1[4] , 
        \wRegInA1[3] , \wRegInA1[2] , \wRegInA1[1] , \wRegInA1[0] }), .Out({
        \wAIn1[31] , \wAIn1[30] , \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , 
        \wAIn1[26] , \wAIn1[25] , \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , 
        \wAIn1[21] , \wAIn1[20] , \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , 
        \wAIn1[16] , \wAIn1[15] , \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , 
        \wAIn1[11] , \wAIn1[10] , \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , 
        \wAIn1[6] , \wAIn1[5] , \wAIn1[4] , \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , 
        \wAIn1[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn83[31] , \wAIn83[30] , \wAIn83[29] , \wAIn83[28] , \wAIn83[27] , 
        \wAIn83[26] , \wAIn83[25] , \wAIn83[24] , \wAIn83[23] , \wAIn83[22] , 
        \wAIn83[21] , \wAIn83[20] , \wAIn83[19] , \wAIn83[18] , \wAIn83[17] , 
        \wAIn83[16] , \wAIn83[15] , \wAIn83[14] , \wAIn83[13] , \wAIn83[12] , 
        \wAIn83[11] , \wAIn83[10] , \wAIn83[9] , \wAIn83[8] , \wAIn83[7] , 
        \wAIn83[6] , \wAIn83[5] , \wAIn83[4] , \wAIn83[3] , \wAIn83[2] , 
        \wAIn83[1] , \wAIn83[0] }), .BIn({\wBIn83[31] , \wBIn83[30] , 
        \wBIn83[29] , \wBIn83[28] , \wBIn83[27] , \wBIn83[26] , \wBIn83[25] , 
        \wBIn83[24] , \wBIn83[23] , \wBIn83[22] , \wBIn83[21] , \wBIn83[20] , 
        \wBIn83[19] , \wBIn83[18] , \wBIn83[17] , \wBIn83[16] , \wBIn83[15] , 
        \wBIn83[14] , \wBIn83[13] , \wBIn83[12] , \wBIn83[11] , \wBIn83[10] , 
        \wBIn83[9] , \wBIn83[8] , \wBIn83[7] , \wBIn83[6] , \wBIn83[5] , 
        \wBIn83[4] , \wBIn83[3] , \wBIn83[2] , \wBIn83[1] , \wBIn83[0] }), 
        .HiOut({\wBMid82[31] , \wBMid82[30] , \wBMid82[29] , \wBMid82[28] , 
        \wBMid82[27] , \wBMid82[26] , \wBMid82[25] , \wBMid82[24] , 
        \wBMid82[23] , \wBMid82[22] , \wBMid82[21] , \wBMid82[20] , 
        \wBMid82[19] , \wBMid82[18] , \wBMid82[17] , \wBMid82[16] , 
        \wBMid82[15] , \wBMid82[14] , \wBMid82[13] , \wBMid82[12] , 
        \wBMid82[11] , \wBMid82[10] , \wBMid82[9] , \wBMid82[8] , \wBMid82[7] , 
        \wBMid82[6] , \wBMid82[5] , \wBMid82[4] , \wBMid82[3] , \wBMid82[2] , 
        \wBMid82[1] , \wBMid82[0] }), .LoOut({\wAMid83[31] , \wAMid83[30] , 
        \wAMid83[29] , \wAMid83[28] , \wAMid83[27] , \wAMid83[26] , 
        \wAMid83[25] , \wAMid83[24] , \wAMid83[23] , \wAMid83[22] , 
        \wAMid83[21] , \wAMid83[20] , \wAMid83[19] , \wAMid83[18] , 
        \wAMid83[17] , \wAMid83[16] , \wAMid83[15] , \wAMid83[14] , 
        \wAMid83[13] , \wAMid83[12] , \wAMid83[11] , \wAMid83[10] , 
        \wAMid83[9] , \wAMid83[8] , \wAMid83[7] , \wAMid83[6] , \wAMid83[5] , 
        \wAMid83[4] , \wAMid83[3] , \wAMid83[2] , \wAMid83[1] , \wAMid83[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid38[31] , \wAMid38[30] , \wAMid38[29] , \wAMid38[28] , 
        \wAMid38[27] , \wAMid38[26] , \wAMid38[25] , \wAMid38[24] , 
        \wAMid38[23] , \wAMid38[22] , \wAMid38[21] , \wAMid38[20] , 
        \wAMid38[19] , \wAMid38[18] , \wAMid38[17] , \wAMid38[16] , 
        \wAMid38[15] , \wAMid38[14] , \wAMid38[13] , \wAMid38[12] , 
        \wAMid38[11] , \wAMid38[10] , \wAMid38[9] , \wAMid38[8] , \wAMid38[7] , 
        \wAMid38[6] , \wAMid38[5] , \wAMid38[4] , \wAMid38[3] , \wAMid38[2] , 
        \wAMid38[1] , \wAMid38[0] }), .BIn({\wBMid38[31] , \wBMid38[30] , 
        \wBMid38[29] , \wBMid38[28] , \wBMid38[27] , \wBMid38[26] , 
        \wBMid38[25] , \wBMid38[24] , \wBMid38[23] , \wBMid38[22] , 
        \wBMid38[21] , \wBMid38[20] , \wBMid38[19] , \wBMid38[18] , 
        \wBMid38[17] , \wBMid38[16] , \wBMid38[15] , \wBMid38[14] , 
        \wBMid38[13] , \wBMid38[12] , \wBMid38[11] , \wBMid38[10] , 
        \wBMid38[9] , \wBMid38[8] , \wBMid38[7] , \wBMid38[6] , \wBMid38[5] , 
        \wBMid38[4] , \wBMid38[3] , \wBMid38[2] , \wBMid38[1] , \wBMid38[0] }), 
        .HiOut({\wRegInB38[31] , \wRegInB38[30] , \wRegInB38[29] , 
        \wRegInB38[28] , \wRegInB38[27] , \wRegInB38[26] , \wRegInB38[25] , 
        \wRegInB38[24] , \wRegInB38[23] , \wRegInB38[22] , \wRegInB38[21] , 
        \wRegInB38[20] , \wRegInB38[19] , \wRegInB38[18] , \wRegInB38[17] , 
        \wRegInB38[16] , \wRegInB38[15] , \wRegInB38[14] , \wRegInB38[13] , 
        \wRegInB38[12] , \wRegInB38[11] , \wRegInB38[10] , \wRegInB38[9] , 
        \wRegInB38[8] , \wRegInB38[7] , \wRegInB38[6] , \wRegInB38[5] , 
        \wRegInB38[4] , \wRegInB38[3] , \wRegInB38[2] , \wRegInB38[1] , 
        \wRegInB38[0] }), .LoOut({\wRegInA39[31] , \wRegInA39[30] , 
        \wRegInA39[29] , \wRegInA39[28] , \wRegInA39[27] , \wRegInA39[26] , 
        \wRegInA39[25] , \wRegInA39[24] , \wRegInA39[23] , \wRegInA39[22] , 
        \wRegInA39[21] , \wRegInA39[20] , \wRegInA39[19] , \wRegInA39[18] , 
        \wRegInA39[17] , \wRegInA39[16] , \wRegInA39[15] , \wRegInA39[14] , 
        \wRegInA39[13] , \wRegInA39[12] , \wRegInA39[11] , \wRegInA39[10] , 
        \wRegInA39[9] , \wRegInA39[8] , \wRegInA39[7] , \wRegInA39[6] , 
        \wRegInA39[5] , \wRegInA39[4] , \wRegInA39[3] , \wRegInA39[2] , 
        \wRegInA39[1] , \wRegInA39[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid56[31] , \wAMid56[30] , \wAMid56[29] , \wAMid56[28] , 
        \wAMid56[27] , \wAMid56[26] , \wAMid56[25] , \wAMid56[24] , 
        \wAMid56[23] , \wAMid56[22] , \wAMid56[21] , \wAMid56[20] , 
        \wAMid56[19] , \wAMid56[18] , \wAMid56[17] , \wAMid56[16] , 
        \wAMid56[15] , \wAMid56[14] , \wAMid56[13] , \wAMid56[12] , 
        \wAMid56[11] , \wAMid56[10] , \wAMid56[9] , \wAMid56[8] , \wAMid56[7] , 
        \wAMid56[6] , \wAMid56[5] , \wAMid56[4] , \wAMid56[3] , \wAMid56[2] , 
        \wAMid56[1] , \wAMid56[0] }), .BIn({\wBMid56[31] , \wBMid56[30] , 
        \wBMid56[29] , \wBMid56[28] , \wBMid56[27] , \wBMid56[26] , 
        \wBMid56[25] , \wBMid56[24] , \wBMid56[23] , \wBMid56[22] , 
        \wBMid56[21] , \wBMid56[20] , \wBMid56[19] , \wBMid56[18] , 
        \wBMid56[17] , \wBMid56[16] , \wBMid56[15] , \wBMid56[14] , 
        \wBMid56[13] , \wBMid56[12] , \wBMid56[11] , \wBMid56[10] , 
        \wBMid56[9] , \wBMid56[8] , \wBMid56[7] , \wBMid56[6] , \wBMid56[5] , 
        \wBMid56[4] , \wBMid56[3] , \wBMid56[2] , \wBMid56[1] , \wBMid56[0] }), 
        .HiOut({\wRegInB56[31] , \wRegInB56[30] , \wRegInB56[29] , 
        \wRegInB56[28] , \wRegInB56[27] , \wRegInB56[26] , \wRegInB56[25] , 
        \wRegInB56[24] , \wRegInB56[23] , \wRegInB56[22] , \wRegInB56[21] , 
        \wRegInB56[20] , \wRegInB56[19] , \wRegInB56[18] , \wRegInB56[17] , 
        \wRegInB56[16] , \wRegInB56[15] , \wRegInB56[14] , \wRegInB56[13] , 
        \wRegInB56[12] , \wRegInB56[11] , \wRegInB56[10] , \wRegInB56[9] , 
        \wRegInB56[8] , \wRegInB56[7] , \wRegInB56[6] , \wRegInB56[5] , 
        \wRegInB56[4] , \wRegInB56[3] , \wRegInB56[2] , \wRegInB56[1] , 
        \wRegInB56[0] }), .LoOut({\wRegInA57[31] , \wRegInA57[30] , 
        \wRegInA57[29] , \wRegInA57[28] , \wRegInA57[27] , \wRegInA57[26] , 
        \wRegInA57[25] , \wRegInA57[24] , \wRegInA57[23] , \wRegInA57[22] , 
        \wRegInA57[21] , \wRegInA57[20] , \wRegInA57[19] , \wRegInA57[18] , 
        \wRegInA57[17] , \wRegInA57[16] , \wRegInA57[15] , \wRegInA57[14] , 
        \wRegInA57[13] , \wRegInA57[12] , \wRegInA57[11] , \wRegInA57[10] , 
        \wRegInA57[9] , \wRegInA57[8] , \wRegInA57[7] , \wRegInA57[6] , 
        \wRegInA57[5] , \wRegInA57[4] , \wRegInA57[3] , \wRegInA57[2] , 
        \wRegInA57[1] , \wRegInA57[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_163 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink164[31] , \ScanLink164[30] , \ScanLink164[29] , 
        \ScanLink164[28] , \ScanLink164[27] , \ScanLink164[26] , 
        \ScanLink164[25] , \ScanLink164[24] , \ScanLink164[23] , 
        \ScanLink164[22] , \ScanLink164[21] , \ScanLink164[20] , 
        \ScanLink164[19] , \ScanLink164[18] , \ScanLink164[17] , 
        \ScanLink164[16] , \ScanLink164[15] , \ScanLink164[14] , 
        \ScanLink164[13] , \ScanLink164[12] , \ScanLink164[11] , 
        \ScanLink164[10] , \ScanLink164[9] , \ScanLink164[8] , 
        \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , \ScanLink164[4] , 
        \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , \ScanLink164[0] 
        }), .ScanOut({\ScanLink163[31] , \ScanLink163[30] , \ScanLink163[29] , 
        \ScanLink163[28] , \ScanLink163[27] , \ScanLink163[26] , 
        \ScanLink163[25] , \ScanLink163[24] , \ScanLink163[23] , 
        \ScanLink163[22] , \ScanLink163[21] , \ScanLink163[20] , 
        \ScanLink163[19] , \ScanLink163[18] , \ScanLink163[17] , 
        \ScanLink163[16] , \ScanLink163[15] , \ScanLink163[14] , 
        \ScanLink163[13] , \ScanLink163[12] , \ScanLink163[11] , 
        \ScanLink163[10] , \ScanLink163[9] , \ScanLink163[8] , 
        \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , \ScanLink163[4] , 
        \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , \ScanLink163[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA46[31] , \wRegInA46[30] , \wRegInA46[29] , 
        \wRegInA46[28] , \wRegInA46[27] , \wRegInA46[26] , \wRegInA46[25] , 
        \wRegInA46[24] , \wRegInA46[23] , \wRegInA46[22] , \wRegInA46[21] , 
        \wRegInA46[20] , \wRegInA46[19] , \wRegInA46[18] , \wRegInA46[17] , 
        \wRegInA46[16] , \wRegInA46[15] , \wRegInA46[14] , \wRegInA46[13] , 
        \wRegInA46[12] , \wRegInA46[11] , \wRegInA46[10] , \wRegInA46[9] , 
        \wRegInA46[8] , \wRegInA46[7] , \wRegInA46[6] , \wRegInA46[5] , 
        \wRegInA46[4] , \wRegInA46[3] , \wRegInA46[2] , \wRegInA46[1] , 
        \wRegInA46[0] }), .Out({\wAIn46[31] , \wAIn46[30] , \wAIn46[29] , 
        \wAIn46[28] , \wAIn46[27] , \wAIn46[26] , \wAIn46[25] , \wAIn46[24] , 
        \wAIn46[23] , \wAIn46[22] , \wAIn46[21] , \wAIn46[20] , \wAIn46[19] , 
        \wAIn46[18] , \wAIn46[17] , \wAIn46[16] , \wAIn46[15] , \wAIn46[14] , 
        \wAIn46[13] , \wAIn46[12] , \wAIn46[11] , \wAIn46[10] , \wAIn46[9] , 
        \wAIn46[8] , \wAIn46[7] , \wAIn46[6] , \wAIn46[5] , \wAIn46[4] , 
        \wAIn46[3] , \wAIn46[2] , \wAIn46[1] , \wAIn46[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_33 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink34[31] , \ScanLink34[30] , \ScanLink34[29] , 
        \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , \ScanLink34[25] , 
        \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , \ScanLink34[21] , 
        \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , \ScanLink34[17] , 
        \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , \ScanLink34[13] , 
        \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , \ScanLink34[9] , 
        \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , \ScanLink34[5] , 
        \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , \ScanLink34[1] , 
        \ScanLink34[0] }), .ScanOut({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA111[31] , \wRegInA111[30] , 
        \wRegInA111[29] , \wRegInA111[28] , \wRegInA111[27] , \wRegInA111[26] , 
        \wRegInA111[25] , \wRegInA111[24] , \wRegInA111[23] , \wRegInA111[22] , 
        \wRegInA111[21] , \wRegInA111[20] , \wRegInA111[19] , \wRegInA111[18] , 
        \wRegInA111[17] , \wRegInA111[16] , \wRegInA111[15] , \wRegInA111[14] , 
        \wRegInA111[13] , \wRegInA111[12] , \wRegInA111[11] , \wRegInA111[10] , 
        \wRegInA111[9] , \wRegInA111[8] , \wRegInA111[7] , \wRegInA111[6] , 
        \wRegInA111[5] , \wRegInA111[4] , \wRegInA111[3] , \wRegInA111[2] , 
        \wRegInA111[1] , \wRegInA111[0] }), .Out({\wAIn111[31] , \wAIn111[30] , 
        \wAIn111[29] , \wAIn111[28] , \wAIn111[27] , \wAIn111[26] , 
        \wAIn111[25] , \wAIn111[24] , \wAIn111[23] , \wAIn111[22] , 
        \wAIn111[21] , \wAIn111[20] , \wAIn111[19] , \wAIn111[18] , 
        \wAIn111[17] , \wAIn111[16] , \wAIn111[15] , \wAIn111[14] , 
        \wAIn111[13] , \wAIn111[12] , \wAIn111[11] , \wAIn111[10] , 
        \wAIn111[9] , \wAIn111[8] , \wAIn111[7] , \wAIn111[6] , \wAIn111[5] , 
        \wAIn111[4] , \wAIn111[3] , \wAIn111[2] , \wAIn111[1] , \wAIn111[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_186 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink187[31] , \ScanLink187[30] , \ScanLink187[29] , 
        \ScanLink187[28] , \ScanLink187[27] , \ScanLink187[26] , 
        \ScanLink187[25] , \ScanLink187[24] , \ScanLink187[23] , 
        \ScanLink187[22] , \ScanLink187[21] , \ScanLink187[20] , 
        \ScanLink187[19] , \ScanLink187[18] , \ScanLink187[17] , 
        \ScanLink187[16] , \ScanLink187[15] , \ScanLink187[14] , 
        \ScanLink187[13] , \ScanLink187[12] , \ScanLink187[11] , 
        \ScanLink187[10] , \ScanLink187[9] , \ScanLink187[8] , 
        \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , \ScanLink187[4] , 
        \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , \ScanLink187[0] 
        }), .ScanOut({\ScanLink186[31] , \ScanLink186[30] , \ScanLink186[29] , 
        \ScanLink186[28] , \ScanLink186[27] , \ScanLink186[26] , 
        \ScanLink186[25] , \ScanLink186[24] , \ScanLink186[23] , 
        \ScanLink186[22] , \ScanLink186[21] , \ScanLink186[20] , 
        \ScanLink186[19] , \ScanLink186[18] , \ScanLink186[17] , 
        \ScanLink186[16] , \ScanLink186[15] , \ScanLink186[14] , 
        \ScanLink186[13] , \ScanLink186[12] , \ScanLink186[11] , 
        \ScanLink186[10] , \ScanLink186[9] , \ScanLink186[8] , 
        \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , \ScanLink186[4] , 
        \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , \ScanLink186[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB34[31] , \wRegInB34[30] , \wRegInB34[29] , 
        \wRegInB34[28] , \wRegInB34[27] , \wRegInB34[26] , \wRegInB34[25] , 
        \wRegInB34[24] , \wRegInB34[23] , \wRegInB34[22] , \wRegInB34[21] , 
        \wRegInB34[20] , \wRegInB34[19] , \wRegInB34[18] , \wRegInB34[17] , 
        \wRegInB34[16] , \wRegInB34[15] , \wRegInB34[14] , \wRegInB34[13] , 
        \wRegInB34[12] , \wRegInB34[11] , \wRegInB34[10] , \wRegInB34[9] , 
        \wRegInB34[8] , \wRegInB34[7] , \wRegInB34[6] , \wRegInB34[5] , 
        \wRegInB34[4] , \wRegInB34[3] , \wRegInB34[2] , \wRegInB34[1] , 
        \wRegInB34[0] }), .Out({\wBIn34[31] , \wBIn34[30] , \wBIn34[29] , 
        \wBIn34[28] , \wBIn34[27] , \wBIn34[26] , \wBIn34[25] , \wBIn34[24] , 
        \wBIn34[23] , \wBIn34[22] , \wBIn34[21] , \wBIn34[20] , \wBIn34[19] , 
        \wBIn34[18] , \wBIn34[17] , \wBIn34[16] , \wBIn34[15] , \wBIn34[14] , 
        \wBIn34[13] , \wBIn34[12] , \wBIn34[11] , \wBIn34[10] , \wBIn34[9] , 
        \wBIn34[8] , \wBIn34[7] , \wBIn34[6] , \wBIn34[5] , \wBIn34[4] , 
        \wBIn34[3] , \wBIn34[2] , \wBIn34[1] , \wBIn34[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid94[31] , \wAMid94[30] , \wAMid94[29] , \wAMid94[28] , 
        \wAMid94[27] , \wAMid94[26] , \wAMid94[25] , \wAMid94[24] , 
        \wAMid94[23] , \wAMid94[22] , \wAMid94[21] , \wAMid94[20] , 
        \wAMid94[19] , \wAMid94[18] , \wAMid94[17] , \wAMid94[16] , 
        \wAMid94[15] , \wAMid94[14] , \wAMid94[13] , \wAMid94[12] , 
        \wAMid94[11] , \wAMid94[10] , \wAMid94[9] , \wAMid94[8] , \wAMid94[7] , 
        \wAMid94[6] , \wAMid94[5] , \wAMid94[4] , \wAMid94[3] , \wAMid94[2] , 
        \wAMid94[1] , \wAMid94[0] }), .BIn({\wBMid94[31] , \wBMid94[30] , 
        \wBMid94[29] , \wBMid94[28] , \wBMid94[27] , \wBMid94[26] , 
        \wBMid94[25] , \wBMid94[24] , \wBMid94[23] , \wBMid94[22] , 
        \wBMid94[21] , \wBMid94[20] , \wBMid94[19] , \wBMid94[18] , 
        \wBMid94[17] , \wBMid94[16] , \wBMid94[15] , \wBMid94[14] , 
        \wBMid94[13] , \wBMid94[12] , \wBMid94[11] , \wBMid94[10] , 
        \wBMid94[9] , \wBMid94[8] , \wBMid94[7] , \wBMid94[6] , \wBMid94[5] , 
        \wBMid94[4] , \wBMid94[3] , \wBMid94[2] , \wBMid94[1] , \wBMid94[0] }), 
        .HiOut({\wRegInB94[31] , \wRegInB94[30] , \wRegInB94[29] , 
        \wRegInB94[28] , \wRegInB94[27] , \wRegInB94[26] , \wRegInB94[25] , 
        \wRegInB94[24] , \wRegInB94[23] , \wRegInB94[22] , \wRegInB94[21] , 
        \wRegInB94[20] , \wRegInB94[19] , \wRegInB94[18] , \wRegInB94[17] , 
        \wRegInB94[16] , \wRegInB94[15] , \wRegInB94[14] , \wRegInB94[13] , 
        \wRegInB94[12] , \wRegInB94[11] , \wRegInB94[10] , \wRegInB94[9] , 
        \wRegInB94[8] , \wRegInB94[7] , \wRegInB94[6] , \wRegInB94[5] , 
        \wRegInB94[4] , \wRegInB94[3] , \wRegInB94[2] , \wRegInB94[1] , 
        \wRegInB94[0] }), .LoOut({\wRegInA95[31] , \wRegInA95[30] , 
        \wRegInA95[29] , \wRegInA95[28] , \wRegInA95[27] , \wRegInA95[26] , 
        \wRegInA95[25] , \wRegInA95[24] , \wRegInA95[23] , \wRegInA95[22] , 
        \wRegInA95[21] , \wRegInA95[20] , \wRegInA95[19] , \wRegInA95[18] , 
        \wRegInA95[17] , \wRegInA95[16] , \wRegInA95[15] , \wRegInA95[14] , 
        \wRegInA95[13] , \wRegInA95[12] , \wRegInA95[11] , \wRegInA95[10] , 
        \wRegInA95[9] , \wRegInA95[8] , \wRegInA95[7] , \wRegInA95[6] , 
        \wRegInA95[5] , \wRegInA95[4] , \wRegInA95[3] , \wRegInA95[2] , 
        \wRegInA95[1] , \wRegInA95[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn7[31] , 
        \wAIn7[30] , \wAIn7[29] , \wAIn7[28] , \wAIn7[27] , \wAIn7[26] , 
        \wAIn7[25] , \wAIn7[24] , \wAIn7[23] , \wAIn7[22] , \wAIn7[21] , 
        \wAIn7[20] , \wAIn7[19] , \wAIn7[18] , \wAIn7[17] , \wAIn7[16] , 
        \wAIn7[15] , \wAIn7[14] , \wAIn7[13] , \wAIn7[12] , \wAIn7[11] , 
        \wAIn7[10] , \wAIn7[9] , \wAIn7[8] , \wAIn7[7] , \wAIn7[6] , 
        \wAIn7[5] , \wAIn7[4] , \wAIn7[3] , \wAIn7[2] , \wAIn7[1] , \wAIn7[0] 
        }), .BIn({\wBIn7[31] , \wBIn7[30] , \wBIn7[29] , \wBIn7[28] , 
        \wBIn7[27] , \wBIn7[26] , \wBIn7[25] , \wBIn7[24] , \wBIn7[23] , 
        \wBIn7[22] , \wBIn7[21] , \wBIn7[20] , \wBIn7[19] , \wBIn7[18] , 
        \wBIn7[17] , \wBIn7[16] , \wBIn7[15] , \wBIn7[14] , \wBIn7[13] , 
        \wBIn7[12] , \wBIn7[11] , \wBIn7[10] , \wBIn7[9] , \wBIn7[8] , 
        \wBIn7[7] , \wBIn7[6] , \wBIn7[5] , \wBIn7[4] , \wBIn7[3] , \wBIn7[2] , 
        \wBIn7[1] , \wBIn7[0] }), .HiOut({\wBMid6[31] , \wBMid6[30] , 
        \wBMid6[29] , \wBMid6[28] , \wBMid6[27] , \wBMid6[26] , \wBMid6[25] , 
        \wBMid6[24] , \wBMid6[23] , \wBMid6[22] , \wBMid6[21] , \wBMid6[20] , 
        \wBMid6[19] , \wBMid6[18] , \wBMid6[17] , \wBMid6[16] , \wBMid6[15] , 
        \wBMid6[14] , \wBMid6[13] , \wBMid6[12] , \wBMid6[11] , \wBMid6[10] , 
        \wBMid6[9] , \wBMid6[8] , \wBMid6[7] , \wBMid6[6] , \wBMid6[5] , 
        \wBMid6[4] , \wBMid6[3] , \wBMid6[2] , \wBMid6[1] , \wBMid6[0] }), 
        .LoOut({\wAMid7[31] , \wAMid7[30] , \wAMid7[29] , \wAMid7[28] , 
        \wAMid7[27] , \wAMid7[26] , \wAMid7[25] , \wAMid7[24] , \wAMid7[23] , 
        \wAMid7[22] , \wAMid7[21] , \wAMid7[20] , \wAMid7[19] , \wAMid7[18] , 
        \wAMid7[17] , \wAMid7[16] , \wAMid7[15] , \wAMid7[14] , \wAMid7[13] , 
        \wAMid7[12] , \wAMid7[11] , \wAMid7[10] , \wAMid7[9] , \wAMid7[8] , 
        \wAMid7[7] , \wAMid7[6] , \wAMid7[5] , \wAMid7[4] , \wAMid7[3] , 
        \wAMid7[2] , \wAMid7[1] , \wAMid7[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn26[31] , \wAIn26[30] , \wAIn26[29] , \wAIn26[28] , \wAIn26[27] , 
        \wAIn26[26] , \wAIn26[25] , \wAIn26[24] , \wAIn26[23] , \wAIn26[22] , 
        \wAIn26[21] , \wAIn26[20] , \wAIn26[19] , \wAIn26[18] , \wAIn26[17] , 
        \wAIn26[16] , \wAIn26[15] , \wAIn26[14] , \wAIn26[13] , \wAIn26[12] , 
        \wAIn26[11] , \wAIn26[10] , \wAIn26[9] , \wAIn26[8] , \wAIn26[7] , 
        \wAIn26[6] , \wAIn26[5] , \wAIn26[4] , \wAIn26[3] , \wAIn26[2] , 
        \wAIn26[1] , \wAIn26[0] }), .BIn({\wBIn26[31] , \wBIn26[30] , 
        \wBIn26[29] , \wBIn26[28] , \wBIn26[27] , \wBIn26[26] , \wBIn26[25] , 
        \wBIn26[24] , \wBIn26[23] , \wBIn26[22] , \wBIn26[21] , \wBIn26[20] , 
        \wBIn26[19] , \wBIn26[18] , \wBIn26[17] , \wBIn26[16] , \wBIn26[15] , 
        \wBIn26[14] , \wBIn26[13] , \wBIn26[12] , \wBIn26[11] , \wBIn26[10] , 
        \wBIn26[9] , \wBIn26[8] , \wBIn26[7] , \wBIn26[6] , \wBIn26[5] , 
        \wBIn26[4] , \wBIn26[3] , \wBIn26[2] , \wBIn26[1] , \wBIn26[0] }), 
        .HiOut({\wBMid25[31] , \wBMid25[30] , \wBMid25[29] , \wBMid25[28] , 
        \wBMid25[27] , \wBMid25[26] , \wBMid25[25] , \wBMid25[24] , 
        \wBMid25[23] , \wBMid25[22] , \wBMid25[21] , \wBMid25[20] , 
        \wBMid25[19] , \wBMid25[18] , \wBMid25[17] , \wBMid25[16] , 
        \wBMid25[15] , \wBMid25[14] , \wBMid25[13] , \wBMid25[12] , 
        \wBMid25[11] , \wBMid25[10] , \wBMid25[9] , \wBMid25[8] , \wBMid25[7] , 
        \wBMid25[6] , \wBMid25[5] , \wBMid25[4] , \wBMid25[3] , \wBMid25[2] , 
        \wBMid25[1] , \wBMid25[0] }), .LoOut({\wAMid26[31] , \wAMid26[30] , 
        \wAMid26[29] , \wAMid26[28] , \wAMid26[27] , \wAMid26[26] , 
        \wAMid26[25] , \wAMid26[24] , \wAMid26[23] , \wAMid26[22] , 
        \wAMid26[21] , \wAMid26[20] , \wAMid26[19] , \wAMid26[18] , 
        \wAMid26[17] , \wAMid26[16] , \wAMid26[15] , \wAMid26[14] , 
        \wAMid26[13] , \wAMid26[12] , \wAMid26[11] , \wAMid26[10] , 
        \wAMid26[9] , \wAMid26[8] , \wAMid26[7] , \wAMid26[6] , \wAMid26[5] , 
        \wAMid26[4] , \wAMid26[3] , \wAMid26[2] , \wAMid26[1] , \wAMid26[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn48[31] , \wAIn48[30] , \wAIn48[29] , \wAIn48[28] , \wAIn48[27] , 
        \wAIn48[26] , \wAIn48[25] , \wAIn48[24] , \wAIn48[23] , \wAIn48[22] , 
        \wAIn48[21] , \wAIn48[20] , \wAIn48[19] , \wAIn48[18] , \wAIn48[17] , 
        \wAIn48[16] , \wAIn48[15] , \wAIn48[14] , \wAIn48[13] , \wAIn48[12] , 
        \wAIn48[11] , \wAIn48[10] , \wAIn48[9] , \wAIn48[8] , \wAIn48[7] , 
        \wAIn48[6] , \wAIn48[5] , \wAIn48[4] , \wAIn48[3] , \wAIn48[2] , 
        \wAIn48[1] , \wAIn48[0] }), .BIn({\wBIn48[31] , \wBIn48[30] , 
        \wBIn48[29] , \wBIn48[28] , \wBIn48[27] , \wBIn48[26] , \wBIn48[25] , 
        \wBIn48[24] , \wBIn48[23] , \wBIn48[22] , \wBIn48[21] , \wBIn48[20] , 
        \wBIn48[19] , \wBIn48[18] , \wBIn48[17] , \wBIn48[16] , \wBIn48[15] , 
        \wBIn48[14] , \wBIn48[13] , \wBIn48[12] , \wBIn48[11] , \wBIn48[10] , 
        \wBIn48[9] , \wBIn48[8] , \wBIn48[7] , \wBIn48[6] , \wBIn48[5] , 
        \wBIn48[4] , \wBIn48[3] , \wBIn48[2] , \wBIn48[1] , \wBIn48[0] }), 
        .HiOut({\wBMid47[31] , \wBMid47[30] , \wBMid47[29] , \wBMid47[28] , 
        \wBMid47[27] , \wBMid47[26] , \wBMid47[25] , \wBMid47[24] , 
        \wBMid47[23] , \wBMid47[22] , \wBMid47[21] , \wBMid47[20] , 
        \wBMid47[19] , \wBMid47[18] , \wBMid47[17] , \wBMid47[16] , 
        \wBMid47[15] , \wBMid47[14] , \wBMid47[13] , \wBMid47[12] , 
        \wBMid47[11] , \wBMid47[10] , \wBMid47[9] , \wBMid47[8] , \wBMid47[7] , 
        \wBMid47[6] , \wBMid47[5] , \wBMid47[4] , \wBMid47[3] , \wBMid47[2] , 
        \wBMid47[1] , \wBMid47[0] }), .LoOut({\wAMid48[31] , \wAMid48[30] , 
        \wAMid48[29] , \wAMid48[28] , \wAMid48[27] , \wAMid48[26] , 
        \wAMid48[25] , \wAMid48[24] , \wAMid48[23] , \wAMid48[22] , 
        \wAMid48[21] , \wAMid48[20] , \wAMid48[19] , \wAMid48[18] , 
        \wAMid48[17] , \wAMid48[16] , \wAMid48[15] , \wAMid48[14] , 
        \wAMid48[13] , \wAMid48[12] , \wAMid48[11] , \wAMid48[10] , 
        \wAMid48[9] , \wAMid48[8] , \wAMid48[7] , \wAMid48[6] , \wAMid48[5] , 
        \wAMid48[4] , \wAMid48[3] , \wAMid48[2] , \wAMid48[1] , \wAMid48[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn53[31] , \wAIn53[30] , \wAIn53[29] , \wAIn53[28] , \wAIn53[27] , 
        \wAIn53[26] , \wAIn53[25] , \wAIn53[24] , \wAIn53[23] , \wAIn53[22] , 
        \wAIn53[21] , \wAIn53[20] , \wAIn53[19] , \wAIn53[18] , \wAIn53[17] , 
        \wAIn53[16] , \wAIn53[15] , \wAIn53[14] , \wAIn53[13] , \wAIn53[12] , 
        \wAIn53[11] , \wAIn53[10] , \wAIn53[9] , \wAIn53[8] , \wAIn53[7] , 
        \wAIn53[6] , \wAIn53[5] , \wAIn53[4] , \wAIn53[3] , \wAIn53[2] , 
        \wAIn53[1] , \wAIn53[0] }), .BIn({\wBIn53[31] , \wBIn53[30] , 
        \wBIn53[29] , \wBIn53[28] , \wBIn53[27] , \wBIn53[26] , \wBIn53[25] , 
        \wBIn53[24] , \wBIn53[23] , \wBIn53[22] , \wBIn53[21] , \wBIn53[20] , 
        \wBIn53[19] , \wBIn53[18] , \wBIn53[17] , \wBIn53[16] , \wBIn53[15] , 
        \wBIn53[14] , \wBIn53[13] , \wBIn53[12] , \wBIn53[11] , \wBIn53[10] , 
        \wBIn53[9] , \wBIn53[8] , \wBIn53[7] , \wBIn53[6] , \wBIn53[5] , 
        \wBIn53[4] , \wBIn53[3] , \wBIn53[2] , \wBIn53[1] , \wBIn53[0] }), 
        .HiOut({\wBMid52[31] , \wBMid52[30] , \wBMid52[29] , \wBMid52[28] , 
        \wBMid52[27] , \wBMid52[26] , \wBMid52[25] , \wBMid52[24] , 
        \wBMid52[23] , \wBMid52[22] , \wBMid52[21] , \wBMid52[20] , 
        \wBMid52[19] , \wBMid52[18] , \wBMid52[17] , \wBMid52[16] , 
        \wBMid52[15] , \wBMid52[14] , \wBMid52[13] , \wBMid52[12] , 
        \wBMid52[11] , \wBMid52[10] , \wBMid52[9] , \wBMid52[8] , \wBMid52[7] , 
        \wBMid52[6] , \wBMid52[5] , \wBMid52[4] , \wBMid52[3] , \wBMid52[2] , 
        \wBMid52[1] , \wBMid52[0] }), .LoOut({\wAMid53[31] , \wAMid53[30] , 
        \wAMid53[29] , \wAMid53[28] , \wAMid53[27] , \wAMid53[26] , 
        \wAMid53[25] , \wAMid53[24] , \wAMid53[23] , \wAMid53[22] , 
        \wAMid53[21] , \wAMid53[20] , \wAMid53[19] , \wAMid53[18] , 
        \wAMid53[17] , \wAMid53[16] , \wAMid53[15] , \wAMid53[14] , 
        \wAMid53[13] , \wAMid53[12] , \wAMid53[11] , \wAMid53[10] , 
        \wAMid53[9] , \wAMid53[8] , \wAMid53[7] , \wAMid53[6] , \wAMid53[5] , 
        \wAMid53[4] , \wAMid53[3] , \wAMid53[2] , \wAMid53[1] , \wAMid53[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn91[31] , \wAIn91[30] , \wAIn91[29] , \wAIn91[28] , \wAIn91[27] , 
        \wAIn91[26] , \wAIn91[25] , \wAIn91[24] , \wAIn91[23] , \wAIn91[22] , 
        \wAIn91[21] , \wAIn91[20] , \wAIn91[19] , \wAIn91[18] , \wAIn91[17] , 
        \wAIn91[16] , \wAIn91[15] , \wAIn91[14] , \wAIn91[13] , \wAIn91[12] , 
        \wAIn91[11] , \wAIn91[10] , \wAIn91[9] , \wAIn91[8] , \wAIn91[7] , 
        \wAIn91[6] , \wAIn91[5] , \wAIn91[4] , \wAIn91[3] , \wAIn91[2] , 
        \wAIn91[1] , \wAIn91[0] }), .BIn({\wBIn91[31] , \wBIn91[30] , 
        \wBIn91[29] , \wBIn91[28] , \wBIn91[27] , \wBIn91[26] , \wBIn91[25] , 
        \wBIn91[24] , \wBIn91[23] , \wBIn91[22] , \wBIn91[21] , \wBIn91[20] , 
        \wBIn91[19] , \wBIn91[18] , \wBIn91[17] , \wBIn91[16] , \wBIn91[15] , 
        \wBIn91[14] , \wBIn91[13] , \wBIn91[12] , \wBIn91[11] , \wBIn91[10] , 
        \wBIn91[9] , \wBIn91[8] , \wBIn91[7] , \wBIn91[6] , \wBIn91[5] , 
        \wBIn91[4] , \wBIn91[3] , \wBIn91[2] , \wBIn91[1] , \wBIn91[0] }), 
        .HiOut({\wBMid90[31] , \wBMid90[30] , \wBMid90[29] , \wBMid90[28] , 
        \wBMid90[27] , \wBMid90[26] , \wBMid90[25] , \wBMid90[24] , 
        \wBMid90[23] , \wBMid90[22] , \wBMid90[21] , \wBMid90[20] , 
        \wBMid90[19] , \wBMid90[18] , \wBMid90[17] , \wBMid90[16] , 
        \wBMid90[15] , \wBMid90[14] , \wBMid90[13] , \wBMid90[12] , 
        \wBMid90[11] , \wBMid90[10] , \wBMid90[9] , \wBMid90[8] , \wBMid90[7] , 
        \wBMid90[6] , \wBMid90[5] , \wBMid90[4] , \wBMid90[3] , \wBMid90[2] , 
        \wBMid90[1] , \wBMid90[0] }), .LoOut({\wAMid91[31] , \wAMid91[30] , 
        \wAMid91[29] , \wAMid91[28] , \wAMid91[27] , \wAMid91[26] , 
        \wAMid91[25] , \wAMid91[24] , \wAMid91[23] , \wAMid91[22] , 
        \wAMid91[21] , \wAMid91[20] , \wAMid91[19] , \wAMid91[18] , 
        \wAMid91[17] , \wAMid91[16] , \wAMid91[15] , \wAMid91[14] , 
        \wAMid91[13] , \wAMid91[12] , \wAMid91[11] , \wAMid91[10] , 
        \wAMid91[9] , \wAMid91[8] , \wAMid91[7] , \wAMid91[6] , \wAMid91[5] , 
        \wAMid91[4] , \wAMid91[3] , \wAMid91[2] , \wAMid91[1] , \wAMid91[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid0[31] , 
        \wAMid0[30] , \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , 
        \wAMid0[25] , \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , 
        \wAMid0[20] , \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , 
        \wAMid0[15] , \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , 
        \wAMid0[10] , \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , 
        \wAMid0[5] , \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , 
        \wAMid0[0] }), .BIn({\wBMid0[31] , \wBMid0[30] , \wBMid0[29] , 
        \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , \wBMid0[24] , 
        \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , \wBMid0[19] , 
        \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , \wBMid0[14] , 
        \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , \wBMid0[9] , 
        \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , \wBMid0[4] , 
        \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), .HiOut({
        \wRegInB0[31] , \wRegInB0[30] , \wRegInB0[29] , \wRegInB0[28] , 
        \wRegInB0[27] , \wRegInB0[26] , \wRegInB0[25] , \wRegInB0[24] , 
        \wRegInB0[23] , \wRegInB0[22] , \wRegInB0[21] , \wRegInB0[20] , 
        \wRegInB0[19] , \wRegInB0[18] , \wRegInB0[17] , \wRegInB0[16] , 
        \wRegInB0[15] , \wRegInB0[14] , \wRegInB0[13] , \wRegInB0[12] , 
        \wRegInB0[11] , \wRegInB0[10] , \wRegInB0[9] , \wRegInB0[8] , 
        \wRegInB0[7] , \wRegInB0[6] , \wRegInB0[5] , \wRegInB0[4] , 
        \wRegInB0[3] , \wRegInB0[2] , \wRegInB0[1] , \wRegInB0[0] }), .LoOut({
        \wRegInA1[31] , \wRegInA1[30] , \wRegInA1[29] , \wRegInA1[28] , 
        \wRegInA1[27] , \wRegInA1[26] , \wRegInA1[25] , \wRegInA1[24] , 
        \wRegInA1[23] , \wRegInA1[22] , \wRegInA1[21] , \wRegInA1[20] , 
        \wRegInA1[19] , \wRegInA1[18] , \wRegInA1[17] , \wRegInA1[16] , 
        \wRegInA1[15] , \wRegInA1[14] , \wRegInA1[13] , \wRegInA1[12] , 
        \wRegInA1[11] , \wRegInA1[10] , \wRegInA1[9] , \wRegInA1[8] , 
        \wRegInA1[7] , \wRegInA1[6] , \wRegInA1[5] , \wRegInA1[4] , 
        \wRegInA1[3] , \wRegInA1[2] , \wRegInA1[1] , \wRegInA1[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_194 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink195[31] , \ScanLink195[30] , \ScanLink195[29] , 
        \ScanLink195[28] , \ScanLink195[27] , \ScanLink195[26] , 
        \ScanLink195[25] , \ScanLink195[24] , \ScanLink195[23] , 
        \ScanLink195[22] , \ScanLink195[21] , \ScanLink195[20] , 
        \ScanLink195[19] , \ScanLink195[18] , \ScanLink195[17] , 
        \ScanLink195[16] , \ScanLink195[15] , \ScanLink195[14] , 
        \ScanLink195[13] , \ScanLink195[12] , \ScanLink195[11] , 
        \ScanLink195[10] , \ScanLink195[9] , \ScanLink195[8] , 
        \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , \ScanLink195[4] , 
        \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , \ScanLink195[0] 
        }), .ScanOut({\ScanLink194[31] , \ScanLink194[30] , \ScanLink194[29] , 
        \ScanLink194[28] , \ScanLink194[27] , \ScanLink194[26] , 
        \ScanLink194[25] , \ScanLink194[24] , \ScanLink194[23] , 
        \ScanLink194[22] , \ScanLink194[21] , \ScanLink194[20] , 
        \ScanLink194[19] , \ScanLink194[18] , \ScanLink194[17] , 
        \ScanLink194[16] , \ScanLink194[15] , \ScanLink194[14] , 
        \ScanLink194[13] , \ScanLink194[12] , \ScanLink194[11] , 
        \ScanLink194[10] , \ScanLink194[9] , \ScanLink194[8] , 
        \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , \ScanLink194[4] , 
        \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , \ScanLink194[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB30[31] , \wRegInB30[30] , \wRegInB30[29] , 
        \wRegInB30[28] , \wRegInB30[27] , \wRegInB30[26] , \wRegInB30[25] , 
        \wRegInB30[24] , \wRegInB30[23] , \wRegInB30[22] , \wRegInB30[21] , 
        \wRegInB30[20] , \wRegInB30[19] , \wRegInB30[18] , \wRegInB30[17] , 
        \wRegInB30[16] , \wRegInB30[15] , \wRegInB30[14] , \wRegInB30[13] , 
        \wRegInB30[12] , \wRegInB30[11] , \wRegInB30[10] , \wRegInB30[9] , 
        \wRegInB30[8] , \wRegInB30[7] , \wRegInB30[6] , \wRegInB30[5] , 
        \wRegInB30[4] , \wRegInB30[3] , \wRegInB30[2] , \wRegInB30[1] , 
        \wRegInB30[0] }), .Out({\wBIn30[31] , \wBIn30[30] , \wBIn30[29] , 
        \wBIn30[28] , \wBIn30[27] , \wBIn30[26] , \wBIn30[25] , \wBIn30[24] , 
        \wBIn30[23] , \wBIn30[22] , \wBIn30[21] , \wBIn30[20] , \wBIn30[19] , 
        \wBIn30[18] , \wBIn30[17] , \wBIn30[16] , \wBIn30[15] , \wBIn30[14] , 
        \wBIn30[13] , \wBIn30[12] , \wBIn30[11] , \wBIn30[10] , \wBIn30[9] , 
        \wBIn30[8] , \wBIn30[7] , \wBIn30[6] , \wBIn30[5] , \wBIn30[4] , 
        \wBIn30[3] , \wBIn30[2] , \wBIn30[1] , \wBIn30[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid86[31] , \wAMid86[30] , \wAMid86[29] , \wAMid86[28] , 
        \wAMid86[27] , \wAMid86[26] , \wAMid86[25] , \wAMid86[24] , 
        \wAMid86[23] , \wAMid86[22] , \wAMid86[21] , \wAMid86[20] , 
        \wAMid86[19] , \wAMid86[18] , \wAMid86[17] , \wAMid86[16] , 
        \wAMid86[15] , \wAMid86[14] , \wAMid86[13] , \wAMid86[12] , 
        \wAMid86[11] , \wAMid86[10] , \wAMid86[9] , \wAMid86[8] , \wAMid86[7] , 
        \wAMid86[6] , \wAMid86[5] , \wAMid86[4] , \wAMid86[3] , \wAMid86[2] , 
        \wAMid86[1] , \wAMid86[0] }), .BIn({\wBMid86[31] , \wBMid86[30] , 
        \wBMid86[29] , \wBMid86[28] , \wBMid86[27] , \wBMid86[26] , 
        \wBMid86[25] , \wBMid86[24] , \wBMid86[23] , \wBMid86[22] , 
        \wBMid86[21] , \wBMid86[20] , \wBMid86[19] , \wBMid86[18] , 
        \wBMid86[17] , \wBMid86[16] , \wBMid86[15] , \wBMid86[14] , 
        \wBMid86[13] , \wBMid86[12] , \wBMid86[11] , \wBMid86[10] , 
        \wBMid86[9] , \wBMid86[8] , \wBMid86[7] , \wBMid86[6] , \wBMid86[5] , 
        \wBMid86[4] , \wBMid86[3] , \wBMid86[2] , \wBMid86[1] , \wBMid86[0] }), 
        .HiOut({\wRegInB86[31] , \wRegInB86[30] , \wRegInB86[29] , 
        \wRegInB86[28] , \wRegInB86[27] , \wRegInB86[26] , \wRegInB86[25] , 
        \wRegInB86[24] , \wRegInB86[23] , \wRegInB86[22] , \wRegInB86[21] , 
        \wRegInB86[20] , \wRegInB86[19] , \wRegInB86[18] , \wRegInB86[17] , 
        \wRegInB86[16] , \wRegInB86[15] , \wRegInB86[14] , \wRegInB86[13] , 
        \wRegInB86[12] , \wRegInB86[11] , \wRegInB86[10] , \wRegInB86[9] , 
        \wRegInB86[8] , \wRegInB86[7] , \wRegInB86[6] , \wRegInB86[5] , 
        \wRegInB86[4] , \wRegInB86[3] , \wRegInB86[2] , \wRegInB86[1] , 
        \wRegInB86[0] }), .LoOut({\wRegInA87[31] , \wRegInA87[30] , 
        \wRegInA87[29] , \wRegInA87[28] , \wRegInA87[27] , \wRegInA87[26] , 
        \wRegInA87[25] , \wRegInA87[24] , \wRegInA87[23] , \wRegInA87[22] , 
        \wRegInA87[21] , \wRegInA87[20] , \wRegInA87[19] , \wRegInA87[18] , 
        \wRegInA87[17] , \wRegInA87[16] , \wRegInA87[15] , \wRegInA87[14] , 
        \wRegInA87[13] , \wRegInA87[12] , \wRegInA87[11] , \wRegInA87[10] , 
        \wRegInA87[9] , \wRegInA87[8] , \wRegInA87[7] , \wRegInA87[6] , 
        \wRegInA87[5] , \wRegInA87[4] , \wRegInA87[3] , \wRegInA87[2] , 
        \wRegInA87[1] , \wRegInA87[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_208 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink209[31] , \ScanLink209[30] , \ScanLink209[29] , 
        \ScanLink209[28] , \ScanLink209[27] , \ScanLink209[26] , 
        \ScanLink209[25] , \ScanLink209[24] , \ScanLink209[23] , 
        \ScanLink209[22] , \ScanLink209[21] , \ScanLink209[20] , 
        \ScanLink209[19] , \ScanLink209[18] , \ScanLink209[17] , 
        \ScanLink209[16] , \ScanLink209[15] , \ScanLink209[14] , 
        \ScanLink209[13] , \ScanLink209[12] , \ScanLink209[11] , 
        \ScanLink209[10] , \ScanLink209[9] , \ScanLink209[8] , 
        \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , \ScanLink209[4] , 
        \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , \ScanLink209[0] 
        }), .ScanOut({\ScanLink208[31] , \ScanLink208[30] , \ScanLink208[29] , 
        \ScanLink208[28] , \ScanLink208[27] , \ScanLink208[26] , 
        \ScanLink208[25] , \ScanLink208[24] , \ScanLink208[23] , 
        \ScanLink208[22] , \ScanLink208[21] , \ScanLink208[20] , 
        \ScanLink208[19] , \ScanLink208[18] , \ScanLink208[17] , 
        \ScanLink208[16] , \ScanLink208[15] , \ScanLink208[14] , 
        \ScanLink208[13] , \ScanLink208[12] , \ScanLink208[11] , 
        \ScanLink208[10] , \ScanLink208[9] , \ScanLink208[8] , 
        \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , \ScanLink208[4] , 
        \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , \ScanLink208[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB23[31] , \wRegInB23[30] , \wRegInB23[29] , 
        \wRegInB23[28] , \wRegInB23[27] , \wRegInB23[26] , \wRegInB23[25] , 
        \wRegInB23[24] , \wRegInB23[23] , \wRegInB23[22] , \wRegInB23[21] , 
        \wRegInB23[20] , \wRegInB23[19] , \wRegInB23[18] , \wRegInB23[17] , 
        \wRegInB23[16] , \wRegInB23[15] , \wRegInB23[14] , \wRegInB23[13] , 
        \wRegInB23[12] , \wRegInB23[11] , \wRegInB23[10] , \wRegInB23[9] , 
        \wRegInB23[8] , \wRegInB23[7] , \wRegInB23[6] , \wRegInB23[5] , 
        \wRegInB23[4] , \wRegInB23[3] , \wRegInB23[2] , \wRegInB23[1] , 
        \wRegInB23[0] }), .Out({\wBIn23[31] , \wBIn23[30] , \wBIn23[29] , 
        \wBIn23[28] , \wBIn23[27] , \wBIn23[26] , \wBIn23[25] , \wBIn23[24] , 
        \wBIn23[23] , \wBIn23[22] , \wBIn23[21] , \wBIn23[20] , \wBIn23[19] , 
        \wBIn23[18] , \wBIn23[17] , \wBIn23[16] , \wBIn23[15] , \wBIn23[14] , 
        \wBIn23[13] , \wBIn23[12] , \wBIn23[11] , \wBIn23[10] , \wBIn23[9] , 
        \wBIn23[8] , \wBIn23[7] , \wBIn23[6] , \wBIn23[5] , \wBIn23[4] , 
        \wBIn23[3] , \wBIn23[2] , \wBIn23[1] , \wBIn23[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_138 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink139[31] , \ScanLink139[30] , \ScanLink139[29] , 
        \ScanLink139[28] , \ScanLink139[27] , \ScanLink139[26] , 
        \ScanLink139[25] , \ScanLink139[24] , \ScanLink139[23] , 
        \ScanLink139[22] , \ScanLink139[21] , \ScanLink139[20] , 
        \ScanLink139[19] , \ScanLink139[18] , \ScanLink139[17] , 
        \ScanLink139[16] , \ScanLink139[15] , \ScanLink139[14] , 
        \ScanLink139[13] , \ScanLink139[12] , \ScanLink139[11] , 
        \ScanLink139[10] , \ScanLink139[9] , \ScanLink139[8] , 
        \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , \ScanLink139[4] , 
        \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , \ScanLink139[0] 
        }), .ScanOut({\ScanLink138[31] , \ScanLink138[30] , \ScanLink138[29] , 
        \ScanLink138[28] , \ScanLink138[27] , \ScanLink138[26] , 
        \ScanLink138[25] , \ScanLink138[24] , \ScanLink138[23] , 
        \ScanLink138[22] , \ScanLink138[21] , \ScanLink138[20] , 
        \ScanLink138[19] , \ScanLink138[18] , \ScanLink138[17] , 
        \ScanLink138[16] , \ScanLink138[15] , \ScanLink138[14] , 
        \ScanLink138[13] , \ScanLink138[12] , \ScanLink138[11] , 
        \ScanLink138[10] , \ScanLink138[9] , \ScanLink138[8] , 
        \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , \ScanLink138[4] , 
        \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , \ScanLink138[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB58[31] , \wRegInB58[30] , \wRegInB58[29] , 
        \wRegInB58[28] , \wRegInB58[27] , \wRegInB58[26] , \wRegInB58[25] , 
        \wRegInB58[24] , \wRegInB58[23] , \wRegInB58[22] , \wRegInB58[21] , 
        \wRegInB58[20] , \wRegInB58[19] , \wRegInB58[18] , \wRegInB58[17] , 
        \wRegInB58[16] , \wRegInB58[15] , \wRegInB58[14] , \wRegInB58[13] , 
        \wRegInB58[12] , \wRegInB58[11] , \wRegInB58[10] , \wRegInB58[9] , 
        \wRegInB58[8] , \wRegInB58[7] , \wRegInB58[6] , \wRegInB58[5] , 
        \wRegInB58[4] , \wRegInB58[3] , \wRegInB58[2] , \wRegInB58[1] , 
        \wRegInB58[0] }), .Out({\wBIn58[31] , \wBIn58[30] , \wBIn58[29] , 
        \wBIn58[28] , \wBIn58[27] , \wBIn58[26] , \wBIn58[25] , \wBIn58[24] , 
        \wBIn58[23] , \wBIn58[22] , \wBIn58[21] , \wBIn58[20] , \wBIn58[19] , 
        \wBIn58[18] , \wBIn58[17] , \wBIn58[16] , \wBIn58[15] , \wBIn58[14] , 
        \wBIn58[13] , \wBIn58[12] , \wBIn58[11] , \wBIn58[10] , \wBIn58[9] , 
        \wBIn58[8] , \wBIn58[7] , \wBIn58[6] , \wBIn58[5] , \wBIn58[4] , 
        \wBIn58[3] , \wBIn58[2] , \wBIn58[1] , \wBIn58[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_68 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink69[31] , \ScanLink69[30] , \ScanLink69[29] , 
        \ScanLink69[28] , \ScanLink69[27] , \ScanLink69[26] , \ScanLink69[25] , 
        \ScanLink69[24] , \ScanLink69[23] , \ScanLink69[22] , \ScanLink69[21] , 
        \ScanLink69[20] , \ScanLink69[19] , \ScanLink69[18] , \ScanLink69[17] , 
        \ScanLink69[16] , \ScanLink69[15] , \ScanLink69[14] , \ScanLink69[13] , 
        \ScanLink69[12] , \ScanLink69[11] , \ScanLink69[10] , \ScanLink69[9] , 
        \ScanLink69[8] , \ScanLink69[7] , \ScanLink69[6] , \ScanLink69[5] , 
        \ScanLink69[4] , \ScanLink69[3] , \ScanLink69[2] , \ScanLink69[1] , 
        \ScanLink69[0] }), .ScanOut({\ScanLink68[31] , \ScanLink68[30] , 
        \ScanLink68[29] , \ScanLink68[28] , \ScanLink68[27] , \ScanLink68[26] , 
        \ScanLink68[25] , \ScanLink68[24] , \ScanLink68[23] , \ScanLink68[22] , 
        \ScanLink68[21] , \ScanLink68[20] , \ScanLink68[19] , \ScanLink68[18] , 
        \ScanLink68[17] , \ScanLink68[16] , \ScanLink68[15] , \ScanLink68[14] , 
        \ScanLink68[13] , \ScanLink68[12] , \ScanLink68[11] , \ScanLink68[10] , 
        \ScanLink68[9] , \ScanLink68[8] , \ScanLink68[7] , \ScanLink68[6] , 
        \ScanLink68[5] , \ScanLink68[4] , \ScanLink68[3] , \ScanLink68[2] , 
        \ScanLink68[1] , \ScanLink68[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB93[31] , \wRegInB93[30] , 
        \wRegInB93[29] , \wRegInB93[28] , \wRegInB93[27] , \wRegInB93[26] , 
        \wRegInB93[25] , \wRegInB93[24] , \wRegInB93[23] , \wRegInB93[22] , 
        \wRegInB93[21] , \wRegInB93[20] , \wRegInB93[19] , \wRegInB93[18] , 
        \wRegInB93[17] , \wRegInB93[16] , \wRegInB93[15] , \wRegInB93[14] , 
        \wRegInB93[13] , \wRegInB93[12] , \wRegInB93[11] , \wRegInB93[10] , 
        \wRegInB93[9] , \wRegInB93[8] , \wRegInB93[7] , \wRegInB93[6] , 
        \wRegInB93[5] , \wRegInB93[4] , \wRegInB93[3] , \wRegInB93[2] , 
        \wRegInB93[1] , \wRegInB93[0] }), .Out({\wBIn93[31] , \wBIn93[30] , 
        \wBIn93[29] , \wBIn93[28] , \wBIn93[27] , \wBIn93[26] , \wBIn93[25] , 
        \wBIn93[24] , \wBIn93[23] , \wBIn93[22] , \wBIn93[21] , \wBIn93[20] , 
        \wBIn93[19] , \wBIn93[18] , \wBIn93[17] , \wBIn93[16] , \wBIn93[15] , 
        \wBIn93[14] , \wBIn93[13] , \wBIn93[12] , \wBIn93[11] , \wBIn93[10] , 
        \wBIn93[9] , \wBIn93[8] , \wBIn93[7] , \wBIn93[6] , \wBIn93[5] , 
        \wBIn93[4] , \wBIn93[3] , \wBIn93[2] , \wBIn93[1] , \wBIn93[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn74[31] , \wAIn74[30] , \wAIn74[29] , \wAIn74[28] , \wAIn74[27] , 
        \wAIn74[26] , \wAIn74[25] , \wAIn74[24] , \wAIn74[23] , \wAIn74[22] , 
        \wAIn74[21] , \wAIn74[20] , \wAIn74[19] , \wAIn74[18] , \wAIn74[17] , 
        \wAIn74[16] , \wAIn74[15] , \wAIn74[14] , \wAIn74[13] , \wAIn74[12] , 
        \wAIn74[11] , \wAIn74[10] , \wAIn74[9] , \wAIn74[8] , \wAIn74[7] , 
        \wAIn74[6] , \wAIn74[5] , \wAIn74[4] , \wAIn74[3] , \wAIn74[2] , 
        \wAIn74[1] , \wAIn74[0] }), .BIn({\wBIn74[31] , \wBIn74[30] , 
        \wBIn74[29] , \wBIn74[28] , \wBIn74[27] , \wBIn74[26] , \wBIn74[25] , 
        \wBIn74[24] , \wBIn74[23] , \wBIn74[22] , \wBIn74[21] , \wBIn74[20] , 
        \wBIn74[19] , \wBIn74[18] , \wBIn74[17] , \wBIn74[16] , \wBIn74[15] , 
        \wBIn74[14] , \wBIn74[13] , \wBIn74[12] , \wBIn74[11] , \wBIn74[10] , 
        \wBIn74[9] , \wBIn74[8] , \wBIn74[7] , \wBIn74[6] , \wBIn74[5] , 
        \wBIn74[4] , \wBIn74[3] , \wBIn74[2] , \wBIn74[1] , \wBIn74[0] }), 
        .HiOut({\wBMid73[31] , \wBMid73[30] , \wBMid73[29] , \wBMid73[28] , 
        \wBMid73[27] , \wBMid73[26] , \wBMid73[25] , \wBMid73[24] , 
        \wBMid73[23] , \wBMid73[22] , \wBMid73[21] , \wBMid73[20] , 
        \wBMid73[19] , \wBMid73[18] , \wBMid73[17] , \wBMid73[16] , 
        \wBMid73[15] , \wBMid73[14] , \wBMid73[13] , \wBMid73[12] , 
        \wBMid73[11] , \wBMid73[10] , \wBMid73[9] , \wBMid73[8] , \wBMid73[7] , 
        \wBMid73[6] , \wBMid73[5] , \wBMid73[4] , \wBMid73[3] , \wBMid73[2] , 
        \wBMid73[1] , \wBMid73[0] }), .LoOut({\wAMid74[31] , \wAMid74[30] , 
        \wAMid74[29] , \wAMid74[28] , \wAMid74[27] , \wAMid74[26] , 
        \wAMid74[25] , \wAMid74[24] , \wAMid74[23] , \wAMid74[22] , 
        \wAMid74[21] , \wAMid74[20] , \wAMid74[19] , \wAMid74[18] , 
        \wAMid74[17] , \wAMid74[16] , \wAMid74[15] , \wAMid74[14] , 
        \wAMid74[13] , \wAMid74[12] , \wAMid74[11] , \wAMid74[10] , 
        \wAMid74[9] , \wAMid74[8] , \wAMid74[7] , \wAMid74[6] , \wAMid74[5] , 
        \wAMid74[4] , \wAMid74[3] , \wAMid74[2] , \wAMid74[1] , \wAMid74[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn104[31] , \wAIn104[30] , \wAIn104[29] , \wAIn104[28] , 
        \wAIn104[27] , \wAIn104[26] , \wAIn104[25] , \wAIn104[24] , 
        \wAIn104[23] , \wAIn104[22] , \wAIn104[21] , \wAIn104[20] , 
        \wAIn104[19] , \wAIn104[18] , \wAIn104[17] , \wAIn104[16] , 
        \wAIn104[15] , \wAIn104[14] , \wAIn104[13] , \wAIn104[12] , 
        \wAIn104[11] , \wAIn104[10] , \wAIn104[9] , \wAIn104[8] , \wAIn104[7] , 
        \wAIn104[6] , \wAIn104[5] , \wAIn104[4] , \wAIn104[3] , \wAIn104[2] , 
        \wAIn104[1] , \wAIn104[0] }), .BIn({\wBIn104[31] , \wBIn104[30] , 
        \wBIn104[29] , \wBIn104[28] , \wBIn104[27] , \wBIn104[26] , 
        \wBIn104[25] , \wBIn104[24] , \wBIn104[23] , \wBIn104[22] , 
        \wBIn104[21] , \wBIn104[20] , \wBIn104[19] , \wBIn104[18] , 
        \wBIn104[17] , \wBIn104[16] , \wBIn104[15] , \wBIn104[14] , 
        \wBIn104[13] , \wBIn104[12] , \wBIn104[11] , \wBIn104[10] , 
        \wBIn104[9] , \wBIn104[8] , \wBIn104[7] , \wBIn104[6] , \wBIn104[5] , 
        \wBIn104[4] , \wBIn104[3] , \wBIn104[2] , \wBIn104[1] , \wBIn104[0] }), 
        .HiOut({\wBMid103[31] , \wBMid103[30] , \wBMid103[29] , \wBMid103[28] , 
        \wBMid103[27] , \wBMid103[26] , \wBMid103[25] , \wBMid103[24] , 
        \wBMid103[23] , \wBMid103[22] , \wBMid103[21] , \wBMid103[20] , 
        \wBMid103[19] , \wBMid103[18] , \wBMid103[17] , \wBMid103[16] , 
        \wBMid103[15] , \wBMid103[14] , \wBMid103[13] , \wBMid103[12] , 
        \wBMid103[11] , \wBMid103[10] , \wBMid103[9] , \wBMid103[8] , 
        \wBMid103[7] , \wBMid103[6] , \wBMid103[5] , \wBMid103[4] , 
        \wBMid103[3] , \wBMid103[2] , \wBMid103[1] , \wBMid103[0] }), .LoOut({
        \wAMid104[31] , \wAMid104[30] , \wAMid104[29] , \wAMid104[28] , 
        \wAMid104[27] , \wAMid104[26] , \wAMid104[25] , \wAMid104[24] , 
        \wAMid104[23] , \wAMid104[22] , \wAMid104[21] , \wAMid104[20] , 
        \wAMid104[19] , \wAMid104[18] , \wAMid104[17] , \wAMid104[16] , 
        \wAMid104[15] , \wAMid104[14] , \wAMid104[13] , \wAMid104[12] , 
        \wAMid104[11] , \wAMid104[10] , \wAMid104[9] , \wAMid104[8] , 
        \wAMid104[7] , \wAMid104[6] , \wAMid104[5] , \wAMid104[4] , 
        \wAMid104[3] , \wAMid104[2] , \wAMid104[1] , \wAMid104[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn123[31] , \wAIn123[30] , \wAIn123[29] , \wAIn123[28] , 
        \wAIn123[27] , \wAIn123[26] , \wAIn123[25] , \wAIn123[24] , 
        \wAIn123[23] , \wAIn123[22] , \wAIn123[21] , \wAIn123[20] , 
        \wAIn123[19] , \wAIn123[18] , \wAIn123[17] , \wAIn123[16] , 
        \wAIn123[15] , \wAIn123[14] , \wAIn123[13] , \wAIn123[12] , 
        \wAIn123[11] , \wAIn123[10] , \wAIn123[9] , \wAIn123[8] , \wAIn123[7] , 
        \wAIn123[6] , \wAIn123[5] , \wAIn123[4] , \wAIn123[3] , \wAIn123[2] , 
        \wAIn123[1] , \wAIn123[0] }), .BIn({\wBIn123[31] , \wBIn123[30] , 
        \wBIn123[29] , \wBIn123[28] , \wBIn123[27] , \wBIn123[26] , 
        \wBIn123[25] , \wBIn123[24] , \wBIn123[23] , \wBIn123[22] , 
        \wBIn123[21] , \wBIn123[20] , \wBIn123[19] , \wBIn123[18] , 
        \wBIn123[17] , \wBIn123[16] , \wBIn123[15] , \wBIn123[14] , 
        \wBIn123[13] , \wBIn123[12] , \wBIn123[11] , \wBIn123[10] , 
        \wBIn123[9] , \wBIn123[8] , \wBIn123[7] , \wBIn123[6] , \wBIn123[5] , 
        \wBIn123[4] , \wBIn123[3] , \wBIn123[2] , \wBIn123[1] , \wBIn123[0] }), 
        .HiOut({\wBMid122[31] , \wBMid122[30] , \wBMid122[29] , \wBMid122[28] , 
        \wBMid122[27] , \wBMid122[26] , \wBMid122[25] , \wBMid122[24] , 
        \wBMid122[23] , \wBMid122[22] , \wBMid122[21] , \wBMid122[20] , 
        \wBMid122[19] , \wBMid122[18] , \wBMid122[17] , \wBMid122[16] , 
        \wBMid122[15] , \wBMid122[14] , \wBMid122[13] , \wBMid122[12] , 
        \wBMid122[11] , \wBMid122[10] , \wBMid122[9] , \wBMid122[8] , 
        \wBMid122[7] , \wBMid122[6] , \wBMid122[5] , \wBMid122[4] , 
        \wBMid122[3] , \wBMid122[2] , \wBMid122[1] , \wBMid122[0] }), .LoOut({
        \wAMid123[31] , \wAMid123[30] , \wAMid123[29] , \wAMid123[28] , 
        \wAMid123[27] , \wAMid123[26] , \wAMid123[25] , \wAMid123[24] , 
        \wAMid123[23] , \wAMid123[22] , \wAMid123[21] , \wAMid123[20] , 
        \wAMid123[19] , \wAMid123[18] , \wAMid123[17] , \wAMid123[16] , 
        \wAMid123[15] , \wAMid123[14] , \wAMid123[13] , \wAMid123[12] , 
        \wAMid123[11] , \wAMid123[10] , \wAMid123[9] , \wAMid123[8] , 
        \wAMid123[7] , \wAMid123[6] , \wAMid123[5] , \wAMid123[4] , 
        \wAMid123[3] , \wAMid123[2] , \wAMid123[1] , \wAMid123[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid63[31] , \wAMid63[30] , \wAMid63[29] , \wAMid63[28] , 
        \wAMid63[27] , \wAMid63[26] , \wAMid63[25] , \wAMid63[24] , 
        \wAMid63[23] , \wAMid63[22] , \wAMid63[21] , \wAMid63[20] , 
        \wAMid63[19] , \wAMid63[18] , \wAMid63[17] , \wAMid63[16] , 
        \wAMid63[15] , \wAMid63[14] , \wAMid63[13] , \wAMid63[12] , 
        \wAMid63[11] , \wAMid63[10] , \wAMid63[9] , \wAMid63[8] , \wAMid63[7] , 
        \wAMid63[6] , \wAMid63[5] , \wAMid63[4] , \wAMid63[3] , \wAMid63[2] , 
        \wAMid63[1] , \wAMid63[0] }), .BIn({\wBMid63[31] , \wBMid63[30] , 
        \wBMid63[29] , \wBMid63[28] , \wBMid63[27] , \wBMid63[26] , 
        \wBMid63[25] , \wBMid63[24] , \wBMid63[23] , \wBMid63[22] , 
        \wBMid63[21] , \wBMid63[20] , \wBMid63[19] , \wBMid63[18] , 
        \wBMid63[17] , \wBMid63[16] , \wBMid63[15] , \wBMid63[14] , 
        \wBMid63[13] , \wBMid63[12] , \wBMid63[11] , \wBMid63[10] , 
        \wBMid63[9] , \wBMid63[8] , \wBMid63[7] , \wBMid63[6] , \wBMid63[5] , 
        \wBMid63[4] , \wBMid63[3] , \wBMid63[2] , \wBMid63[1] , \wBMid63[0] }), 
        .HiOut({\wRegInB63[31] , \wRegInB63[30] , \wRegInB63[29] , 
        \wRegInB63[28] , \wRegInB63[27] , \wRegInB63[26] , \wRegInB63[25] , 
        \wRegInB63[24] , \wRegInB63[23] , \wRegInB63[22] , \wRegInB63[21] , 
        \wRegInB63[20] , \wRegInB63[19] , \wRegInB63[18] , \wRegInB63[17] , 
        \wRegInB63[16] , \wRegInB63[15] , \wRegInB63[14] , \wRegInB63[13] , 
        \wRegInB63[12] , \wRegInB63[11] , \wRegInB63[10] , \wRegInB63[9] , 
        \wRegInB63[8] , \wRegInB63[7] , \wRegInB63[6] , \wRegInB63[5] , 
        \wRegInB63[4] , \wRegInB63[3] , \wRegInB63[2] , \wRegInB63[1] , 
        \wRegInB63[0] }), .LoOut({\wRegInA64[31] , \wRegInA64[30] , 
        \wRegInA64[29] , \wRegInA64[28] , \wRegInA64[27] , \wRegInA64[26] , 
        \wRegInA64[25] , \wRegInA64[24] , \wRegInA64[23] , \wRegInA64[22] , 
        \wRegInA64[21] , \wRegInA64[20] , \wRegInA64[19] , \wRegInA64[18] , 
        \wRegInA64[17] , \wRegInA64[16] , \wRegInA64[15] , \wRegInA64[14] , 
        \wRegInA64[13] , \wRegInA64[12] , \wRegInA64[11] , \wRegInA64[10] , 
        \wRegInA64[9] , \wRegInA64[8] , \wRegInA64[7] , \wRegInA64[6] , 
        \wRegInA64[5] , \wRegInA64[4] , \wRegInA64[3] , \wRegInA64[2] , 
        \wRegInA64[1] , \wRegInA64[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_156 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink157[31] , \ScanLink157[30] , \ScanLink157[29] , 
        \ScanLink157[28] , \ScanLink157[27] , \ScanLink157[26] , 
        \ScanLink157[25] , \ScanLink157[24] , \ScanLink157[23] , 
        \ScanLink157[22] , \ScanLink157[21] , \ScanLink157[20] , 
        \ScanLink157[19] , \ScanLink157[18] , \ScanLink157[17] , 
        \ScanLink157[16] , \ScanLink157[15] , \ScanLink157[14] , 
        \ScanLink157[13] , \ScanLink157[12] , \ScanLink157[11] , 
        \ScanLink157[10] , \ScanLink157[9] , \ScanLink157[8] , 
        \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , \ScanLink157[4] , 
        \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , \ScanLink157[0] 
        }), .ScanOut({\ScanLink156[31] , \ScanLink156[30] , \ScanLink156[29] , 
        \ScanLink156[28] , \ScanLink156[27] , \ScanLink156[26] , 
        \ScanLink156[25] , \ScanLink156[24] , \ScanLink156[23] , 
        \ScanLink156[22] , \ScanLink156[21] , \ScanLink156[20] , 
        \ScanLink156[19] , \ScanLink156[18] , \ScanLink156[17] , 
        \ScanLink156[16] , \ScanLink156[15] , \ScanLink156[14] , 
        \ScanLink156[13] , \ScanLink156[12] , \ScanLink156[11] , 
        \ScanLink156[10] , \ScanLink156[9] , \ScanLink156[8] , 
        \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , \ScanLink156[4] , 
        \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , \ScanLink156[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB49[31] , \wRegInB49[30] , \wRegInB49[29] , 
        \wRegInB49[28] , \wRegInB49[27] , \wRegInB49[26] , \wRegInB49[25] , 
        \wRegInB49[24] , \wRegInB49[23] , \wRegInB49[22] , \wRegInB49[21] , 
        \wRegInB49[20] , \wRegInB49[19] , \wRegInB49[18] , \wRegInB49[17] , 
        \wRegInB49[16] , \wRegInB49[15] , \wRegInB49[14] , \wRegInB49[13] , 
        \wRegInB49[12] , \wRegInB49[11] , \wRegInB49[10] , \wRegInB49[9] , 
        \wRegInB49[8] , \wRegInB49[7] , \wRegInB49[6] , \wRegInB49[5] , 
        \wRegInB49[4] , \wRegInB49[3] , \wRegInB49[2] , \wRegInB49[1] , 
        \wRegInB49[0] }), .Out({\wBIn49[31] , \wBIn49[30] , \wBIn49[29] , 
        \wBIn49[28] , \wBIn49[27] , \wBIn49[26] , \wBIn49[25] , \wBIn49[24] , 
        \wBIn49[23] , \wBIn49[22] , \wBIn49[21] , \wBIn49[20] , \wBIn49[19] , 
        \wBIn49[18] , \wBIn49[17] , \wBIn49[16] , \wBIn49[15] , \wBIn49[14] , 
        \wBIn49[13] , \wBIn49[12] , \wBIn49[11] , \wBIn49[10] , \wBIn49[9] , 
        \wBIn49[8] , \wBIn49[7] , \wBIn49[6] , \wBIn49[5] , \wBIn49[4] , 
        \wBIn49[3] , \wBIn49[2] , \wBIn49[1] , \wBIn49[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_241 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink242[31] , \ScanLink242[30] , \ScanLink242[29] , 
        \ScanLink242[28] , \ScanLink242[27] , \ScanLink242[26] , 
        \ScanLink242[25] , \ScanLink242[24] , \ScanLink242[23] , 
        \ScanLink242[22] , \ScanLink242[21] , \ScanLink242[20] , 
        \ScanLink242[19] , \ScanLink242[18] , \ScanLink242[17] , 
        \ScanLink242[16] , \ScanLink242[15] , \ScanLink242[14] , 
        \ScanLink242[13] , \ScanLink242[12] , \ScanLink242[11] , 
        \ScanLink242[10] , \ScanLink242[9] , \ScanLink242[8] , 
        \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , \ScanLink242[4] , 
        \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , \ScanLink242[0] 
        }), .ScanOut({\ScanLink241[31] , \ScanLink241[30] , \ScanLink241[29] , 
        \ScanLink241[28] , \ScanLink241[27] , \ScanLink241[26] , 
        \ScanLink241[25] , \ScanLink241[24] , \ScanLink241[23] , 
        \ScanLink241[22] , \ScanLink241[21] , \ScanLink241[20] , 
        \ScanLink241[19] , \ScanLink241[18] , \ScanLink241[17] , 
        \ScanLink241[16] , \ScanLink241[15] , \ScanLink241[14] , 
        \ScanLink241[13] , \ScanLink241[12] , \ScanLink241[11] , 
        \ScanLink241[10] , \ScanLink241[9] , \ScanLink241[8] , 
        \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , \ScanLink241[4] , 
        \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , \ScanLink241[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA7[31] , \wRegInA7[30] , \wRegInA7[29] , \wRegInA7[28] , 
        \wRegInA7[27] , \wRegInA7[26] , \wRegInA7[25] , \wRegInA7[24] , 
        \wRegInA7[23] , \wRegInA7[22] , \wRegInA7[21] , \wRegInA7[20] , 
        \wRegInA7[19] , \wRegInA7[18] , \wRegInA7[17] , \wRegInA7[16] , 
        \wRegInA7[15] , \wRegInA7[14] , \wRegInA7[13] , \wRegInA7[12] , 
        \wRegInA7[11] , \wRegInA7[10] , \wRegInA7[9] , \wRegInA7[8] , 
        \wRegInA7[7] , \wRegInA7[6] , \wRegInA7[5] , \wRegInA7[4] , 
        \wRegInA7[3] , \wRegInA7[2] , \wRegInA7[1] , \wRegInA7[0] }), .Out({
        \wAIn7[31] , \wAIn7[30] , \wAIn7[29] , \wAIn7[28] , \wAIn7[27] , 
        \wAIn7[26] , \wAIn7[25] , \wAIn7[24] , \wAIn7[23] , \wAIn7[22] , 
        \wAIn7[21] , \wAIn7[20] , \wAIn7[19] , \wAIn7[18] , \wAIn7[17] , 
        \wAIn7[16] , \wAIn7[15] , \wAIn7[14] , \wAIn7[13] , \wAIn7[12] , 
        \wAIn7[11] , \wAIn7[10] , \wAIn7[9] , \wAIn7[8] , \wAIn7[7] , 
        \wAIn7[6] , \wAIn7[5] , \wAIn7[4] , \wAIn7[3] , \wAIn7[2] , \wAIn7[1] , 
        \wAIn7[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid44[31] , \wAMid44[30] , \wAMid44[29] , \wAMid44[28] , 
        \wAMid44[27] , \wAMid44[26] , \wAMid44[25] , \wAMid44[24] , 
        \wAMid44[23] , \wAMid44[22] , \wAMid44[21] , \wAMid44[20] , 
        \wAMid44[19] , \wAMid44[18] , \wAMid44[17] , \wAMid44[16] , 
        \wAMid44[15] , \wAMid44[14] , \wAMid44[13] , \wAMid44[12] , 
        \wAMid44[11] , \wAMid44[10] , \wAMid44[9] , \wAMid44[8] , \wAMid44[7] , 
        \wAMid44[6] , \wAMid44[5] , \wAMid44[4] , \wAMid44[3] , \wAMid44[2] , 
        \wAMid44[1] , \wAMid44[0] }), .BIn({\wBMid44[31] , \wBMid44[30] , 
        \wBMid44[29] , \wBMid44[28] , \wBMid44[27] , \wBMid44[26] , 
        \wBMid44[25] , \wBMid44[24] , \wBMid44[23] , \wBMid44[22] , 
        \wBMid44[21] , \wBMid44[20] , \wBMid44[19] , \wBMid44[18] , 
        \wBMid44[17] , \wBMid44[16] , \wBMid44[15] , \wBMid44[14] , 
        \wBMid44[13] , \wBMid44[12] , \wBMid44[11] , \wBMid44[10] , 
        \wBMid44[9] , \wBMid44[8] , \wBMid44[7] , \wBMid44[6] , \wBMid44[5] , 
        \wBMid44[4] , \wBMid44[3] , \wBMid44[2] , \wBMid44[1] , \wBMid44[0] }), 
        .HiOut({\wRegInB44[31] , \wRegInB44[30] , \wRegInB44[29] , 
        \wRegInB44[28] , \wRegInB44[27] , \wRegInB44[26] , \wRegInB44[25] , 
        \wRegInB44[24] , \wRegInB44[23] , \wRegInB44[22] , \wRegInB44[21] , 
        \wRegInB44[20] , \wRegInB44[19] , \wRegInB44[18] , \wRegInB44[17] , 
        \wRegInB44[16] , \wRegInB44[15] , \wRegInB44[14] , \wRegInB44[13] , 
        \wRegInB44[12] , \wRegInB44[11] , \wRegInB44[10] , \wRegInB44[9] , 
        \wRegInB44[8] , \wRegInB44[7] , \wRegInB44[6] , \wRegInB44[5] , 
        \wRegInB44[4] , \wRegInB44[3] , \wRegInB44[2] , \wRegInB44[1] , 
        \wRegInB44[0] }), .LoOut({\wRegInA45[31] , \wRegInA45[30] , 
        \wRegInA45[29] , \wRegInA45[28] , \wRegInA45[27] , \wRegInA45[26] , 
        \wRegInA45[25] , \wRegInA45[24] , \wRegInA45[23] , \wRegInA45[22] , 
        \wRegInA45[21] , \wRegInA45[20] , \wRegInA45[19] , \wRegInA45[18] , 
        \wRegInA45[17] , \wRegInA45[16] , \wRegInA45[15] , \wRegInA45[14] , 
        \wRegInA45[13] , \wRegInA45[12] , \wRegInA45[11] , \wRegInA45[10] , 
        \wRegInA45[9] , \wRegInA45[8] , \wRegInA45[7] , \wRegInA45[6] , 
        \wRegInA45[5] , \wRegInA45[4] , \wRegInA45[3] , \wRegInA45[2] , 
        \wRegInA45[1] , \wRegInA45[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid78[31] , \wAMid78[30] , \wAMid78[29] , \wAMid78[28] , 
        \wAMid78[27] , \wAMid78[26] , \wAMid78[25] , \wAMid78[24] , 
        \wAMid78[23] , \wAMid78[22] , \wAMid78[21] , \wAMid78[20] , 
        \wAMid78[19] , \wAMid78[18] , \wAMid78[17] , \wAMid78[16] , 
        \wAMid78[15] , \wAMid78[14] , \wAMid78[13] , \wAMid78[12] , 
        \wAMid78[11] , \wAMid78[10] , \wAMid78[9] , \wAMid78[8] , \wAMid78[7] , 
        \wAMid78[6] , \wAMid78[5] , \wAMid78[4] , \wAMid78[3] , \wAMid78[2] , 
        \wAMid78[1] , \wAMid78[0] }), .BIn({\wBMid78[31] , \wBMid78[30] , 
        \wBMid78[29] , \wBMid78[28] , \wBMid78[27] , \wBMid78[26] , 
        \wBMid78[25] , \wBMid78[24] , \wBMid78[23] , \wBMid78[22] , 
        \wBMid78[21] , \wBMid78[20] , \wBMid78[19] , \wBMid78[18] , 
        \wBMid78[17] , \wBMid78[16] , \wBMid78[15] , \wBMid78[14] , 
        \wBMid78[13] , \wBMid78[12] , \wBMid78[11] , \wBMid78[10] , 
        \wBMid78[9] , \wBMid78[8] , \wBMid78[7] , \wBMid78[6] , \wBMid78[5] , 
        \wBMid78[4] , \wBMid78[3] , \wBMid78[2] , \wBMid78[1] , \wBMid78[0] }), 
        .HiOut({\wRegInB78[31] , \wRegInB78[30] , \wRegInB78[29] , 
        \wRegInB78[28] , \wRegInB78[27] , \wRegInB78[26] , \wRegInB78[25] , 
        \wRegInB78[24] , \wRegInB78[23] , \wRegInB78[22] , \wRegInB78[21] , 
        \wRegInB78[20] , \wRegInB78[19] , \wRegInB78[18] , \wRegInB78[17] , 
        \wRegInB78[16] , \wRegInB78[15] , \wRegInB78[14] , \wRegInB78[13] , 
        \wRegInB78[12] , \wRegInB78[11] , \wRegInB78[10] , \wRegInB78[9] , 
        \wRegInB78[8] , \wRegInB78[7] , \wRegInB78[6] , \wRegInB78[5] , 
        \wRegInB78[4] , \wRegInB78[3] , \wRegInB78[2] , \wRegInB78[1] , 
        \wRegInB78[0] }), .LoOut({\wRegInA79[31] , \wRegInA79[30] , 
        \wRegInA79[29] , \wRegInA79[28] , \wRegInA79[27] , \wRegInA79[26] , 
        \wRegInA79[25] , \wRegInA79[24] , \wRegInA79[23] , \wRegInA79[22] , 
        \wRegInA79[21] , \wRegInA79[20] , \wRegInA79[19] , \wRegInA79[18] , 
        \wRegInA79[17] , \wRegInA79[16] , \wRegInA79[15] , \wRegInA79[14] , 
        \wRegInA79[13] , \wRegInA79[12] , \wRegInA79[11] , \wRegInA79[10] , 
        \wRegInA79[9] , \wRegInA79[8] , \wRegInA79[7] , \wRegInA79[6] , 
        \wRegInA79[5] , \wRegInA79[4] , \wRegInA79[3] , \wRegInA79[2] , 
        \wRegInA79[1] , \wRegInA79[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid115[31] , \wAMid115[30] , \wAMid115[29] , \wAMid115[28] , 
        \wAMid115[27] , \wAMid115[26] , \wAMid115[25] , \wAMid115[24] , 
        \wAMid115[23] , \wAMid115[22] , \wAMid115[21] , \wAMid115[20] , 
        \wAMid115[19] , \wAMid115[18] , \wAMid115[17] , \wAMid115[16] , 
        \wAMid115[15] , \wAMid115[14] , \wAMid115[13] , \wAMid115[12] , 
        \wAMid115[11] , \wAMid115[10] , \wAMid115[9] , \wAMid115[8] , 
        \wAMid115[7] , \wAMid115[6] , \wAMid115[5] , \wAMid115[4] , 
        \wAMid115[3] , \wAMid115[2] , \wAMid115[1] , \wAMid115[0] }), .BIn({
        \wBMid115[31] , \wBMid115[30] , \wBMid115[29] , \wBMid115[28] , 
        \wBMid115[27] , \wBMid115[26] , \wBMid115[25] , \wBMid115[24] , 
        \wBMid115[23] , \wBMid115[22] , \wBMid115[21] , \wBMid115[20] , 
        \wBMid115[19] , \wBMid115[18] , \wBMid115[17] , \wBMid115[16] , 
        \wBMid115[15] , \wBMid115[14] , \wBMid115[13] , \wBMid115[12] , 
        \wBMid115[11] , \wBMid115[10] , \wBMid115[9] , \wBMid115[8] , 
        \wBMid115[7] , \wBMid115[6] , \wBMid115[5] , \wBMid115[4] , 
        \wBMid115[3] , \wBMid115[2] , \wBMid115[1] , \wBMid115[0] }), .HiOut({
        \wRegInB115[31] , \wRegInB115[30] , \wRegInB115[29] , \wRegInB115[28] , 
        \wRegInB115[27] , \wRegInB115[26] , \wRegInB115[25] , \wRegInB115[24] , 
        \wRegInB115[23] , \wRegInB115[22] , \wRegInB115[21] , \wRegInB115[20] , 
        \wRegInB115[19] , \wRegInB115[18] , \wRegInB115[17] , \wRegInB115[16] , 
        \wRegInB115[15] , \wRegInB115[14] , \wRegInB115[13] , \wRegInB115[12] , 
        \wRegInB115[11] , \wRegInB115[10] , \wRegInB115[9] , \wRegInB115[8] , 
        \wRegInB115[7] , \wRegInB115[6] , \wRegInB115[5] , \wRegInB115[4] , 
        \wRegInB115[3] , \wRegInB115[2] , \wRegInB115[1] , \wRegInB115[0] }), 
        .LoOut({\wRegInA116[31] , \wRegInA116[30] , \wRegInA116[29] , 
        \wRegInA116[28] , \wRegInA116[27] , \wRegInA116[26] , \wRegInA116[25] , 
        \wRegInA116[24] , \wRegInA116[23] , \wRegInA116[22] , \wRegInA116[21] , 
        \wRegInA116[20] , \wRegInA116[19] , \wRegInA116[18] , \wRegInA116[17] , 
        \wRegInA116[16] , \wRegInA116[15] , \wRegInA116[14] , \wRegInA116[13] , 
        \wRegInA116[12] , \wRegInA116[11] , \wRegInA116[10] , \wRegInA116[9] , 
        \wRegInA116[8] , \wRegInA116[7] , \wRegInA116[6] , \wRegInA116[5] , 
        \wRegInA116[4] , \wRegInA116[3] , \wRegInA116[2] , \wRegInA116[1] , 
        \wRegInA116[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_171 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink172[31] , \ScanLink172[30] , \ScanLink172[29] , 
        \ScanLink172[28] , \ScanLink172[27] , \ScanLink172[26] , 
        \ScanLink172[25] , \ScanLink172[24] , \ScanLink172[23] , 
        \ScanLink172[22] , \ScanLink172[21] , \ScanLink172[20] , 
        \ScanLink172[19] , \ScanLink172[18] , \ScanLink172[17] , 
        \ScanLink172[16] , \ScanLink172[15] , \ScanLink172[14] , 
        \ScanLink172[13] , \ScanLink172[12] , \ScanLink172[11] , 
        \ScanLink172[10] , \ScanLink172[9] , \ScanLink172[8] , 
        \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , \ScanLink172[4] , 
        \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , \ScanLink172[0] 
        }), .ScanOut({\ScanLink171[31] , \ScanLink171[30] , \ScanLink171[29] , 
        \ScanLink171[28] , \ScanLink171[27] , \ScanLink171[26] , 
        \ScanLink171[25] , \ScanLink171[24] , \ScanLink171[23] , 
        \ScanLink171[22] , \ScanLink171[21] , \ScanLink171[20] , 
        \ScanLink171[19] , \ScanLink171[18] , \ScanLink171[17] , 
        \ScanLink171[16] , \ScanLink171[15] , \ScanLink171[14] , 
        \ScanLink171[13] , \ScanLink171[12] , \ScanLink171[11] , 
        \ScanLink171[10] , \ScanLink171[9] , \ScanLink171[8] , 
        \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , \ScanLink171[4] , 
        \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , \ScanLink171[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA42[31] , \wRegInA42[30] , \wRegInA42[29] , 
        \wRegInA42[28] , \wRegInA42[27] , \wRegInA42[26] , \wRegInA42[25] , 
        \wRegInA42[24] , \wRegInA42[23] , \wRegInA42[22] , \wRegInA42[21] , 
        \wRegInA42[20] , \wRegInA42[19] , \wRegInA42[18] , \wRegInA42[17] , 
        \wRegInA42[16] , \wRegInA42[15] , \wRegInA42[14] , \wRegInA42[13] , 
        \wRegInA42[12] , \wRegInA42[11] , \wRegInA42[10] , \wRegInA42[9] , 
        \wRegInA42[8] , \wRegInA42[7] , \wRegInA42[6] , \wRegInA42[5] , 
        \wRegInA42[4] , \wRegInA42[3] , \wRegInA42[2] , \wRegInA42[1] , 
        \wRegInA42[0] }), .Out({\wAIn42[31] , \wAIn42[30] , \wAIn42[29] , 
        \wAIn42[28] , \wAIn42[27] , \wAIn42[26] , \wAIn42[25] , \wAIn42[24] , 
        \wAIn42[23] , \wAIn42[22] , \wAIn42[21] , \wAIn42[20] , \wAIn42[19] , 
        \wAIn42[18] , \wAIn42[17] , \wAIn42[16] , \wAIn42[15] , \wAIn42[14] , 
        \wAIn42[13] , \wAIn42[12] , \wAIn42[11] , \wAIn42[10] , \wAIn42[9] , 
        \wAIn42[8] , \wAIn42[7] , \wAIn42[6] , \wAIn42[5] , \wAIn42[4] , 
        \wAIn42[3] , \wAIn42[2] , \wAIn42[1] , \wAIn42[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_21 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink22[31] , \ScanLink22[30] , \ScanLink22[29] , 
        \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , \ScanLink22[25] , 
        \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , \ScanLink22[21] , 
        \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , \ScanLink22[17] , 
        \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , \ScanLink22[13] , 
        \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , \ScanLink22[9] , 
        \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , \ScanLink22[5] , 
        \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , \ScanLink22[1] , 
        \ScanLink22[0] }), .ScanOut({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA117[31] , \wRegInA117[30] , 
        \wRegInA117[29] , \wRegInA117[28] , \wRegInA117[27] , \wRegInA117[26] , 
        \wRegInA117[25] , \wRegInA117[24] , \wRegInA117[23] , \wRegInA117[22] , 
        \wRegInA117[21] , \wRegInA117[20] , \wRegInA117[19] , \wRegInA117[18] , 
        \wRegInA117[17] , \wRegInA117[16] , \wRegInA117[15] , \wRegInA117[14] , 
        \wRegInA117[13] , \wRegInA117[12] , \wRegInA117[11] , \wRegInA117[10] , 
        \wRegInA117[9] , \wRegInA117[8] , \wRegInA117[7] , \wRegInA117[6] , 
        \wRegInA117[5] , \wRegInA117[4] , \wRegInA117[3] , \wRegInA117[2] , 
        \wRegInA117[1] , \wRegInA117[0] }), .Out({\wAIn117[31] , \wAIn117[30] , 
        \wAIn117[29] , \wAIn117[28] , \wAIn117[27] , \wAIn117[26] , 
        \wAIn117[25] , \wAIn117[24] , \wAIn117[23] , \wAIn117[22] , 
        \wAIn117[21] , \wAIn117[20] , \wAIn117[19] , \wAIn117[18] , 
        \wAIn117[17] , \wAIn117[16] , \wAIn117[15] , \wAIn117[14] , 
        \wAIn117[13] , \wAIn117[12] , \wAIn117[11] , \wAIn117[10] , 
        \wAIn117[9] , \wAIn117[8] , \wAIn117[7] , \wAIn117[6] , \wAIn117[5] , 
        \wAIn117[4] , \wAIn117[3] , \wAIn117[2] , \wAIn117[1] , \wAIn117[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_96 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink97[31] , \ScanLink97[30] , \ScanLink97[29] , 
        \ScanLink97[28] , \ScanLink97[27] , \ScanLink97[26] , \ScanLink97[25] , 
        \ScanLink97[24] , \ScanLink97[23] , \ScanLink97[22] , \ScanLink97[21] , 
        \ScanLink97[20] , \ScanLink97[19] , \ScanLink97[18] , \ScanLink97[17] , 
        \ScanLink97[16] , \ScanLink97[15] , \ScanLink97[14] , \ScanLink97[13] , 
        \ScanLink97[12] , \ScanLink97[11] , \ScanLink97[10] , \ScanLink97[9] , 
        \ScanLink97[8] , \ScanLink97[7] , \ScanLink97[6] , \ScanLink97[5] , 
        \ScanLink97[4] , \ScanLink97[3] , \ScanLink97[2] , \ScanLink97[1] , 
        \ScanLink97[0] }), .ScanOut({\ScanLink96[31] , \ScanLink96[30] , 
        \ScanLink96[29] , \ScanLink96[28] , \ScanLink96[27] , \ScanLink96[26] , 
        \ScanLink96[25] , \ScanLink96[24] , \ScanLink96[23] , \ScanLink96[22] , 
        \ScanLink96[21] , \ScanLink96[20] , \ScanLink96[19] , \ScanLink96[18] , 
        \ScanLink96[17] , \ScanLink96[16] , \ScanLink96[15] , \ScanLink96[14] , 
        \ScanLink96[13] , \ScanLink96[12] , \ScanLink96[11] , \ScanLink96[10] , 
        \ScanLink96[9] , \ScanLink96[8] , \ScanLink96[7] , \ScanLink96[6] , 
        \ScanLink96[5] , \ScanLink96[4] , \ScanLink96[3] , \ScanLink96[2] , 
        \ScanLink96[1] , \ScanLink96[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB79[31] , \wRegInB79[30] , 
        \wRegInB79[29] , \wRegInB79[28] , \wRegInB79[27] , \wRegInB79[26] , 
        \wRegInB79[25] , \wRegInB79[24] , \wRegInB79[23] , \wRegInB79[22] , 
        \wRegInB79[21] , \wRegInB79[20] , \wRegInB79[19] , \wRegInB79[18] , 
        \wRegInB79[17] , \wRegInB79[16] , \wRegInB79[15] , \wRegInB79[14] , 
        \wRegInB79[13] , \wRegInB79[12] , \wRegInB79[11] , \wRegInB79[10] , 
        \wRegInB79[9] , \wRegInB79[8] , \wRegInB79[7] , \wRegInB79[6] , 
        \wRegInB79[5] , \wRegInB79[4] , \wRegInB79[3] , \wRegInB79[2] , 
        \wRegInB79[1] , \wRegInB79[0] }), .Out({\wBIn79[31] , \wBIn79[30] , 
        \wBIn79[29] , \wBIn79[28] , \wBIn79[27] , \wBIn79[26] , \wBIn79[25] , 
        \wBIn79[24] , \wBIn79[23] , \wBIn79[22] , \wBIn79[21] , \wBIn79[20] , 
        \wBIn79[19] , \wBIn79[18] , \wBIn79[17] , \wBIn79[16] , \wBIn79[15] , 
        \wBIn79[14] , \wBIn79[13] , \wBIn79[12] , \wBIn79[11] , \wBIn79[10] , 
        \wBIn79[9] , \wBIn79[8] , \wBIn79[7] , \wBIn79[6] , \wBIn79[5] , 
        \wBIn79[4] , \wBIn79[3] , \wBIn79[2] , \wBIn79[1] , \wBIn79[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid16[31] , \wAMid16[30] , \wAMid16[29] , \wAMid16[28] , 
        \wAMid16[27] , \wAMid16[26] , \wAMid16[25] , \wAMid16[24] , 
        \wAMid16[23] , \wAMid16[22] , \wAMid16[21] , \wAMid16[20] , 
        \wAMid16[19] , \wAMid16[18] , \wAMid16[17] , \wAMid16[16] , 
        \wAMid16[15] , \wAMid16[14] , \wAMid16[13] , \wAMid16[12] , 
        \wAMid16[11] , \wAMid16[10] , \wAMid16[9] , \wAMid16[8] , \wAMid16[7] , 
        \wAMid16[6] , \wAMid16[5] , \wAMid16[4] , \wAMid16[3] , \wAMid16[2] , 
        \wAMid16[1] , \wAMid16[0] }), .BIn({\wBMid16[31] , \wBMid16[30] , 
        \wBMid16[29] , \wBMid16[28] , \wBMid16[27] , \wBMid16[26] , 
        \wBMid16[25] , \wBMid16[24] , \wBMid16[23] , \wBMid16[22] , 
        \wBMid16[21] , \wBMid16[20] , \wBMid16[19] , \wBMid16[18] , 
        \wBMid16[17] , \wBMid16[16] , \wBMid16[15] , \wBMid16[14] , 
        \wBMid16[13] , \wBMid16[12] , \wBMid16[11] , \wBMid16[10] , 
        \wBMid16[9] , \wBMid16[8] , \wBMid16[7] , \wBMid16[6] , \wBMid16[5] , 
        \wBMid16[4] , \wBMid16[3] , \wBMid16[2] , \wBMid16[1] , \wBMid16[0] }), 
        .HiOut({\wRegInB16[31] , \wRegInB16[30] , \wRegInB16[29] , 
        \wRegInB16[28] , \wRegInB16[27] , \wRegInB16[26] , \wRegInB16[25] , 
        \wRegInB16[24] , \wRegInB16[23] , \wRegInB16[22] , \wRegInB16[21] , 
        \wRegInB16[20] , \wRegInB16[19] , \wRegInB16[18] , \wRegInB16[17] , 
        \wRegInB16[16] , \wRegInB16[15] , \wRegInB16[14] , \wRegInB16[13] , 
        \wRegInB16[12] , \wRegInB16[11] , \wRegInB16[10] , \wRegInB16[9] , 
        \wRegInB16[8] , \wRegInB16[7] , \wRegInB16[6] , \wRegInB16[5] , 
        \wRegInB16[4] , \wRegInB16[3] , \wRegInB16[2] , \wRegInB16[1] , 
        \wRegInB16[0] }), .LoOut({\wRegInA17[31] , \wRegInA17[30] , 
        \wRegInA17[29] , \wRegInA17[28] , \wRegInA17[27] , \wRegInA17[26] , 
        \wRegInA17[25] , \wRegInA17[24] , \wRegInA17[23] , \wRegInA17[22] , 
        \wRegInA17[21] , \wRegInA17[20] , \wRegInA17[19] , \wRegInA17[18] , 
        \wRegInA17[17] , \wRegInA17[16] , \wRegInA17[15] , \wRegInA17[14] , 
        \wRegInA17[13] , \wRegInA17[12] , \wRegInA17[11] , \wRegInA17[10] , 
        \wRegInA17[9] , \wRegInA17[8] , \wRegInA17[7] , \wRegInA17[6] , 
        \wRegInA17[5] , \wRegInA17[4] , \wRegInA17[3] , \wRegInA17[2] , 
        \wRegInA17[1] , \wRegInA17[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_213 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink214[31] , \ScanLink214[30] , \ScanLink214[29] , 
        \ScanLink214[28] , \ScanLink214[27] , \ScanLink214[26] , 
        \ScanLink214[25] , \ScanLink214[24] , \ScanLink214[23] , 
        \ScanLink214[22] , \ScanLink214[21] , \ScanLink214[20] , 
        \ScanLink214[19] , \ScanLink214[18] , \ScanLink214[17] , 
        \ScanLink214[16] , \ScanLink214[15] , \ScanLink214[14] , 
        \ScanLink214[13] , \ScanLink214[12] , \ScanLink214[11] , 
        \ScanLink214[10] , \ScanLink214[9] , \ScanLink214[8] , 
        \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , \ScanLink214[4] , 
        \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , \ScanLink214[0] 
        }), .ScanOut({\ScanLink213[31] , \ScanLink213[30] , \ScanLink213[29] , 
        \ScanLink213[28] , \ScanLink213[27] , \ScanLink213[26] , 
        \ScanLink213[25] , \ScanLink213[24] , \ScanLink213[23] , 
        \ScanLink213[22] , \ScanLink213[21] , \ScanLink213[20] , 
        \ScanLink213[19] , \ScanLink213[18] , \ScanLink213[17] , 
        \ScanLink213[16] , \ScanLink213[15] , \ScanLink213[14] , 
        \ScanLink213[13] , \ScanLink213[12] , \ScanLink213[11] , 
        \ScanLink213[10] , \ScanLink213[9] , \ScanLink213[8] , 
        \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , \ScanLink213[4] , 
        \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , \ScanLink213[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA21[31] , \wRegInA21[30] , \wRegInA21[29] , 
        \wRegInA21[28] , \wRegInA21[27] , \wRegInA21[26] , \wRegInA21[25] , 
        \wRegInA21[24] , \wRegInA21[23] , \wRegInA21[22] , \wRegInA21[21] , 
        \wRegInA21[20] , \wRegInA21[19] , \wRegInA21[18] , \wRegInA21[17] , 
        \wRegInA21[16] , \wRegInA21[15] , \wRegInA21[14] , \wRegInA21[13] , 
        \wRegInA21[12] , \wRegInA21[11] , \wRegInA21[10] , \wRegInA21[9] , 
        \wRegInA21[8] , \wRegInA21[7] , \wRegInA21[6] , \wRegInA21[5] , 
        \wRegInA21[4] , \wRegInA21[3] , \wRegInA21[2] , \wRegInA21[1] , 
        \wRegInA21[0] }), .Out({\wAIn21[31] , \wAIn21[30] , \wAIn21[29] , 
        \wAIn21[28] , \wAIn21[27] , \wAIn21[26] , \wAIn21[25] , \wAIn21[24] , 
        \wAIn21[23] , \wAIn21[22] , \wAIn21[21] , \wAIn21[20] , \wAIn21[19] , 
        \wAIn21[18] , \wAIn21[17] , \wAIn21[16] , \wAIn21[15] , \wAIn21[14] , 
        \wAIn21[13] , \wAIn21[12] , \wAIn21[11] , \wAIn21[10] , \wAIn21[9] , 
        \wAIn21[8] , \wAIn21[7] , \wAIn21[6] , \wAIn21[5] , \wAIn21[4] , 
        \wAIn21[3] , \wAIn21[2] , \wAIn21[1] , \wAIn21[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_73 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink74[31] , \ScanLink74[30] , \ScanLink74[29] , 
        \ScanLink74[28] , \ScanLink74[27] , \ScanLink74[26] , \ScanLink74[25] , 
        \ScanLink74[24] , \ScanLink74[23] , \ScanLink74[22] , \ScanLink74[21] , 
        \ScanLink74[20] , \ScanLink74[19] , \ScanLink74[18] , \ScanLink74[17] , 
        \ScanLink74[16] , \ScanLink74[15] , \ScanLink74[14] , \ScanLink74[13] , 
        \ScanLink74[12] , \ScanLink74[11] , \ScanLink74[10] , \ScanLink74[9] , 
        \ScanLink74[8] , \ScanLink74[7] , \ScanLink74[6] , \ScanLink74[5] , 
        \ScanLink74[4] , \ScanLink74[3] , \ScanLink74[2] , \ScanLink74[1] , 
        \ScanLink74[0] }), .ScanOut({\ScanLink73[31] , \ScanLink73[30] , 
        \ScanLink73[29] , \ScanLink73[28] , \ScanLink73[27] , \ScanLink73[26] , 
        \ScanLink73[25] , \ScanLink73[24] , \ScanLink73[23] , \ScanLink73[22] , 
        \ScanLink73[21] , \ScanLink73[20] , \ScanLink73[19] , \ScanLink73[18] , 
        \ScanLink73[17] , \ScanLink73[16] , \ScanLink73[15] , \ScanLink73[14] , 
        \ScanLink73[13] , \ScanLink73[12] , \ScanLink73[11] , \ScanLink73[10] , 
        \ScanLink73[9] , \ScanLink73[8] , \ScanLink73[7] , \ScanLink73[6] , 
        \ScanLink73[5] , \ScanLink73[4] , \ScanLink73[3] , \ScanLink73[2] , 
        \ScanLink73[1] , \ScanLink73[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA91[31] , \wRegInA91[30] , 
        \wRegInA91[29] , \wRegInA91[28] , \wRegInA91[27] , \wRegInA91[26] , 
        \wRegInA91[25] , \wRegInA91[24] , \wRegInA91[23] , \wRegInA91[22] , 
        \wRegInA91[21] , \wRegInA91[20] , \wRegInA91[19] , \wRegInA91[18] , 
        \wRegInA91[17] , \wRegInA91[16] , \wRegInA91[15] , \wRegInA91[14] , 
        \wRegInA91[13] , \wRegInA91[12] , \wRegInA91[11] , \wRegInA91[10] , 
        \wRegInA91[9] , \wRegInA91[8] , \wRegInA91[7] , \wRegInA91[6] , 
        \wRegInA91[5] , \wRegInA91[4] , \wRegInA91[3] , \wRegInA91[2] , 
        \wRegInA91[1] , \wRegInA91[0] }), .Out({\wAIn91[31] , \wAIn91[30] , 
        \wAIn91[29] , \wAIn91[28] , \wAIn91[27] , \wAIn91[26] , \wAIn91[25] , 
        \wAIn91[24] , \wAIn91[23] , \wAIn91[22] , \wAIn91[21] , \wAIn91[20] , 
        \wAIn91[19] , \wAIn91[18] , \wAIn91[17] , \wAIn91[16] , \wAIn91[15] , 
        \wAIn91[14] , \wAIn91[13] , \wAIn91[12] , \wAIn91[11] , \wAIn91[10] , 
        \wAIn91[9] , \wAIn91[8] , \wAIn91[7] , \wAIn91[6] , \wAIn91[5] , 
        \wAIn91[4] , \wAIn91[3] , \wAIn91[2] , \wAIn91[1] , \wAIn91[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_123 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink124[31] , \ScanLink124[30] , \ScanLink124[29] , 
        \ScanLink124[28] , \ScanLink124[27] , \ScanLink124[26] , 
        \ScanLink124[25] , \ScanLink124[24] , \ScanLink124[23] , 
        \ScanLink124[22] , \ScanLink124[21] , \ScanLink124[20] , 
        \ScanLink124[19] , \ScanLink124[18] , \ScanLink124[17] , 
        \ScanLink124[16] , \ScanLink124[15] , \ScanLink124[14] , 
        \ScanLink124[13] , \ScanLink124[12] , \ScanLink124[11] , 
        \ScanLink124[10] , \ScanLink124[9] , \ScanLink124[8] , 
        \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , \ScanLink124[4] , 
        \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , \ScanLink124[0] 
        }), .ScanOut({\ScanLink123[31] , \ScanLink123[30] , \ScanLink123[29] , 
        \ScanLink123[28] , \ScanLink123[27] , \ScanLink123[26] , 
        \ScanLink123[25] , \ScanLink123[24] , \ScanLink123[23] , 
        \ScanLink123[22] , \ScanLink123[21] , \ScanLink123[20] , 
        \ScanLink123[19] , \ScanLink123[18] , \ScanLink123[17] , 
        \ScanLink123[16] , \ScanLink123[15] , \ScanLink123[14] , 
        \ScanLink123[13] , \ScanLink123[12] , \ScanLink123[11] , 
        \ScanLink123[10] , \ScanLink123[9] , \ScanLink123[8] , 
        \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , \ScanLink123[4] , 
        \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , \ScanLink123[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA66[31] , \wRegInA66[30] , \wRegInA66[29] , 
        \wRegInA66[28] , \wRegInA66[27] , \wRegInA66[26] , \wRegInA66[25] , 
        \wRegInA66[24] , \wRegInA66[23] , \wRegInA66[22] , \wRegInA66[21] , 
        \wRegInA66[20] , \wRegInA66[19] , \wRegInA66[18] , \wRegInA66[17] , 
        \wRegInA66[16] , \wRegInA66[15] , \wRegInA66[14] , \wRegInA66[13] , 
        \wRegInA66[12] , \wRegInA66[11] , \wRegInA66[10] , \wRegInA66[9] , 
        \wRegInA66[8] , \wRegInA66[7] , \wRegInA66[6] , \wRegInA66[5] , 
        \wRegInA66[4] , \wRegInA66[3] , \wRegInA66[2] , \wRegInA66[1] , 
        \wRegInA66[0] }), .Out({\wAIn66[31] , \wAIn66[30] , \wAIn66[29] , 
        \wAIn66[28] , \wAIn66[27] , \wAIn66[26] , \wAIn66[25] , \wAIn66[24] , 
        \wAIn66[23] , \wAIn66[22] , \wAIn66[21] , \wAIn66[20] , \wAIn66[19] , 
        \wAIn66[18] , \wAIn66[17] , \wAIn66[16] , \wAIn66[15] , \wAIn66[14] , 
        \wAIn66[13] , \wAIn66[12] , \wAIn66[11] , \wAIn66[10] , \wAIn66[9] , 
        \wAIn66[8] , \wAIn66[7] , \wAIn66[6] , \wAIn66[5] , \wAIn66[4] , 
        \wAIn66[3] , \wAIn66[2] , \wAIn66[1] , \wAIn66[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid31[31] , \wAMid31[30] , \wAMid31[29] , \wAMid31[28] , 
        \wAMid31[27] , \wAMid31[26] , \wAMid31[25] , \wAMid31[24] , 
        \wAMid31[23] , \wAMid31[22] , \wAMid31[21] , \wAMid31[20] , 
        \wAMid31[19] , \wAMid31[18] , \wAMid31[17] , \wAMid31[16] , 
        \wAMid31[15] , \wAMid31[14] , \wAMid31[13] , \wAMid31[12] , 
        \wAMid31[11] , \wAMid31[10] , \wAMid31[9] , \wAMid31[8] , \wAMid31[7] , 
        \wAMid31[6] , \wAMid31[5] , \wAMid31[4] , \wAMid31[3] , \wAMid31[2] , 
        \wAMid31[1] , \wAMid31[0] }), .BIn({\wBMid31[31] , \wBMid31[30] , 
        \wBMid31[29] , \wBMid31[28] , \wBMid31[27] , \wBMid31[26] , 
        \wBMid31[25] , \wBMid31[24] , \wBMid31[23] , \wBMid31[22] , 
        \wBMid31[21] , \wBMid31[20] , \wBMid31[19] , \wBMid31[18] , 
        \wBMid31[17] , \wBMid31[16] , \wBMid31[15] , \wBMid31[14] , 
        \wBMid31[13] , \wBMid31[12] , \wBMid31[11] , \wBMid31[10] , 
        \wBMid31[9] , \wBMid31[8] , \wBMid31[7] , \wBMid31[6] , \wBMid31[5] , 
        \wBMid31[4] , \wBMid31[3] , \wBMid31[2] , \wBMid31[1] , \wBMid31[0] }), 
        .HiOut({\wRegInB31[31] , \wRegInB31[30] , \wRegInB31[29] , 
        \wRegInB31[28] , \wRegInB31[27] , \wRegInB31[26] , \wRegInB31[25] , 
        \wRegInB31[24] , \wRegInB31[23] , \wRegInB31[22] , \wRegInB31[21] , 
        \wRegInB31[20] , \wRegInB31[19] , \wRegInB31[18] , \wRegInB31[17] , 
        \wRegInB31[16] , \wRegInB31[15] , \wRegInB31[14] , \wRegInB31[13] , 
        \wRegInB31[12] , \wRegInB31[11] , \wRegInB31[10] , \wRegInB31[9] , 
        \wRegInB31[8] , \wRegInB31[7] , \wRegInB31[6] , \wRegInB31[5] , 
        \wRegInB31[4] , \wRegInB31[3] , \wRegInB31[2] , \wRegInB31[1] , 
        \wRegInB31[0] }), .LoOut({\wRegInA32[31] , \wRegInA32[30] , 
        \wRegInA32[29] , \wRegInA32[28] , \wRegInA32[27] , \wRegInA32[26] , 
        \wRegInA32[25] , \wRegInA32[24] , \wRegInA32[23] , \wRegInA32[22] , 
        \wRegInA32[21] , \wRegInA32[20] , \wRegInA32[19] , \wRegInA32[18] , 
        \wRegInA32[17] , \wRegInA32[16] , \wRegInA32[15] , \wRegInA32[14] , 
        \wRegInA32[13] , \wRegInA32[12] , \wRegInA32[11] , \wRegInA32[10] , 
        \wRegInA32[9] , \wRegInA32[8] , \wRegInA32[7] , \wRegInA32[6] , 
        \wRegInA32[5] , \wRegInA32[4] , \wRegInA32[3] , \wRegInA32[2] , 
        \wRegInA32[1] , \wRegInA32[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_234 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink235[31] , \ScanLink235[30] , \ScanLink235[29] , 
        \ScanLink235[28] , \ScanLink235[27] , \ScanLink235[26] , 
        \ScanLink235[25] , \ScanLink235[24] , \ScanLink235[23] , 
        \ScanLink235[22] , \ScanLink235[21] , \ScanLink235[20] , 
        \ScanLink235[19] , \ScanLink235[18] , \ScanLink235[17] , 
        \ScanLink235[16] , \ScanLink235[15] , \ScanLink235[14] , 
        \ScanLink235[13] , \ScanLink235[12] , \ScanLink235[11] , 
        \ScanLink235[10] , \ScanLink235[9] , \ScanLink235[8] , 
        \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , \ScanLink235[4] , 
        \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , \ScanLink235[0] 
        }), .ScanOut({\ScanLink234[31] , \ScanLink234[30] , \ScanLink234[29] , 
        \ScanLink234[28] , \ScanLink234[27] , \ScanLink234[26] , 
        \ScanLink234[25] , \ScanLink234[24] , \ScanLink234[23] , 
        \ScanLink234[22] , \ScanLink234[21] , \ScanLink234[20] , 
        \ScanLink234[19] , \ScanLink234[18] , \ScanLink234[17] , 
        \ScanLink234[16] , \ScanLink234[15] , \ScanLink234[14] , 
        \ScanLink234[13] , \ScanLink234[12] , \ScanLink234[11] , 
        \ScanLink234[10] , \ScanLink234[9] , \ScanLink234[8] , 
        \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , \ScanLink234[4] , 
        \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , \ScanLink234[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB10[31] , \wRegInB10[30] , \wRegInB10[29] , 
        \wRegInB10[28] , \wRegInB10[27] , \wRegInB10[26] , \wRegInB10[25] , 
        \wRegInB10[24] , \wRegInB10[23] , \wRegInB10[22] , \wRegInB10[21] , 
        \wRegInB10[20] , \wRegInB10[19] , \wRegInB10[18] , \wRegInB10[17] , 
        \wRegInB10[16] , \wRegInB10[15] , \wRegInB10[14] , \wRegInB10[13] , 
        \wRegInB10[12] , \wRegInB10[11] , \wRegInB10[10] , \wRegInB10[9] , 
        \wRegInB10[8] , \wRegInB10[7] , \wRegInB10[6] , \wRegInB10[5] , 
        \wRegInB10[4] , \wRegInB10[3] , \wRegInB10[2] , \wRegInB10[1] , 
        \wRegInB10[0] }), .Out({\wBIn10[31] , \wBIn10[30] , \wBIn10[29] , 
        \wBIn10[28] , \wBIn10[27] , \wBIn10[26] , \wBIn10[25] , \wBIn10[24] , 
        \wBIn10[23] , \wBIn10[22] , \wBIn10[21] , \wBIn10[20] , \wBIn10[19] , 
        \wBIn10[18] , \wBIn10[17] , \wBIn10[16] , \wBIn10[15] , \wBIn10[14] , 
        \wBIn10[13] , \wBIn10[12] , \wBIn10[11] , \wBIn10[10] , \wBIn10[9] , 
        \wBIn10[8] , \wBIn10[7] , \wBIn10[6] , \wBIn10[5] , \wBIn10[4] , 
        \wBIn10[3] , \wBIn10[2] , \wBIn10[1] , \wBIn10[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_104 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink105[31] , \ScanLink105[30] , \ScanLink105[29] , 
        \ScanLink105[28] , \ScanLink105[27] , \ScanLink105[26] , 
        \ScanLink105[25] , \ScanLink105[24] , \ScanLink105[23] , 
        \ScanLink105[22] , \ScanLink105[21] , \ScanLink105[20] , 
        \ScanLink105[19] , \ScanLink105[18] , \ScanLink105[17] , 
        \ScanLink105[16] , \ScanLink105[15] , \ScanLink105[14] , 
        \ScanLink105[13] , \ScanLink105[12] , \ScanLink105[11] , 
        \ScanLink105[10] , \ScanLink105[9] , \ScanLink105[8] , 
        \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , \ScanLink105[4] , 
        \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , \ScanLink105[0] 
        }), .ScanOut({\ScanLink104[31] , \ScanLink104[30] , \ScanLink104[29] , 
        \ScanLink104[28] , \ScanLink104[27] , \ScanLink104[26] , 
        \ScanLink104[25] , \ScanLink104[24] , \ScanLink104[23] , 
        \ScanLink104[22] , \ScanLink104[21] , \ScanLink104[20] , 
        \ScanLink104[19] , \ScanLink104[18] , \ScanLink104[17] , 
        \ScanLink104[16] , \ScanLink104[15] , \ScanLink104[14] , 
        \ScanLink104[13] , \ScanLink104[12] , \ScanLink104[11] , 
        \ScanLink104[10] , \ScanLink104[9] , \ScanLink104[8] , 
        \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , \ScanLink104[4] , 
        \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , \ScanLink104[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB75[31] , \wRegInB75[30] , \wRegInB75[29] , 
        \wRegInB75[28] , \wRegInB75[27] , \wRegInB75[26] , \wRegInB75[25] , 
        \wRegInB75[24] , \wRegInB75[23] , \wRegInB75[22] , \wRegInB75[21] , 
        \wRegInB75[20] , \wRegInB75[19] , \wRegInB75[18] , \wRegInB75[17] , 
        \wRegInB75[16] , \wRegInB75[15] , \wRegInB75[14] , \wRegInB75[13] , 
        \wRegInB75[12] , \wRegInB75[11] , \wRegInB75[10] , \wRegInB75[9] , 
        \wRegInB75[8] , \wRegInB75[7] , \wRegInB75[6] , \wRegInB75[5] , 
        \wRegInB75[4] , \wRegInB75[3] , \wRegInB75[2] , \wRegInB75[1] , 
        \wRegInB75[0] }), .Out({\wBIn75[31] , \wBIn75[30] , \wBIn75[29] , 
        \wBIn75[28] , \wBIn75[27] , \wBIn75[26] , \wBIn75[25] , \wBIn75[24] , 
        \wBIn75[23] , \wBIn75[22] , \wBIn75[21] , \wBIn75[20] , \wBIn75[19] , 
        \wBIn75[18] , \wBIn75[17] , \wBIn75[16] , \wBIn75[15] , \wBIn75[14] , 
        \wBIn75[13] , \wBIn75[12] , \wBIn75[11] , \wBIn75[10] , \wBIn75[9] , 
        \wBIn75[8] , \wBIn75[7] , \wBIn75[6] , \wBIn75[5] , \wBIn75[4] , 
        \wBIn75[3] , \wBIn75[2] , \wBIn75[1] , \wBIn75[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_54 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink55[31] , \ScanLink55[30] , \ScanLink55[29] , 
        \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , \ScanLink55[25] , 
        \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , \ScanLink55[21] , 
        \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , \ScanLink55[17] , 
        \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , \ScanLink55[13] , 
        \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , \ScanLink55[9] , 
        \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , \ScanLink55[5] , 
        \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , \ScanLink55[1] , 
        \ScanLink55[0] }), .ScanOut({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB100[31] , \wRegInB100[30] , 
        \wRegInB100[29] , \wRegInB100[28] , \wRegInB100[27] , \wRegInB100[26] , 
        \wRegInB100[25] , \wRegInB100[24] , \wRegInB100[23] , \wRegInB100[22] , 
        \wRegInB100[21] , \wRegInB100[20] , \wRegInB100[19] , \wRegInB100[18] , 
        \wRegInB100[17] , \wRegInB100[16] , \wRegInB100[15] , \wRegInB100[14] , 
        \wRegInB100[13] , \wRegInB100[12] , \wRegInB100[11] , \wRegInB100[10] , 
        \wRegInB100[9] , \wRegInB100[8] , \wRegInB100[7] , \wRegInB100[6] , 
        \wRegInB100[5] , \wRegInB100[4] , \wRegInB100[3] , \wRegInB100[2] , 
        \wRegInB100[1] , \wRegInB100[0] }), .Out({\wBIn100[31] , \wBIn100[30] , 
        \wBIn100[29] , \wBIn100[28] , \wBIn100[27] , \wBIn100[26] , 
        \wBIn100[25] , \wBIn100[24] , \wBIn100[23] , \wBIn100[22] , 
        \wBIn100[21] , \wBIn100[20] , \wBIn100[19] , \wBIn100[18] , 
        \wBIn100[17] , \wBIn100[16] , \wBIn100[15] , \wBIn100[14] , 
        \wBIn100[13] , \wBIn100[12] , \wBIn100[11] , \wBIn100[10] , 
        \wBIn100[9] , \wBIn100[8] , \wBIn100[7] , \wBIn100[6] , \wBIn100[5] , 
        \wBIn100[4] , \wBIn100[3] , \wBIn100[2] , \wBIn100[1] , \wBIn100[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn9[31] , 
        \wAIn9[30] , \wAIn9[29] , \wAIn9[28] , \wAIn9[27] , \wAIn9[26] , 
        \wAIn9[25] , \wAIn9[24] , \wAIn9[23] , \wAIn9[22] , \wAIn9[21] , 
        \wAIn9[20] , \wAIn9[19] , \wAIn9[18] , \wAIn9[17] , \wAIn9[16] , 
        \wAIn9[15] , \wAIn9[14] , \wAIn9[13] , \wAIn9[12] , \wAIn9[11] , 
        \wAIn9[10] , \wAIn9[9] , \wAIn9[8] , \wAIn9[7] , \wAIn9[6] , 
        \wAIn9[5] , \wAIn9[4] , \wAIn9[3] , \wAIn9[2] , \wAIn9[1] , \wAIn9[0] 
        }), .BIn({\wBIn9[31] , \wBIn9[30] , \wBIn9[29] , \wBIn9[28] , 
        \wBIn9[27] , \wBIn9[26] , \wBIn9[25] , \wBIn9[24] , \wBIn9[23] , 
        \wBIn9[22] , \wBIn9[21] , \wBIn9[20] , \wBIn9[19] , \wBIn9[18] , 
        \wBIn9[17] , \wBIn9[16] , \wBIn9[15] , \wBIn9[14] , \wBIn9[13] , 
        \wBIn9[12] , \wBIn9[11] , \wBIn9[10] , \wBIn9[9] , \wBIn9[8] , 
        \wBIn9[7] , \wBIn9[6] , \wBIn9[5] , \wBIn9[4] , \wBIn9[3] , \wBIn9[2] , 
        \wBIn9[1] , \wBIn9[0] }), .HiOut({\wBMid8[31] , \wBMid8[30] , 
        \wBMid8[29] , \wBMid8[28] , \wBMid8[27] , \wBMid8[26] , \wBMid8[25] , 
        \wBMid8[24] , \wBMid8[23] , \wBMid8[22] , \wBMid8[21] , \wBMid8[20] , 
        \wBMid8[19] , \wBMid8[18] , \wBMid8[17] , \wBMid8[16] , \wBMid8[15] , 
        \wBMid8[14] , \wBMid8[13] , \wBMid8[12] , \wBMid8[11] , \wBMid8[10] , 
        \wBMid8[9] , \wBMid8[8] , \wBMid8[7] , \wBMid8[6] , \wBMid8[5] , 
        \wBMid8[4] , \wBMid8[3] , \wBMid8[2] , \wBMid8[1] , \wBMid8[0] }), 
        .LoOut({\wAMid9[31] , \wAMid9[30] , \wAMid9[29] , \wAMid9[28] , 
        \wAMid9[27] , \wAMid9[26] , \wAMid9[25] , \wAMid9[24] , \wAMid9[23] , 
        \wAMid9[22] , \wAMid9[21] , \wAMid9[20] , \wAMid9[19] , \wAMid9[18] , 
        \wAMid9[17] , \wAMid9[16] , \wAMid9[15] , \wAMid9[14] , \wAMid9[13] , 
        \wAMid9[12] , \wAMid9[11] , \wAMid9[10] , \wAMid9[9] , \wAMid9[8] , 
        \wAMid9[7] , \wAMid9[6] , \wAMid9[5] , \wAMid9[4] , \wAMid9[3] , 
        \wAMid9[2] , \wAMid9[1] , \wAMid9[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn11[31] , \wAIn11[30] , \wAIn11[29] , \wAIn11[28] , \wAIn11[27] , 
        \wAIn11[26] , \wAIn11[25] , \wAIn11[24] , \wAIn11[23] , \wAIn11[22] , 
        \wAIn11[21] , \wAIn11[20] , \wAIn11[19] , \wAIn11[18] , \wAIn11[17] , 
        \wAIn11[16] , \wAIn11[15] , \wAIn11[14] , \wAIn11[13] , \wAIn11[12] , 
        \wAIn11[11] , \wAIn11[10] , \wAIn11[9] , \wAIn11[8] , \wAIn11[7] , 
        \wAIn11[6] , \wAIn11[5] , \wAIn11[4] , \wAIn11[3] , \wAIn11[2] , 
        \wAIn11[1] , \wAIn11[0] }), .BIn({\wBIn11[31] , \wBIn11[30] , 
        \wBIn11[29] , \wBIn11[28] , \wBIn11[27] , \wBIn11[26] , \wBIn11[25] , 
        \wBIn11[24] , \wBIn11[23] , \wBIn11[22] , \wBIn11[21] , \wBIn11[20] , 
        \wBIn11[19] , \wBIn11[18] , \wBIn11[17] , \wBIn11[16] , \wBIn11[15] , 
        \wBIn11[14] , \wBIn11[13] , \wBIn11[12] , \wBIn11[11] , \wBIn11[10] , 
        \wBIn11[9] , \wBIn11[8] , \wBIn11[7] , \wBIn11[6] , \wBIn11[5] , 
        \wBIn11[4] , \wBIn11[3] , \wBIn11[2] , \wBIn11[1] , \wBIn11[0] }), 
        .HiOut({\wBMid10[31] , \wBMid10[30] , \wBMid10[29] , \wBMid10[28] , 
        \wBMid10[27] , \wBMid10[26] , \wBMid10[25] , \wBMid10[24] , 
        \wBMid10[23] , \wBMid10[22] , \wBMid10[21] , \wBMid10[20] , 
        \wBMid10[19] , \wBMid10[18] , \wBMid10[17] , \wBMid10[16] , 
        \wBMid10[15] , \wBMid10[14] , \wBMid10[13] , \wBMid10[12] , 
        \wBMid10[11] , \wBMid10[10] , \wBMid10[9] , \wBMid10[8] , \wBMid10[7] , 
        \wBMid10[6] , \wBMid10[5] , \wBMid10[4] , \wBMid10[3] , \wBMid10[2] , 
        \wBMid10[1] , \wBMid10[0] }), .LoOut({\wAMid11[31] , \wAMid11[30] , 
        \wAMid11[29] , \wAMid11[28] , \wAMid11[27] , \wAMid11[26] , 
        \wAMid11[25] , \wAMid11[24] , \wAMid11[23] , \wAMid11[22] , 
        \wAMid11[21] , \wAMid11[20] , \wAMid11[19] , \wAMid11[18] , 
        \wAMid11[17] , \wAMid11[16] , \wAMid11[15] , \wAMid11[14] , 
        \wAMid11[13] , \wAMid11[12] , \wAMid11[11] , \wAMid11[10] , 
        \wAMid11[9] , \wAMid11[8] , \wAMid11[7] , \wAMid11[6] , \wAMid11[5] , 
        \wAMid11[4] , \wAMid11[3] , \wAMid11[2] , \wAMid11[1] , \wAMid11[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn43[31] , \wAIn43[30] , \wAIn43[29] , \wAIn43[28] , \wAIn43[27] , 
        \wAIn43[26] , \wAIn43[25] , \wAIn43[24] , \wAIn43[23] , \wAIn43[22] , 
        \wAIn43[21] , \wAIn43[20] , \wAIn43[19] , \wAIn43[18] , \wAIn43[17] , 
        \wAIn43[16] , \wAIn43[15] , \wAIn43[14] , \wAIn43[13] , \wAIn43[12] , 
        \wAIn43[11] , \wAIn43[10] , \wAIn43[9] , \wAIn43[8] , \wAIn43[7] , 
        \wAIn43[6] , \wAIn43[5] , \wAIn43[4] , \wAIn43[3] , \wAIn43[2] , 
        \wAIn43[1] , \wAIn43[0] }), .BIn({\wBIn43[31] , \wBIn43[30] , 
        \wBIn43[29] , \wBIn43[28] , \wBIn43[27] , \wBIn43[26] , \wBIn43[25] , 
        \wBIn43[24] , \wBIn43[23] , \wBIn43[22] , \wBIn43[21] , \wBIn43[20] , 
        \wBIn43[19] , \wBIn43[18] , \wBIn43[17] , \wBIn43[16] , \wBIn43[15] , 
        \wBIn43[14] , \wBIn43[13] , \wBIn43[12] , \wBIn43[11] , \wBIn43[10] , 
        \wBIn43[9] , \wBIn43[8] , \wBIn43[7] , \wBIn43[6] , \wBIn43[5] , 
        \wBIn43[4] , \wBIn43[3] , \wBIn43[2] , \wBIn43[1] , \wBIn43[0] }), 
        .HiOut({\wBMid42[31] , \wBMid42[30] , \wBMid42[29] , \wBMid42[28] , 
        \wBMid42[27] , \wBMid42[26] , \wBMid42[25] , \wBMid42[24] , 
        \wBMid42[23] , \wBMid42[22] , \wBMid42[21] , \wBMid42[20] , 
        \wBMid42[19] , \wBMid42[18] , \wBMid42[17] , \wBMid42[16] , 
        \wBMid42[15] , \wBMid42[14] , \wBMid42[13] , \wBMid42[12] , 
        \wBMid42[11] , \wBMid42[10] , \wBMid42[9] , \wBMid42[8] , \wBMid42[7] , 
        \wBMid42[6] , \wBMid42[5] , \wBMid42[4] , \wBMid42[3] , \wBMid42[2] , 
        \wBMid42[1] , \wBMid42[0] }), .LoOut({\wAMid43[31] , \wAMid43[30] , 
        \wAMid43[29] , \wAMid43[28] , \wAMid43[27] , \wAMid43[26] , 
        \wAMid43[25] , \wAMid43[24] , \wAMid43[23] , \wAMid43[22] , 
        \wAMid43[21] , \wAMid43[20] , \wAMid43[19] , \wAMid43[18] , 
        \wAMid43[17] , \wAMid43[16] , \wAMid43[15] , \wAMid43[14] , 
        \wAMid43[13] , \wAMid43[12] , \wAMid43[11] , \wAMid43[10] , 
        \wAMid43[9] , \wAMid43[8] , \wAMid43[7] , \wAMid43[6] , \wAMid43[5] , 
        \wAMid43[4] , \wAMid43[3] , \wAMid43[2] , \wAMid43[1] , \wAMid43[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn64[31] , \wAIn64[30] , \wAIn64[29] , \wAIn64[28] , \wAIn64[27] , 
        \wAIn64[26] , \wAIn64[25] , \wAIn64[24] , \wAIn64[23] , \wAIn64[22] , 
        \wAIn64[21] , \wAIn64[20] , \wAIn64[19] , \wAIn64[18] , \wAIn64[17] , 
        \wAIn64[16] , \wAIn64[15] , \wAIn64[14] , \wAIn64[13] , \wAIn64[12] , 
        \wAIn64[11] , \wAIn64[10] , \wAIn64[9] , \wAIn64[8] , \wAIn64[7] , 
        \wAIn64[6] , \wAIn64[5] , \wAIn64[4] , \wAIn64[3] , \wAIn64[2] , 
        \wAIn64[1] , \wAIn64[0] }), .BIn({\wBIn64[31] , \wBIn64[30] , 
        \wBIn64[29] , \wBIn64[28] , \wBIn64[27] , \wBIn64[26] , \wBIn64[25] , 
        \wBIn64[24] , \wBIn64[23] , \wBIn64[22] , \wBIn64[21] , \wBIn64[20] , 
        \wBIn64[19] , \wBIn64[18] , \wBIn64[17] , \wBIn64[16] , \wBIn64[15] , 
        \wBIn64[14] , \wBIn64[13] , \wBIn64[12] , \wBIn64[11] , \wBIn64[10] , 
        \wBIn64[9] , \wBIn64[8] , \wBIn64[7] , \wBIn64[6] , \wBIn64[5] , 
        \wBIn64[4] , \wBIn64[3] , \wBIn64[2] , \wBIn64[1] , \wBIn64[0] }), 
        .HiOut({\wBMid63[31] , \wBMid63[30] , \wBMid63[29] , \wBMid63[28] , 
        \wBMid63[27] , \wBMid63[26] , \wBMid63[25] , \wBMid63[24] , 
        \wBMid63[23] , \wBMid63[22] , \wBMid63[21] , \wBMid63[20] , 
        \wBMid63[19] , \wBMid63[18] , \wBMid63[17] , \wBMid63[16] , 
        \wBMid63[15] , \wBMid63[14] , \wBMid63[13] , \wBMid63[12] , 
        \wBMid63[11] , \wBMid63[10] , \wBMid63[9] , \wBMid63[8] , \wBMid63[7] , 
        \wBMid63[6] , \wBMid63[5] , \wBMid63[4] , \wBMid63[3] , \wBMid63[2] , 
        \wBMid63[1] , \wBMid63[0] }), .LoOut({\wAMid64[31] , \wAMid64[30] , 
        \wAMid64[29] , \wAMid64[28] , \wAMid64[27] , \wAMid64[26] , 
        \wAMid64[25] , \wAMid64[24] , \wAMid64[23] , \wAMid64[22] , 
        \wAMid64[21] , \wAMid64[20] , \wAMid64[19] , \wAMid64[18] , 
        \wAMid64[17] , \wAMid64[16] , \wAMid64[15] , \wAMid64[14] , 
        \wAMid64[13] , \wAMid64[12] , \wAMid64[11] , \wAMid64[10] , 
        \wAMid64[9] , \wAMid64[8] , \wAMid64[7] , \wAMid64[6] , \wAMid64[5] , 
        \wAMid64[4] , \wAMid64[3] , \wAMid64[2] , \wAMid64[1] , \wAMid64[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn81[31] , \wAIn81[30] , \wAIn81[29] , \wAIn81[28] , \wAIn81[27] , 
        \wAIn81[26] , \wAIn81[25] , \wAIn81[24] , \wAIn81[23] , \wAIn81[22] , 
        \wAIn81[21] , \wAIn81[20] , \wAIn81[19] , \wAIn81[18] , \wAIn81[17] , 
        \wAIn81[16] , \wAIn81[15] , \wAIn81[14] , \wAIn81[13] , \wAIn81[12] , 
        \wAIn81[11] , \wAIn81[10] , \wAIn81[9] , \wAIn81[8] , \wAIn81[7] , 
        \wAIn81[6] , \wAIn81[5] , \wAIn81[4] , \wAIn81[3] , \wAIn81[2] , 
        \wAIn81[1] , \wAIn81[0] }), .BIn({\wBIn81[31] , \wBIn81[30] , 
        \wBIn81[29] , \wBIn81[28] , \wBIn81[27] , \wBIn81[26] , \wBIn81[25] , 
        \wBIn81[24] , \wBIn81[23] , \wBIn81[22] , \wBIn81[21] , \wBIn81[20] , 
        \wBIn81[19] , \wBIn81[18] , \wBIn81[17] , \wBIn81[16] , \wBIn81[15] , 
        \wBIn81[14] , \wBIn81[13] , \wBIn81[12] , \wBIn81[11] , \wBIn81[10] , 
        \wBIn81[9] , \wBIn81[8] , \wBIn81[7] , \wBIn81[6] , \wBIn81[5] , 
        \wBIn81[4] , \wBIn81[3] , \wBIn81[2] , \wBIn81[1] , \wBIn81[0] }), 
        .HiOut({\wBMid80[31] , \wBMid80[30] , \wBMid80[29] , \wBMid80[28] , 
        \wBMid80[27] , \wBMid80[26] , \wBMid80[25] , \wBMid80[24] , 
        \wBMid80[23] , \wBMid80[22] , \wBMid80[21] , \wBMid80[20] , 
        \wBMid80[19] , \wBMid80[18] , \wBMid80[17] , \wBMid80[16] , 
        \wBMid80[15] , \wBMid80[14] , \wBMid80[13] , \wBMid80[12] , 
        \wBMid80[11] , \wBMid80[10] , \wBMid80[9] , \wBMid80[8] , \wBMid80[7] , 
        \wBMid80[6] , \wBMid80[5] , \wBMid80[4] , \wBMid80[3] , \wBMid80[2] , 
        \wBMid80[1] , \wBMid80[0] }), .LoOut({\wAMid81[31] , \wAMid81[30] , 
        \wAMid81[29] , \wAMid81[28] , \wAMid81[27] , \wAMid81[26] , 
        \wAMid81[25] , \wAMid81[24] , \wAMid81[23] , \wAMid81[22] , 
        \wAMid81[21] , \wAMid81[20] , \wAMid81[19] , \wAMid81[18] , 
        \wAMid81[17] , \wAMid81[16] , \wAMid81[15] , \wAMid81[14] , 
        \wAMid81[13] , \wAMid81[12] , \wAMid81[11] , \wAMid81[10] , 
        \wAMid81[9] , \wAMid81[8] , \wAMid81[7] , \wAMid81[6] , \wAMid81[5] , 
        \wAMid81[4] , \wAMid81[3] , \wAMid81[2] , \wAMid81[1] , \wAMid81[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid96[31] , \wAMid96[30] , \wAMid96[29] , \wAMid96[28] , 
        \wAMid96[27] , \wAMid96[26] , \wAMid96[25] , \wAMid96[24] , 
        \wAMid96[23] , \wAMid96[22] , \wAMid96[21] , \wAMid96[20] , 
        \wAMid96[19] , \wAMid96[18] , \wAMid96[17] , \wAMid96[16] , 
        \wAMid96[15] , \wAMid96[14] , \wAMid96[13] , \wAMid96[12] , 
        \wAMid96[11] , \wAMid96[10] , \wAMid96[9] , \wAMid96[8] , \wAMid96[7] , 
        \wAMid96[6] , \wAMid96[5] , \wAMid96[4] , \wAMid96[3] , \wAMid96[2] , 
        \wAMid96[1] , \wAMid96[0] }), .BIn({\wBMid96[31] , \wBMid96[30] , 
        \wBMid96[29] , \wBMid96[28] , \wBMid96[27] , \wBMid96[26] , 
        \wBMid96[25] , \wBMid96[24] , \wBMid96[23] , \wBMid96[22] , 
        \wBMid96[21] , \wBMid96[20] , \wBMid96[19] , \wBMid96[18] , 
        \wBMid96[17] , \wBMid96[16] , \wBMid96[15] , \wBMid96[14] , 
        \wBMid96[13] , \wBMid96[12] , \wBMid96[11] , \wBMid96[10] , 
        \wBMid96[9] , \wBMid96[8] , \wBMid96[7] , \wBMid96[6] , \wBMid96[5] , 
        \wBMid96[4] , \wBMid96[3] , \wBMid96[2] , \wBMid96[1] , \wBMid96[0] }), 
        .HiOut({\wRegInB96[31] , \wRegInB96[30] , \wRegInB96[29] , 
        \wRegInB96[28] , \wRegInB96[27] , \wRegInB96[26] , \wRegInB96[25] , 
        \wRegInB96[24] , \wRegInB96[23] , \wRegInB96[22] , \wRegInB96[21] , 
        \wRegInB96[20] , \wRegInB96[19] , \wRegInB96[18] , \wRegInB96[17] , 
        \wRegInB96[16] , \wRegInB96[15] , \wRegInB96[14] , \wRegInB96[13] , 
        \wRegInB96[12] , \wRegInB96[11] , \wRegInB96[10] , \wRegInB96[9] , 
        \wRegInB96[8] , \wRegInB96[7] , \wRegInB96[6] , \wRegInB96[5] , 
        \wRegInB96[4] , \wRegInB96[3] , \wRegInB96[2] , \wRegInB96[1] , 
        \wRegInB96[0] }), .LoOut({\wRegInA97[31] , \wRegInA97[30] , 
        \wRegInA97[29] , \wRegInA97[28] , \wRegInA97[27] , \wRegInA97[26] , 
        \wRegInA97[25] , \wRegInA97[24] , \wRegInA97[23] , \wRegInA97[22] , 
        \wRegInA97[21] , \wRegInA97[20] , \wRegInA97[19] , \wRegInA97[18] , 
        \wRegInA97[17] , \wRegInA97[16] , \wRegInA97[15] , \wRegInA97[14] , 
        \wRegInA97[13] , \wRegInA97[12] , \wRegInA97[11] , \wRegInA97[10] , 
        \wRegInA97[9] , \wRegInA97[8] , \wRegInA97[7] , \wRegInA97[6] , 
        \wRegInA97[5] , \wRegInA97[4] , \wRegInA97[3] , \wRegInA97[2] , 
        \wRegInA97[1] , \wRegInA97[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn114[31] , \wAIn114[30] , \wAIn114[29] , \wAIn114[28] , 
        \wAIn114[27] , \wAIn114[26] , \wAIn114[25] , \wAIn114[24] , 
        \wAIn114[23] , \wAIn114[22] , \wAIn114[21] , \wAIn114[20] , 
        \wAIn114[19] , \wAIn114[18] , \wAIn114[17] , \wAIn114[16] , 
        \wAIn114[15] , \wAIn114[14] , \wAIn114[13] , \wAIn114[12] , 
        \wAIn114[11] , \wAIn114[10] , \wAIn114[9] , \wAIn114[8] , \wAIn114[7] , 
        \wAIn114[6] , \wAIn114[5] , \wAIn114[4] , \wAIn114[3] , \wAIn114[2] , 
        \wAIn114[1] , \wAIn114[0] }), .BIn({\wBIn114[31] , \wBIn114[30] , 
        \wBIn114[29] , \wBIn114[28] , \wBIn114[27] , \wBIn114[26] , 
        \wBIn114[25] , \wBIn114[24] , \wBIn114[23] , \wBIn114[22] , 
        \wBIn114[21] , \wBIn114[20] , \wBIn114[19] , \wBIn114[18] , 
        \wBIn114[17] , \wBIn114[16] , \wBIn114[15] , \wBIn114[14] , 
        \wBIn114[13] , \wBIn114[12] , \wBIn114[11] , \wBIn114[10] , 
        \wBIn114[9] , \wBIn114[8] , \wBIn114[7] , \wBIn114[6] , \wBIn114[5] , 
        \wBIn114[4] , \wBIn114[3] , \wBIn114[2] , \wBIn114[1] , \wBIn114[0] }), 
        .HiOut({\wBMid113[31] , \wBMid113[30] , \wBMid113[29] , \wBMid113[28] , 
        \wBMid113[27] , \wBMid113[26] , \wBMid113[25] , \wBMid113[24] , 
        \wBMid113[23] , \wBMid113[22] , \wBMid113[21] , \wBMid113[20] , 
        \wBMid113[19] , \wBMid113[18] , \wBMid113[17] , \wBMid113[16] , 
        \wBMid113[15] , \wBMid113[14] , \wBMid113[13] , \wBMid113[12] , 
        \wBMid113[11] , \wBMid113[10] , \wBMid113[9] , \wBMid113[8] , 
        \wBMid113[7] , \wBMid113[6] , \wBMid113[5] , \wBMid113[4] , 
        \wBMid113[3] , \wBMid113[2] , \wBMid113[1] , \wBMid113[0] }), .LoOut({
        \wAMid114[31] , \wAMid114[30] , \wAMid114[29] , \wAMid114[28] , 
        \wAMid114[27] , \wAMid114[26] , \wAMid114[25] , \wAMid114[24] , 
        \wAMid114[23] , \wAMid114[22] , \wAMid114[21] , \wAMid114[20] , 
        \wAMid114[19] , \wAMid114[18] , \wAMid114[17] , \wAMid114[16] , 
        \wAMid114[15] , \wAMid114[14] , \wAMid114[13] , \wAMid114[12] , 
        \wAMid114[11] , \wAMid114[10] , \wAMid114[9] , \wAMid114[8] , 
        \wAMid114[7] , \wAMid114[6] , \wAMid114[5] , \wAMid114[4] , 
        \wAMid114[3] , \wAMid114[2] , \wAMid114[1] , \wAMid114[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_251 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink252[31] , \ScanLink252[30] , \ScanLink252[29] , 
        \ScanLink252[28] , \ScanLink252[27] , \ScanLink252[26] , 
        \ScanLink252[25] , \ScanLink252[24] , \ScanLink252[23] , 
        \ScanLink252[22] , \ScanLink252[21] , \ScanLink252[20] , 
        \ScanLink252[19] , \ScanLink252[18] , \ScanLink252[17] , 
        \ScanLink252[16] , \ScanLink252[15] , \ScanLink252[14] , 
        \ScanLink252[13] , \ScanLink252[12] , \ScanLink252[11] , 
        \ScanLink252[10] , \ScanLink252[9] , \ScanLink252[8] , 
        \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , \ScanLink252[4] , 
        \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , \ScanLink252[0] 
        }), .ScanOut({\ScanLink251[31] , \ScanLink251[30] , \ScanLink251[29] , 
        \ScanLink251[28] , \ScanLink251[27] , \ScanLink251[26] , 
        \ScanLink251[25] , \ScanLink251[24] , \ScanLink251[23] , 
        \ScanLink251[22] , \ScanLink251[21] , \ScanLink251[20] , 
        \ScanLink251[19] , \ScanLink251[18] , \ScanLink251[17] , 
        \ScanLink251[16] , \ScanLink251[15] , \ScanLink251[14] , 
        \ScanLink251[13] , \ScanLink251[12] , \ScanLink251[11] , 
        \ScanLink251[10] , \ScanLink251[9] , \ScanLink251[8] , 
        \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , \ScanLink251[4] , 
        \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , \ScanLink251[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA2[31] , \wRegInA2[30] , \wRegInA2[29] , \wRegInA2[28] , 
        \wRegInA2[27] , \wRegInA2[26] , \wRegInA2[25] , \wRegInA2[24] , 
        \wRegInA2[23] , \wRegInA2[22] , \wRegInA2[21] , \wRegInA2[20] , 
        \wRegInA2[19] , \wRegInA2[18] , \wRegInA2[17] , \wRegInA2[16] , 
        \wRegInA2[15] , \wRegInA2[14] , \wRegInA2[13] , \wRegInA2[12] , 
        \wRegInA2[11] , \wRegInA2[10] , \wRegInA2[9] , \wRegInA2[8] , 
        \wRegInA2[7] , \wRegInA2[6] , \wRegInA2[5] , \wRegInA2[4] , 
        \wRegInA2[3] , \wRegInA2[2] , \wRegInA2[1] , \wRegInA2[0] }), .Out({
        \wAIn2[31] , \wAIn2[30] , \wAIn2[29] , \wAIn2[28] , \wAIn2[27] , 
        \wAIn2[26] , \wAIn2[25] , \wAIn2[24] , \wAIn2[23] , \wAIn2[22] , 
        \wAIn2[21] , \wAIn2[20] , \wAIn2[19] , \wAIn2[18] , \wAIn2[17] , 
        \wAIn2[16] , \wAIn2[15] , \wAIn2[14] , \wAIn2[13] , \wAIn2[12] , 
        \wAIn2[11] , \wAIn2[10] , \wAIn2[9] , \wAIn2[8] , \wAIn2[7] , 
        \wAIn2[6] , \wAIn2[5] , \wAIn2[4] , \wAIn2[3] , \wAIn2[2] , \wAIn2[1] , 
        \wAIn2[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_218 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink219[31] , \ScanLink219[30] , \ScanLink219[29] , 
        \ScanLink219[28] , \ScanLink219[27] , \ScanLink219[26] , 
        \ScanLink219[25] , \ScanLink219[24] , \ScanLink219[23] , 
        \ScanLink219[22] , \ScanLink219[21] , \ScanLink219[20] , 
        \ScanLink219[19] , \ScanLink219[18] , \ScanLink219[17] , 
        \ScanLink219[16] , \ScanLink219[15] , \ScanLink219[14] , 
        \ScanLink219[13] , \ScanLink219[12] , \ScanLink219[11] , 
        \ScanLink219[10] , \ScanLink219[9] , \ScanLink219[8] , 
        \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , \ScanLink219[4] , 
        \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , \ScanLink219[0] 
        }), .ScanOut({\ScanLink218[31] , \ScanLink218[30] , \ScanLink218[29] , 
        \ScanLink218[28] , \ScanLink218[27] , \ScanLink218[26] , 
        \ScanLink218[25] , \ScanLink218[24] , \ScanLink218[23] , 
        \ScanLink218[22] , \ScanLink218[21] , \ScanLink218[20] , 
        \ScanLink218[19] , \ScanLink218[18] , \ScanLink218[17] , 
        \ScanLink218[16] , \ScanLink218[15] , \ScanLink218[14] , 
        \ScanLink218[13] , \ScanLink218[12] , \ScanLink218[11] , 
        \ScanLink218[10] , \ScanLink218[9] , \ScanLink218[8] , 
        \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , \ScanLink218[4] , 
        \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , \ScanLink218[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB18[31] , \wRegInB18[30] , \wRegInB18[29] , 
        \wRegInB18[28] , \wRegInB18[27] , \wRegInB18[26] , \wRegInB18[25] , 
        \wRegInB18[24] , \wRegInB18[23] , \wRegInB18[22] , \wRegInB18[21] , 
        \wRegInB18[20] , \wRegInB18[19] , \wRegInB18[18] , \wRegInB18[17] , 
        \wRegInB18[16] , \wRegInB18[15] , \wRegInB18[14] , \wRegInB18[13] , 
        \wRegInB18[12] , \wRegInB18[11] , \wRegInB18[10] , \wRegInB18[9] , 
        \wRegInB18[8] , \wRegInB18[7] , \wRegInB18[6] , \wRegInB18[5] , 
        \wRegInB18[4] , \wRegInB18[3] , \wRegInB18[2] , \wRegInB18[1] , 
        \wRegInB18[0] }), .Out({\wBIn18[31] , \wBIn18[30] , \wBIn18[29] , 
        \wBIn18[28] , \wBIn18[27] , \wBIn18[26] , \wBIn18[25] , \wBIn18[24] , 
        \wBIn18[23] , \wBIn18[22] , \wBIn18[21] , \wBIn18[20] , \wBIn18[19] , 
        \wBIn18[18] , \wBIn18[17] , \wBIn18[16] , \wBIn18[15] , \wBIn18[14] , 
        \wBIn18[13] , \wBIn18[12] , \wBIn18[11] , \wBIn18[10] , \wBIn18[9] , 
        \wBIn18[8] , \wBIn18[7] , \wBIn18[6] , \wBIn18[5] , \wBIn18[4] , 
        \wBIn18[3] , \wBIn18[2] , \wBIn18[1] , \wBIn18[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_184 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink185[31] , \ScanLink185[30] , \ScanLink185[29] , 
        \ScanLink185[28] , \ScanLink185[27] , \ScanLink185[26] , 
        \ScanLink185[25] , \ScanLink185[24] , \ScanLink185[23] , 
        \ScanLink185[22] , \ScanLink185[21] , \ScanLink185[20] , 
        \ScanLink185[19] , \ScanLink185[18] , \ScanLink185[17] , 
        \ScanLink185[16] , \ScanLink185[15] , \ScanLink185[14] , 
        \ScanLink185[13] , \ScanLink185[12] , \ScanLink185[11] , 
        \ScanLink185[10] , \ScanLink185[9] , \ScanLink185[8] , 
        \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , \ScanLink185[4] , 
        \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , \ScanLink185[0] 
        }), .ScanOut({\ScanLink184[31] , \ScanLink184[30] , \ScanLink184[29] , 
        \ScanLink184[28] , \ScanLink184[27] , \ScanLink184[26] , 
        \ScanLink184[25] , \ScanLink184[24] , \ScanLink184[23] , 
        \ScanLink184[22] , \ScanLink184[21] , \ScanLink184[20] , 
        \ScanLink184[19] , \ScanLink184[18] , \ScanLink184[17] , 
        \ScanLink184[16] , \ScanLink184[15] , \ScanLink184[14] , 
        \ScanLink184[13] , \ScanLink184[12] , \ScanLink184[11] , 
        \ScanLink184[10] , \ScanLink184[9] , \ScanLink184[8] , 
        \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , \ScanLink184[4] , 
        \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , \ScanLink184[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB35[31] , \wRegInB35[30] , \wRegInB35[29] , 
        \wRegInB35[28] , \wRegInB35[27] , \wRegInB35[26] , \wRegInB35[25] , 
        \wRegInB35[24] , \wRegInB35[23] , \wRegInB35[22] , \wRegInB35[21] , 
        \wRegInB35[20] , \wRegInB35[19] , \wRegInB35[18] , \wRegInB35[17] , 
        \wRegInB35[16] , \wRegInB35[15] , \wRegInB35[14] , \wRegInB35[13] , 
        \wRegInB35[12] , \wRegInB35[11] , \wRegInB35[10] , \wRegInB35[9] , 
        \wRegInB35[8] , \wRegInB35[7] , \wRegInB35[6] , \wRegInB35[5] , 
        \wRegInB35[4] , \wRegInB35[3] , \wRegInB35[2] , \wRegInB35[1] , 
        \wRegInB35[0] }), .Out({\wBIn35[31] , \wBIn35[30] , \wBIn35[29] , 
        \wBIn35[28] , \wBIn35[27] , \wBIn35[26] , \wBIn35[25] , \wBIn35[24] , 
        \wBIn35[23] , \wBIn35[22] , \wBIn35[21] , \wBIn35[20] , \wBIn35[19] , 
        \wBIn35[18] , \wBIn35[17] , \wBIn35[16] , \wBIn35[15] , \wBIn35[14] , 
        \wBIn35[13] , \wBIn35[12] , \wBIn35[11] , \wBIn35[10] , \wBIn35[9] , 
        \wBIn35[8] , \wBIn35[7] , \wBIn35[6] , \wBIn35[5] , \wBIn35[4] , 
        \wBIn35[3] , \wBIn35[2] , \wBIn35[1] , \wBIn35[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_128 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink129[31] , \ScanLink129[30] , \ScanLink129[29] , 
        \ScanLink129[28] , \ScanLink129[27] , \ScanLink129[26] , 
        \ScanLink129[25] , \ScanLink129[24] , \ScanLink129[23] , 
        \ScanLink129[22] , \ScanLink129[21] , \ScanLink129[20] , 
        \ScanLink129[19] , \ScanLink129[18] , \ScanLink129[17] , 
        \ScanLink129[16] , \ScanLink129[15] , \ScanLink129[14] , 
        \ScanLink129[13] , \ScanLink129[12] , \ScanLink129[11] , 
        \ScanLink129[10] , \ScanLink129[9] , \ScanLink129[8] , 
        \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , \ScanLink129[4] , 
        \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , \ScanLink129[0] 
        }), .ScanOut({\ScanLink128[31] , \ScanLink128[30] , \ScanLink128[29] , 
        \ScanLink128[28] , \ScanLink128[27] , \ScanLink128[26] , 
        \ScanLink128[25] , \ScanLink128[24] , \ScanLink128[23] , 
        \ScanLink128[22] , \ScanLink128[21] , \ScanLink128[20] , 
        \ScanLink128[19] , \ScanLink128[18] , \ScanLink128[17] , 
        \ScanLink128[16] , \ScanLink128[15] , \ScanLink128[14] , 
        \ScanLink128[13] , \ScanLink128[12] , \ScanLink128[11] , 
        \ScanLink128[10] , \ScanLink128[9] , \ScanLink128[8] , 
        \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , \ScanLink128[4] , 
        \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , \ScanLink128[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB63[31] , \wRegInB63[30] , \wRegInB63[29] , 
        \wRegInB63[28] , \wRegInB63[27] , \wRegInB63[26] , \wRegInB63[25] , 
        \wRegInB63[24] , \wRegInB63[23] , \wRegInB63[22] , \wRegInB63[21] , 
        \wRegInB63[20] , \wRegInB63[19] , \wRegInB63[18] , \wRegInB63[17] , 
        \wRegInB63[16] , \wRegInB63[15] , \wRegInB63[14] , \wRegInB63[13] , 
        \wRegInB63[12] , \wRegInB63[11] , \wRegInB63[10] , \wRegInB63[9] , 
        \wRegInB63[8] , \wRegInB63[7] , \wRegInB63[6] , \wRegInB63[5] , 
        \wRegInB63[4] , \wRegInB63[3] , \wRegInB63[2] , \wRegInB63[1] , 
        \wRegInB63[0] }), .Out({\wBIn63[31] , \wBIn63[30] , \wBIn63[29] , 
        \wBIn63[28] , \wBIn63[27] , \wBIn63[26] , \wBIn63[25] , \wBIn63[24] , 
        \wBIn63[23] , \wBIn63[22] , \wBIn63[21] , \wBIn63[20] , \wBIn63[19] , 
        \wBIn63[18] , \wBIn63[17] , \wBIn63[16] , \wBIn63[15] , \wBIn63[14] , 
        \wBIn63[13] , \wBIn63[12] , \wBIn63[11] , \wBIn63[10] , \wBIn63[9] , 
        \wBIn63[8] , \wBIn63[7] , \wBIn63[6] , \wBIn63[5] , \wBIn63[4] , 
        \wBIn63[3] , \wBIn63[2] , \wBIn63[1] , \wBIn63[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_78 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink79[31] , \ScanLink79[30] , \ScanLink79[29] , 
        \ScanLink79[28] , \ScanLink79[27] , \ScanLink79[26] , \ScanLink79[25] , 
        \ScanLink79[24] , \ScanLink79[23] , \ScanLink79[22] , \ScanLink79[21] , 
        \ScanLink79[20] , \ScanLink79[19] , \ScanLink79[18] , \ScanLink79[17] , 
        \ScanLink79[16] , \ScanLink79[15] , \ScanLink79[14] , \ScanLink79[13] , 
        \ScanLink79[12] , \ScanLink79[11] , \ScanLink79[10] , \ScanLink79[9] , 
        \ScanLink79[8] , \ScanLink79[7] , \ScanLink79[6] , \ScanLink79[5] , 
        \ScanLink79[4] , \ScanLink79[3] , \ScanLink79[2] , \ScanLink79[1] , 
        \ScanLink79[0] }), .ScanOut({\ScanLink78[31] , \ScanLink78[30] , 
        \ScanLink78[29] , \ScanLink78[28] , \ScanLink78[27] , \ScanLink78[26] , 
        \ScanLink78[25] , \ScanLink78[24] , \ScanLink78[23] , \ScanLink78[22] , 
        \ScanLink78[21] , \ScanLink78[20] , \ScanLink78[19] , \ScanLink78[18] , 
        \ScanLink78[17] , \ScanLink78[16] , \ScanLink78[15] , \ScanLink78[14] , 
        \ScanLink78[13] , \ScanLink78[12] , \ScanLink78[11] , \ScanLink78[10] , 
        \ScanLink78[9] , \ScanLink78[8] , \ScanLink78[7] , \ScanLink78[6] , 
        \ScanLink78[5] , \ScanLink78[4] , \ScanLink78[3] , \ScanLink78[2] , 
        \ScanLink78[1] , \ScanLink78[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB88[31] , \wRegInB88[30] , 
        \wRegInB88[29] , \wRegInB88[28] , \wRegInB88[27] , \wRegInB88[26] , 
        \wRegInB88[25] , \wRegInB88[24] , \wRegInB88[23] , \wRegInB88[22] , 
        \wRegInB88[21] , \wRegInB88[20] , \wRegInB88[19] , \wRegInB88[18] , 
        \wRegInB88[17] , \wRegInB88[16] , \wRegInB88[15] , \wRegInB88[14] , 
        \wRegInB88[13] , \wRegInB88[12] , \wRegInB88[11] , \wRegInB88[10] , 
        \wRegInB88[9] , \wRegInB88[8] , \wRegInB88[7] , \wRegInB88[6] , 
        \wRegInB88[5] , \wRegInB88[4] , \wRegInB88[3] , \wRegInB88[2] , 
        \wRegInB88[1] , \wRegInB88[0] }), .Out({\wBIn88[31] , \wBIn88[30] , 
        \wBIn88[29] , \wBIn88[28] , \wBIn88[27] , \wBIn88[26] , \wBIn88[25] , 
        \wBIn88[24] , \wBIn88[23] , \wBIn88[22] , \wBIn88[21] , \wBIn88[20] , 
        \wBIn88[19] , \wBIn88[18] , \wBIn88[17] , \wBIn88[16] , \wBIn88[15] , 
        \wBIn88[14] , \wBIn88[13] , \wBIn88[12] , \wBIn88[11] , \wBIn88[10] , 
        \wBIn88[9] , \wBIn88[8] , \wBIn88[7] , \wBIn88[6] , \wBIn88[5] , 
        \wBIn88[4] , \wBIn88[3] , \wBIn88[2] , \wBIn88[1] , \wBIn88[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid54[31] , \wAMid54[30] , \wAMid54[29] , \wAMid54[28] , 
        \wAMid54[27] , \wAMid54[26] , \wAMid54[25] , \wAMid54[24] , 
        \wAMid54[23] , \wAMid54[22] , \wAMid54[21] , \wAMid54[20] , 
        \wAMid54[19] , \wAMid54[18] , \wAMid54[17] , \wAMid54[16] , 
        \wAMid54[15] , \wAMid54[14] , \wAMid54[13] , \wAMid54[12] , 
        \wAMid54[11] , \wAMid54[10] , \wAMid54[9] , \wAMid54[8] , \wAMid54[7] , 
        \wAMid54[6] , \wAMid54[5] , \wAMid54[4] , \wAMid54[3] , \wAMid54[2] , 
        \wAMid54[1] , \wAMid54[0] }), .BIn({\wBMid54[31] , \wBMid54[30] , 
        \wBMid54[29] , \wBMid54[28] , \wBMid54[27] , \wBMid54[26] , 
        \wBMid54[25] , \wBMid54[24] , \wBMid54[23] , \wBMid54[22] , 
        \wBMid54[21] , \wBMid54[20] , \wBMid54[19] , \wBMid54[18] , 
        \wBMid54[17] , \wBMid54[16] , \wBMid54[15] , \wBMid54[14] , 
        \wBMid54[13] , \wBMid54[12] , \wBMid54[11] , \wBMid54[10] , 
        \wBMid54[9] , \wBMid54[8] , \wBMid54[7] , \wBMid54[6] , \wBMid54[5] , 
        \wBMid54[4] , \wBMid54[3] , \wBMid54[2] , \wBMid54[1] , \wBMid54[0] }), 
        .HiOut({\wRegInB54[31] , \wRegInB54[30] , \wRegInB54[29] , 
        \wRegInB54[28] , \wRegInB54[27] , \wRegInB54[26] , \wRegInB54[25] , 
        \wRegInB54[24] , \wRegInB54[23] , \wRegInB54[22] , \wRegInB54[21] , 
        \wRegInB54[20] , \wRegInB54[19] , \wRegInB54[18] , \wRegInB54[17] , 
        \wRegInB54[16] , \wRegInB54[15] , \wRegInB54[14] , \wRegInB54[13] , 
        \wRegInB54[12] , \wRegInB54[11] , \wRegInB54[10] , \wRegInB54[9] , 
        \wRegInB54[8] , \wRegInB54[7] , \wRegInB54[6] , \wRegInB54[5] , 
        \wRegInB54[4] , \wRegInB54[3] , \wRegInB54[2] , \wRegInB54[1] , 
        \wRegInB54[0] }), .LoOut({\wRegInA55[31] , \wRegInA55[30] , 
        \wRegInA55[29] , \wRegInA55[28] , \wRegInA55[27] , \wRegInA55[26] , 
        \wRegInA55[25] , \wRegInA55[24] , \wRegInA55[23] , \wRegInA55[22] , 
        \wRegInA55[21] , \wRegInA55[20] , \wRegInA55[19] , \wRegInA55[18] , 
        \wRegInA55[17] , \wRegInA55[16] , \wRegInA55[15] , \wRegInA55[14] , 
        \wRegInA55[13] , \wRegInA55[12] , \wRegInA55[11] , \wRegInA55[10] , 
        \wRegInA55[9] , \wRegInA55[8] , \wRegInA55[7] , \wRegInA55[6] , 
        \wRegInA55[5] , \wRegInA55[4] , \wRegInA55[3] , \wRegInA55[2] , 
        \wRegInA55[1] , \wRegInA55[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_31 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink32[31] , \ScanLink32[30] , \ScanLink32[29] , 
        \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , \ScanLink32[25] , 
        \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , \ScanLink32[21] , 
        \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , \ScanLink32[17] , 
        \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , \ScanLink32[13] , 
        \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , \ScanLink32[9] , 
        \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , \ScanLink32[5] , 
        \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , \ScanLink32[1] , 
        \ScanLink32[0] }), .ScanOut({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA112[31] , \wRegInA112[30] , 
        \wRegInA112[29] , \wRegInA112[28] , \wRegInA112[27] , \wRegInA112[26] , 
        \wRegInA112[25] , \wRegInA112[24] , \wRegInA112[23] , \wRegInA112[22] , 
        \wRegInA112[21] , \wRegInA112[20] , \wRegInA112[19] , \wRegInA112[18] , 
        \wRegInA112[17] , \wRegInA112[16] , \wRegInA112[15] , \wRegInA112[14] , 
        \wRegInA112[13] , \wRegInA112[12] , \wRegInA112[11] , \wRegInA112[10] , 
        \wRegInA112[9] , \wRegInA112[8] , \wRegInA112[7] , \wRegInA112[6] , 
        \wRegInA112[5] , \wRegInA112[4] , \wRegInA112[3] , \wRegInA112[2] , 
        \wRegInA112[1] , \wRegInA112[0] }), .Out({\wAIn112[31] , \wAIn112[30] , 
        \wAIn112[29] , \wAIn112[28] , \wAIn112[27] , \wAIn112[26] , 
        \wAIn112[25] , \wAIn112[24] , \wAIn112[23] , \wAIn112[22] , 
        \wAIn112[21] , \wAIn112[20] , \wAIn112[19] , \wAIn112[18] , 
        \wAIn112[17] , \wAIn112[16] , \wAIn112[15] , \wAIn112[14] , 
        \wAIn112[13] , \wAIn112[12] , \wAIn112[11] , \wAIn112[10] , 
        \wAIn112[9] , \wAIn112[8] , \wAIn112[7] , \wAIn112[6] , \wAIn112[5] , 
        \wAIn112[4] , \wAIn112[3] , \wAIn112[2] , \wAIn112[1] , \wAIn112[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_161 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink162[31] , \ScanLink162[30] , \ScanLink162[29] , 
        \ScanLink162[28] , \ScanLink162[27] , \ScanLink162[26] , 
        \ScanLink162[25] , \ScanLink162[24] , \ScanLink162[23] , 
        \ScanLink162[22] , \ScanLink162[21] , \ScanLink162[20] , 
        \ScanLink162[19] , \ScanLink162[18] , \ScanLink162[17] , 
        \ScanLink162[16] , \ScanLink162[15] , \ScanLink162[14] , 
        \ScanLink162[13] , \ScanLink162[12] , \ScanLink162[11] , 
        \ScanLink162[10] , \ScanLink162[9] , \ScanLink162[8] , 
        \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , \ScanLink162[4] , 
        \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , \ScanLink162[0] 
        }), .ScanOut({\ScanLink161[31] , \ScanLink161[30] , \ScanLink161[29] , 
        \ScanLink161[28] , \ScanLink161[27] , \ScanLink161[26] , 
        \ScanLink161[25] , \ScanLink161[24] , \ScanLink161[23] , 
        \ScanLink161[22] , \ScanLink161[21] , \ScanLink161[20] , 
        \ScanLink161[19] , \ScanLink161[18] , \ScanLink161[17] , 
        \ScanLink161[16] , \ScanLink161[15] , \ScanLink161[14] , 
        \ScanLink161[13] , \ScanLink161[12] , \ScanLink161[11] , 
        \ScanLink161[10] , \ScanLink161[9] , \ScanLink161[8] , 
        \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , \ScanLink161[4] , 
        \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , \ScanLink161[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA47[31] , \wRegInA47[30] , \wRegInA47[29] , 
        \wRegInA47[28] , \wRegInA47[27] , \wRegInA47[26] , \wRegInA47[25] , 
        \wRegInA47[24] , \wRegInA47[23] , \wRegInA47[22] , \wRegInA47[21] , 
        \wRegInA47[20] , \wRegInA47[19] , \wRegInA47[18] , \wRegInA47[17] , 
        \wRegInA47[16] , \wRegInA47[15] , \wRegInA47[14] , \wRegInA47[13] , 
        \wRegInA47[12] , \wRegInA47[11] , \wRegInA47[10] , \wRegInA47[9] , 
        \wRegInA47[8] , \wRegInA47[7] , \wRegInA47[6] , \wRegInA47[5] , 
        \wRegInA47[4] , \wRegInA47[3] , \wRegInA47[2] , \wRegInA47[1] , 
        \wRegInA47[0] }), .Out({\wAIn47[31] , \wAIn47[30] , \wAIn47[29] , 
        \wAIn47[28] , \wAIn47[27] , \wAIn47[26] , \wAIn47[25] , \wAIn47[24] , 
        \wAIn47[23] , \wAIn47[22] , \wAIn47[21] , \wAIn47[20] , \wAIn47[19] , 
        \wAIn47[18] , \wAIn47[17] , \wAIn47[16] , \wAIn47[15] , \wAIn47[14] , 
        \wAIn47[13] , \wAIn47[12] , \wAIn47[11] , \wAIn47[10] , \wAIn47[9] , 
        \wAIn47[8] , \wAIn47[7] , \wAIn47[6] , \wAIn47[5] , \wAIn47[4] , 
        \wAIn47[3] , \wAIn47[2] , \wAIn47[1] , \wAIn47[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid73[31] , \wAMid73[30] , \wAMid73[29] , \wAMid73[28] , 
        \wAMid73[27] , \wAMid73[26] , \wAMid73[25] , \wAMid73[24] , 
        \wAMid73[23] , \wAMid73[22] , \wAMid73[21] , \wAMid73[20] , 
        \wAMid73[19] , \wAMid73[18] , \wAMid73[17] , \wAMid73[16] , 
        \wAMid73[15] , \wAMid73[14] , \wAMid73[13] , \wAMid73[12] , 
        \wAMid73[11] , \wAMid73[10] , \wAMid73[9] , \wAMid73[8] , \wAMid73[7] , 
        \wAMid73[6] , \wAMid73[5] , \wAMid73[4] , \wAMid73[3] , \wAMid73[2] , 
        \wAMid73[1] , \wAMid73[0] }), .BIn({\wBMid73[31] , \wBMid73[30] , 
        \wBMid73[29] , \wBMid73[28] , \wBMid73[27] , \wBMid73[26] , 
        \wBMid73[25] , \wBMid73[24] , \wBMid73[23] , \wBMid73[22] , 
        \wBMid73[21] , \wBMid73[20] , \wBMid73[19] , \wBMid73[18] , 
        \wBMid73[17] , \wBMid73[16] , \wBMid73[15] , \wBMid73[14] , 
        \wBMid73[13] , \wBMid73[12] , \wBMid73[11] , \wBMid73[10] , 
        \wBMid73[9] , \wBMid73[8] , \wBMid73[7] , \wBMid73[6] , \wBMid73[5] , 
        \wBMid73[4] , \wBMid73[3] , \wBMid73[2] , \wBMid73[1] , \wBMid73[0] }), 
        .HiOut({\wRegInB73[31] , \wRegInB73[30] , \wRegInB73[29] , 
        \wRegInB73[28] , \wRegInB73[27] , \wRegInB73[26] , \wRegInB73[25] , 
        \wRegInB73[24] , \wRegInB73[23] , \wRegInB73[22] , \wRegInB73[21] , 
        \wRegInB73[20] , \wRegInB73[19] , \wRegInB73[18] , \wRegInB73[17] , 
        \wRegInB73[16] , \wRegInB73[15] , \wRegInB73[14] , \wRegInB73[13] , 
        \wRegInB73[12] , \wRegInB73[11] , \wRegInB73[10] , \wRegInB73[9] , 
        \wRegInB73[8] , \wRegInB73[7] , \wRegInB73[6] , \wRegInB73[5] , 
        \wRegInB73[4] , \wRegInB73[3] , \wRegInB73[2] , \wRegInB73[1] , 
        \wRegInB73[0] }), .LoOut({\wRegInA74[31] , \wRegInA74[30] , 
        \wRegInA74[29] , \wRegInA74[28] , \wRegInA74[27] , \wRegInA74[26] , 
        \wRegInA74[25] , \wRegInA74[24] , \wRegInA74[23] , \wRegInA74[22] , 
        \wRegInA74[21] , \wRegInA74[20] , \wRegInA74[19] , \wRegInA74[18] , 
        \wRegInA74[17] , \wRegInA74[16] , \wRegInA74[15] , \wRegInA74[14] , 
        \wRegInA74[13] , \wRegInA74[12] , \wRegInA74[11] , \wRegInA74[10] , 
        \wRegInA74[9] , \wRegInA74[8] , \wRegInA74[7] , \wRegInA74[6] , 
        \wRegInA74[5] , \wRegInA74[4] , \wRegInA74[3] , \wRegInA74[2] , 
        \wRegInA74[1] , \wRegInA74[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_146 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink147[31] , \ScanLink147[30] , \ScanLink147[29] , 
        \ScanLink147[28] , \ScanLink147[27] , \ScanLink147[26] , 
        \ScanLink147[25] , \ScanLink147[24] , \ScanLink147[23] , 
        \ScanLink147[22] , \ScanLink147[21] , \ScanLink147[20] , 
        \ScanLink147[19] , \ScanLink147[18] , \ScanLink147[17] , 
        \ScanLink147[16] , \ScanLink147[15] , \ScanLink147[14] , 
        \ScanLink147[13] , \ScanLink147[12] , \ScanLink147[11] , 
        \ScanLink147[10] , \ScanLink147[9] , \ScanLink147[8] , 
        \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , \ScanLink147[4] , 
        \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , \ScanLink147[0] 
        }), .ScanOut({\ScanLink146[31] , \ScanLink146[30] , \ScanLink146[29] , 
        \ScanLink146[28] , \ScanLink146[27] , \ScanLink146[26] , 
        \ScanLink146[25] , \ScanLink146[24] , \ScanLink146[23] , 
        \ScanLink146[22] , \ScanLink146[21] , \ScanLink146[20] , 
        \ScanLink146[19] , \ScanLink146[18] , \ScanLink146[17] , 
        \ScanLink146[16] , \ScanLink146[15] , \ScanLink146[14] , 
        \ScanLink146[13] , \ScanLink146[12] , \ScanLink146[11] , 
        \ScanLink146[10] , \ScanLink146[9] , \ScanLink146[8] , 
        \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , \ScanLink146[4] , 
        \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , \ScanLink146[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB54[31] , \wRegInB54[30] , \wRegInB54[29] , 
        \wRegInB54[28] , \wRegInB54[27] , \wRegInB54[26] , \wRegInB54[25] , 
        \wRegInB54[24] , \wRegInB54[23] , \wRegInB54[22] , \wRegInB54[21] , 
        \wRegInB54[20] , \wRegInB54[19] , \wRegInB54[18] , \wRegInB54[17] , 
        \wRegInB54[16] , \wRegInB54[15] , \wRegInB54[14] , \wRegInB54[13] , 
        \wRegInB54[12] , \wRegInB54[11] , \wRegInB54[10] , \wRegInB54[9] , 
        \wRegInB54[8] , \wRegInB54[7] , \wRegInB54[6] , \wRegInB54[5] , 
        \wRegInB54[4] , \wRegInB54[3] , \wRegInB54[2] , \wRegInB54[1] , 
        \wRegInB54[0] }), .Out({\wBIn54[31] , \wBIn54[30] , \wBIn54[29] , 
        \wBIn54[28] , \wBIn54[27] , \wBIn54[26] , \wBIn54[25] , \wBIn54[24] , 
        \wBIn54[23] , \wBIn54[22] , \wBIn54[21] , \wBIn54[20] , \wBIn54[19] , 
        \wBIn54[18] , \wBIn54[17] , \wBIn54[16] , \wBIn54[15] , \wBIn54[14] , 
        \wBIn54[13] , \wBIn54[12] , \wBIn54[11] , \wBIn54[10] , \wBIn54[9] , 
        \wBIn54[8] , \wBIn54[7] , \wBIn54[6] , \wBIn54[5] , \wBIn54[4] , 
        \wBIn54[3] , \wBIn54[2] , \wBIn54[1] , \wBIn54[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_16 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink17[31] , \ScanLink17[30] , \ScanLink17[29] , 
        \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , \ScanLink17[25] , 
        \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , \ScanLink17[21] , 
        \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , \ScanLink17[17] , 
        \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , \ScanLink17[13] , 
        \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , \ScanLink17[9] , 
        \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , \ScanLink17[5] , 
        \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , \ScanLink17[1] , 
        \ScanLink17[0] }), .ScanOut({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB119[31] , \wRegInB119[30] , 
        \wRegInB119[29] , \wRegInB119[28] , \wRegInB119[27] , \wRegInB119[26] , 
        \wRegInB119[25] , \wRegInB119[24] , \wRegInB119[23] , \wRegInB119[22] , 
        \wRegInB119[21] , \wRegInB119[20] , \wRegInB119[19] , \wRegInB119[18] , 
        \wRegInB119[17] , \wRegInB119[16] , \wRegInB119[15] , \wRegInB119[14] , 
        \wRegInB119[13] , \wRegInB119[12] , \wRegInB119[11] , \wRegInB119[10] , 
        \wRegInB119[9] , \wRegInB119[8] , \wRegInB119[7] , \wRegInB119[6] , 
        \wRegInB119[5] , \wRegInB119[4] , \wRegInB119[3] , \wRegInB119[2] , 
        \wRegInB119[1] , \wRegInB119[0] }), .Out({\wBIn119[31] , \wBIn119[30] , 
        \wBIn119[29] , \wBIn119[28] , \wBIn119[27] , \wBIn119[26] , 
        \wBIn119[25] , \wBIn119[24] , \wBIn119[23] , \wBIn119[22] , 
        \wBIn119[21] , \wBIn119[20] , \wBIn119[19] , \wBIn119[18] , 
        \wBIn119[17] , \wBIn119[16] , \wBIn119[15] , \wBIn119[14] , 
        \wBIn119[13] , \wBIn119[12] , \wBIn119[11] , \wBIn119[10] , 
        \wBIn119[9] , \wBIn119[8] , \wBIn119[7] , \wBIn119[6] , \wBIn119[5] , 
        \wBIn119[4] , \wBIn119[3] , \wBIn119[2] , \wBIn119[1] , \wBIn119[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn58[31] , \wAIn58[30] , \wAIn58[29] , \wAIn58[28] , \wAIn58[27] , 
        \wAIn58[26] , \wAIn58[25] , \wAIn58[24] , \wAIn58[23] , \wAIn58[22] , 
        \wAIn58[21] , \wAIn58[20] , \wAIn58[19] , \wAIn58[18] , \wAIn58[17] , 
        \wAIn58[16] , \wAIn58[15] , \wAIn58[14] , \wAIn58[13] , \wAIn58[12] , 
        \wAIn58[11] , \wAIn58[10] , \wAIn58[9] , \wAIn58[8] , \wAIn58[7] , 
        \wAIn58[6] , \wAIn58[5] , \wAIn58[4] , \wAIn58[3] , \wAIn58[2] , 
        \wAIn58[1] , \wAIn58[0] }), .BIn({\wBIn58[31] , \wBIn58[30] , 
        \wBIn58[29] , \wBIn58[28] , \wBIn58[27] , \wBIn58[26] , \wBIn58[25] , 
        \wBIn58[24] , \wBIn58[23] , \wBIn58[22] , \wBIn58[21] , \wBIn58[20] , 
        \wBIn58[19] , \wBIn58[18] , \wBIn58[17] , \wBIn58[16] , \wBIn58[15] , 
        \wBIn58[14] , \wBIn58[13] , \wBIn58[12] , \wBIn58[11] , \wBIn58[10] , 
        \wBIn58[9] , \wBIn58[8] , \wBIn58[7] , \wBIn58[6] , \wBIn58[5] , 
        \wBIn58[4] , \wBIn58[3] , \wBIn58[2] , \wBIn58[1] , \wBIn58[0] }), 
        .HiOut({\wBMid57[31] , \wBMid57[30] , \wBMid57[29] , \wBMid57[28] , 
        \wBMid57[27] , \wBMid57[26] , \wBMid57[25] , \wBMid57[24] , 
        \wBMid57[23] , \wBMid57[22] , \wBMid57[21] , \wBMid57[20] , 
        \wBMid57[19] , \wBMid57[18] , \wBMid57[17] , \wBMid57[16] , 
        \wBMid57[15] , \wBMid57[14] , \wBMid57[13] , \wBMid57[12] , 
        \wBMid57[11] , \wBMid57[10] , \wBMid57[9] , \wBMid57[8] , \wBMid57[7] , 
        \wBMid57[6] , \wBMid57[5] , \wBMid57[4] , \wBMid57[3] , \wBMid57[2] , 
        \wBMid57[1] , \wBMid57[0] }), .LoOut({\wAMid58[31] , \wAMid58[30] , 
        \wAMid58[29] , \wAMid58[28] , \wAMid58[27] , \wAMid58[26] , 
        \wAMid58[25] , \wAMid58[24] , \wAMid58[23] , \wAMid58[22] , 
        \wAMid58[21] , \wAMid58[20] , \wAMid58[19] , \wAMid58[18] , 
        \wAMid58[17] , \wAMid58[16] , \wAMid58[15] , \wAMid58[14] , 
        \wAMid58[13] , \wAMid58[12] , \wAMid58[11] , \wAMid58[10] , 
        \wAMid58[9] , \wAMid58[8] , \wAMid58[7] , \wAMid58[6] , \wAMid58[5] , 
        \wAMid58[4] , \wAMid58[3] , \wAMid58[2] , \wAMid58[1] , \wAMid58[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid105[31] , \wAMid105[30] , \wAMid105[29] , \wAMid105[28] , 
        \wAMid105[27] , \wAMid105[26] , \wAMid105[25] , \wAMid105[24] , 
        \wAMid105[23] , \wAMid105[22] , \wAMid105[21] , \wAMid105[20] , 
        \wAMid105[19] , \wAMid105[18] , \wAMid105[17] , \wAMid105[16] , 
        \wAMid105[15] , \wAMid105[14] , \wAMid105[13] , \wAMid105[12] , 
        \wAMid105[11] , \wAMid105[10] , \wAMid105[9] , \wAMid105[8] , 
        \wAMid105[7] , \wAMid105[6] , \wAMid105[5] , \wAMid105[4] , 
        \wAMid105[3] , \wAMid105[2] , \wAMid105[1] , \wAMid105[0] }), .BIn({
        \wBMid105[31] , \wBMid105[30] , \wBMid105[29] , \wBMid105[28] , 
        \wBMid105[27] , \wBMid105[26] , \wBMid105[25] , \wBMid105[24] , 
        \wBMid105[23] , \wBMid105[22] , \wBMid105[21] , \wBMid105[20] , 
        \wBMid105[19] , \wBMid105[18] , \wBMid105[17] , \wBMid105[16] , 
        \wBMid105[15] , \wBMid105[14] , \wBMid105[13] , \wBMid105[12] , 
        \wBMid105[11] , \wBMid105[10] , \wBMid105[9] , \wBMid105[8] , 
        \wBMid105[7] , \wBMid105[6] , \wBMid105[5] , \wBMid105[4] , 
        \wBMid105[3] , \wBMid105[2] , \wBMid105[1] , \wBMid105[0] }), .HiOut({
        \wRegInB105[31] , \wRegInB105[30] , \wRegInB105[29] , \wRegInB105[28] , 
        \wRegInB105[27] , \wRegInB105[26] , \wRegInB105[25] , \wRegInB105[24] , 
        \wRegInB105[23] , \wRegInB105[22] , \wRegInB105[21] , \wRegInB105[20] , 
        \wRegInB105[19] , \wRegInB105[18] , \wRegInB105[17] , \wRegInB105[16] , 
        \wRegInB105[15] , \wRegInB105[14] , \wRegInB105[13] , \wRegInB105[12] , 
        \wRegInB105[11] , \wRegInB105[10] , \wRegInB105[9] , \wRegInB105[8] , 
        \wRegInB105[7] , \wRegInB105[6] , \wRegInB105[5] , \wRegInB105[4] , 
        \wRegInB105[3] , \wRegInB105[2] , \wRegInB105[1] , \wRegInB105[0] }), 
        .LoOut({\wRegInA106[31] , \wRegInA106[30] , \wRegInA106[29] , 
        \wRegInA106[28] , \wRegInA106[27] , \wRegInA106[26] , \wRegInA106[25] , 
        \wRegInA106[24] , \wRegInA106[23] , \wRegInA106[22] , \wRegInA106[21] , 
        \wRegInA106[20] , \wRegInA106[19] , \wRegInA106[18] , \wRegInA106[17] , 
        \wRegInA106[16] , \wRegInA106[15] , \wRegInA106[14] , \wRegInA106[13] , 
        \wRegInA106[12] , \wRegInA106[11] , \wRegInA106[10] , \wRegInA106[9] , 
        \wRegInA106[8] , \wRegInA106[7] , \wRegInA106[6] , \wRegInA106[5] , 
        \wRegInA106[4] , \wRegInA106[3] , \wRegInA106[2] , \wRegInA106[1] , 
        \wRegInA106[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid122[31] , \wAMid122[30] , \wAMid122[29] , \wAMid122[28] , 
        \wAMid122[27] , \wAMid122[26] , \wAMid122[25] , \wAMid122[24] , 
        \wAMid122[23] , \wAMid122[22] , \wAMid122[21] , \wAMid122[20] , 
        \wAMid122[19] , \wAMid122[18] , \wAMid122[17] , \wAMid122[16] , 
        \wAMid122[15] , \wAMid122[14] , \wAMid122[13] , \wAMid122[12] , 
        \wAMid122[11] , \wAMid122[10] , \wAMid122[9] , \wAMid122[8] , 
        \wAMid122[7] , \wAMid122[6] , \wAMid122[5] , \wAMid122[4] , 
        \wAMid122[3] , \wAMid122[2] , \wAMid122[1] , \wAMid122[0] }), .BIn({
        \wBMid122[31] , \wBMid122[30] , \wBMid122[29] , \wBMid122[28] , 
        \wBMid122[27] , \wBMid122[26] , \wBMid122[25] , \wBMid122[24] , 
        \wBMid122[23] , \wBMid122[22] , \wBMid122[21] , \wBMid122[20] , 
        \wBMid122[19] , \wBMid122[18] , \wBMid122[17] , \wBMid122[16] , 
        \wBMid122[15] , \wBMid122[14] , \wBMid122[13] , \wBMid122[12] , 
        \wBMid122[11] , \wBMid122[10] , \wBMid122[9] , \wBMid122[8] , 
        \wBMid122[7] , \wBMid122[6] , \wBMid122[5] , \wBMid122[4] , 
        \wBMid122[3] , \wBMid122[2] , \wBMid122[1] , \wBMid122[0] }), .HiOut({
        \wRegInB122[31] , \wRegInB122[30] , \wRegInB122[29] , \wRegInB122[28] , 
        \wRegInB122[27] , \wRegInB122[26] , \wRegInB122[25] , \wRegInB122[24] , 
        \wRegInB122[23] , \wRegInB122[22] , \wRegInB122[21] , \wRegInB122[20] , 
        \wRegInB122[19] , \wRegInB122[18] , \wRegInB122[17] , \wRegInB122[16] , 
        \wRegInB122[15] , \wRegInB122[14] , \wRegInB122[13] , \wRegInB122[12] , 
        \wRegInB122[11] , \wRegInB122[10] , \wRegInB122[9] , \wRegInB122[8] , 
        \wRegInB122[7] , \wRegInB122[6] , \wRegInB122[5] , \wRegInB122[4] , 
        \wRegInB122[3] , \wRegInB122[2] , \wRegInB122[1] , \wRegInB122[0] }), 
        .LoOut({\wRegInA123[31] , \wRegInA123[30] , \wRegInA123[29] , 
        \wRegInA123[28] , \wRegInA123[27] , \wRegInA123[26] , \wRegInA123[25] , 
        \wRegInA123[24] , \wRegInA123[23] , \wRegInA123[22] , \wRegInA123[21] , 
        \wRegInA123[20] , \wRegInA123[19] , \wRegInA123[18] , \wRegInA123[17] , 
        \wRegInA123[16] , \wRegInA123[15] , \wRegInA123[14] , \wRegInA123[13] , 
        \wRegInA123[12] , \wRegInA123[11] , \wRegInA123[10] , \wRegInA123[9] , 
        \wRegInA123[8] , \wRegInA123[7] , \wRegInA123[6] , \wRegInA123[5] , 
        \wRegInA123[4] , \wRegInA123[3] , \wRegInA123[2] , \wRegInA123[1] , 
        \wRegInA123[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_86 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink87[31] , \ScanLink87[30] , \ScanLink87[29] , 
        \ScanLink87[28] , \ScanLink87[27] , \ScanLink87[26] , \ScanLink87[25] , 
        \ScanLink87[24] , \ScanLink87[23] , \ScanLink87[22] , \ScanLink87[21] , 
        \ScanLink87[20] , \ScanLink87[19] , \ScanLink87[18] , \ScanLink87[17] , 
        \ScanLink87[16] , \ScanLink87[15] , \ScanLink87[14] , \ScanLink87[13] , 
        \ScanLink87[12] , \ScanLink87[11] , \ScanLink87[10] , \ScanLink87[9] , 
        \ScanLink87[8] , \ScanLink87[7] , \ScanLink87[6] , \ScanLink87[5] , 
        \ScanLink87[4] , \ScanLink87[3] , \ScanLink87[2] , \ScanLink87[1] , 
        \ScanLink87[0] }), .ScanOut({\ScanLink86[31] , \ScanLink86[30] , 
        \ScanLink86[29] , \ScanLink86[28] , \ScanLink86[27] , \ScanLink86[26] , 
        \ScanLink86[25] , \ScanLink86[24] , \ScanLink86[23] , \ScanLink86[22] , 
        \ScanLink86[21] , \ScanLink86[20] , \ScanLink86[19] , \ScanLink86[18] , 
        \ScanLink86[17] , \ScanLink86[16] , \ScanLink86[15] , \ScanLink86[14] , 
        \ScanLink86[13] , \ScanLink86[12] , \ScanLink86[11] , \ScanLink86[10] , 
        \ScanLink86[9] , \ScanLink86[8] , \ScanLink86[7] , \ScanLink86[6] , 
        \ScanLink86[5] , \ScanLink86[4] , \ScanLink86[3] , \ScanLink86[2] , 
        \ScanLink86[1] , \ScanLink86[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB84[31] , \wRegInB84[30] , 
        \wRegInB84[29] , \wRegInB84[28] , \wRegInB84[27] , \wRegInB84[26] , 
        \wRegInB84[25] , \wRegInB84[24] , \wRegInB84[23] , \wRegInB84[22] , 
        \wRegInB84[21] , \wRegInB84[20] , \wRegInB84[19] , \wRegInB84[18] , 
        \wRegInB84[17] , \wRegInB84[16] , \wRegInB84[15] , \wRegInB84[14] , 
        \wRegInB84[13] , \wRegInB84[12] , \wRegInB84[11] , \wRegInB84[10] , 
        \wRegInB84[9] , \wRegInB84[8] , \wRegInB84[7] , \wRegInB84[6] , 
        \wRegInB84[5] , \wRegInB84[4] , \wRegInB84[3] , \wRegInB84[2] , 
        \wRegInB84[1] , \wRegInB84[0] }), .Out({\wBIn84[31] , \wBIn84[30] , 
        \wBIn84[29] , \wBIn84[28] , \wBIn84[27] , \wBIn84[26] , \wBIn84[25] , 
        \wBIn84[24] , \wBIn84[23] , \wBIn84[22] , \wBIn84[21] , \wBIn84[20] , 
        \wBIn84[19] , \wBIn84[18] , \wBIn84[17] , \wBIn84[16] , \wBIn84[15] , 
        \wBIn84[14] , \wBIn84[13] , \wBIn84[12] , \wBIn84[11] , \wBIn84[10] , 
        \wBIn84[9] , \wBIn84[8] , \wBIn84[7] , \wBIn84[6] , \wBIn84[5] , 
        \wBIn84[4] , \wBIn84[3] , \wBIn84[2] , \wBIn84[1] , \wBIn84[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid68[31] , \wAMid68[30] , \wAMid68[29] , \wAMid68[28] , 
        \wAMid68[27] , \wAMid68[26] , \wAMid68[25] , \wAMid68[24] , 
        \wAMid68[23] , \wAMid68[22] , \wAMid68[21] , \wAMid68[20] , 
        \wAMid68[19] , \wAMid68[18] , \wAMid68[17] , \wAMid68[16] , 
        \wAMid68[15] , \wAMid68[14] , \wAMid68[13] , \wAMid68[12] , 
        \wAMid68[11] , \wAMid68[10] , \wAMid68[9] , \wAMid68[8] , \wAMid68[7] , 
        \wAMid68[6] , \wAMid68[5] , \wAMid68[4] , \wAMid68[3] , \wAMid68[2] , 
        \wAMid68[1] , \wAMid68[0] }), .BIn({\wBMid68[31] , \wBMid68[30] , 
        \wBMid68[29] , \wBMid68[28] , \wBMid68[27] , \wBMid68[26] , 
        \wBMid68[25] , \wBMid68[24] , \wBMid68[23] , \wBMid68[22] , 
        \wBMid68[21] , \wBMid68[20] , \wBMid68[19] , \wBMid68[18] , 
        \wBMid68[17] , \wBMid68[16] , \wBMid68[15] , \wBMid68[14] , 
        \wBMid68[13] , \wBMid68[12] , \wBMid68[11] , \wBMid68[10] , 
        \wBMid68[9] , \wBMid68[8] , \wBMid68[7] , \wBMid68[6] , \wBMid68[5] , 
        \wBMid68[4] , \wBMid68[3] , \wBMid68[2] , \wBMid68[1] , \wBMid68[0] }), 
        .HiOut({\wRegInB68[31] , \wRegInB68[30] , \wRegInB68[29] , 
        \wRegInB68[28] , \wRegInB68[27] , \wRegInB68[26] , \wRegInB68[25] , 
        \wRegInB68[24] , \wRegInB68[23] , \wRegInB68[22] , \wRegInB68[21] , 
        \wRegInB68[20] , \wRegInB68[19] , \wRegInB68[18] , \wRegInB68[17] , 
        \wRegInB68[16] , \wRegInB68[15] , \wRegInB68[14] , \wRegInB68[13] , 
        \wRegInB68[12] , \wRegInB68[11] , \wRegInB68[10] , \wRegInB68[9] , 
        \wRegInB68[8] , \wRegInB68[7] , \wRegInB68[6] , \wRegInB68[5] , 
        \wRegInB68[4] , \wRegInB68[3] , \wRegInB68[2] , \wRegInB68[1] , 
        \wRegInB68[0] }), .LoOut({\wRegInA69[31] , \wRegInA69[30] , 
        \wRegInA69[29] , \wRegInA69[28] , \wRegInA69[27] , \wRegInA69[26] , 
        \wRegInA69[25] , \wRegInA69[24] , \wRegInA69[23] , \wRegInA69[22] , 
        \wRegInA69[21] , \wRegInA69[20] , \wRegInA69[19] , \wRegInA69[18] , 
        \wRegInA69[17] , \wRegInA69[16] , \wRegInA69[15] , \wRegInA69[14] , 
        \wRegInA69[13] , \wRegInA69[12] , \wRegInA69[11] , \wRegInA69[10] , 
        \wRegInA69[9] , \wRegInA69[8] , \wRegInA69[7] , \wRegInA69[6] , 
        \wRegInA69[5] , \wRegInA69[4] , \wRegInA69[3] , \wRegInA69[2] , 
        \wRegInA69[1] , \wRegInA69[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn18[31] , \wAIn18[30] , \wAIn18[29] , \wAIn18[28] , \wAIn18[27] , 
        \wAIn18[26] , \wAIn18[25] , \wAIn18[24] , \wAIn18[23] , \wAIn18[22] , 
        \wAIn18[21] , \wAIn18[20] , \wAIn18[19] , \wAIn18[18] , \wAIn18[17] , 
        \wAIn18[16] , \wAIn18[15] , \wAIn18[14] , \wAIn18[13] , \wAIn18[12] , 
        \wAIn18[11] , \wAIn18[10] , \wAIn18[9] , \wAIn18[8] , \wAIn18[7] , 
        \wAIn18[6] , \wAIn18[5] , \wAIn18[4] , \wAIn18[3] , \wAIn18[2] , 
        \wAIn18[1] , \wAIn18[0] }), .BIn({\wBIn18[31] , \wBIn18[30] , 
        \wBIn18[29] , \wBIn18[28] , \wBIn18[27] , \wBIn18[26] , \wBIn18[25] , 
        \wBIn18[24] , \wBIn18[23] , \wBIn18[22] , \wBIn18[21] , \wBIn18[20] , 
        \wBIn18[19] , \wBIn18[18] , \wBIn18[17] , \wBIn18[16] , \wBIn18[15] , 
        \wBIn18[14] , \wBIn18[13] , \wBIn18[12] , \wBIn18[11] , \wBIn18[10] , 
        \wBIn18[9] , \wBIn18[8] , \wBIn18[7] , \wBIn18[6] , \wBIn18[5] , 
        \wBIn18[4] , \wBIn18[3] , \wBIn18[2] , \wBIn18[1] , \wBIn18[0] }), 
        .HiOut({\wBMid17[31] , \wBMid17[30] , \wBMid17[29] , \wBMid17[28] , 
        \wBMid17[27] , \wBMid17[26] , \wBMid17[25] , \wBMid17[24] , 
        \wBMid17[23] , \wBMid17[22] , \wBMid17[21] , \wBMid17[20] , 
        \wBMid17[19] , \wBMid17[18] , \wBMid17[17] , \wBMid17[16] , 
        \wBMid17[15] , \wBMid17[14] , \wBMid17[13] , \wBMid17[12] , 
        \wBMid17[11] , \wBMid17[10] , \wBMid17[9] , \wBMid17[8] , \wBMid17[7] , 
        \wBMid17[6] , \wBMid17[5] , \wBMid17[4] , \wBMid17[3] , \wBMid17[2] , 
        \wBMid17[1] , \wBMid17[0] }), .LoOut({\wAMid18[31] , \wAMid18[30] , 
        \wAMid18[29] , \wAMid18[28] , \wAMid18[27] , \wAMid18[26] , 
        \wAMid18[25] , \wAMid18[24] , \wAMid18[23] , \wAMid18[22] , 
        \wAMid18[21] , \wAMid18[20] , \wAMid18[19] , \wAMid18[18] , 
        \wAMid18[17] , \wAMid18[16] , \wAMid18[15] , \wAMid18[14] , 
        \wAMid18[13] , \wAMid18[12] , \wAMid18[11] , \wAMid18[10] , 
        \wAMid18[9] , \wAMid18[8] , \wAMid18[7] , \wAMid18[6] , \wAMid18[5] , 
        \wAMid18[4] , \wAMid18[3] , \wAMid18[2] , \wAMid18[1] , \wAMid18[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn24[31] , \wAIn24[30] , \wAIn24[29] , \wAIn24[28] , \wAIn24[27] , 
        \wAIn24[26] , \wAIn24[25] , \wAIn24[24] , \wAIn24[23] , \wAIn24[22] , 
        \wAIn24[21] , \wAIn24[20] , \wAIn24[19] , \wAIn24[18] , \wAIn24[17] , 
        \wAIn24[16] , \wAIn24[15] , \wAIn24[14] , \wAIn24[13] , \wAIn24[12] , 
        \wAIn24[11] , \wAIn24[10] , \wAIn24[9] , \wAIn24[8] , \wAIn24[7] , 
        \wAIn24[6] , \wAIn24[5] , \wAIn24[4] , \wAIn24[3] , \wAIn24[2] , 
        \wAIn24[1] , \wAIn24[0] }), .BIn({\wBIn24[31] , \wBIn24[30] , 
        \wBIn24[29] , \wBIn24[28] , \wBIn24[27] , \wBIn24[26] , \wBIn24[25] , 
        \wBIn24[24] , \wBIn24[23] , \wBIn24[22] , \wBIn24[21] , \wBIn24[20] , 
        \wBIn24[19] , \wBIn24[18] , \wBIn24[17] , \wBIn24[16] , \wBIn24[15] , 
        \wBIn24[14] , \wBIn24[13] , \wBIn24[12] , \wBIn24[11] , \wBIn24[10] , 
        \wBIn24[9] , \wBIn24[8] , \wBIn24[7] , \wBIn24[6] , \wBIn24[5] , 
        \wBIn24[4] , \wBIn24[3] , \wBIn24[2] , \wBIn24[1] , \wBIn24[0] }), 
        .HiOut({\wBMid23[31] , \wBMid23[30] , \wBMid23[29] , \wBMid23[28] , 
        \wBMid23[27] , \wBMid23[26] , \wBMid23[25] , \wBMid23[24] , 
        \wBMid23[23] , \wBMid23[22] , \wBMid23[21] , \wBMid23[20] , 
        \wBMid23[19] , \wBMid23[18] , \wBMid23[17] , \wBMid23[16] , 
        \wBMid23[15] , \wBMid23[14] , \wBMid23[13] , \wBMid23[12] , 
        \wBMid23[11] , \wBMid23[10] , \wBMid23[9] , \wBMid23[8] , \wBMid23[7] , 
        \wBMid23[6] , \wBMid23[5] , \wBMid23[4] , \wBMid23[3] , \wBMid23[2] , 
        \wBMid23[1] , \wBMid23[0] }), .LoOut({\wAMid24[31] , \wAMid24[30] , 
        \wAMid24[29] , \wAMid24[28] , \wAMid24[27] , \wAMid24[26] , 
        \wAMid24[25] , \wAMid24[24] , \wAMid24[23] , \wAMid24[22] , 
        \wAMid24[21] , \wAMid24[20] , \wAMid24[19] , \wAMid24[18] , 
        \wAMid24[17] , \wAMid24[16] , \wAMid24[15] , \wAMid24[14] , 
        \wAMid24[13] , \wAMid24[12] , \wAMid24[11] , \wAMid24[10] , 
        \wAMid24[9] , \wAMid24[8] , \wAMid24[7] , \wAMid24[6] , \wAMid24[5] , 
        \wAMid24[4] , \wAMid24[3] , \wAMid24[2] , \wAMid24[1] , \wAMid24[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn36[31] , \wAIn36[30] , \wAIn36[29] , \wAIn36[28] , \wAIn36[27] , 
        \wAIn36[26] , \wAIn36[25] , \wAIn36[24] , \wAIn36[23] , \wAIn36[22] , 
        \wAIn36[21] , \wAIn36[20] , \wAIn36[19] , \wAIn36[18] , \wAIn36[17] , 
        \wAIn36[16] , \wAIn36[15] , \wAIn36[14] , \wAIn36[13] , \wAIn36[12] , 
        \wAIn36[11] , \wAIn36[10] , \wAIn36[9] , \wAIn36[8] , \wAIn36[7] , 
        \wAIn36[6] , \wAIn36[5] , \wAIn36[4] , \wAIn36[3] , \wAIn36[2] , 
        \wAIn36[1] , \wAIn36[0] }), .BIn({\wBIn36[31] , \wBIn36[30] , 
        \wBIn36[29] , \wBIn36[28] , \wBIn36[27] , \wBIn36[26] , \wBIn36[25] , 
        \wBIn36[24] , \wBIn36[23] , \wBIn36[22] , \wBIn36[21] , \wBIn36[20] , 
        \wBIn36[19] , \wBIn36[18] , \wBIn36[17] , \wBIn36[16] , \wBIn36[15] , 
        \wBIn36[14] , \wBIn36[13] , \wBIn36[12] , \wBIn36[11] , \wBIn36[10] , 
        \wBIn36[9] , \wBIn36[8] , \wBIn36[7] , \wBIn36[6] , \wBIn36[5] , 
        \wBIn36[4] , \wBIn36[3] , \wBIn36[2] , \wBIn36[1] , \wBIn36[0] }), 
        .HiOut({\wBMid35[31] , \wBMid35[30] , \wBMid35[29] , \wBMid35[28] , 
        \wBMid35[27] , \wBMid35[26] , \wBMid35[25] , \wBMid35[24] , 
        \wBMid35[23] , \wBMid35[22] , \wBMid35[21] , \wBMid35[20] , 
        \wBMid35[19] , \wBMid35[18] , \wBMid35[17] , \wBMid35[16] , 
        \wBMid35[15] , \wBMid35[14] , \wBMid35[13] , \wBMid35[12] , 
        \wBMid35[11] , \wBMid35[10] , \wBMid35[9] , \wBMid35[8] , \wBMid35[7] , 
        \wBMid35[6] , \wBMid35[5] , \wBMid35[4] , \wBMid35[3] , \wBMid35[2] , 
        \wBMid35[1] , \wBMid35[0] }), .LoOut({\wAMid36[31] , \wAMid36[30] , 
        \wAMid36[29] , \wAMid36[28] , \wAMid36[27] , \wAMid36[26] , 
        \wAMid36[25] , \wAMid36[24] , \wAMid36[23] , \wAMid36[22] , 
        \wAMid36[21] , \wAMid36[20] , \wAMid36[19] , \wAMid36[18] , 
        \wAMid36[17] , \wAMid36[16] , \wAMid36[15] , \wAMid36[14] , 
        \wAMid36[13] , \wAMid36[12] , \wAMid36[11] , \wAMid36[10] , 
        \wAMid36[9] , \wAMid36[8] , \wAMid36[7] , \wAMid36[6] , \wAMid36[5] , 
        \wAMid36[4] , \wAMid36[3] , \wAMid36[2] , \wAMid36[1] , \wAMid36[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid21[31] , \wAMid21[30] , \wAMid21[29] , \wAMid21[28] , 
        \wAMid21[27] , \wAMid21[26] , \wAMid21[25] , \wAMid21[24] , 
        \wAMid21[23] , \wAMid21[22] , \wAMid21[21] , \wAMid21[20] , 
        \wAMid21[19] , \wAMid21[18] , \wAMid21[17] , \wAMid21[16] , 
        \wAMid21[15] , \wAMid21[14] , \wAMid21[13] , \wAMid21[12] , 
        \wAMid21[11] , \wAMid21[10] , \wAMid21[9] , \wAMid21[8] , \wAMid21[7] , 
        \wAMid21[6] , \wAMid21[5] , \wAMid21[4] , \wAMid21[3] , \wAMid21[2] , 
        \wAMid21[1] , \wAMid21[0] }), .BIn({\wBMid21[31] , \wBMid21[30] , 
        \wBMid21[29] , \wBMid21[28] , \wBMid21[27] , \wBMid21[26] , 
        \wBMid21[25] , \wBMid21[24] , \wBMid21[23] , \wBMid21[22] , 
        \wBMid21[21] , \wBMid21[20] , \wBMid21[19] , \wBMid21[18] , 
        \wBMid21[17] , \wBMid21[16] , \wBMid21[15] , \wBMid21[14] , 
        \wBMid21[13] , \wBMid21[12] , \wBMid21[11] , \wBMid21[10] , 
        \wBMid21[9] , \wBMid21[8] , \wBMid21[7] , \wBMid21[6] , \wBMid21[5] , 
        \wBMid21[4] , \wBMid21[3] , \wBMid21[2] , \wBMid21[1] , \wBMid21[0] }), 
        .HiOut({\wRegInB21[31] , \wRegInB21[30] , \wRegInB21[29] , 
        \wRegInB21[28] , \wRegInB21[27] , \wRegInB21[26] , \wRegInB21[25] , 
        \wRegInB21[24] , \wRegInB21[23] , \wRegInB21[22] , \wRegInB21[21] , 
        \wRegInB21[20] , \wRegInB21[19] , \wRegInB21[18] , \wRegInB21[17] , 
        \wRegInB21[16] , \wRegInB21[15] , \wRegInB21[14] , \wRegInB21[13] , 
        \wRegInB21[12] , \wRegInB21[11] , \wRegInB21[10] , \wRegInB21[9] , 
        \wRegInB21[8] , \wRegInB21[7] , \wRegInB21[6] , \wRegInB21[5] , 
        \wRegInB21[4] , \wRegInB21[3] , \wRegInB21[2] , \wRegInB21[1] , 
        \wRegInB21[0] }), .LoOut({\wRegInA22[31] , \wRegInA22[30] , 
        \wRegInA22[29] , \wRegInA22[28] , \wRegInA22[27] , \wRegInA22[26] , 
        \wRegInA22[25] , \wRegInA22[24] , \wRegInA22[23] , \wRegInA22[22] , 
        \wRegInA22[21] , \wRegInA22[20] , \wRegInA22[19] , \wRegInA22[18] , 
        \wRegInA22[17] , \wRegInA22[16] , \wRegInA22[15] , \wRegInA22[14] , 
        \wRegInA22[13] , \wRegInA22[12] , \wRegInA22[11] , \wRegInA22[10] , 
        \wRegInA22[9] , \wRegInA22[8] , \wRegInA22[7] , \wRegInA22[6] , 
        \wRegInA22[5] , \wRegInA22[4] , \wRegInA22[3] , \wRegInA22[2] , 
        \wRegInA22[1] , \wRegInA22[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_44 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink45[31] , \ScanLink45[30] , \ScanLink45[29] , 
        \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , \ScanLink45[25] , 
        \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , \ScanLink45[21] , 
        \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , \ScanLink45[17] , 
        \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , \ScanLink45[13] , 
        \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , \ScanLink45[9] , 
        \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , \ScanLink45[5] , 
        \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , \ScanLink45[1] , 
        \ScanLink45[0] }), .ScanOut({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB105[31] , \wRegInB105[30] , 
        \wRegInB105[29] , \wRegInB105[28] , \wRegInB105[27] , \wRegInB105[26] , 
        \wRegInB105[25] , \wRegInB105[24] , \wRegInB105[23] , \wRegInB105[22] , 
        \wRegInB105[21] , \wRegInB105[20] , \wRegInB105[19] , \wRegInB105[18] , 
        \wRegInB105[17] , \wRegInB105[16] , \wRegInB105[15] , \wRegInB105[14] , 
        \wRegInB105[13] , \wRegInB105[12] , \wRegInB105[11] , \wRegInB105[10] , 
        \wRegInB105[9] , \wRegInB105[8] , \wRegInB105[7] , \wRegInB105[6] , 
        \wRegInB105[5] , \wRegInB105[4] , \wRegInB105[3] , \wRegInB105[2] , 
        \wRegInB105[1] , \wRegInB105[0] }), .Out({\wBIn105[31] , \wBIn105[30] , 
        \wBIn105[29] , \wBIn105[28] , \wBIn105[27] , \wBIn105[26] , 
        \wBIn105[25] , \wBIn105[24] , \wBIn105[23] , \wBIn105[22] , 
        \wBIn105[21] , \wBIn105[20] , \wBIn105[19] , \wBIn105[18] , 
        \wBIn105[17] , \wBIn105[16] , \wBIn105[15] , \wBIn105[14] , 
        \wBIn105[13] , \wBIn105[12] , \wBIn105[11] , \wBIn105[10] , 
        \wBIn105[9] , \wBIn105[8] , \wBIn105[7] , \wBIn105[6] , \wBIn105[5] , 
        \wBIn105[4] , \wBIn105[3] , \wBIn105[2] , \wBIn105[1] , \wBIn105[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_224 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink225[31] , \ScanLink225[30] , \ScanLink225[29] , 
        \ScanLink225[28] , \ScanLink225[27] , \ScanLink225[26] , 
        \ScanLink225[25] , \ScanLink225[24] , \ScanLink225[23] , 
        \ScanLink225[22] , \ScanLink225[21] , \ScanLink225[20] , 
        \ScanLink225[19] , \ScanLink225[18] , \ScanLink225[17] , 
        \ScanLink225[16] , \ScanLink225[15] , \ScanLink225[14] , 
        \ScanLink225[13] , \ScanLink225[12] , \ScanLink225[11] , 
        \ScanLink225[10] , \ScanLink225[9] , \ScanLink225[8] , 
        \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , \ScanLink225[4] , 
        \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , \ScanLink225[0] 
        }), .ScanOut({\ScanLink224[31] , \ScanLink224[30] , \ScanLink224[29] , 
        \ScanLink224[28] , \ScanLink224[27] , \ScanLink224[26] , 
        \ScanLink224[25] , \ScanLink224[24] , \ScanLink224[23] , 
        \ScanLink224[22] , \ScanLink224[21] , \ScanLink224[20] , 
        \ScanLink224[19] , \ScanLink224[18] , \ScanLink224[17] , 
        \ScanLink224[16] , \ScanLink224[15] , \ScanLink224[14] , 
        \ScanLink224[13] , \ScanLink224[12] , \ScanLink224[11] , 
        \ScanLink224[10] , \ScanLink224[9] , \ScanLink224[8] , 
        \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , \ScanLink224[4] , 
        \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , \ScanLink224[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB15[31] , \wRegInB15[30] , \wRegInB15[29] , 
        \wRegInB15[28] , \wRegInB15[27] , \wRegInB15[26] , \wRegInB15[25] , 
        \wRegInB15[24] , \wRegInB15[23] , \wRegInB15[22] , \wRegInB15[21] , 
        \wRegInB15[20] , \wRegInB15[19] , \wRegInB15[18] , \wRegInB15[17] , 
        \wRegInB15[16] , \wRegInB15[15] , \wRegInB15[14] , \wRegInB15[13] , 
        \wRegInB15[12] , \wRegInB15[11] , \wRegInB15[10] , \wRegInB15[9] , 
        \wRegInB15[8] , \wRegInB15[7] , \wRegInB15[6] , \wRegInB15[5] , 
        \wRegInB15[4] , \wRegInB15[3] , \wRegInB15[2] , \wRegInB15[1] , 
        \wRegInB15[0] }), .Out({\wBIn15[31] , \wBIn15[30] , \wBIn15[29] , 
        \wBIn15[28] , \wBIn15[27] , \wBIn15[26] , \wBIn15[25] , \wBIn15[24] , 
        \wBIn15[23] , \wBIn15[22] , \wBIn15[21] , \wBIn15[20] , \wBIn15[19] , 
        \wBIn15[18] , \wBIn15[17] , \wBIn15[16] , \wBIn15[15] , \wBIn15[14] , 
        \wBIn15[13] , \wBIn15[12] , \wBIn15[11] , \wBIn15[10] , \wBIn15[9] , 
        \wBIn15[8] , \wBIn15[7] , \wBIn15[6] , \wBIn15[5] , \wBIn15[4] , 
        \wBIn15[3] , \wBIn15[2] , \wBIn15[1] , \wBIn15[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_114 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink115[31] , \ScanLink115[30] , \ScanLink115[29] , 
        \ScanLink115[28] , \ScanLink115[27] , \ScanLink115[26] , 
        \ScanLink115[25] , \ScanLink115[24] , \ScanLink115[23] , 
        \ScanLink115[22] , \ScanLink115[21] , \ScanLink115[20] , 
        \ScanLink115[19] , \ScanLink115[18] , \ScanLink115[17] , 
        \ScanLink115[16] , \ScanLink115[15] , \ScanLink115[14] , 
        \ScanLink115[13] , \ScanLink115[12] , \ScanLink115[11] , 
        \ScanLink115[10] , \ScanLink115[9] , \ScanLink115[8] , 
        \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , \ScanLink115[4] , 
        \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , \ScanLink115[0] 
        }), .ScanOut({\ScanLink114[31] , \ScanLink114[30] , \ScanLink114[29] , 
        \ScanLink114[28] , \ScanLink114[27] , \ScanLink114[26] , 
        \ScanLink114[25] , \ScanLink114[24] , \ScanLink114[23] , 
        \ScanLink114[22] , \ScanLink114[21] , \ScanLink114[20] , 
        \ScanLink114[19] , \ScanLink114[18] , \ScanLink114[17] , 
        \ScanLink114[16] , \ScanLink114[15] , \ScanLink114[14] , 
        \ScanLink114[13] , \ScanLink114[12] , \ScanLink114[11] , 
        \ScanLink114[10] , \ScanLink114[9] , \ScanLink114[8] , 
        \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , \ScanLink114[4] , 
        \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , \ScanLink114[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB70[31] , \wRegInB70[30] , \wRegInB70[29] , 
        \wRegInB70[28] , \wRegInB70[27] , \wRegInB70[26] , \wRegInB70[25] , 
        \wRegInB70[24] , \wRegInB70[23] , \wRegInB70[22] , \wRegInB70[21] , 
        \wRegInB70[20] , \wRegInB70[19] , \wRegInB70[18] , \wRegInB70[17] , 
        \wRegInB70[16] , \wRegInB70[15] , \wRegInB70[14] , \wRegInB70[13] , 
        \wRegInB70[12] , \wRegInB70[11] , \wRegInB70[10] , \wRegInB70[9] , 
        \wRegInB70[8] , \wRegInB70[7] , \wRegInB70[6] , \wRegInB70[5] , 
        \wRegInB70[4] , \wRegInB70[3] , \wRegInB70[2] , \wRegInB70[1] , 
        \wRegInB70[0] }), .Out({\wBIn70[31] , \wBIn70[30] , \wBIn70[29] , 
        \wBIn70[28] , \wBIn70[27] , \wBIn70[26] , \wBIn70[25] , \wBIn70[24] , 
        \wBIn70[23] , \wBIn70[22] , \wBIn70[21] , \wBIn70[20] , \wBIn70[19] , 
        \wBIn70[18] , \wBIn70[17] , \wBIn70[16] , \wBIn70[15] , \wBIn70[14] , 
        \wBIn70[13] , \wBIn70[12] , \wBIn70[11] , \wBIn70[10] , \wBIn70[9] , 
        \wBIn70[8] , \wBIn70[7] , \wBIn70[6] , \wBIn70[5] , \wBIn70[4] , 
        \wBIn70[3] , \wBIn70[2] , \wBIn70[1] , \wBIn70[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_203 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink204[31] , \ScanLink204[30] , \ScanLink204[29] , 
        \ScanLink204[28] , \ScanLink204[27] , \ScanLink204[26] , 
        \ScanLink204[25] , \ScanLink204[24] , \ScanLink204[23] , 
        \ScanLink204[22] , \ScanLink204[21] , \ScanLink204[20] , 
        \ScanLink204[19] , \ScanLink204[18] , \ScanLink204[17] , 
        \ScanLink204[16] , \ScanLink204[15] , \ScanLink204[14] , 
        \ScanLink204[13] , \ScanLink204[12] , \ScanLink204[11] , 
        \ScanLink204[10] , \ScanLink204[9] , \ScanLink204[8] , 
        \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , \ScanLink204[4] , 
        \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , \ScanLink204[0] 
        }), .ScanOut({\ScanLink203[31] , \ScanLink203[30] , \ScanLink203[29] , 
        \ScanLink203[28] , \ScanLink203[27] , \ScanLink203[26] , 
        \ScanLink203[25] , \ScanLink203[24] , \ScanLink203[23] , 
        \ScanLink203[22] , \ScanLink203[21] , \ScanLink203[20] , 
        \ScanLink203[19] , \ScanLink203[18] , \ScanLink203[17] , 
        \ScanLink203[16] , \ScanLink203[15] , \ScanLink203[14] , 
        \ScanLink203[13] , \ScanLink203[12] , \ScanLink203[11] , 
        \ScanLink203[10] , \ScanLink203[9] , \ScanLink203[8] , 
        \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , \ScanLink203[4] , 
        \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , \ScanLink203[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA26[31] , \wRegInA26[30] , \wRegInA26[29] , 
        \wRegInA26[28] , \wRegInA26[27] , \wRegInA26[26] , \wRegInA26[25] , 
        \wRegInA26[24] , \wRegInA26[23] , \wRegInA26[22] , \wRegInA26[21] , 
        \wRegInA26[20] , \wRegInA26[19] , \wRegInA26[18] , \wRegInA26[17] , 
        \wRegInA26[16] , \wRegInA26[15] , \wRegInA26[14] , \wRegInA26[13] , 
        \wRegInA26[12] , \wRegInA26[11] , \wRegInA26[10] , \wRegInA26[9] , 
        \wRegInA26[8] , \wRegInA26[7] , \wRegInA26[6] , \wRegInA26[5] , 
        \wRegInA26[4] , \wRegInA26[3] , \wRegInA26[2] , \wRegInA26[1] , 
        \wRegInA26[0] }), .Out({\wAIn26[31] , \wAIn26[30] , \wAIn26[29] , 
        \wAIn26[28] , \wAIn26[27] , \wAIn26[26] , \wAIn26[25] , \wAIn26[24] , 
        \wAIn26[23] , \wAIn26[22] , \wAIn26[21] , \wAIn26[20] , \wAIn26[19] , 
        \wAIn26[18] , \wAIn26[17] , \wAIn26[16] , \wAIn26[15] , \wAIn26[14] , 
        \wAIn26[13] , \wAIn26[12] , \wAIn26[11] , \wAIn26[10] , \wAIn26[9] , 
        \wAIn26[8] , \wAIn26[7] , \wAIn26[6] , \wAIn26[5] , \wAIn26[4] , 
        \wAIn26[3] , \wAIn26[2] , \wAIn26[1] , \wAIn26[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_7 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[31] , \ScanLink8[30] , \ScanLink8[29] , 
        \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , \ScanLink8[25] , 
        \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , \ScanLink8[21] , 
        \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , \ScanLink8[17] , 
        \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , \ScanLink8[13] , 
        \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , \ScanLink8[9] , 
        \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA124[31] , \wRegInA124[30] , 
        \wRegInA124[29] , \wRegInA124[28] , \wRegInA124[27] , \wRegInA124[26] , 
        \wRegInA124[25] , \wRegInA124[24] , \wRegInA124[23] , \wRegInA124[22] , 
        \wRegInA124[21] , \wRegInA124[20] , \wRegInA124[19] , \wRegInA124[18] , 
        \wRegInA124[17] , \wRegInA124[16] , \wRegInA124[15] , \wRegInA124[14] , 
        \wRegInA124[13] , \wRegInA124[12] , \wRegInA124[11] , \wRegInA124[10] , 
        \wRegInA124[9] , \wRegInA124[8] , \wRegInA124[7] , \wRegInA124[6] , 
        \wRegInA124[5] , \wRegInA124[4] , \wRegInA124[3] , \wRegInA124[2] , 
        \wRegInA124[1] , \wRegInA124[0] }), .Out({\wAIn124[31] , \wAIn124[30] , 
        \wAIn124[29] , \wAIn124[28] , \wAIn124[27] , \wAIn124[26] , 
        \wAIn124[25] , \wAIn124[24] , \wAIn124[23] , \wAIn124[22] , 
        \wAIn124[21] , \wAIn124[20] , \wAIn124[19] , \wAIn124[18] , 
        \wAIn124[17] , \wAIn124[16] , \wAIn124[15] , \wAIn124[14] , 
        \wAIn124[13] , \wAIn124[12] , \wAIn124[11] , \wAIn124[10] , 
        \wAIn124[9] , \wAIn124[8] , \wAIn124[7] , \wAIn124[6] , \wAIn124[5] , 
        \wAIn124[4] , \wAIn124[3] , \wAIn124[2] , \wAIn124[1] , \wAIn124[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn88[31] , \wAIn88[30] , \wAIn88[29] , \wAIn88[28] , \wAIn88[27] , 
        \wAIn88[26] , \wAIn88[25] , \wAIn88[24] , \wAIn88[23] , \wAIn88[22] , 
        \wAIn88[21] , \wAIn88[20] , \wAIn88[19] , \wAIn88[18] , \wAIn88[17] , 
        \wAIn88[16] , \wAIn88[15] , \wAIn88[14] , \wAIn88[13] , \wAIn88[12] , 
        \wAIn88[11] , \wAIn88[10] , \wAIn88[9] , \wAIn88[8] , \wAIn88[7] , 
        \wAIn88[6] , \wAIn88[5] , \wAIn88[4] , \wAIn88[3] , \wAIn88[2] , 
        \wAIn88[1] , \wAIn88[0] }), .BIn({\wBIn88[31] , \wBIn88[30] , 
        \wBIn88[29] , \wBIn88[28] , \wBIn88[27] , \wBIn88[26] , \wBIn88[25] , 
        \wBIn88[24] , \wBIn88[23] , \wBIn88[22] , \wBIn88[21] , \wBIn88[20] , 
        \wBIn88[19] , \wBIn88[18] , \wBIn88[17] , \wBIn88[16] , \wBIn88[15] , 
        \wBIn88[14] , \wBIn88[13] , \wBIn88[12] , \wBIn88[11] , \wBIn88[10] , 
        \wBIn88[9] , \wBIn88[8] , \wBIn88[7] , \wBIn88[6] , \wBIn88[5] , 
        \wBIn88[4] , \wBIn88[3] , \wBIn88[2] , \wBIn88[1] , \wBIn88[0] }), 
        .HiOut({\wBMid87[31] , \wBMid87[30] , \wBMid87[29] , \wBMid87[28] , 
        \wBMid87[27] , \wBMid87[26] , \wBMid87[25] , \wBMid87[24] , 
        \wBMid87[23] , \wBMid87[22] , \wBMid87[21] , \wBMid87[20] , 
        \wBMid87[19] , \wBMid87[18] , \wBMid87[17] , \wBMid87[16] , 
        \wBMid87[15] , \wBMid87[14] , \wBMid87[13] , \wBMid87[12] , 
        \wBMid87[11] , \wBMid87[10] , \wBMid87[9] , \wBMid87[8] , \wBMid87[7] , 
        \wBMid87[6] , \wBMid87[5] , \wBMid87[4] , \wBMid87[3] , \wBMid87[2] , 
        \wBMid87[1] , \wBMid87[0] }), .LoOut({\wAMid88[31] , \wAMid88[30] , 
        \wAMid88[29] , \wAMid88[28] , \wAMid88[27] , \wAMid88[26] , 
        \wAMid88[25] , \wAMid88[24] , \wAMid88[23] , \wAMid88[22] , 
        \wAMid88[21] , \wAMid88[20] , \wAMid88[19] , \wAMid88[18] , 
        \wAMid88[17] , \wAMid88[16] , \wAMid88[15] , \wAMid88[14] , 
        \wAMid88[13] , \wAMid88[12] , \wAMid88[11] , \wAMid88[10] , 
        \wAMid88[9] , \wAMid88[8] , \wAMid88[7] , \wAMid88[6] , \wAMid88[5] , 
        \wAMid88[4] , \wAMid88[3] , \wAMid88[2] , \wAMid88[1] , \wAMid88[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_133 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink134[31] , \ScanLink134[30] , \ScanLink134[29] , 
        \ScanLink134[28] , \ScanLink134[27] , \ScanLink134[26] , 
        \ScanLink134[25] , \ScanLink134[24] , \ScanLink134[23] , 
        \ScanLink134[22] , \ScanLink134[21] , \ScanLink134[20] , 
        \ScanLink134[19] , \ScanLink134[18] , \ScanLink134[17] , 
        \ScanLink134[16] , \ScanLink134[15] , \ScanLink134[14] , 
        \ScanLink134[13] , \ScanLink134[12] , \ScanLink134[11] , 
        \ScanLink134[10] , \ScanLink134[9] , \ScanLink134[8] , 
        \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , \ScanLink134[4] , 
        \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , \ScanLink134[0] 
        }), .ScanOut({\ScanLink133[31] , \ScanLink133[30] , \ScanLink133[29] , 
        \ScanLink133[28] , \ScanLink133[27] , \ScanLink133[26] , 
        \ScanLink133[25] , \ScanLink133[24] , \ScanLink133[23] , 
        \ScanLink133[22] , \ScanLink133[21] , \ScanLink133[20] , 
        \ScanLink133[19] , \ScanLink133[18] , \ScanLink133[17] , 
        \ScanLink133[16] , \ScanLink133[15] , \ScanLink133[14] , 
        \ScanLink133[13] , \ScanLink133[12] , \ScanLink133[11] , 
        \ScanLink133[10] , \ScanLink133[9] , \ScanLink133[8] , 
        \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , \ScanLink133[4] , 
        \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , \ScanLink133[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA61[31] , \wRegInA61[30] , \wRegInA61[29] , 
        \wRegInA61[28] , \wRegInA61[27] , \wRegInA61[26] , \wRegInA61[25] , 
        \wRegInA61[24] , \wRegInA61[23] , \wRegInA61[22] , \wRegInA61[21] , 
        \wRegInA61[20] , \wRegInA61[19] , \wRegInA61[18] , \wRegInA61[17] , 
        \wRegInA61[16] , \wRegInA61[15] , \wRegInA61[14] , \wRegInA61[13] , 
        \wRegInA61[12] , \wRegInA61[11] , \wRegInA61[10] , \wRegInA61[9] , 
        \wRegInA61[8] , \wRegInA61[7] , \wRegInA61[6] , \wRegInA61[5] , 
        \wRegInA61[4] , \wRegInA61[3] , \wRegInA61[2] , \wRegInA61[1] , 
        \wRegInA61[0] }), .Out({\wAIn61[31] , \wAIn61[30] , \wAIn61[29] , 
        \wAIn61[28] , \wAIn61[27] , \wAIn61[26] , \wAIn61[25] , \wAIn61[24] , 
        \wAIn61[23] , \wAIn61[22] , \wAIn61[21] , \wAIn61[20] , \wAIn61[19] , 
        \wAIn61[18] , \wAIn61[17] , \wAIn61[16] , \wAIn61[15] , \wAIn61[14] , 
        \wAIn61[13] , \wAIn61[12] , \wAIn61[11] , \wAIn61[10] , \wAIn61[9] , 
        \wAIn61[8] , \wAIn61[7] , \wAIn61[6] , \wAIn61[5] , \wAIn61[4] , 
        \wAIn61[3] , \wAIn61[2] , \wAIn61[1] , \wAIn61[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_63 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink64[31] , \ScanLink64[30] , \ScanLink64[29] , 
        \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , \ScanLink64[25] , 
        \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , \ScanLink64[21] , 
        \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , \ScanLink64[17] , 
        \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , \ScanLink64[13] , 
        \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , \ScanLink64[9] , 
        \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , \ScanLink64[5] , 
        \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , \ScanLink64[1] , 
        \ScanLink64[0] }), .ScanOut({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA96[31] , \wRegInA96[30] , 
        \wRegInA96[29] , \wRegInA96[28] , \wRegInA96[27] , \wRegInA96[26] , 
        \wRegInA96[25] , \wRegInA96[24] , \wRegInA96[23] , \wRegInA96[22] , 
        \wRegInA96[21] , \wRegInA96[20] , \wRegInA96[19] , \wRegInA96[18] , 
        \wRegInA96[17] , \wRegInA96[16] , \wRegInA96[15] , \wRegInA96[14] , 
        \wRegInA96[13] , \wRegInA96[12] , \wRegInA96[11] , \wRegInA96[10] , 
        \wRegInA96[9] , \wRegInA96[8] , \wRegInA96[7] , \wRegInA96[6] , 
        \wRegInA96[5] , \wRegInA96[4] , \wRegInA96[3] , \wRegInA96[2] , 
        \wRegInA96[1] , \wRegInA96[0] }), .Out({\wAIn96[31] , \wAIn96[30] , 
        \wAIn96[29] , \wAIn96[28] , \wAIn96[27] , \wAIn96[26] , \wAIn96[25] , 
        \wAIn96[24] , \wAIn96[23] , \wAIn96[22] , \wAIn96[21] , \wAIn96[20] , 
        \wAIn96[19] , \wAIn96[18] , \wAIn96[17] , \wAIn96[16] , \wAIn96[15] , 
        \wAIn96[14] , \wAIn96[13] , \wAIn96[12] , \wAIn96[11] , \wAIn96[10] , 
        \wAIn96[9] , \wAIn96[8] , \wAIn96[7] , \wAIn96[6] , \wAIn96[5] , 
        \wAIn96[4] , \wAIn96[3] , \wAIn96[2] , \wAIn96[1] , \wAIn96[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid33[31] , \wAMid33[30] , \wAMid33[29] , \wAMid33[28] , 
        \wAMid33[27] , \wAMid33[26] , \wAMid33[25] , \wAMid33[24] , 
        \wAMid33[23] , \wAMid33[22] , \wAMid33[21] , \wAMid33[20] , 
        \wAMid33[19] , \wAMid33[18] , \wAMid33[17] , \wAMid33[16] , 
        \wAMid33[15] , \wAMid33[14] , \wAMid33[13] , \wAMid33[12] , 
        \wAMid33[11] , \wAMid33[10] , \wAMid33[9] , \wAMid33[8] , \wAMid33[7] , 
        \wAMid33[6] , \wAMid33[5] , \wAMid33[4] , \wAMid33[3] , \wAMid33[2] , 
        \wAMid33[1] , \wAMid33[0] }), .BIn({\wBMid33[31] , \wBMid33[30] , 
        \wBMid33[29] , \wBMid33[28] , \wBMid33[27] , \wBMid33[26] , 
        \wBMid33[25] , \wBMid33[24] , \wBMid33[23] , \wBMid33[22] , 
        \wBMid33[21] , \wBMid33[20] , \wBMid33[19] , \wBMid33[18] , 
        \wBMid33[17] , \wBMid33[16] , \wBMid33[15] , \wBMid33[14] , 
        \wBMid33[13] , \wBMid33[12] , \wBMid33[11] , \wBMid33[10] , 
        \wBMid33[9] , \wBMid33[8] , \wBMid33[7] , \wBMid33[6] , \wBMid33[5] , 
        \wBMid33[4] , \wBMid33[3] , \wBMid33[2] , \wBMid33[1] , \wBMid33[0] }), 
        .HiOut({\wRegInB33[31] , \wRegInB33[30] , \wRegInB33[29] , 
        \wRegInB33[28] , \wRegInB33[27] , \wRegInB33[26] , \wRegInB33[25] , 
        \wRegInB33[24] , \wRegInB33[23] , \wRegInB33[22] , \wRegInB33[21] , 
        \wRegInB33[20] , \wRegInB33[19] , \wRegInB33[18] , \wRegInB33[17] , 
        \wRegInB33[16] , \wRegInB33[15] , \wRegInB33[14] , \wRegInB33[13] , 
        \wRegInB33[12] , \wRegInB33[11] , \wRegInB33[10] , \wRegInB33[9] , 
        \wRegInB33[8] , \wRegInB33[7] , \wRegInB33[6] , \wRegInB33[5] , 
        \wRegInB33[4] , \wRegInB33[3] , \wRegInB33[2] , \wRegInB33[1] , 
        \wRegInB33[0] }), .LoOut({\wRegInA34[31] , \wRegInA34[30] , 
        \wRegInA34[29] , \wRegInA34[28] , \wRegInA34[27] , \wRegInA34[26] , 
        \wRegInA34[25] , \wRegInA34[24] , \wRegInA34[23] , \wRegInA34[22] , 
        \wRegInA34[21] , \wRegInA34[20] , \wRegInA34[19] , \wRegInA34[18] , 
        \wRegInA34[17] , \wRegInA34[16] , \wRegInA34[15] , \wRegInA34[14] , 
        \wRegInA34[13] , \wRegInA34[12] , \wRegInA34[11] , \wRegInA34[10] , 
        \wRegInA34[9] , \wRegInA34[8] , \wRegInA34[7] , \wRegInA34[6] , 
        \wRegInA34[5] , \wRegInA34[4] , \wRegInA34[3] , \wRegInA34[2] , 
        \wRegInA34[1] , \wRegInA34[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_106 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink107[31] , \ScanLink107[30] , \ScanLink107[29] , 
        \ScanLink107[28] , \ScanLink107[27] , \ScanLink107[26] , 
        \ScanLink107[25] , \ScanLink107[24] , \ScanLink107[23] , 
        \ScanLink107[22] , \ScanLink107[21] , \ScanLink107[20] , 
        \ScanLink107[19] , \ScanLink107[18] , \ScanLink107[17] , 
        \ScanLink107[16] , \ScanLink107[15] , \ScanLink107[14] , 
        \ScanLink107[13] , \ScanLink107[12] , \ScanLink107[11] , 
        \ScanLink107[10] , \ScanLink107[9] , \ScanLink107[8] , 
        \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , \ScanLink107[4] , 
        \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , \ScanLink107[0] 
        }), .ScanOut({\ScanLink106[31] , \ScanLink106[30] , \ScanLink106[29] , 
        \ScanLink106[28] , \ScanLink106[27] , \ScanLink106[26] , 
        \ScanLink106[25] , \ScanLink106[24] , \ScanLink106[23] , 
        \ScanLink106[22] , \ScanLink106[21] , \ScanLink106[20] , 
        \ScanLink106[19] , \ScanLink106[18] , \ScanLink106[17] , 
        \ScanLink106[16] , \ScanLink106[15] , \ScanLink106[14] , 
        \ScanLink106[13] , \ScanLink106[12] , \ScanLink106[11] , 
        \ScanLink106[10] , \ScanLink106[9] , \ScanLink106[8] , 
        \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , \ScanLink106[4] , 
        \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , \ScanLink106[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB74[31] , \wRegInB74[30] , \wRegInB74[29] , 
        \wRegInB74[28] , \wRegInB74[27] , \wRegInB74[26] , \wRegInB74[25] , 
        \wRegInB74[24] , \wRegInB74[23] , \wRegInB74[22] , \wRegInB74[21] , 
        \wRegInB74[20] , \wRegInB74[19] , \wRegInB74[18] , \wRegInB74[17] , 
        \wRegInB74[16] , \wRegInB74[15] , \wRegInB74[14] , \wRegInB74[13] , 
        \wRegInB74[12] , \wRegInB74[11] , \wRegInB74[10] , \wRegInB74[9] , 
        \wRegInB74[8] , \wRegInB74[7] , \wRegInB74[6] , \wRegInB74[5] , 
        \wRegInB74[4] , \wRegInB74[3] , \wRegInB74[2] , \wRegInB74[1] , 
        \wRegInB74[0] }), .Out({\wBIn74[31] , \wBIn74[30] , \wBIn74[29] , 
        \wBIn74[28] , \wBIn74[27] , \wBIn74[26] , \wBIn74[25] , \wBIn74[24] , 
        \wBIn74[23] , \wBIn74[22] , \wBIn74[21] , \wBIn74[20] , \wBIn74[19] , 
        \wBIn74[18] , \wBIn74[17] , \wBIn74[16] , \wBIn74[15] , \wBIn74[14] , 
        \wBIn74[13] , \wBIn74[12] , \wBIn74[11] , \wBIn74[10] , \wBIn74[9] , 
        \wBIn74[8] , \wBIn74[7] , \wBIn74[6] , \wBIn74[5] , \wBIn74[4] , 
        \wBIn74[3] , \wBIn74[2] , \wBIn74[1] , \wBIn74[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_56 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink57[31] , \ScanLink57[30] , \ScanLink57[29] , 
        \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , \ScanLink57[25] , 
        \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , \ScanLink57[21] , 
        \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , \ScanLink57[17] , 
        \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , \ScanLink57[13] , 
        \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , \ScanLink57[9] , 
        \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , \ScanLink57[5] , 
        \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , \ScanLink57[1] , 
        \ScanLink57[0] }), .ScanOut({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB99[31] , \wRegInB99[30] , 
        \wRegInB99[29] , \wRegInB99[28] , \wRegInB99[27] , \wRegInB99[26] , 
        \wRegInB99[25] , \wRegInB99[24] , \wRegInB99[23] , \wRegInB99[22] , 
        \wRegInB99[21] , \wRegInB99[20] , \wRegInB99[19] , \wRegInB99[18] , 
        \wRegInB99[17] , \wRegInB99[16] , \wRegInB99[15] , \wRegInB99[14] , 
        \wRegInB99[13] , \wRegInB99[12] , \wRegInB99[11] , \wRegInB99[10] , 
        \wRegInB99[9] , \wRegInB99[8] , \wRegInB99[7] , \wRegInB99[6] , 
        \wRegInB99[5] , \wRegInB99[4] , \wRegInB99[3] , \wRegInB99[2] , 
        \wRegInB99[1] , \wRegInB99[0] }), .Out({\wBIn99[31] , \wBIn99[30] , 
        \wBIn99[29] , \wBIn99[28] , \wBIn99[27] , \wBIn99[26] , \wBIn99[25] , 
        \wBIn99[24] , \wBIn99[23] , \wBIn99[22] , \wBIn99[21] , \wBIn99[20] , 
        \wBIn99[19] , \wBIn99[18] , \wBIn99[17] , \wBIn99[16] , \wBIn99[15] , 
        \wBIn99[14] , \wBIn99[13] , \wBIn99[12] , \wBIn99[11] , \wBIn99[10] , 
        \wBIn99[9] , \wBIn99[8] , \wBIn99[7] , \wBIn99[6] , \wBIn99[5] , 
        \wBIn99[4] , \wBIn99[3] , \wBIn99[2] , \wBIn99[1] , \wBIn99[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_236 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink237[31] , \ScanLink237[30] , \ScanLink237[29] , 
        \ScanLink237[28] , \ScanLink237[27] , \ScanLink237[26] , 
        \ScanLink237[25] , \ScanLink237[24] , \ScanLink237[23] , 
        \ScanLink237[22] , \ScanLink237[21] , \ScanLink237[20] , 
        \ScanLink237[19] , \ScanLink237[18] , \ScanLink237[17] , 
        \ScanLink237[16] , \ScanLink237[15] , \ScanLink237[14] , 
        \ScanLink237[13] , \ScanLink237[12] , \ScanLink237[11] , 
        \ScanLink237[10] , \ScanLink237[9] , \ScanLink237[8] , 
        \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , \ScanLink237[4] , 
        \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , \ScanLink237[0] 
        }), .ScanOut({\ScanLink236[31] , \ScanLink236[30] , \ScanLink236[29] , 
        \ScanLink236[28] , \ScanLink236[27] , \ScanLink236[26] , 
        \ScanLink236[25] , \ScanLink236[24] , \ScanLink236[23] , 
        \ScanLink236[22] , \ScanLink236[21] , \ScanLink236[20] , 
        \ScanLink236[19] , \ScanLink236[18] , \ScanLink236[17] , 
        \ScanLink236[16] , \ScanLink236[15] , \ScanLink236[14] , 
        \ScanLink236[13] , \ScanLink236[12] , \ScanLink236[11] , 
        \ScanLink236[10] , \ScanLink236[9] , \ScanLink236[8] , 
        \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , \ScanLink236[4] , 
        \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , \ScanLink236[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB9[31] , \wRegInB9[30] , \wRegInB9[29] , \wRegInB9[28] , 
        \wRegInB9[27] , \wRegInB9[26] , \wRegInB9[25] , \wRegInB9[24] , 
        \wRegInB9[23] , \wRegInB9[22] , \wRegInB9[21] , \wRegInB9[20] , 
        \wRegInB9[19] , \wRegInB9[18] , \wRegInB9[17] , \wRegInB9[16] , 
        \wRegInB9[15] , \wRegInB9[14] , \wRegInB9[13] , \wRegInB9[12] , 
        \wRegInB9[11] , \wRegInB9[10] , \wRegInB9[9] , \wRegInB9[8] , 
        \wRegInB9[7] , \wRegInB9[6] , \wRegInB9[5] , \wRegInB9[4] , 
        \wRegInB9[3] , \wRegInB9[2] , \wRegInB9[1] , \wRegInB9[0] }), .Out({
        \wBIn9[31] , \wBIn9[30] , \wBIn9[29] , \wBIn9[28] , \wBIn9[27] , 
        \wBIn9[26] , \wBIn9[25] , \wBIn9[24] , \wBIn9[23] , \wBIn9[22] , 
        \wBIn9[21] , \wBIn9[20] , \wBIn9[19] , \wBIn9[18] , \wBIn9[17] , 
        \wBIn9[16] , \wBIn9[15] , \wBIn9[14] , \wBIn9[13] , \wBIn9[12] , 
        \wBIn9[11] , \wBIn9[10] , \wBIn9[9] , \wBIn9[8] , \wBIn9[7] , 
        \wBIn9[6] , \wBIn9[5] , \wBIn9[4] , \wBIn9[3] , \wBIn9[2] , \wBIn9[1] , 
        \wBIn9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_211 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink212[31] , \ScanLink212[30] , \ScanLink212[29] , 
        \ScanLink212[28] , \ScanLink212[27] , \ScanLink212[26] , 
        \ScanLink212[25] , \ScanLink212[24] , \ScanLink212[23] , 
        \ScanLink212[22] , \ScanLink212[21] , \ScanLink212[20] , 
        \ScanLink212[19] , \ScanLink212[18] , \ScanLink212[17] , 
        \ScanLink212[16] , \ScanLink212[15] , \ScanLink212[14] , 
        \ScanLink212[13] , \ScanLink212[12] , \ScanLink212[11] , 
        \ScanLink212[10] , \ScanLink212[9] , \ScanLink212[8] , 
        \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , \ScanLink212[4] , 
        \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , \ScanLink212[0] 
        }), .ScanOut({\ScanLink211[31] , \ScanLink211[30] , \ScanLink211[29] , 
        \ScanLink211[28] , \ScanLink211[27] , \ScanLink211[26] , 
        \ScanLink211[25] , \ScanLink211[24] , \ScanLink211[23] , 
        \ScanLink211[22] , \ScanLink211[21] , \ScanLink211[20] , 
        \ScanLink211[19] , \ScanLink211[18] , \ScanLink211[17] , 
        \ScanLink211[16] , \ScanLink211[15] , \ScanLink211[14] , 
        \ScanLink211[13] , \ScanLink211[12] , \ScanLink211[11] , 
        \ScanLink211[10] , \ScanLink211[9] , \ScanLink211[8] , 
        \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , \ScanLink211[4] , 
        \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , \ScanLink211[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA22[31] , \wRegInA22[30] , \wRegInA22[29] , 
        \wRegInA22[28] , \wRegInA22[27] , \wRegInA22[26] , \wRegInA22[25] , 
        \wRegInA22[24] , \wRegInA22[23] , \wRegInA22[22] , \wRegInA22[21] , 
        \wRegInA22[20] , \wRegInA22[19] , \wRegInA22[18] , \wRegInA22[17] , 
        \wRegInA22[16] , \wRegInA22[15] , \wRegInA22[14] , \wRegInA22[13] , 
        \wRegInA22[12] , \wRegInA22[11] , \wRegInA22[10] , \wRegInA22[9] , 
        \wRegInA22[8] , \wRegInA22[7] , \wRegInA22[6] , \wRegInA22[5] , 
        \wRegInA22[4] , \wRegInA22[3] , \wRegInA22[2] , \wRegInA22[1] , 
        \wRegInA22[0] }), .Out({\wAIn22[31] , \wAIn22[30] , \wAIn22[29] , 
        \wAIn22[28] , \wAIn22[27] , \wAIn22[26] , \wAIn22[25] , \wAIn22[24] , 
        \wAIn22[23] , \wAIn22[22] , \wAIn22[21] , \wAIn22[20] , \wAIn22[19] , 
        \wAIn22[18] , \wAIn22[17] , \wAIn22[16] , \wAIn22[15] , \wAIn22[14] , 
        \wAIn22[13] , \wAIn22[12] , \wAIn22[11] , \wAIn22[10] , \wAIn22[9] , 
        \wAIn22[8] , \wAIn22[7] , \wAIn22[6] , \wAIn22[5] , \wAIn22[4] , 
        \wAIn22[3] , \wAIn22[2] , \wAIn22[1] , \wAIn22[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn51[31] , \wAIn51[30] , \wAIn51[29] , \wAIn51[28] , \wAIn51[27] , 
        \wAIn51[26] , \wAIn51[25] , \wAIn51[24] , \wAIn51[23] , \wAIn51[22] , 
        \wAIn51[21] , \wAIn51[20] , \wAIn51[19] , \wAIn51[18] , \wAIn51[17] , 
        \wAIn51[16] , \wAIn51[15] , \wAIn51[14] , \wAIn51[13] , \wAIn51[12] , 
        \wAIn51[11] , \wAIn51[10] , \wAIn51[9] , \wAIn51[8] , \wAIn51[7] , 
        \wAIn51[6] , \wAIn51[5] , \wAIn51[4] , \wAIn51[3] , \wAIn51[2] , 
        \wAIn51[1] , \wAIn51[0] }), .BIn({\wBIn51[31] , \wBIn51[30] , 
        \wBIn51[29] , \wBIn51[28] , \wBIn51[27] , \wBIn51[26] , \wBIn51[25] , 
        \wBIn51[24] , \wBIn51[23] , \wBIn51[22] , \wBIn51[21] , \wBIn51[20] , 
        \wBIn51[19] , \wBIn51[18] , \wBIn51[17] , \wBIn51[16] , \wBIn51[15] , 
        \wBIn51[14] , \wBIn51[13] , \wBIn51[12] , \wBIn51[11] , \wBIn51[10] , 
        \wBIn51[9] , \wBIn51[8] , \wBIn51[7] , \wBIn51[6] , \wBIn51[5] , 
        \wBIn51[4] , \wBIn51[3] , \wBIn51[2] , \wBIn51[1] , \wBIn51[0] }), 
        .HiOut({\wBMid50[31] , \wBMid50[30] , \wBMid50[29] , \wBMid50[28] , 
        \wBMid50[27] , \wBMid50[26] , \wBMid50[25] , \wBMid50[24] , 
        \wBMid50[23] , \wBMid50[22] , \wBMid50[21] , \wBMid50[20] , 
        \wBMid50[19] , \wBMid50[18] , \wBMid50[17] , \wBMid50[16] , 
        \wBMid50[15] , \wBMid50[14] , \wBMid50[13] , \wBMid50[12] , 
        \wBMid50[11] , \wBMid50[10] , \wBMid50[9] , \wBMid50[8] , \wBMid50[7] , 
        \wBMid50[6] , \wBMid50[5] , \wBMid50[4] , \wBMid50[3] , \wBMid50[2] , 
        \wBMid50[1] , \wBMid50[0] }), .LoOut({\wAMid51[31] , \wAMid51[30] , 
        \wAMid51[29] , \wAMid51[28] , \wAMid51[27] , \wAMid51[26] , 
        \wAMid51[25] , \wAMid51[24] , \wAMid51[23] , \wAMid51[22] , 
        \wAMid51[21] , \wAMid51[20] , \wAMid51[19] , \wAMid51[18] , 
        \wAMid51[17] , \wAMid51[16] , \wAMid51[15] , \wAMid51[14] , 
        \wAMid51[13] , \wAMid51[12] , \wAMid51[11] , \wAMid51[10] , 
        \wAMid51[9] , \wAMid51[8] , \wAMid51[7] , \wAMid51[6] , \wAMid51[5] , 
        \wAMid51[4] , \wAMid51[3] , \wAMid51[2] , \wAMid51[1] , \wAMid51[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn76[31] , \wAIn76[30] , \wAIn76[29] , \wAIn76[28] , \wAIn76[27] , 
        \wAIn76[26] , \wAIn76[25] , \wAIn76[24] , \wAIn76[23] , \wAIn76[22] , 
        \wAIn76[21] , \wAIn76[20] , \wAIn76[19] , \wAIn76[18] , \wAIn76[17] , 
        \wAIn76[16] , \wAIn76[15] , \wAIn76[14] , \wAIn76[13] , \wAIn76[12] , 
        \wAIn76[11] , \wAIn76[10] , \wAIn76[9] , \wAIn76[8] , \wAIn76[7] , 
        \wAIn76[6] , \wAIn76[5] , \wAIn76[4] , \wAIn76[3] , \wAIn76[2] , 
        \wAIn76[1] , \wAIn76[0] }), .BIn({\wBIn76[31] , \wBIn76[30] , 
        \wBIn76[29] , \wBIn76[28] , \wBIn76[27] , \wBIn76[26] , \wBIn76[25] , 
        \wBIn76[24] , \wBIn76[23] , \wBIn76[22] , \wBIn76[21] , \wBIn76[20] , 
        \wBIn76[19] , \wBIn76[18] , \wBIn76[17] , \wBIn76[16] , \wBIn76[15] , 
        \wBIn76[14] , \wBIn76[13] , \wBIn76[12] , \wBIn76[11] , \wBIn76[10] , 
        \wBIn76[9] , \wBIn76[8] , \wBIn76[7] , \wBIn76[6] , \wBIn76[5] , 
        \wBIn76[4] , \wBIn76[3] , \wBIn76[2] , \wBIn76[1] , \wBIn76[0] }), 
        .HiOut({\wBMid75[31] , \wBMid75[30] , \wBMid75[29] , \wBMid75[28] , 
        \wBMid75[27] , \wBMid75[26] , \wBMid75[25] , \wBMid75[24] , 
        \wBMid75[23] , \wBMid75[22] , \wBMid75[21] , \wBMid75[20] , 
        \wBMid75[19] , \wBMid75[18] , \wBMid75[17] , \wBMid75[16] , 
        \wBMid75[15] , \wBMid75[14] , \wBMid75[13] , \wBMid75[12] , 
        \wBMid75[11] , \wBMid75[10] , \wBMid75[9] , \wBMid75[8] , \wBMid75[7] , 
        \wBMid75[6] , \wBMid75[5] , \wBMid75[4] , \wBMid75[3] , \wBMid75[2] , 
        \wBMid75[1] , \wBMid75[0] }), .LoOut({\wAMid76[31] , \wAMid76[30] , 
        \wAMid76[29] , \wAMid76[28] , \wAMid76[27] , \wAMid76[26] , 
        \wAMid76[25] , \wAMid76[24] , \wAMid76[23] , \wAMid76[22] , 
        \wAMid76[21] , \wAMid76[20] , \wAMid76[19] , \wAMid76[18] , 
        \wAMid76[17] , \wAMid76[16] , \wAMid76[15] , \wAMid76[14] , 
        \wAMid76[13] , \wAMid76[12] , \wAMid76[11] , \wAMid76[10] , 
        \wAMid76[9] , \wAMid76[8] , \wAMid76[7] , \wAMid76[6] , \wAMid76[5] , 
        \wAMid76[4] , \wAMid76[3] , \wAMid76[2] , \wAMid76[1] , \wAMid76[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn106[31] , \wAIn106[30] , \wAIn106[29] , \wAIn106[28] , 
        \wAIn106[27] , \wAIn106[26] , \wAIn106[25] , \wAIn106[24] , 
        \wAIn106[23] , \wAIn106[22] , \wAIn106[21] , \wAIn106[20] , 
        \wAIn106[19] , \wAIn106[18] , \wAIn106[17] , \wAIn106[16] , 
        \wAIn106[15] , \wAIn106[14] , \wAIn106[13] , \wAIn106[12] , 
        \wAIn106[11] , \wAIn106[10] , \wAIn106[9] , \wAIn106[8] , \wAIn106[7] , 
        \wAIn106[6] , \wAIn106[5] , \wAIn106[4] , \wAIn106[3] , \wAIn106[2] , 
        \wAIn106[1] , \wAIn106[0] }), .BIn({\wBIn106[31] , \wBIn106[30] , 
        \wBIn106[29] , \wBIn106[28] , \wBIn106[27] , \wBIn106[26] , 
        \wBIn106[25] , \wBIn106[24] , \wBIn106[23] , \wBIn106[22] , 
        \wBIn106[21] , \wBIn106[20] , \wBIn106[19] , \wBIn106[18] , 
        \wBIn106[17] , \wBIn106[16] , \wBIn106[15] , \wBIn106[14] , 
        \wBIn106[13] , \wBIn106[12] , \wBIn106[11] , \wBIn106[10] , 
        \wBIn106[9] , \wBIn106[8] , \wBIn106[7] , \wBIn106[6] , \wBIn106[5] , 
        \wBIn106[4] , \wBIn106[3] , \wBIn106[2] , \wBIn106[1] , \wBIn106[0] }), 
        .HiOut({\wBMid105[31] , \wBMid105[30] , \wBMid105[29] , \wBMid105[28] , 
        \wBMid105[27] , \wBMid105[26] , \wBMid105[25] , \wBMid105[24] , 
        \wBMid105[23] , \wBMid105[22] , \wBMid105[21] , \wBMid105[20] , 
        \wBMid105[19] , \wBMid105[18] , \wBMid105[17] , \wBMid105[16] , 
        \wBMid105[15] , \wBMid105[14] , \wBMid105[13] , \wBMid105[12] , 
        \wBMid105[11] , \wBMid105[10] , \wBMid105[9] , \wBMid105[8] , 
        \wBMid105[7] , \wBMid105[6] , \wBMid105[5] , \wBMid105[4] , 
        \wBMid105[3] , \wBMid105[2] , \wBMid105[1] , \wBMid105[0] }), .LoOut({
        \wAMid106[31] , \wAMid106[30] , \wAMid106[29] , \wAMid106[28] , 
        \wAMid106[27] , \wAMid106[26] , \wAMid106[25] , \wAMid106[24] , 
        \wAMid106[23] , \wAMid106[22] , \wAMid106[21] , \wAMid106[20] , 
        \wAMid106[19] , \wAMid106[18] , \wAMid106[17] , \wAMid106[16] , 
        \wAMid106[15] , \wAMid106[14] , \wAMid106[13] , \wAMid106[12] , 
        \wAMid106[11] , \wAMid106[10] , \wAMid106[9] , \wAMid106[8] , 
        \wAMid106[7] , \wAMid106[6] , \wAMid106[5] , \wAMid106[4] , 
        \wAMid106[3] , \wAMid106[2] , \wAMid106[1] , \wAMid106[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid14[31] , \wAMid14[30] , \wAMid14[29] , \wAMid14[28] , 
        \wAMid14[27] , \wAMid14[26] , \wAMid14[25] , \wAMid14[24] , 
        \wAMid14[23] , \wAMid14[22] , \wAMid14[21] , \wAMid14[20] , 
        \wAMid14[19] , \wAMid14[18] , \wAMid14[17] , \wAMid14[16] , 
        \wAMid14[15] , \wAMid14[14] , \wAMid14[13] , \wAMid14[12] , 
        \wAMid14[11] , \wAMid14[10] , \wAMid14[9] , \wAMid14[8] , \wAMid14[7] , 
        \wAMid14[6] , \wAMid14[5] , \wAMid14[4] , \wAMid14[3] , \wAMid14[2] , 
        \wAMid14[1] , \wAMid14[0] }), .BIn({\wBMid14[31] , \wBMid14[30] , 
        \wBMid14[29] , \wBMid14[28] , \wBMid14[27] , \wBMid14[26] , 
        \wBMid14[25] , \wBMid14[24] , \wBMid14[23] , \wBMid14[22] , 
        \wBMid14[21] , \wBMid14[20] , \wBMid14[19] , \wBMid14[18] , 
        \wBMid14[17] , \wBMid14[16] , \wBMid14[15] , \wBMid14[14] , 
        \wBMid14[13] , \wBMid14[12] , \wBMid14[11] , \wBMid14[10] , 
        \wBMid14[9] , \wBMid14[8] , \wBMid14[7] , \wBMid14[6] , \wBMid14[5] , 
        \wBMid14[4] , \wBMid14[3] , \wBMid14[2] , \wBMid14[1] , \wBMid14[0] }), 
        .HiOut({\wRegInB14[31] , \wRegInB14[30] , \wRegInB14[29] , 
        \wRegInB14[28] , \wRegInB14[27] , \wRegInB14[26] , \wRegInB14[25] , 
        \wRegInB14[24] , \wRegInB14[23] , \wRegInB14[22] , \wRegInB14[21] , 
        \wRegInB14[20] , \wRegInB14[19] , \wRegInB14[18] , \wRegInB14[17] , 
        \wRegInB14[16] , \wRegInB14[15] , \wRegInB14[14] , \wRegInB14[13] , 
        \wRegInB14[12] , \wRegInB14[11] , \wRegInB14[10] , \wRegInB14[9] , 
        \wRegInB14[8] , \wRegInB14[7] , \wRegInB14[6] , \wRegInB14[5] , 
        \wRegInB14[4] , \wRegInB14[3] , \wRegInB14[2] , \wRegInB14[1] , 
        \wRegInB14[0] }), .LoOut({\wRegInA15[31] , \wRegInA15[30] , 
        \wRegInA15[29] , \wRegInA15[28] , \wRegInA15[27] , \wRegInA15[26] , 
        \wRegInA15[25] , \wRegInA15[24] , \wRegInA15[23] , \wRegInA15[22] , 
        \wRegInA15[21] , \wRegInA15[20] , \wRegInA15[19] , \wRegInA15[18] , 
        \wRegInA15[17] , \wRegInA15[16] , \wRegInA15[15] , \wRegInA15[14] , 
        \wRegInA15[13] , \wRegInA15[12] , \wRegInA15[11] , \wRegInA15[10] , 
        \wRegInA15[9] , \wRegInA15[8] , \wRegInA15[7] , \wRegInA15[6] , 
        \wRegInA15[5] , \wRegInA15[4] , \wRegInA15[3] , \wRegInA15[2] , 
        \wRegInA15[1] , \wRegInA15[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_121 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink122[31] , \ScanLink122[30] , \ScanLink122[29] , 
        \ScanLink122[28] , \ScanLink122[27] , \ScanLink122[26] , 
        \ScanLink122[25] , \ScanLink122[24] , \ScanLink122[23] , 
        \ScanLink122[22] , \ScanLink122[21] , \ScanLink122[20] , 
        \ScanLink122[19] , \ScanLink122[18] , \ScanLink122[17] , 
        \ScanLink122[16] , \ScanLink122[15] , \ScanLink122[14] , 
        \ScanLink122[13] , \ScanLink122[12] , \ScanLink122[11] , 
        \ScanLink122[10] , \ScanLink122[9] , \ScanLink122[8] , 
        \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , \ScanLink122[4] , 
        \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , \ScanLink122[0] 
        }), .ScanOut({\ScanLink121[31] , \ScanLink121[30] , \ScanLink121[29] , 
        \ScanLink121[28] , \ScanLink121[27] , \ScanLink121[26] , 
        \ScanLink121[25] , \ScanLink121[24] , \ScanLink121[23] , 
        \ScanLink121[22] , \ScanLink121[21] , \ScanLink121[20] , 
        \ScanLink121[19] , \ScanLink121[18] , \ScanLink121[17] , 
        \ScanLink121[16] , \ScanLink121[15] , \ScanLink121[14] , 
        \ScanLink121[13] , \ScanLink121[12] , \ScanLink121[11] , 
        \ScanLink121[10] , \ScanLink121[9] , \ScanLink121[8] , 
        \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , \ScanLink121[4] , 
        \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , \ScanLink121[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA67[31] , \wRegInA67[30] , \wRegInA67[29] , 
        \wRegInA67[28] , \wRegInA67[27] , \wRegInA67[26] , \wRegInA67[25] , 
        \wRegInA67[24] , \wRegInA67[23] , \wRegInA67[22] , \wRegInA67[21] , 
        \wRegInA67[20] , \wRegInA67[19] , \wRegInA67[18] , \wRegInA67[17] , 
        \wRegInA67[16] , \wRegInA67[15] , \wRegInA67[14] , \wRegInA67[13] , 
        \wRegInA67[12] , \wRegInA67[11] , \wRegInA67[10] , \wRegInA67[9] , 
        \wRegInA67[8] , \wRegInA67[7] , \wRegInA67[6] , \wRegInA67[5] , 
        \wRegInA67[4] , \wRegInA67[3] , \wRegInA67[2] , \wRegInA67[1] , 
        \wRegInA67[0] }), .Out({\wAIn67[31] , \wAIn67[30] , \wAIn67[29] , 
        \wAIn67[28] , \wAIn67[27] , \wAIn67[26] , \wAIn67[25] , \wAIn67[24] , 
        \wAIn67[23] , \wAIn67[22] , \wAIn67[21] , \wAIn67[20] , \wAIn67[19] , 
        \wAIn67[18] , \wAIn67[17] , \wAIn67[16] , \wAIn67[15] , \wAIn67[14] , 
        \wAIn67[13] , \wAIn67[12] , \wAIn67[11] , \wAIn67[10] , \wAIn67[9] , 
        \wAIn67[8] , \wAIn67[7] , \wAIn67[6] , \wAIn67[5] , \wAIn67[4] , 
        \wAIn67[3] , \wAIn67[2] , \wAIn67[1] , \wAIn67[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid117[31] , \wAMid117[30] , \wAMid117[29] , \wAMid117[28] , 
        \wAMid117[27] , \wAMid117[26] , \wAMid117[25] , \wAMid117[24] , 
        \wAMid117[23] , \wAMid117[22] , \wAMid117[21] , \wAMid117[20] , 
        \wAMid117[19] , \wAMid117[18] , \wAMid117[17] , \wAMid117[16] , 
        \wAMid117[15] , \wAMid117[14] , \wAMid117[13] , \wAMid117[12] , 
        \wAMid117[11] , \wAMid117[10] , \wAMid117[9] , \wAMid117[8] , 
        \wAMid117[7] , \wAMid117[6] , \wAMid117[5] , \wAMid117[4] , 
        \wAMid117[3] , \wAMid117[2] , \wAMid117[1] , \wAMid117[0] }), .BIn({
        \wBMid117[31] , \wBMid117[30] , \wBMid117[29] , \wBMid117[28] , 
        \wBMid117[27] , \wBMid117[26] , \wBMid117[25] , \wBMid117[24] , 
        \wBMid117[23] , \wBMid117[22] , \wBMid117[21] , \wBMid117[20] , 
        \wBMid117[19] , \wBMid117[18] , \wBMid117[17] , \wBMid117[16] , 
        \wBMid117[15] , \wBMid117[14] , \wBMid117[13] , \wBMid117[12] , 
        \wBMid117[11] , \wBMid117[10] , \wBMid117[9] , \wBMid117[8] , 
        \wBMid117[7] , \wBMid117[6] , \wBMid117[5] , \wBMid117[4] , 
        \wBMid117[3] , \wBMid117[2] , \wBMid117[1] , \wBMid117[0] }), .HiOut({
        \wRegInB117[31] , \wRegInB117[30] , \wRegInB117[29] , \wRegInB117[28] , 
        \wRegInB117[27] , \wRegInB117[26] , \wRegInB117[25] , \wRegInB117[24] , 
        \wRegInB117[23] , \wRegInB117[22] , \wRegInB117[21] , \wRegInB117[20] , 
        \wRegInB117[19] , \wRegInB117[18] , \wRegInB117[17] , \wRegInB117[16] , 
        \wRegInB117[15] , \wRegInB117[14] , \wRegInB117[13] , \wRegInB117[12] , 
        \wRegInB117[11] , \wRegInB117[10] , \wRegInB117[9] , \wRegInB117[8] , 
        \wRegInB117[7] , \wRegInB117[6] , \wRegInB117[5] , \wRegInB117[4] , 
        \wRegInB117[3] , \wRegInB117[2] , \wRegInB117[1] , \wRegInB117[0] }), 
        .LoOut({\wRegInA118[31] , \wRegInA118[30] , \wRegInA118[29] , 
        \wRegInA118[28] , \wRegInA118[27] , \wRegInA118[26] , \wRegInA118[25] , 
        \wRegInA118[24] , \wRegInA118[23] , \wRegInA118[22] , \wRegInA118[21] , 
        \wRegInA118[20] , \wRegInA118[19] , \wRegInA118[18] , \wRegInA118[17] , 
        \wRegInA118[16] , \wRegInA118[15] , \wRegInA118[14] , \wRegInA118[13] , 
        \wRegInA118[12] , \wRegInA118[11] , \wRegInA118[10] , \wRegInA118[9] , 
        \wRegInA118[8] , \wRegInA118[7] , \wRegInA118[6] , \wRegInA118[5] , 
        \wRegInA118[4] , \wRegInA118[3] , \wRegInA118[2] , \wRegInA118[1] , 
        \wRegInA118[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_168 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink169[31] , \ScanLink169[30] , \ScanLink169[29] , 
        \ScanLink169[28] , \ScanLink169[27] , \ScanLink169[26] , 
        \ScanLink169[25] , \ScanLink169[24] , \ScanLink169[23] , 
        \ScanLink169[22] , \ScanLink169[21] , \ScanLink169[20] , 
        \ScanLink169[19] , \ScanLink169[18] , \ScanLink169[17] , 
        \ScanLink169[16] , \ScanLink169[15] , \ScanLink169[14] , 
        \ScanLink169[13] , \ScanLink169[12] , \ScanLink169[11] , 
        \ScanLink169[10] , \ScanLink169[9] , \ScanLink169[8] , 
        \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , \ScanLink169[4] , 
        \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , \ScanLink169[0] 
        }), .ScanOut({\ScanLink168[31] , \ScanLink168[30] , \ScanLink168[29] , 
        \ScanLink168[28] , \ScanLink168[27] , \ScanLink168[26] , 
        \ScanLink168[25] , \ScanLink168[24] , \ScanLink168[23] , 
        \ScanLink168[22] , \ScanLink168[21] , \ScanLink168[20] , 
        \ScanLink168[19] , \ScanLink168[18] , \ScanLink168[17] , 
        \ScanLink168[16] , \ScanLink168[15] , \ScanLink168[14] , 
        \ScanLink168[13] , \ScanLink168[12] , \ScanLink168[11] , 
        \ScanLink168[10] , \ScanLink168[9] , \ScanLink168[8] , 
        \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , \ScanLink168[4] , 
        \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , \ScanLink168[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB43[31] , \wRegInB43[30] , \wRegInB43[29] , 
        \wRegInB43[28] , \wRegInB43[27] , \wRegInB43[26] , \wRegInB43[25] , 
        \wRegInB43[24] , \wRegInB43[23] , \wRegInB43[22] , \wRegInB43[21] , 
        \wRegInB43[20] , \wRegInB43[19] , \wRegInB43[18] , \wRegInB43[17] , 
        \wRegInB43[16] , \wRegInB43[15] , \wRegInB43[14] , \wRegInB43[13] , 
        \wRegInB43[12] , \wRegInB43[11] , \wRegInB43[10] , \wRegInB43[9] , 
        \wRegInB43[8] , \wRegInB43[7] , \wRegInB43[6] , \wRegInB43[5] , 
        \wRegInB43[4] , \wRegInB43[3] , \wRegInB43[2] , \wRegInB43[1] , 
        \wRegInB43[0] }), .Out({\wBIn43[31] , \wBIn43[30] , \wBIn43[29] , 
        \wBIn43[28] , \wBIn43[27] , \wBIn43[26] , \wBIn43[25] , \wBIn43[24] , 
        \wBIn43[23] , \wBIn43[22] , \wBIn43[21] , \wBIn43[20] , \wBIn43[19] , 
        \wBIn43[18] , \wBIn43[17] , \wBIn43[16] , \wBIn43[15] , \wBIn43[14] , 
        \wBIn43[13] , \wBIn43[12] , \wBIn43[11] , \wBIn43[10] , \wBIn43[9] , 
        \wBIn43[8] , \wBIn43[7] , \wBIn43[6] , \wBIn43[5] , \wBIn43[4] , 
        \wBIn43[3] , \wBIn43[2] , \wBIn43[1] , \wBIn43[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_71 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink72[31] , \ScanLink72[30] , \ScanLink72[29] , 
        \ScanLink72[28] , \ScanLink72[27] , \ScanLink72[26] , \ScanLink72[25] , 
        \ScanLink72[24] , \ScanLink72[23] , \ScanLink72[22] , \ScanLink72[21] , 
        \ScanLink72[20] , \ScanLink72[19] , \ScanLink72[18] , \ScanLink72[17] , 
        \ScanLink72[16] , \ScanLink72[15] , \ScanLink72[14] , \ScanLink72[13] , 
        \ScanLink72[12] , \ScanLink72[11] , \ScanLink72[10] , \ScanLink72[9] , 
        \ScanLink72[8] , \ScanLink72[7] , \ScanLink72[6] , \ScanLink72[5] , 
        \ScanLink72[4] , \ScanLink72[3] , \ScanLink72[2] , \ScanLink72[1] , 
        \ScanLink72[0] }), .ScanOut({\ScanLink71[31] , \ScanLink71[30] , 
        \ScanLink71[29] , \ScanLink71[28] , \ScanLink71[27] , \ScanLink71[26] , 
        \ScanLink71[25] , \ScanLink71[24] , \ScanLink71[23] , \ScanLink71[22] , 
        \ScanLink71[21] , \ScanLink71[20] , \ScanLink71[19] , \ScanLink71[18] , 
        \ScanLink71[17] , \ScanLink71[16] , \ScanLink71[15] , \ScanLink71[14] , 
        \ScanLink71[13] , \ScanLink71[12] , \ScanLink71[11] , \ScanLink71[10] , 
        \ScanLink71[9] , \ScanLink71[8] , \ScanLink71[7] , \ScanLink71[6] , 
        \ScanLink71[5] , \ScanLink71[4] , \ScanLink71[3] , \ScanLink71[2] , 
        \ScanLink71[1] , \ScanLink71[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA92[31] , \wRegInA92[30] , 
        \wRegInA92[29] , \wRegInA92[28] , \wRegInA92[27] , \wRegInA92[26] , 
        \wRegInA92[25] , \wRegInA92[24] , \wRegInA92[23] , \wRegInA92[22] , 
        \wRegInA92[21] , \wRegInA92[20] , \wRegInA92[19] , \wRegInA92[18] , 
        \wRegInA92[17] , \wRegInA92[16] , \wRegInA92[15] , \wRegInA92[14] , 
        \wRegInA92[13] , \wRegInA92[12] , \wRegInA92[11] , \wRegInA92[10] , 
        \wRegInA92[9] , \wRegInA92[8] , \wRegInA92[7] , \wRegInA92[6] , 
        \wRegInA92[5] , \wRegInA92[4] , \wRegInA92[3] , \wRegInA92[2] , 
        \wRegInA92[1] , \wRegInA92[0] }), .Out({\wAIn92[31] , \wAIn92[30] , 
        \wAIn92[29] , \wAIn92[28] , \wAIn92[27] , \wAIn92[26] , \wAIn92[25] , 
        \wAIn92[24] , \wAIn92[23] , \wAIn92[22] , \wAIn92[21] , \wAIn92[20] , 
        \wAIn92[19] , \wAIn92[18] , \wAIn92[17] , \wAIn92[16] , \wAIn92[15] , 
        \wAIn92[14] , \wAIn92[13] , \wAIn92[12] , \wAIn92[11] , \wAIn92[10] , 
        \wAIn92[9] , \wAIn92[8] , \wAIn92[7] , \wAIn92[6] , \wAIn92[5] , 
        \wAIn92[4] , \wAIn92[3] , \wAIn92[2] , \wAIn92[1] , \wAIn92[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_38 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink39[31] , \ScanLink39[30] , \ScanLink39[29] , 
        \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , \ScanLink39[25] , 
        \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , \ScanLink39[21] , 
        \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , \ScanLink39[17] , 
        \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , \ScanLink39[13] , 
        \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , \ScanLink39[9] , 
        \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , \ScanLink39[5] , 
        \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , \ScanLink39[1] , 
        \ScanLink39[0] }), .ScanOut({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB108[31] , \wRegInB108[30] , 
        \wRegInB108[29] , \wRegInB108[28] , \wRegInB108[27] , \wRegInB108[26] , 
        \wRegInB108[25] , \wRegInB108[24] , \wRegInB108[23] , \wRegInB108[22] , 
        \wRegInB108[21] , \wRegInB108[20] , \wRegInB108[19] , \wRegInB108[18] , 
        \wRegInB108[17] , \wRegInB108[16] , \wRegInB108[15] , \wRegInB108[14] , 
        \wRegInB108[13] , \wRegInB108[12] , \wRegInB108[11] , \wRegInB108[10] , 
        \wRegInB108[9] , \wRegInB108[8] , \wRegInB108[7] , \wRegInB108[6] , 
        \wRegInB108[5] , \wRegInB108[4] , \wRegInB108[3] , \wRegInB108[2] , 
        \wRegInB108[1] , \wRegInB108[0] }), .Out({\wBIn108[31] , \wBIn108[30] , 
        \wBIn108[29] , \wBIn108[28] , \wBIn108[27] , \wBIn108[26] , 
        \wBIn108[25] , \wBIn108[24] , \wBIn108[23] , \wBIn108[22] , 
        \wBIn108[21] , \wBIn108[20] , \wBIn108[19] , \wBIn108[18] , 
        \wBIn108[17] , \wBIn108[16] , \wBIn108[15] , \wBIn108[14] , 
        \wBIn108[13] , \wBIn108[12] , \wBIn108[11] , \wBIn108[10] , 
        \wBIn108[9] , \wBIn108[8] , \wBIn108[7] , \wBIn108[6] , \wBIn108[5] , 
        \wBIn108[4] , \wBIn108[3] , \wBIn108[2] , \wBIn108[1] , \wBIn108[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_94 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink95[31] , \ScanLink95[30] , \ScanLink95[29] , 
        \ScanLink95[28] , \ScanLink95[27] , \ScanLink95[26] , \ScanLink95[25] , 
        \ScanLink95[24] , \ScanLink95[23] , \ScanLink95[22] , \ScanLink95[21] , 
        \ScanLink95[20] , \ScanLink95[19] , \ScanLink95[18] , \ScanLink95[17] , 
        \ScanLink95[16] , \ScanLink95[15] , \ScanLink95[14] , \ScanLink95[13] , 
        \ScanLink95[12] , \ScanLink95[11] , \ScanLink95[10] , \ScanLink95[9] , 
        \ScanLink95[8] , \ScanLink95[7] , \ScanLink95[6] , \ScanLink95[5] , 
        \ScanLink95[4] , \ScanLink95[3] , \ScanLink95[2] , \ScanLink95[1] , 
        \ScanLink95[0] }), .ScanOut({\ScanLink94[31] , \ScanLink94[30] , 
        \ScanLink94[29] , \ScanLink94[28] , \ScanLink94[27] , \ScanLink94[26] , 
        \ScanLink94[25] , \ScanLink94[24] , \ScanLink94[23] , \ScanLink94[22] , 
        \ScanLink94[21] , \ScanLink94[20] , \ScanLink94[19] , \ScanLink94[18] , 
        \ScanLink94[17] , \ScanLink94[16] , \ScanLink94[15] , \ScanLink94[14] , 
        \ScanLink94[13] , \ScanLink94[12] , \ScanLink94[11] , \ScanLink94[10] , 
        \ScanLink94[9] , \ScanLink94[8] , \ScanLink94[7] , \ScanLink94[6] , 
        \ScanLink94[5] , \ScanLink94[4] , \ScanLink94[3] , \ScanLink94[2] , 
        \ScanLink94[1] , \ScanLink94[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB80[31] , \wRegInB80[30] , 
        \wRegInB80[29] , \wRegInB80[28] , \wRegInB80[27] , \wRegInB80[26] , 
        \wRegInB80[25] , \wRegInB80[24] , \wRegInB80[23] , \wRegInB80[22] , 
        \wRegInB80[21] , \wRegInB80[20] , \wRegInB80[19] , \wRegInB80[18] , 
        \wRegInB80[17] , \wRegInB80[16] , \wRegInB80[15] , \wRegInB80[14] , 
        \wRegInB80[13] , \wRegInB80[12] , \wRegInB80[11] , \wRegInB80[10] , 
        \wRegInB80[9] , \wRegInB80[8] , \wRegInB80[7] , \wRegInB80[6] , 
        \wRegInB80[5] , \wRegInB80[4] , \wRegInB80[3] , \wRegInB80[2] , 
        \wRegInB80[1] , \wRegInB80[0] }), .Out({\wBIn80[31] , \wBIn80[30] , 
        \wBIn80[29] , \wBIn80[28] , \wBIn80[27] , \wBIn80[26] , \wBIn80[25] , 
        \wBIn80[24] , \wBIn80[23] , \wBIn80[22] , \wBIn80[21] , \wBIn80[20] , 
        \wBIn80[19] , \wBIn80[18] , \wBIn80[17] , \wBIn80[16] , \wBIn80[15] , 
        \wBIn80[14] , \wBIn80[13] , \wBIn80[12] , \wBIn80[11] , \wBIn80[10] , 
        \wBIn80[9] , \wBIn80[8] , \wBIn80[7] , \wBIn80[6] , \wBIn80[5] , 
        \wBIn80[4] , \wBIn80[3] , \wBIn80[2] , \wBIn80[1] , \wBIn80[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_243 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink244[31] , \ScanLink244[30] , \ScanLink244[29] , 
        \ScanLink244[28] , \ScanLink244[27] , \ScanLink244[26] , 
        \ScanLink244[25] , \ScanLink244[24] , \ScanLink244[23] , 
        \ScanLink244[22] , \ScanLink244[21] , \ScanLink244[20] , 
        \ScanLink244[19] , \ScanLink244[18] , \ScanLink244[17] , 
        \ScanLink244[16] , \ScanLink244[15] , \ScanLink244[14] , 
        \ScanLink244[13] , \ScanLink244[12] , \ScanLink244[11] , 
        \ScanLink244[10] , \ScanLink244[9] , \ScanLink244[8] , 
        \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , \ScanLink244[4] , 
        \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , \ScanLink244[0] 
        }), .ScanOut({\ScanLink243[31] , \ScanLink243[30] , \ScanLink243[29] , 
        \ScanLink243[28] , \ScanLink243[27] , \ScanLink243[26] , 
        \ScanLink243[25] , \ScanLink243[24] , \ScanLink243[23] , 
        \ScanLink243[22] , \ScanLink243[21] , \ScanLink243[20] , 
        \ScanLink243[19] , \ScanLink243[18] , \ScanLink243[17] , 
        \ScanLink243[16] , \ScanLink243[15] , \ScanLink243[14] , 
        \ScanLink243[13] , \ScanLink243[12] , \ScanLink243[11] , 
        \ScanLink243[10] , \ScanLink243[9] , \ScanLink243[8] , 
        \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , \ScanLink243[4] , 
        \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , \ScanLink243[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA6[31] , \wRegInA6[30] , \wRegInA6[29] , \wRegInA6[28] , 
        \wRegInA6[27] , \wRegInA6[26] , \wRegInA6[25] , \wRegInA6[24] , 
        \wRegInA6[23] , \wRegInA6[22] , \wRegInA6[21] , \wRegInA6[20] , 
        \wRegInA6[19] , \wRegInA6[18] , \wRegInA6[17] , \wRegInA6[16] , 
        \wRegInA6[15] , \wRegInA6[14] , \wRegInA6[13] , \wRegInA6[12] , 
        \wRegInA6[11] , \wRegInA6[10] , \wRegInA6[9] , \wRegInA6[8] , 
        \wRegInA6[7] , \wRegInA6[6] , \wRegInA6[5] , \wRegInA6[4] , 
        \wRegInA6[3] , \wRegInA6[2] , \wRegInA6[1] , \wRegInA6[0] }), .Out({
        \wAIn6[31] , \wAIn6[30] , \wAIn6[29] , \wAIn6[28] , \wAIn6[27] , 
        \wAIn6[26] , \wAIn6[25] , \wAIn6[24] , \wAIn6[23] , \wAIn6[22] , 
        \wAIn6[21] , \wAIn6[20] , \wAIn6[19] , \wAIn6[18] , \wAIn6[17] , 
        \wAIn6[16] , \wAIn6[15] , \wAIn6[14] , \wAIn6[13] , \wAIn6[12] , 
        \wAIn6[11] , \wAIn6[10] , \wAIn6[9] , \wAIn6[8] , \wAIn6[7] , 
        \wAIn6[6] , \wAIn6[5] , \wAIn6[4] , \wAIn6[3] , \wAIn6[2] , \wAIn6[1] , 
        \wAIn6[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid46[31] , \wAMid46[30] , \wAMid46[29] , \wAMid46[28] , 
        \wAMid46[27] , \wAMid46[26] , \wAMid46[25] , \wAMid46[24] , 
        \wAMid46[23] , \wAMid46[22] , \wAMid46[21] , \wAMid46[20] , 
        \wAMid46[19] , \wAMid46[18] , \wAMid46[17] , \wAMid46[16] , 
        \wAMid46[15] , \wAMid46[14] , \wAMid46[13] , \wAMid46[12] , 
        \wAMid46[11] , \wAMid46[10] , \wAMid46[9] , \wAMid46[8] , \wAMid46[7] , 
        \wAMid46[6] , \wAMid46[5] , \wAMid46[4] , \wAMid46[3] , \wAMid46[2] , 
        \wAMid46[1] , \wAMid46[0] }), .BIn({\wBMid46[31] , \wBMid46[30] , 
        \wBMid46[29] , \wBMid46[28] , \wBMid46[27] , \wBMid46[26] , 
        \wBMid46[25] , \wBMid46[24] , \wBMid46[23] , \wBMid46[22] , 
        \wBMid46[21] , \wBMid46[20] , \wBMid46[19] , \wBMid46[18] , 
        \wBMid46[17] , \wBMid46[16] , \wBMid46[15] , \wBMid46[14] , 
        \wBMid46[13] , \wBMid46[12] , \wBMid46[11] , \wBMid46[10] , 
        \wBMid46[9] , \wBMid46[8] , \wBMid46[7] , \wBMid46[6] , \wBMid46[5] , 
        \wBMid46[4] , \wBMid46[3] , \wBMid46[2] , \wBMid46[1] , \wBMid46[0] }), 
        .HiOut({\wRegInB46[31] , \wRegInB46[30] , \wRegInB46[29] , 
        \wRegInB46[28] , \wRegInB46[27] , \wRegInB46[26] , \wRegInB46[25] , 
        \wRegInB46[24] , \wRegInB46[23] , \wRegInB46[22] , \wRegInB46[21] , 
        \wRegInB46[20] , \wRegInB46[19] , \wRegInB46[18] , \wRegInB46[17] , 
        \wRegInB46[16] , \wRegInB46[15] , \wRegInB46[14] , \wRegInB46[13] , 
        \wRegInB46[12] , \wRegInB46[11] , \wRegInB46[10] , \wRegInB46[9] , 
        \wRegInB46[8] , \wRegInB46[7] , \wRegInB46[6] , \wRegInB46[5] , 
        \wRegInB46[4] , \wRegInB46[3] , \wRegInB46[2] , \wRegInB46[1] , 
        \wRegInB46[0] }), .LoOut({\wRegInA47[31] , \wRegInA47[30] , 
        \wRegInA47[29] , \wRegInA47[28] , \wRegInA47[27] , \wRegInA47[26] , 
        \wRegInA47[25] , \wRegInA47[24] , \wRegInA47[23] , \wRegInA47[22] , 
        \wRegInA47[21] , \wRegInA47[20] , \wRegInA47[19] , \wRegInA47[18] , 
        \wRegInA47[17] , \wRegInA47[16] , \wRegInA47[15] , \wRegInA47[14] , 
        \wRegInA47[13] , \wRegInA47[12] , \wRegInA47[11] , \wRegInA47[10] , 
        \wRegInA47[9] , \wRegInA47[8] , \wRegInA47[7] , \wRegInA47[6] , 
        \wRegInA47[5] , \wRegInA47[4] , \wRegInA47[3] , \wRegInA47[2] , 
        \wRegInA47[1] , \wRegInA47[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_173 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink174[31] , \ScanLink174[30] , \ScanLink174[29] , 
        \ScanLink174[28] , \ScanLink174[27] , \ScanLink174[26] , 
        \ScanLink174[25] , \ScanLink174[24] , \ScanLink174[23] , 
        \ScanLink174[22] , \ScanLink174[21] , \ScanLink174[20] , 
        \ScanLink174[19] , \ScanLink174[18] , \ScanLink174[17] , 
        \ScanLink174[16] , \ScanLink174[15] , \ScanLink174[14] , 
        \ScanLink174[13] , \ScanLink174[12] , \ScanLink174[11] , 
        \ScanLink174[10] , \ScanLink174[9] , \ScanLink174[8] , 
        \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , \ScanLink174[4] , 
        \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , \ScanLink174[0] 
        }), .ScanOut({\ScanLink173[31] , \ScanLink173[30] , \ScanLink173[29] , 
        \ScanLink173[28] , \ScanLink173[27] , \ScanLink173[26] , 
        \ScanLink173[25] , \ScanLink173[24] , \ScanLink173[23] , 
        \ScanLink173[22] , \ScanLink173[21] , \ScanLink173[20] , 
        \ScanLink173[19] , \ScanLink173[18] , \ScanLink173[17] , 
        \ScanLink173[16] , \ScanLink173[15] , \ScanLink173[14] , 
        \ScanLink173[13] , \ScanLink173[12] , \ScanLink173[11] , 
        \ScanLink173[10] , \ScanLink173[9] , \ScanLink173[8] , 
        \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , \ScanLink173[4] , 
        \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , \ScanLink173[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA41[31] , \wRegInA41[30] , \wRegInA41[29] , 
        \wRegInA41[28] , \wRegInA41[27] , \wRegInA41[26] , \wRegInA41[25] , 
        \wRegInA41[24] , \wRegInA41[23] , \wRegInA41[22] , \wRegInA41[21] , 
        \wRegInA41[20] , \wRegInA41[19] , \wRegInA41[18] , \wRegInA41[17] , 
        \wRegInA41[16] , \wRegInA41[15] , \wRegInA41[14] , \wRegInA41[13] , 
        \wRegInA41[12] , \wRegInA41[11] , \wRegInA41[10] , \wRegInA41[9] , 
        \wRegInA41[8] , \wRegInA41[7] , \wRegInA41[6] , \wRegInA41[5] , 
        \wRegInA41[4] , \wRegInA41[3] , \wRegInA41[2] , \wRegInA41[1] , 
        \wRegInA41[0] }), .Out({\wAIn41[31] , \wAIn41[30] , \wAIn41[29] , 
        \wAIn41[28] , \wAIn41[27] , \wAIn41[26] , \wAIn41[25] , \wAIn41[24] , 
        \wAIn41[23] , \wAIn41[22] , \wAIn41[21] , \wAIn41[20] , \wAIn41[19] , 
        \wAIn41[18] , \wAIn41[17] , \wAIn41[16] , \wAIn41[15] , \wAIn41[14] , 
        \wAIn41[13] , \wAIn41[12] , \wAIn41[11] , \wAIn41[10] , \wAIn41[9] , 
        \wAIn41[8] , \wAIn41[7] , \wAIn41[6] , \wAIn41[5] , \wAIn41[4] , 
        \wAIn41[3] , \wAIn41[2] , \wAIn41[1] , \wAIn41[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_23 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink24[31] , \ScanLink24[30] , \ScanLink24[29] , 
        \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , \ScanLink24[25] , 
        \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , \ScanLink24[21] , 
        \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , \ScanLink24[17] , 
        \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , \ScanLink24[13] , 
        \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , \ScanLink24[9] , 
        \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , \ScanLink24[5] , 
        \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , \ScanLink24[1] , 
        \ScanLink24[0] }), .ScanOut({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA116[31] , \wRegInA116[30] , 
        \wRegInA116[29] , \wRegInA116[28] , \wRegInA116[27] , \wRegInA116[26] , 
        \wRegInA116[25] , \wRegInA116[24] , \wRegInA116[23] , \wRegInA116[22] , 
        \wRegInA116[21] , \wRegInA116[20] , \wRegInA116[19] , \wRegInA116[18] , 
        \wRegInA116[17] , \wRegInA116[16] , \wRegInA116[15] , \wRegInA116[14] , 
        \wRegInA116[13] , \wRegInA116[12] , \wRegInA116[11] , \wRegInA116[10] , 
        \wRegInA116[9] , \wRegInA116[8] , \wRegInA116[7] , \wRegInA116[6] , 
        \wRegInA116[5] , \wRegInA116[4] , \wRegInA116[3] , \wRegInA116[2] , 
        \wRegInA116[1] , \wRegInA116[0] }), .Out({\wAIn116[31] , \wAIn116[30] , 
        \wAIn116[29] , \wAIn116[28] , \wAIn116[27] , \wAIn116[26] , 
        \wAIn116[25] , \wAIn116[24] , \wAIn116[23] , \wAIn116[22] , 
        \wAIn116[21] , \wAIn116[20] , \wAIn116[19] , \wAIn116[18] , 
        \wAIn116[17] , \wAIn116[16] , \wAIn116[15] , \wAIn116[14] , 
        \wAIn116[13] , \wAIn116[12] , \wAIn116[11] , \wAIn116[10] , 
        \wAIn116[9] , \wAIn116[8] , \wAIn116[7] , \wAIn116[6] , \wAIn116[5] , 
        \wAIn116[4] , \wAIn116[3] , \wAIn116[2] , \wAIn116[1] , \wAIn116[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid61[31] , \wAMid61[30] , \wAMid61[29] , \wAMid61[28] , 
        \wAMid61[27] , \wAMid61[26] , \wAMid61[25] , \wAMid61[24] , 
        \wAMid61[23] , \wAMid61[22] , \wAMid61[21] , \wAMid61[20] , 
        \wAMid61[19] , \wAMid61[18] , \wAMid61[17] , \wAMid61[16] , 
        \wAMid61[15] , \wAMid61[14] , \wAMid61[13] , \wAMid61[12] , 
        \wAMid61[11] , \wAMid61[10] , \wAMid61[9] , \wAMid61[8] , \wAMid61[7] , 
        \wAMid61[6] , \wAMid61[5] , \wAMid61[4] , \wAMid61[3] , \wAMid61[2] , 
        \wAMid61[1] , \wAMid61[0] }), .BIn({\wBMid61[31] , \wBMid61[30] , 
        \wBMid61[29] , \wBMid61[28] , \wBMid61[27] , \wBMid61[26] , 
        \wBMid61[25] , \wBMid61[24] , \wBMid61[23] , \wBMid61[22] , 
        \wBMid61[21] , \wBMid61[20] , \wBMid61[19] , \wBMid61[18] , 
        \wBMid61[17] , \wBMid61[16] , \wBMid61[15] , \wBMid61[14] , 
        \wBMid61[13] , \wBMid61[12] , \wBMid61[11] , \wBMid61[10] , 
        \wBMid61[9] , \wBMid61[8] , \wBMid61[7] , \wBMid61[6] , \wBMid61[5] , 
        \wBMid61[4] , \wBMid61[3] , \wBMid61[2] , \wBMid61[1] , \wBMid61[0] }), 
        .HiOut({\wRegInB61[31] , \wRegInB61[30] , \wRegInB61[29] , 
        \wRegInB61[28] , \wRegInB61[27] , \wRegInB61[26] , \wRegInB61[25] , 
        \wRegInB61[24] , \wRegInB61[23] , \wRegInB61[22] , \wRegInB61[21] , 
        \wRegInB61[20] , \wRegInB61[19] , \wRegInB61[18] , \wRegInB61[17] , 
        \wRegInB61[16] , \wRegInB61[15] , \wRegInB61[14] , \wRegInB61[13] , 
        \wRegInB61[12] , \wRegInB61[11] , \wRegInB61[10] , \wRegInB61[9] , 
        \wRegInB61[8] , \wRegInB61[7] , \wRegInB61[6] , \wRegInB61[5] , 
        \wRegInB61[4] , \wRegInB61[3] , \wRegInB61[2] , \wRegInB61[1] , 
        \wRegInB61[0] }), .LoOut({\wRegInA62[31] , \wRegInA62[30] , 
        \wRegInA62[29] , \wRegInA62[28] , \wRegInA62[27] , \wRegInA62[26] , 
        \wRegInA62[25] , \wRegInA62[24] , \wRegInA62[23] , \wRegInA62[22] , 
        \wRegInA62[21] , \wRegInA62[20] , \wRegInA62[19] , \wRegInA62[18] , 
        \wRegInA62[17] , \wRegInA62[16] , \wRegInA62[15] , \wRegInA62[14] , 
        \wRegInA62[13] , \wRegInA62[12] , \wRegInA62[11] , \wRegInA62[10] , 
        \wRegInA62[9] , \wRegInA62[8] , \wRegInA62[7] , \wRegInA62[6] , 
        \wRegInA62[5] , \wRegInA62[4] , \wRegInA62[3] , \wRegInA62[2] , 
        \wRegInA62[1] , \wRegInA62[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_154 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink155[31] , \ScanLink155[30] , \ScanLink155[29] , 
        \ScanLink155[28] , \ScanLink155[27] , \ScanLink155[26] , 
        \ScanLink155[25] , \ScanLink155[24] , \ScanLink155[23] , 
        \ScanLink155[22] , \ScanLink155[21] , \ScanLink155[20] , 
        \ScanLink155[19] , \ScanLink155[18] , \ScanLink155[17] , 
        \ScanLink155[16] , \ScanLink155[15] , \ScanLink155[14] , 
        \ScanLink155[13] , \ScanLink155[12] , \ScanLink155[11] , 
        \ScanLink155[10] , \ScanLink155[9] , \ScanLink155[8] , 
        \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , \ScanLink155[4] , 
        \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , \ScanLink155[0] 
        }), .ScanOut({\ScanLink154[31] , \ScanLink154[30] , \ScanLink154[29] , 
        \ScanLink154[28] , \ScanLink154[27] , \ScanLink154[26] , 
        \ScanLink154[25] , \ScanLink154[24] , \ScanLink154[23] , 
        \ScanLink154[22] , \ScanLink154[21] , \ScanLink154[20] , 
        \ScanLink154[19] , \ScanLink154[18] , \ScanLink154[17] , 
        \ScanLink154[16] , \ScanLink154[15] , \ScanLink154[14] , 
        \ScanLink154[13] , \ScanLink154[12] , \ScanLink154[11] , 
        \ScanLink154[10] , \ScanLink154[9] , \ScanLink154[8] , 
        \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , \ScanLink154[4] , 
        \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , \ScanLink154[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB50[31] , \wRegInB50[30] , \wRegInB50[29] , 
        \wRegInB50[28] , \wRegInB50[27] , \wRegInB50[26] , \wRegInB50[25] , 
        \wRegInB50[24] , \wRegInB50[23] , \wRegInB50[22] , \wRegInB50[21] , 
        \wRegInB50[20] , \wRegInB50[19] , \wRegInB50[18] , \wRegInB50[17] , 
        \wRegInB50[16] , \wRegInB50[15] , \wRegInB50[14] , \wRegInB50[13] , 
        \wRegInB50[12] , \wRegInB50[11] , \wRegInB50[10] , \wRegInB50[9] , 
        \wRegInB50[8] , \wRegInB50[7] , \wRegInB50[6] , \wRegInB50[5] , 
        \wRegInB50[4] , \wRegInB50[3] , \wRegInB50[2] , \wRegInB50[1] , 
        \wRegInB50[0] }), .Out({\wBIn50[31] , \wBIn50[30] , \wBIn50[29] , 
        \wBIn50[28] , \wBIn50[27] , \wBIn50[26] , \wBIn50[25] , \wBIn50[24] , 
        \wBIn50[23] , \wBIn50[22] , \wBIn50[21] , \wBIn50[20] , \wBIn50[19] , 
        \wBIn50[18] , \wBIn50[17] , \wBIn50[16] , \wBIn50[15] , \wBIn50[14] , 
        \wBIn50[13] , \wBIn50[12] , \wBIn50[11] , \wBIn50[10] , \wBIn50[9] , 
        \wBIn50[8] , \wBIn50[7] , \wBIn50[6] , \wBIn50[5] , \wBIn50[4] , 
        \wBIn50[3] , \wBIn50[2] , \wBIn50[1] , \wBIn50[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn121[31] , \wAIn121[30] , \wAIn121[29] , \wAIn121[28] , 
        \wAIn121[27] , \wAIn121[26] , \wAIn121[25] , \wAIn121[24] , 
        \wAIn121[23] , \wAIn121[22] , \wAIn121[21] , \wAIn121[20] , 
        \wAIn121[19] , \wAIn121[18] , \wAIn121[17] , \wAIn121[16] , 
        \wAIn121[15] , \wAIn121[14] , \wAIn121[13] , \wAIn121[12] , 
        \wAIn121[11] , \wAIn121[10] , \wAIn121[9] , \wAIn121[8] , \wAIn121[7] , 
        \wAIn121[6] , \wAIn121[5] , \wAIn121[4] , \wAIn121[3] , \wAIn121[2] , 
        \wAIn121[1] , \wAIn121[0] }), .BIn({\wBIn121[31] , \wBIn121[30] , 
        \wBIn121[29] , \wBIn121[28] , \wBIn121[27] , \wBIn121[26] , 
        \wBIn121[25] , \wBIn121[24] , \wBIn121[23] , \wBIn121[22] , 
        \wBIn121[21] , \wBIn121[20] , \wBIn121[19] , \wBIn121[18] , 
        \wBIn121[17] , \wBIn121[16] , \wBIn121[15] , \wBIn121[14] , 
        \wBIn121[13] , \wBIn121[12] , \wBIn121[11] , \wBIn121[10] , 
        \wBIn121[9] , \wBIn121[8] , \wBIn121[7] , \wBIn121[6] , \wBIn121[5] , 
        \wBIn121[4] , \wBIn121[3] , \wBIn121[2] , \wBIn121[1] , \wBIn121[0] }), 
        .HiOut({\wBMid120[31] , \wBMid120[30] , \wBMid120[29] , \wBMid120[28] , 
        \wBMid120[27] , \wBMid120[26] , \wBMid120[25] , \wBMid120[24] , 
        \wBMid120[23] , \wBMid120[22] , \wBMid120[21] , \wBMid120[20] , 
        \wBMid120[19] , \wBMid120[18] , \wBMid120[17] , \wBMid120[16] , 
        \wBMid120[15] , \wBMid120[14] , \wBMid120[13] , \wBMid120[12] , 
        \wBMid120[11] , \wBMid120[10] , \wBMid120[9] , \wBMid120[8] , 
        \wBMid120[7] , \wBMid120[6] , \wBMid120[5] , \wBMid120[4] , 
        \wBMid120[3] , \wBMid120[2] , \wBMid120[1] , \wBMid120[0] }), .LoOut({
        \wAMid121[31] , \wAMid121[30] , \wAMid121[29] , \wAMid121[28] , 
        \wAMid121[27] , \wAMid121[26] , \wAMid121[25] , \wAMid121[24] , 
        \wAMid121[23] , \wAMid121[22] , \wAMid121[21] , \wAMid121[20] , 
        \wAMid121[19] , \wAMid121[18] , \wAMid121[17] , \wAMid121[16] , 
        \wAMid121[15] , \wAMid121[14] , \wAMid121[13] , \wAMid121[12] , 
        \wAMid121[11] , \wAMid121[10] , \wAMid121[9] , \wAMid121[8] , 
        \wAMid121[7] , \wAMid121[6] , \wAMid121[5] , \wAMid121[4] , 
        \wAMid121[3] , \wAMid121[2] , \wAMid121[1] , \wAMid121[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid28[31] , \wAMid28[30] , \wAMid28[29] , \wAMid28[28] , 
        \wAMid28[27] , \wAMid28[26] , \wAMid28[25] , \wAMid28[24] , 
        \wAMid28[23] , \wAMid28[22] , \wAMid28[21] , \wAMid28[20] , 
        \wAMid28[19] , \wAMid28[18] , \wAMid28[17] , \wAMid28[16] , 
        \wAMid28[15] , \wAMid28[14] , \wAMid28[13] , \wAMid28[12] , 
        \wAMid28[11] , \wAMid28[10] , \wAMid28[9] , \wAMid28[8] , \wAMid28[7] , 
        \wAMid28[6] , \wAMid28[5] , \wAMid28[4] , \wAMid28[3] , \wAMid28[2] , 
        \wAMid28[1] , \wAMid28[0] }), .BIn({\wBMid28[31] , \wBMid28[30] , 
        \wBMid28[29] , \wBMid28[28] , \wBMid28[27] , \wBMid28[26] , 
        \wBMid28[25] , \wBMid28[24] , \wBMid28[23] , \wBMid28[22] , 
        \wBMid28[21] , \wBMid28[20] , \wBMid28[19] , \wBMid28[18] , 
        \wBMid28[17] , \wBMid28[16] , \wBMid28[15] , \wBMid28[14] , 
        \wBMid28[13] , \wBMid28[12] , \wBMid28[11] , \wBMid28[10] , 
        \wBMid28[9] , \wBMid28[8] , \wBMid28[7] , \wBMid28[6] , \wBMid28[5] , 
        \wBMid28[4] , \wBMid28[3] , \wBMid28[2] , \wBMid28[1] , \wBMid28[0] }), 
        .HiOut({\wRegInB28[31] , \wRegInB28[30] , \wRegInB28[29] , 
        \wRegInB28[28] , \wRegInB28[27] , \wRegInB28[26] , \wRegInB28[25] , 
        \wRegInB28[24] , \wRegInB28[23] , \wRegInB28[22] , \wRegInB28[21] , 
        \wRegInB28[20] , \wRegInB28[19] , \wRegInB28[18] , \wRegInB28[17] , 
        \wRegInB28[16] , \wRegInB28[15] , \wRegInB28[14] , \wRegInB28[13] , 
        \wRegInB28[12] , \wRegInB28[11] , \wRegInB28[10] , \wRegInB28[9] , 
        \wRegInB28[8] , \wRegInB28[7] , \wRegInB28[6] , \wRegInB28[5] , 
        \wRegInB28[4] , \wRegInB28[3] , \wRegInB28[2] , \wRegInB28[1] , 
        \wRegInB28[0] }), .LoOut({\wRegInA29[31] , \wRegInA29[30] , 
        \wRegInA29[29] , \wRegInA29[28] , \wRegInA29[27] , \wRegInA29[26] , 
        \wRegInA29[25] , \wRegInA29[24] , \wRegInA29[23] , \wRegInA29[22] , 
        \wRegInA29[21] , \wRegInA29[20] , \wRegInA29[19] , \wRegInA29[18] , 
        \wRegInA29[17] , \wRegInA29[16] , \wRegInA29[15] , \wRegInA29[14] , 
        \wRegInA29[13] , \wRegInA29[12] , \wRegInA29[11] , \wRegInA29[10] , 
        \wRegInA29[9] , \wRegInA29[8] , \wRegInA29[7] , \wRegInA29[6] , 
        \wRegInA29[5] , \wRegInA29[4] , \wRegInA29[3] , \wRegInA29[2] , 
        \wRegInA29[1] , \wRegInA29[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn38[31] , \wAIn38[30] , \wAIn38[29] , \wAIn38[28] , \wAIn38[27] , 
        \wAIn38[26] , \wAIn38[25] , \wAIn38[24] , \wAIn38[23] , \wAIn38[22] , 
        \wAIn38[21] , \wAIn38[20] , \wAIn38[19] , \wAIn38[18] , \wAIn38[17] , 
        \wAIn38[16] , \wAIn38[15] , \wAIn38[14] , \wAIn38[13] , \wAIn38[12] , 
        \wAIn38[11] , \wAIn38[10] , \wAIn38[9] , \wAIn38[8] , \wAIn38[7] , 
        \wAIn38[6] , \wAIn38[5] , \wAIn38[4] , \wAIn38[3] , \wAIn38[2] , 
        \wAIn38[1] , \wAIn38[0] }), .BIn({\wBIn38[31] , \wBIn38[30] , 
        \wBIn38[29] , \wBIn38[28] , \wBIn38[27] , \wBIn38[26] , \wBIn38[25] , 
        \wBIn38[24] , \wBIn38[23] , \wBIn38[22] , \wBIn38[21] , \wBIn38[20] , 
        \wBIn38[19] , \wBIn38[18] , \wBIn38[17] , \wBIn38[16] , \wBIn38[15] , 
        \wBIn38[14] , \wBIn38[13] , \wBIn38[12] , \wBIn38[11] , \wBIn38[10] , 
        \wBIn38[9] , \wBIn38[8] , \wBIn38[7] , \wBIn38[6] , \wBIn38[5] , 
        \wBIn38[4] , \wBIn38[3] , \wBIn38[2] , \wBIn38[1] , \wBIn38[0] }), 
        .HiOut({\wBMid37[31] , \wBMid37[30] , \wBMid37[29] , \wBMid37[28] , 
        \wBMid37[27] , \wBMid37[26] , \wBMid37[25] , \wBMid37[24] , 
        \wBMid37[23] , \wBMid37[22] , \wBMid37[21] , \wBMid37[20] , 
        \wBMid37[19] , \wBMid37[18] , \wBMid37[17] , \wBMid37[16] , 
        \wBMid37[15] , \wBMid37[14] , \wBMid37[13] , \wBMid37[12] , 
        \wBMid37[11] , \wBMid37[10] , \wBMid37[9] , \wBMid37[8] , \wBMid37[7] , 
        \wBMid37[6] , \wBMid37[5] , \wBMid37[4] , \wBMid37[3] , \wBMid37[2] , 
        \wBMid37[1] , \wBMid37[0] }), .LoOut({\wAMid38[31] , \wAMid38[30] , 
        \wAMid38[29] , \wAMid38[28] , \wAMid38[27] , \wAMid38[26] , 
        \wAMid38[25] , \wAMid38[24] , \wAMid38[23] , \wAMid38[22] , 
        \wAMid38[21] , \wAMid38[20] , \wAMid38[19] , \wAMid38[18] , 
        \wAMid38[17] , \wAMid38[16] , \wAMid38[15] , \wAMid38[14] , 
        \wAMid38[13] , \wAMid38[12] , \wAMid38[11] , \wAMid38[10] , 
        \wAMid38[9] , \wAMid38[8] , \wAMid38[7] , \wAMid38[6] , \wAMid38[5] , 
        \wAMid38[4] , \wAMid38[3] , \wAMid38[2] , \wAMid38[1] , \wAMid38[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn93[31] , \wAIn93[30] , \wAIn93[29] , \wAIn93[28] , \wAIn93[27] , 
        \wAIn93[26] , \wAIn93[25] , \wAIn93[24] , \wAIn93[23] , \wAIn93[22] , 
        \wAIn93[21] , \wAIn93[20] , \wAIn93[19] , \wAIn93[18] , \wAIn93[17] , 
        \wAIn93[16] , \wAIn93[15] , \wAIn93[14] , \wAIn93[13] , \wAIn93[12] , 
        \wAIn93[11] , \wAIn93[10] , \wAIn93[9] , \wAIn93[8] , \wAIn93[7] , 
        \wAIn93[6] , \wAIn93[5] , \wAIn93[4] , \wAIn93[3] , \wAIn93[2] , 
        \wAIn93[1] , \wAIn93[0] }), .BIn({\wBIn93[31] , \wBIn93[30] , 
        \wBIn93[29] , \wBIn93[28] , \wBIn93[27] , \wBIn93[26] , \wBIn93[25] , 
        \wBIn93[24] , \wBIn93[23] , \wBIn93[22] , \wBIn93[21] , \wBIn93[20] , 
        \wBIn93[19] , \wBIn93[18] , \wBIn93[17] , \wBIn93[16] , \wBIn93[15] , 
        \wBIn93[14] , \wBIn93[13] , \wBIn93[12] , \wBIn93[11] , \wBIn93[10] , 
        \wBIn93[9] , \wBIn93[8] , \wBIn93[7] , \wBIn93[6] , \wBIn93[5] , 
        \wBIn93[4] , \wBIn93[3] , \wBIn93[2] , \wBIn93[1] , \wBIn93[0] }), 
        .HiOut({\wBMid92[31] , \wBMid92[30] , \wBMid92[29] , \wBMid92[28] , 
        \wBMid92[27] , \wBMid92[26] , \wBMid92[25] , \wBMid92[24] , 
        \wBMid92[23] , \wBMid92[22] , \wBMid92[21] , \wBMid92[20] , 
        \wBMid92[19] , \wBMid92[18] , \wBMid92[17] , \wBMid92[16] , 
        \wBMid92[15] , \wBMid92[14] , \wBMid92[13] , \wBMid92[12] , 
        \wBMid92[11] , \wBMid92[10] , \wBMid92[9] , \wBMid92[8] , \wBMid92[7] , 
        \wBMid92[6] , \wBMid92[5] , \wBMid92[4] , \wBMid92[3] , \wBMid92[2] , 
        \wBMid92[1] , \wBMid92[0] }), .LoOut({\wAMid93[31] , \wAMid93[30] , 
        \wAMid93[29] , \wAMid93[28] , \wAMid93[27] , \wAMid93[26] , 
        \wAMid93[25] , \wAMid93[24] , \wAMid93[23] , \wAMid93[22] , 
        \wAMid93[21] , \wAMid93[20] , \wAMid93[19] , \wAMid93[18] , 
        \wAMid93[17] , \wAMid93[16] , \wAMid93[15] , \wAMid93[14] , 
        \wAMid93[13] , \wAMid93[12] , \wAMid93[11] , \wAMid93[10] , 
        \wAMid93[9] , \wAMid93[8] , \wAMid93[7] , \wAMid93[6] , \wAMid93[5] , 
        \wAMid93[4] , \wAMid93[3] , \wAMid93[2] , \wAMid93[1] , \wAMid93[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid2[31] , 
        \wAMid2[30] , \wAMid2[29] , \wAMid2[28] , \wAMid2[27] , \wAMid2[26] , 
        \wAMid2[25] , \wAMid2[24] , \wAMid2[23] , \wAMid2[22] , \wAMid2[21] , 
        \wAMid2[20] , \wAMid2[19] , \wAMid2[18] , \wAMid2[17] , \wAMid2[16] , 
        \wAMid2[15] , \wAMid2[14] , \wAMid2[13] , \wAMid2[12] , \wAMid2[11] , 
        \wAMid2[10] , \wAMid2[9] , \wAMid2[8] , \wAMid2[7] , \wAMid2[6] , 
        \wAMid2[5] , \wAMid2[4] , \wAMid2[3] , \wAMid2[2] , \wAMid2[1] , 
        \wAMid2[0] }), .BIn({\wBMid2[31] , \wBMid2[30] , \wBMid2[29] , 
        \wBMid2[28] , \wBMid2[27] , \wBMid2[26] , \wBMid2[25] , \wBMid2[24] , 
        \wBMid2[23] , \wBMid2[22] , \wBMid2[21] , \wBMid2[20] , \wBMid2[19] , 
        \wBMid2[18] , \wBMid2[17] , \wBMid2[16] , \wBMid2[15] , \wBMid2[14] , 
        \wBMid2[13] , \wBMid2[12] , \wBMid2[11] , \wBMid2[10] , \wBMid2[9] , 
        \wBMid2[8] , \wBMid2[7] , \wBMid2[6] , \wBMid2[5] , \wBMid2[4] , 
        \wBMid2[3] , \wBMid2[2] , \wBMid2[1] , \wBMid2[0] }), .HiOut({
        \wRegInB2[31] , \wRegInB2[30] , \wRegInB2[29] , \wRegInB2[28] , 
        \wRegInB2[27] , \wRegInB2[26] , \wRegInB2[25] , \wRegInB2[24] , 
        \wRegInB2[23] , \wRegInB2[22] , \wRegInB2[21] , \wRegInB2[20] , 
        \wRegInB2[19] , \wRegInB2[18] , \wRegInB2[17] , \wRegInB2[16] , 
        \wRegInB2[15] , \wRegInB2[14] , \wRegInB2[13] , \wRegInB2[12] , 
        \wRegInB2[11] , \wRegInB2[10] , \wRegInB2[9] , \wRegInB2[8] , 
        \wRegInB2[7] , \wRegInB2[6] , \wRegInB2[5] , \wRegInB2[4] , 
        \wRegInB2[3] , \wRegInB2[2] , \wRegInB2[1] , \wRegInB2[0] }), .LoOut({
        \wRegInA3[31] , \wRegInA3[30] , \wRegInA3[29] , \wRegInA3[28] , 
        \wRegInA3[27] , \wRegInA3[26] , \wRegInA3[25] , \wRegInA3[24] , 
        \wRegInA3[23] , \wRegInA3[22] , \wRegInA3[21] , \wRegInA3[20] , 
        \wRegInA3[19] , \wRegInA3[18] , \wRegInA3[17] , \wRegInA3[16] , 
        \wRegInA3[15] , \wRegInA3[14] , \wRegInA3[13] , \wRegInA3[12] , 
        \wRegInA3[11] , \wRegInA3[10] , \wRegInA3[9] , \wRegInA3[8] , 
        \wRegInA3[7] , \wRegInA3[6] , \wRegInA3[5] , \wRegInA3[4] , 
        \wRegInA3[3] , \wRegInA3[2] , \wRegInA3[1] , \wRegInA3[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid84[31] , \wAMid84[30] , \wAMid84[29] , \wAMid84[28] , 
        \wAMid84[27] , \wAMid84[26] , \wAMid84[25] , \wAMid84[24] , 
        \wAMid84[23] , \wAMid84[22] , \wAMid84[21] , \wAMid84[20] , 
        \wAMid84[19] , \wAMid84[18] , \wAMid84[17] , \wAMid84[16] , 
        \wAMid84[15] , \wAMid84[14] , \wAMid84[13] , \wAMid84[12] , 
        \wAMid84[11] , \wAMid84[10] , \wAMid84[9] , \wAMid84[8] , \wAMid84[7] , 
        \wAMid84[6] , \wAMid84[5] , \wAMid84[4] , \wAMid84[3] , \wAMid84[2] , 
        \wAMid84[1] , \wAMid84[0] }), .BIn({\wBMid84[31] , \wBMid84[30] , 
        \wBMid84[29] , \wBMid84[28] , \wBMid84[27] , \wBMid84[26] , 
        \wBMid84[25] , \wBMid84[24] , \wBMid84[23] , \wBMid84[22] , 
        \wBMid84[21] , \wBMid84[20] , \wBMid84[19] , \wBMid84[18] , 
        \wBMid84[17] , \wBMid84[16] , \wBMid84[15] , \wBMid84[14] , 
        \wBMid84[13] , \wBMid84[12] , \wBMid84[11] , \wBMid84[10] , 
        \wBMid84[9] , \wBMid84[8] , \wBMid84[7] , \wBMid84[6] , \wBMid84[5] , 
        \wBMid84[4] , \wBMid84[3] , \wBMid84[2] , \wBMid84[1] , \wBMid84[0] }), 
        .HiOut({\wRegInB84[31] , \wRegInB84[30] , \wRegInB84[29] , 
        \wRegInB84[28] , \wRegInB84[27] , \wRegInB84[26] , \wRegInB84[25] , 
        \wRegInB84[24] , \wRegInB84[23] , \wRegInB84[22] , \wRegInB84[21] , 
        \wRegInB84[20] , \wRegInB84[19] , \wRegInB84[18] , \wRegInB84[17] , 
        \wRegInB84[16] , \wRegInB84[15] , \wRegInB84[14] , \wRegInB84[13] , 
        \wRegInB84[12] , \wRegInB84[11] , \wRegInB84[10] , \wRegInB84[9] , 
        \wRegInB84[8] , \wRegInB84[7] , \wRegInB84[6] , \wRegInB84[5] , 
        \wRegInB84[4] , \wRegInB84[3] , \wRegInB84[2] , \wRegInB84[1] , 
        \wRegInB84[0] }), .LoOut({\wRegInA85[31] , \wRegInA85[30] , 
        \wRegInA85[29] , \wRegInA85[28] , \wRegInA85[27] , \wRegInA85[26] , 
        \wRegInA85[25] , \wRegInA85[24] , \wRegInA85[23] , \wRegInA85[22] , 
        \wRegInA85[21] , \wRegInA85[20] , \wRegInA85[19] , \wRegInA85[18] , 
        \wRegInA85[17] , \wRegInA85[16] , \wRegInA85[15] , \wRegInA85[14] , 
        \wRegInA85[13] , \wRegInA85[12] , \wRegInA85[11] , \wRegInA85[10] , 
        \wRegInA85[9] , \wRegInA85[8] , \wRegInA85[7] , \wRegInA85[6] , 
        \wRegInA85[5] , \wRegInA85[4] , \wRegInA85[3] , \wRegInA85[2] , 
        \wRegInA85[1] , \wRegInA85[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_196 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink197[31] , \ScanLink197[30] , \ScanLink197[29] , 
        \ScanLink197[28] , \ScanLink197[27] , \ScanLink197[26] , 
        \ScanLink197[25] , \ScanLink197[24] , \ScanLink197[23] , 
        \ScanLink197[22] , \ScanLink197[21] , \ScanLink197[20] , 
        \ScanLink197[19] , \ScanLink197[18] , \ScanLink197[17] , 
        \ScanLink197[16] , \ScanLink197[15] , \ScanLink197[14] , 
        \ScanLink197[13] , \ScanLink197[12] , \ScanLink197[11] , 
        \ScanLink197[10] , \ScanLink197[9] , \ScanLink197[8] , 
        \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , \ScanLink197[4] , 
        \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , \ScanLink197[0] 
        }), .ScanOut({\ScanLink196[31] , \ScanLink196[30] , \ScanLink196[29] , 
        \ScanLink196[28] , \ScanLink196[27] , \ScanLink196[26] , 
        \ScanLink196[25] , \ScanLink196[24] , \ScanLink196[23] , 
        \ScanLink196[22] , \ScanLink196[21] , \ScanLink196[20] , 
        \ScanLink196[19] , \ScanLink196[18] , \ScanLink196[17] , 
        \ScanLink196[16] , \ScanLink196[15] , \ScanLink196[14] , 
        \ScanLink196[13] , \ScanLink196[12] , \ScanLink196[11] , 
        \ScanLink196[10] , \ScanLink196[9] , \ScanLink196[8] , 
        \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , \ScanLink196[4] , 
        \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , \ScanLink196[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB29[31] , \wRegInB29[30] , \wRegInB29[29] , 
        \wRegInB29[28] , \wRegInB29[27] , \wRegInB29[26] , \wRegInB29[25] , 
        \wRegInB29[24] , \wRegInB29[23] , \wRegInB29[22] , \wRegInB29[21] , 
        \wRegInB29[20] , \wRegInB29[19] , \wRegInB29[18] , \wRegInB29[17] , 
        \wRegInB29[16] , \wRegInB29[15] , \wRegInB29[14] , \wRegInB29[13] , 
        \wRegInB29[12] , \wRegInB29[11] , \wRegInB29[10] , \wRegInB29[9] , 
        \wRegInB29[8] , \wRegInB29[7] , \wRegInB29[6] , \wRegInB29[5] , 
        \wRegInB29[4] , \wRegInB29[3] , \wRegInB29[2] , \wRegInB29[1] , 
        \wRegInB29[0] }), .Out({\wBIn29[31] , \wBIn29[30] , \wBIn29[29] , 
        \wBIn29[28] , \wBIn29[27] , \wBIn29[26] , \wBIn29[25] , \wBIn29[24] , 
        \wBIn29[23] , \wBIn29[22] , \wBIn29[21] , \wBIn29[20] , \wBIn29[19] , 
        \wBIn29[18] , \wBIn29[17] , \wBIn29[16] , \wBIn29[15] , \wBIn29[14] , 
        \wBIn29[13] , \wBIn29[12] , \wBIn29[11] , \wBIn29[10] , \wBIn29[9] , 
        \wBIn29[8] , \wBIn29[7] , \wBIn29[6] , \wBIn29[5] , \wBIn29[4] , 
        \wBIn29[3] , \wBIn29[2] , \wBIn29[1] , \wBIn29[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_9 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[31] , \ScanLink10[30] , \ScanLink10[29] , 
        \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , \ScanLink10[25] , 
        \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , \ScanLink10[21] , 
        \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , \ScanLink10[17] , 
        \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , \ScanLink10[13] , 
        \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , \ScanLink10[9] , 
        \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA123[31] , \wRegInA123[30] , 
        \wRegInA123[29] , \wRegInA123[28] , \wRegInA123[27] , \wRegInA123[26] , 
        \wRegInA123[25] , \wRegInA123[24] , \wRegInA123[23] , \wRegInA123[22] , 
        \wRegInA123[21] , \wRegInA123[20] , \wRegInA123[19] , \wRegInA123[18] , 
        \wRegInA123[17] , \wRegInA123[16] , \wRegInA123[15] , \wRegInA123[14] , 
        \wRegInA123[13] , \wRegInA123[12] , \wRegInA123[11] , \wRegInA123[10] , 
        \wRegInA123[9] , \wRegInA123[8] , \wRegInA123[7] , \wRegInA123[6] , 
        \wRegInA123[5] , \wRegInA123[4] , \wRegInA123[3] , \wRegInA123[2] , 
        \wRegInA123[1] , \wRegInA123[0] }), .Out({\wAIn123[31] , \wAIn123[30] , 
        \wAIn123[29] , \wAIn123[28] , \wAIn123[27] , \wAIn123[26] , 
        \wAIn123[25] , \wAIn123[24] , \wAIn123[23] , \wAIn123[22] , 
        \wAIn123[21] , \wAIn123[20] , \wAIn123[19] , \wAIn123[18] , 
        \wAIn123[17] , \wAIn123[16] , \wAIn123[15] , \wAIn123[14] , 
        \wAIn123[13] , \wAIn123[12] , \wAIn123[11] , \wAIn123[10] , 
        \wAIn123[9] , \wAIn123[8] , \wAIn123[7] , \wAIn123[6] , \wAIn123[5] , 
        \wAIn123[4] , \wAIn123[3] , \wAIn123[2] , \wAIn123[1] , \wAIn123[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn56[31] , \wAIn56[30] , \wAIn56[29] , \wAIn56[28] , \wAIn56[27] , 
        \wAIn56[26] , \wAIn56[25] , \wAIn56[24] , \wAIn56[23] , \wAIn56[22] , 
        \wAIn56[21] , \wAIn56[20] , \wAIn56[19] , \wAIn56[18] , \wAIn56[17] , 
        \wAIn56[16] , \wAIn56[15] , \wAIn56[14] , \wAIn56[13] , \wAIn56[12] , 
        \wAIn56[11] , \wAIn56[10] , \wAIn56[9] , \wAIn56[8] , \wAIn56[7] , 
        \wAIn56[6] , \wAIn56[5] , \wAIn56[4] , \wAIn56[3] , \wAIn56[2] , 
        \wAIn56[1] , \wAIn56[0] }), .BIn({\wBIn56[31] , \wBIn56[30] , 
        \wBIn56[29] , \wBIn56[28] , \wBIn56[27] , \wBIn56[26] , \wBIn56[25] , 
        \wBIn56[24] , \wBIn56[23] , \wBIn56[22] , \wBIn56[21] , \wBIn56[20] , 
        \wBIn56[19] , \wBIn56[18] , \wBIn56[17] , \wBIn56[16] , \wBIn56[15] , 
        \wBIn56[14] , \wBIn56[13] , \wBIn56[12] , \wBIn56[11] , \wBIn56[10] , 
        \wBIn56[9] , \wBIn56[8] , \wBIn56[7] , \wBIn56[6] , \wBIn56[5] , 
        \wBIn56[4] , \wBIn56[3] , \wBIn56[2] , \wBIn56[1] , \wBIn56[0] }), 
        .HiOut({\wBMid55[31] , \wBMid55[30] , \wBMid55[29] , \wBMid55[28] , 
        \wBMid55[27] , \wBMid55[26] , \wBMid55[25] , \wBMid55[24] , 
        \wBMid55[23] , \wBMid55[22] , \wBMid55[21] , \wBMid55[20] , 
        \wBMid55[19] , \wBMid55[18] , \wBMid55[17] , \wBMid55[16] , 
        \wBMid55[15] , \wBMid55[14] , \wBMid55[13] , \wBMid55[12] , 
        \wBMid55[11] , \wBMid55[10] , \wBMid55[9] , \wBMid55[8] , \wBMid55[7] , 
        \wBMid55[6] , \wBMid55[5] , \wBMid55[4] , \wBMid55[3] , \wBMid55[2] , 
        \wBMid55[1] , \wBMid55[0] }), .LoOut({\wAMid56[31] , \wAMid56[30] , 
        \wAMid56[29] , \wAMid56[28] , \wAMid56[27] , \wAMid56[26] , 
        \wAMid56[25] , \wAMid56[24] , \wAMid56[23] , \wAMid56[22] , 
        \wAMid56[21] , \wAMid56[20] , \wAMid56[19] , \wAMid56[18] , 
        \wAMid56[17] , \wAMid56[16] , \wAMid56[15] , \wAMid56[14] , 
        \wAMid56[13] , \wAMid56[12] , \wAMid56[11] , \wAMid56[10] , 
        \wAMid56[9] , \wAMid56[8] , \wAMid56[7] , \wAMid56[6] , \wAMid56[5] , 
        \wAMid56[4] , \wAMid56[3] , \wAMid56[2] , \wAMid56[1] , \wAMid56[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn94[31] , \wAIn94[30] , \wAIn94[29] , \wAIn94[28] , \wAIn94[27] , 
        \wAIn94[26] , \wAIn94[25] , \wAIn94[24] , \wAIn94[23] , \wAIn94[22] , 
        \wAIn94[21] , \wAIn94[20] , \wAIn94[19] , \wAIn94[18] , \wAIn94[17] , 
        \wAIn94[16] , \wAIn94[15] , \wAIn94[14] , \wAIn94[13] , \wAIn94[12] , 
        \wAIn94[11] , \wAIn94[10] , \wAIn94[9] , \wAIn94[8] , \wAIn94[7] , 
        \wAIn94[6] , \wAIn94[5] , \wAIn94[4] , \wAIn94[3] , \wAIn94[2] , 
        \wAIn94[1] , \wAIn94[0] }), .BIn({\wBIn94[31] , \wBIn94[30] , 
        \wBIn94[29] , \wBIn94[28] , \wBIn94[27] , \wBIn94[26] , \wBIn94[25] , 
        \wBIn94[24] , \wBIn94[23] , \wBIn94[22] , \wBIn94[21] , \wBIn94[20] , 
        \wBIn94[19] , \wBIn94[18] , \wBIn94[17] , \wBIn94[16] , \wBIn94[15] , 
        \wBIn94[14] , \wBIn94[13] , \wBIn94[12] , \wBIn94[11] , \wBIn94[10] , 
        \wBIn94[9] , \wBIn94[8] , \wBIn94[7] , \wBIn94[6] , \wBIn94[5] , 
        \wBIn94[4] , \wBIn94[3] , \wBIn94[2] , \wBIn94[1] , \wBIn94[0] }), 
        .HiOut({\wBMid93[31] , \wBMid93[30] , \wBMid93[29] , \wBMid93[28] , 
        \wBMid93[27] , \wBMid93[26] , \wBMid93[25] , \wBMid93[24] , 
        \wBMid93[23] , \wBMid93[22] , \wBMid93[21] , \wBMid93[20] , 
        \wBMid93[19] , \wBMid93[18] , \wBMid93[17] , \wBMid93[16] , 
        \wBMid93[15] , \wBMid93[14] , \wBMid93[13] , \wBMid93[12] , 
        \wBMid93[11] , \wBMid93[10] , \wBMid93[9] , \wBMid93[8] , \wBMid93[7] , 
        \wBMid93[6] , \wBMid93[5] , \wBMid93[4] , \wBMid93[3] , \wBMid93[2] , 
        \wBMid93[1] , \wBMid93[0] }), .LoOut({\wAMid94[31] , \wAMid94[30] , 
        \wAMid94[29] , \wAMid94[28] , \wAMid94[27] , \wAMid94[26] , 
        \wAMid94[25] , \wAMid94[24] , \wAMid94[23] , \wAMid94[22] , 
        \wAMid94[21] , \wAMid94[20] , \wAMid94[19] , \wAMid94[18] , 
        \wAMid94[17] , \wAMid94[16] , \wAMid94[15] , \wAMid94[14] , 
        \wAMid94[13] , \wAMid94[12] , \wAMid94[11] , \wAMid94[10] , 
        \wAMid94[9] , \wAMid94[8] , \wAMid94[7] , \wAMid94[6] , \wAMid94[5] , 
        \wAMid94[4] , \wAMid94[3] , \wAMid94[2] , \wAMid94[1] , \wAMid94[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_191 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink192[31] , \ScanLink192[30] , \ScanLink192[29] , 
        \ScanLink192[28] , \ScanLink192[27] , \ScanLink192[26] , 
        \ScanLink192[25] , \ScanLink192[24] , \ScanLink192[23] , 
        \ScanLink192[22] , \ScanLink192[21] , \ScanLink192[20] , 
        \ScanLink192[19] , \ScanLink192[18] , \ScanLink192[17] , 
        \ScanLink192[16] , \ScanLink192[15] , \ScanLink192[14] , 
        \ScanLink192[13] , \ScanLink192[12] , \ScanLink192[11] , 
        \ScanLink192[10] , \ScanLink192[9] , \ScanLink192[8] , 
        \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , \ScanLink192[4] , 
        \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , \ScanLink192[0] 
        }), .ScanOut({\ScanLink191[31] , \ScanLink191[30] , \ScanLink191[29] , 
        \ScanLink191[28] , \ScanLink191[27] , \ScanLink191[26] , 
        \ScanLink191[25] , \ScanLink191[24] , \ScanLink191[23] , 
        \ScanLink191[22] , \ScanLink191[21] , \ScanLink191[20] , 
        \ScanLink191[19] , \ScanLink191[18] , \ScanLink191[17] , 
        \ScanLink191[16] , \ScanLink191[15] , \ScanLink191[14] , 
        \ScanLink191[13] , \ScanLink191[12] , \ScanLink191[11] , 
        \ScanLink191[10] , \ScanLink191[9] , \ScanLink191[8] , 
        \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , \ScanLink191[4] , 
        \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , \ScanLink191[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA32[31] , \wRegInA32[30] , \wRegInA32[29] , 
        \wRegInA32[28] , \wRegInA32[27] , \wRegInA32[26] , \wRegInA32[25] , 
        \wRegInA32[24] , \wRegInA32[23] , \wRegInA32[22] , \wRegInA32[21] , 
        \wRegInA32[20] , \wRegInA32[19] , \wRegInA32[18] , \wRegInA32[17] , 
        \wRegInA32[16] , \wRegInA32[15] , \wRegInA32[14] , \wRegInA32[13] , 
        \wRegInA32[12] , \wRegInA32[11] , \wRegInA32[10] , \wRegInA32[9] , 
        \wRegInA32[8] , \wRegInA32[7] , \wRegInA32[6] , \wRegInA32[5] , 
        \wRegInA32[4] , \wRegInA32[3] , \wRegInA32[2] , \wRegInA32[1] , 
        \wRegInA32[0] }), .Out({\wAIn32[31] , \wAIn32[30] , \wAIn32[29] , 
        \wAIn32[28] , \wAIn32[27] , \wAIn32[26] , \wAIn32[25] , \wAIn32[24] , 
        \wAIn32[23] , \wAIn32[22] , \wAIn32[21] , \wAIn32[20] , \wAIn32[19] , 
        \wAIn32[18] , \wAIn32[17] , \wAIn32[16] , \wAIn32[15] , \wAIn32[14] , 
        \wAIn32[13] , \wAIn32[12] , \wAIn32[11] , \wAIn32[10] , \wAIn32[9] , 
        \wAIn32[8] , \wAIn32[7] , \wAIn32[6] , \wAIn32[5] , \wAIn32[4] , 
        \wAIn32[3] , \wAIn32[2] , \wAIn32[1] , \wAIn32[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn126[31] , \wAIn126[30] , \wAIn126[29] , \wAIn126[28] , 
        \wAIn126[27] , \wAIn126[26] , \wAIn126[25] , \wAIn126[24] , 
        \wAIn126[23] , \wAIn126[22] , \wAIn126[21] , \wAIn126[20] , 
        \wAIn126[19] , \wAIn126[18] , \wAIn126[17] , \wAIn126[16] , 
        \wAIn126[15] , \wAIn126[14] , \wAIn126[13] , \wAIn126[12] , 
        \wAIn126[11] , \wAIn126[10] , \wAIn126[9] , \wAIn126[8] , \wAIn126[7] , 
        \wAIn126[6] , \wAIn126[5] , \wAIn126[4] , \wAIn126[3] , \wAIn126[2] , 
        \wAIn126[1] , \wAIn126[0] }), .BIn({\wBIn126[31] , \wBIn126[30] , 
        \wBIn126[29] , \wBIn126[28] , \wBIn126[27] , \wBIn126[26] , 
        \wBIn126[25] , \wBIn126[24] , \wBIn126[23] , \wBIn126[22] , 
        \wBIn126[21] , \wBIn126[20] , \wBIn126[19] , \wBIn126[18] , 
        \wBIn126[17] , \wBIn126[16] , \wBIn126[15] , \wBIn126[14] , 
        \wBIn126[13] , \wBIn126[12] , \wBIn126[11] , \wBIn126[10] , 
        \wBIn126[9] , \wBIn126[8] , \wBIn126[7] , \wBIn126[6] , \wBIn126[5] , 
        \wBIn126[4] , \wBIn126[3] , \wBIn126[2] , \wBIn126[1] , \wBIn126[0] }), 
        .HiOut({\wBMid125[31] , \wBMid125[30] , \wBMid125[29] , \wBMid125[28] , 
        \wBMid125[27] , \wBMid125[26] , \wBMid125[25] , \wBMid125[24] , 
        \wBMid125[23] , \wBMid125[22] , \wBMid125[21] , \wBMid125[20] , 
        \wBMid125[19] , \wBMid125[18] , \wBMid125[17] , \wBMid125[16] , 
        \wBMid125[15] , \wBMid125[14] , \wBMid125[13] , \wBMid125[12] , 
        \wBMid125[11] , \wBMid125[10] , \wBMid125[9] , \wBMid125[8] , 
        \wBMid125[7] , \wBMid125[6] , \wBMid125[5] , \wBMid125[4] , 
        \wBMid125[3] , \wBMid125[2] , \wBMid125[1] , \wBMid125[0] }), .LoOut({
        \wAMid126[31] , \wAMid126[30] , \wAMid126[29] , \wAMid126[28] , 
        \wAMid126[27] , \wAMid126[26] , \wAMid126[25] , \wAMid126[24] , 
        \wAMid126[23] , \wAMid126[22] , \wAMid126[21] , \wAMid126[20] , 
        \wAMid126[19] , \wAMid126[18] , \wAMid126[17] , \wAMid126[16] , 
        \wAMid126[15] , \wAMid126[14] , \wAMid126[13] , \wAMid126[12] , 
        \wAMid126[11] , \wAMid126[10] , \wAMid126[9] , \wAMid126[8] , 
        \wAMid126[7] , \wAMid126[6] , \wAMid126[5] , \wAMid126[4] , 
        \wAMid126[3] , \wAMid126[2] , \wAMid126[1] , \wAMid126[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid5[31] , 
        \wAMid5[30] , \wAMid5[29] , \wAMid5[28] , \wAMid5[27] , \wAMid5[26] , 
        \wAMid5[25] , \wAMid5[24] , \wAMid5[23] , \wAMid5[22] , \wAMid5[21] , 
        \wAMid5[20] , \wAMid5[19] , \wAMid5[18] , \wAMid5[17] , \wAMid5[16] , 
        \wAMid5[15] , \wAMid5[14] , \wAMid5[13] , \wAMid5[12] , \wAMid5[11] , 
        \wAMid5[10] , \wAMid5[9] , \wAMid5[8] , \wAMid5[7] , \wAMid5[6] , 
        \wAMid5[5] , \wAMid5[4] , \wAMid5[3] , \wAMid5[2] , \wAMid5[1] , 
        \wAMid5[0] }), .BIn({\wBMid5[31] , \wBMid5[30] , \wBMid5[29] , 
        \wBMid5[28] , \wBMid5[27] , \wBMid5[26] , \wBMid5[25] , \wBMid5[24] , 
        \wBMid5[23] , \wBMid5[22] , \wBMid5[21] , \wBMid5[20] , \wBMid5[19] , 
        \wBMid5[18] , \wBMid5[17] , \wBMid5[16] , \wBMid5[15] , \wBMid5[14] , 
        \wBMid5[13] , \wBMid5[12] , \wBMid5[11] , \wBMid5[10] , \wBMid5[9] , 
        \wBMid5[8] , \wBMid5[7] , \wBMid5[6] , \wBMid5[5] , \wBMid5[4] , 
        \wBMid5[3] , \wBMid5[2] , \wBMid5[1] , \wBMid5[0] }), .HiOut({
        \wRegInB5[31] , \wRegInB5[30] , \wRegInB5[29] , \wRegInB5[28] , 
        \wRegInB5[27] , \wRegInB5[26] , \wRegInB5[25] , \wRegInB5[24] , 
        \wRegInB5[23] , \wRegInB5[22] , \wRegInB5[21] , \wRegInB5[20] , 
        \wRegInB5[19] , \wRegInB5[18] , \wRegInB5[17] , \wRegInB5[16] , 
        \wRegInB5[15] , \wRegInB5[14] , \wRegInB5[13] , \wRegInB5[12] , 
        \wRegInB5[11] , \wRegInB5[10] , \wRegInB5[9] , \wRegInB5[8] , 
        \wRegInB5[7] , \wRegInB5[6] , \wRegInB5[5] , \wRegInB5[4] , 
        \wRegInB5[3] , \wRegInB5[2] , \wRegInB5[1] , \wRegInB5[0] }), .LoOut({
        \wRegInA6[31] , \wRegInA6[30] , \wRegInA6[29] , \wRegInA6[28] , 
        \wRegInA6[27] , \wRegInA6[26] , \wRegInA6[25] , \wRegInA6[24] , 
        \wRegInA6[23] , \wRegInA6[22] , \wRegInA6[21] , \wRegInA6[20] , 
        \wRegInA6[19] , \wRegInA6[18] , \wRegInA6[17] , \wRegInA6[16] , 
        \wRegInA6[15] , \wRegInA6[14] , \wRegInA6[13] , \wRegInA6[12] , 
        \wRegInA6[11] , \wRegInA6[10] , \wRegInA6[9] , \wRegInA6[8] , 
        \wRegInA6[7] , \wRegInA6[6] , \wRegInA6[5] , \wRegInA6[4] , 
        \wRegInA6[3] , \wRegInA6[2] , \wRegInA6[1] , \wRegInA6[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid83[31] , \wAMid83[30] , \wAMid83[29] , \wAMid83[28] , 
        \wAMid83[27] , \wAMid83[26] , \wAMid83[25] , \wAMid83[24] , 
        \wAMid83[23] , \wAMid83[22] , \wAMid83[21] , \wAMid83[20] , 
        \wAMid83[19] , \wAMid83[18] , \wAMid83[17] , \wAMid83[16] , 
        \wAMid83[15] , \wAMid83[14] , \wAMid83[13] , \wAMid83[12] , 
        \wAMid83[11] , \wAMid83[10] , \wAMid83[9] , \wAMid83[8] , \wAMid83[7] , 
        \wAMid83[6] , \wAMid83[5] , \wAMid83[4] , \wAMid83[3] , \wAMid83[2] , 
        \wAMid83[1] , \wAMid83[0] }), .BIn({\wBMid83[31] , \wBMid83[30] , 
        \wBMid83[29] , \wBMid83[28] , \wBMid83[27] , \wBMid83[26] , 
        \wBMid83[25] , \wBMid83[24] , \wBMid83[23] , \wBMid83[22] , 
        \wBMid83[21] , \wBMid83[20] , \wBMid83[19] , \wBMid83[18] , 
        \wBMid83[17] , \wBMid83[16] , \wBMid83[15] , \wBMid83[14] , 
        \wBMid83[13] , \wBMid83[12] , \wBMid83[11] , \wBMid83[10] , 
        \wBMid83[9] , \wBMid83[8] , \wBMid83[7] , \wBMid83[6] , \wBMid83[5] , 
        \wBMid83[4] , \wBMid83[3] , \wBMid83[2] , \wBMid83[1] , \wBMid83[0] }), 
        .HiOut({\wRegInB83[31] , \wRegInB83[30] , \wRegInB83[29] , 
        \wRegInB83[28] , \wRegInB83[27] , \wRegInB83[26] , \wRegInB83[25] , 
        \wRegInB83[24] , \wRegInB83[23] , \wRegInB83[22] , \wRegInB83[21] , 
        \wRegInB83[20] , \wRegInB83[19] , \wRegInB83[18] , \wRegInB83[17] , 
        \wRegInB83[16] , \wRegInB83[15] , \wRegInB83[14] , \wRegInB83[13] , 
        \wRegInB83[12] , \wRegInB83[11] , \wRegInB83[10] , \wRegInB83[9] , 
        \wRegInB83[8] , \wRegInB83[7] , \wRegInB83[6] , \wRegInB83[5] , 
        \wRegInB83[4] , \wRegInB83[3] , \wRegInB83[2] , \wRegInB83[1] , 
        \wRegInB83[0] }), .LoOut({\wRegInA84[31] , \wRegInA84[30] , 
        \wRegInA84[29] , \wRegInA84[28] , \wRegInA84[27] , \wRegInA84[26] , 
        \wRegInA84[25] , \wRegInA84[24] , \wRegInA84[23] , \wRegInA84[22] , 
        \wRegInA84[21] , \wRegInA84[20] , \wRegInA84[19] , \wRegInA84[18] , 
        \wRegInA84[17] , \wRegInA84[16] , \wRegInA84[15] , \wRegInA84[14] , 
        \wRegInA84[13] , \wRegInA84[12] , \wRegInA84[11] , \wRegInA84[10] , 
        \wRegInA84[9] , \wRegInA84[8] , \wRegInA84[7] , \wRegInA84[6] , 
        \wRegInA84[5] , \wRegInA84[4] , \wRegInA84[3] , \wRegInA84[2] , 
        \wRegInA84[1] , \wRegInA84[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_88 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink89[31] , \ScanLink89[30] , \ScanLink89[29] , 
        \ScanLink89[28] , \ScanLink89[27] , \ScanLink89[26] , \ScanLink89[25] , 
        \ScanLink89[24] , \ScanLink89[23] , \ScanLink89[22] , \ScanLink89[21] , 
        \ScanLink89[20] , \ScanLink89[19] , \ScanLink89[18] , \ScanLink89[17] , 
        \ScanLink89[16] , \ScanLink89[15] , \ScanLink89[14] , \ScanLink89[13] , 
        \ScanLink89[12] , \ScanLink89[11] , \ScanLink89[10] , \ScanLink89[9] , 
        \ScanLink89[8] , \ScanLink89[7] , \ScanLink89[6] , \ScanLink89[5] , 
        \ScanLink89[4] , \ScanLink89[3] , \ScanLink89[2] , \ScanLink89[1] , 
        \ScanLink89[0] }), .ScanOut({\ScanLink88[31] , \ScanLink88[30] , 
        \ScanLink88[29] , \ScanLink88[28] , \ScanLink88[27] , \ScanLink88[26] , 
        \ScanLink88[25] , \ScanLink88[24] , \ScanLink88[23] , \ScanLink88[22] , 
        \ScanLink88[21] , \ScanLink88[20] , \ScanLink88[19] , \ScanLink88[18] , 
        \ScanLink88[17] , \ScanLink88[16] , \ScanLink88[15] , \ScanLink88[14] , 
        \ScanLink88[13] , \ScanLink88[12] , \ScanLink88[11] , \ScanLink88[10] , 
        \ScanLink88[9] , \ScanLink88[8] , \ScanLink88[7] , \ScanLink88[6] , 
        \ScanLink88[5] , \ScanLink88[4] , \ScanLink88[3] , \ScanLink88[2] , 
        \ScanLink88[1] , \ScanLink88[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB83[31] , \wRegInB83[30] , 
        \wRegInB83[29] , \wRegInB83[28] , \wRegInB83[27] , \wRegInB83[26] , 
        \wRegInB83[25] , \wRegInB83[24] , \wRegInB83[23] , \wRegInB83[22] , 
        \wRegInB83[21] , \wRegInB83[20] , \wRegInB83[19] , \wRegInB83[18] , 
        \wRegInB83[17] , \wRegInB83[16] , \wRegInB83[15] , \wRegInB83[14] , 
        \wRegInB83[13] , \wRegInB83[12] , \wRegInB83[11] , \wRegInB83[10] , 
        \wRegInB83[9] , \wRegInB83[8] , \wRegInB83[7] , \wRegInB83[6] , 
        \wRegInB83[5] , \wRegInB83[4] , \wRegInB83[3] , \wRegInB83[2] , 
        \wRegInB83[1] , \wRegInB83[0] }), .Out({\wBIn83[31] , \wBIn83[30] , 
        \wBIn83[29] , \wBIn83[28] , \wBIn83[27] , \wBIn83[26] , \wBIn83[25] , 
        \wBIn83[24] , \wBIn83[23] , \wBIn83[22] , \wBIn83[21] , \wBIn83[20] , 
        \wBIn83[19] , \wBIn83[18] , \wBIn83[17] , \wBIn83[16] , \wBIn83[15] , 
        \wBIn83[14] , \wBIn83[13] , \wBIn83[12] , \wBIn83[11] , \wBIn83[10] , 
        \wBIn83[9] , \wBIn83[8] , \wBIn83[7] , \wBIn83[6] , \wBIn83[5] , 
        \wBIn83[4] , \wBIn83[3] , \wBIn83[2] , \wBIn83[1] , \wBIn83[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn71[31] , \wAIn71[30] , \wAIn71[29] , \wAIn71[28] , \wAIn71[27] , 
        \wAIn71[26] , \wAIn71[25] , \wAIn71[24] , \wAIn71[23] , \wAIn71[22] , 
        \wAIn71[21] , \wAIn71[20] , \wAIn71[19] , \wAIn71[18] , \wAIn71[17] , 
        \wAIn71[16] , \wAIn71[15] , \wAIn71[14] , \wAIn71[13] , \wAIn71[12] , 
        \wAIn71[11] , \wAIn71[10] , \wAIn71[9] , \wAIn71[8] , \wAIn71[7] , 
        \wAIn71[6] , \wAIn71[5] , \wAIn71[4] , \wAIn71[3] , \wAIn71[2] , 
        \wAIn71[1] , \wAIn71[0] }), .BIn({\wBIn71[31] , \wBIn71[30] , 
        \wBIn71[29] , \wBIn71[28] , \wBIn71[27] , \wBIn71[26] , \wBIn71[25] , 
        \wBIn71[24] , \wBIn71[23] , \wBIn71[22] , \wBIn71[21] , \wBIn71[20] , 
        \wBIn71[19] , \wBIn71[18] , \wBIn71[17] , \wBIn71[16] , \wBIn71[15] , 
        \wBIn71[14] , \wBIn71[13] , \wBIn71[12] , \wBIn71[11] , \wBIn71[10] , 
        \wBIn71[9] , \wBIn71[8] , \wBIn71[7] , \wBIn71[6] , \wBIn71[5] , 
        \wBIn71[4] , \wBIn71[3] , \wBIn71[2] , \wBIn71[1] , \wBIn71[0] }), 
        .HiOut({\wBMid70[31] , \wBMid70[30] , \wBMid70[29] , \wBMid70[28] , 
        \wBMid70[27] , \wBMid70[26] , \wBMid70[25] , \wBMid70[24] , 
        \wBMid70[23] , \wBMid70[22] , \wBMid70[21] , \wBMid70[20] , 
        \wBMid70[19] , \wBMid70[18] , \wBMid70[17] , \wBMid70[16] , 
        \wBMid70[15] , \wBMid70[14] , \wBMid70[13] , \wBMid70[12] , 
        \wBMid70[11] , \wBMid70[10] , \wBMid70[9] , \wBMid70[8] , \wBMid70[7] , 
        \wBMid70[6] , \wBMid70[5] , \wBMid70[4] , \wBMid70[3] , \wBMid70[2] , 
        \wBMid70[1] , \wBMid70[0] }), .LoOut({\wAMid71[31] , \wAMid71[30] , 
        \wAMid71[29] , \wAMid71[28] , \wAMid71[27] , \wAMid71[26] , 
        \wAMid71[25] , \wAMid71[24] , \wAMid71[23] , \wAMid71[22] , 
        \wAMid71[21] , \wAMid71[20] , \wAMid71[19] , \wAMid71[18] , 
        \wAMid71[17] , \wAMid71[16] , \wAMid71[15] , \wAMid71[14] , 
        \wAMid71[13] , \wAMid71[12] , \wAMid71[11] , \wAMid71[10] , 
        \wAMid71[9] , \wAMid71[8] , \wAMid71[7] , \wAMid71[6] , \wAMid71[5] , 
        \wAMid71[4] , \wAMid71[3] , \wAMid71[2] , \wAMid71[1] , \wAMid71[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid66[31] , \wAMid66[30] , \wAMid66[29] , \wAMid66[28] , 
        \wAMid66[27] , \wAMid66[26] , \wAMid66[25] , \wAMid66[24] , 
        \wAMid66[23] , \wAMid66[22] , \wAMid66[21] , \wAMid66[20] , 
        \wAMid66[19] , \wAMid66[18] , \wAMid66[17] , \wAMid66[16] , 
        \wAMid66[15] , \wAMid66[14] , \wAMid66[13] , \wAMid66[12] , 
        \wAMid66[11] , \wAMid66[10] , \wAMid66[9] , \wAMid66[8] , \wAMid66[7] , 
        \wAMid66[6] , \wAMid66[5] , \wAMid66[4] , \wAMid66[3] , \wAMid66[2] , 
        \wAMid66[1] , \wAMid66[0] }), .BIn({\wBMid66[31] , \wBMid66[30] , 
        \wBMid66[29] , \wBMid66[28] , \wBMid66[27] , \wBMid66[26] , 
        \wBMid66[25] , \wBMid66[24] , \wBMid66[23] , \wBMid66[22] , 
        \wBMid66[21] , \wBMid66[20] , \wBMid66[19] , \wBMid66[18] , 
        \wBMid66[17] , \wBMid66[16] , \wBMid66[15] , \wBMid66[14] , 
        \wBMid66[13] , \wBMid66[12] , \wBMid66[11] , \wBMid66[10] , 
        \wBMid66[9] , \wBMid66[8] , \wBMid66[7] , \wBMid66[6] , \wBMid66[5] , 
        \wBMid66[4] , \wBMid66[3] , \wBMid66[2] , \wBMid66[1] , \wBMid66[0] }), 
        .HiOut({\wRegInB66[31] , \wRegInB66[30] , \wRegInB66[29] , 
        \wRegInB66[28] , \wRegInB66[27] , \wRegInB66[26] , \wRegInB66[25] , 
        \wRegInB66[24] , \wRegInB66[23] , \wRegInB66[22] , \wRegInB66[21] , 
        \wRegInB66[20] , \wRegInB66[19] , \wRegInB66[18] , \wRegInB66[17] , 
        \wRegInB66[16] , \wRegInB66[15] , \wRegInB66[14] , \wRegInB66[13] , 
        \wRegInB66[12] , \wRegInB66[11] , \wRegInB66[10] , \wRegInB66[9] , 
        \wRegInB66[8] , \wRegInB66[7] , \wRegInB66[6] , \wRegInB66[5] , 
        \wRegInB66[4] , \wRegInB66[3] , \wRegInB66[2] , \wRegInB66[1] , 
        \wRegInB66[0] }), .LoOut({\wRegInA67[31] , \wRegInA67[30] , 
        \wRegInA67[29] , \wRegInA67[28] , \wRegInA67[27] , \wRegInA67[26] , 
        \wRegInA67[25] , \wRegInA67[24] , \wRegInA67[23] , \wRegInA67[22] , 
        \wRegInA67[21] , \wRegInA67[20] , \wRegInA67[19] , \wRegInA67[18] , 
        \wRegInA67[17] , \wRegInA67[16] , \wRegInA67[15] , \wRegInA67[14] , 
        \wRegInA67[13] , \wRegInA67[12] , \wRegInA67[11] , \wRegInA67[10] , 
        \wRegInA67[9] , \wRegInA67[8] , \wRegInA67[7] , \wRegInA67[6] , 
        \wRegInA67[5] , \wRegInA67[4] , \wRegInA67[3] , \wRegInA67[2] , 
        \wRegInA67[1] , \wRegInA67[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_153 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink154[31] , \ScanLink154[30] , \ScanLink154[29] , 
        \ScanLink154[28] , \ScanLink154[27] , \ScanLink154[26] , 
        \ScanLink154[25] , \ScanLink154[24] , \ScanLink154[23] , 
        \ScanLink154[22] , \ScanLink154[21] , \ScanLink154[20] , 
        \ScanLink154[19] , \ScanLink154[18] , \ScanLink154[17] , 
        \ScanLink154[16] , \ScanLink154[15] , \ScanLink154[14] , 
        \ScanLink154[13] , \ScanLink154[12] , \ScanLink154[11] , 
        \ScanLink154[10] , \ScanLink154[9] , \ScanLink154[8] , 
        \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , \ScanLink154[4] , 
        \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , \ScanLink154[0] 
        }), .ScanOut({\ScanLink153[31] , \ScanLink153[30] , \ScanLink153[29] , 
        \ScanLink153[28] , \ScanLink153[27] , \ScanLink153[26] , 
        \ScanLink153[25] , \ScanLink153[24] , \ScanLink153[23] , 
        \ScanLink153[22] , \ScanLink153[21] , \ScanLink153[20] , 
        \ScanLink153[19] , \ScanLink153[18] , \ScanLink153[17] , 
        \ScanLink153[16] , \ScanLink153[15] , \ScanLink153[14] , 
        \ScanLink153[13] , \ScanLink153[12] , \ScanLink153[11] , 
        \ScanLink153[10] , \ScanLink153[9] , \ScanLink153[8] , 
        \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , \ScanLink153[4] , 
        \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , \ScanLink153[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA51[31] , \wRegInA51[30] , \wRegInA51[29] , 
        \wRegInA51[28] , \wRegInA51[27] , \wRegInA51[26] , \wRegInA51[25] , 
        \wRegInA51[24] , \wRegInA51[23] , \wRegInA51[22] , \wRegInA51[21] , 
        \wRegInA51[20] , \wRegInA51[19] , \wRegInA51[18] , \wRegInA51[17] , 
        \wRegInA51[16] , \wRegInA51[15] , \wRegInA51[14] , \wRegInA51[13] , 
        \wRegInA51[12] , \wRegInA51[11] , \wRegInA51[10] , \wRegInA51[9] , 
        \wRegInA51[8] , \wRegInA51[7] , \wRegInA51[6] , \wRegInA51[5] , 
        \wRegInA51[4] , \wRegInA51[3] , \wRegInA51[2] , \wRegInA51[1] , 
        \wRegInA51[0] }), .Out({\wAIn51[31] , \wAIn51[30] , \wAIn51[29] , 
        \wAIn51[28] , \wAIn51[27] , \wAIn51[26] , \wAIn51[25] , \wAIn51[24] , 
        \wAIn51[23] , \wAIn51[22] , \wAIn51[21] , \wAIn51[20] , \wAIn51[19] , 
        \wAIn51[18] , \wAIn51[17] , \wAIn51[16] , \wAIn51[15] , \wAIn51[14] , 
        \wAIn51[13] , \wAIn51[12] , \wAIn51[11] , \wAIn51[10] , \wAIn51[9] , 
        \wAIn51[8] , \wAIn51[7] , \wAIn51[6] , \wAIn51[5] , \wAIn51[4] , 
        \wAIn51[3] , \wAIn51[2] , \wAIn51[1] , \wAIn51[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn101[31] , \wAIn101[30] , \wAIn101[29] , \wAIn101[28] , 
        \wAIn101[27] , \wAIn101[26] , \wAIn101[25] , \wAIn101[24] , 
        \wAIn101[23] , \wAIn101[22] , \wAIn101[21] , \wAIn101[20] , 
        \wAIn101[19] , \wAIn101[18] , \wAIn101[17] , \wAIn101[16] , 
        \wAIn101[15] , \wAIn101[14] , \wAIn101[13] , \wAIn101[12] , 
        \wAIn101[11] , \wAIn101[10] , \wAIn101[9] , \wAIn101[8] , \wAIn101[7] , 
        \wAIn101[6] , \wAIn101[5] , \wAIn101[4] , \wAIn101[3] , \wAIn101[2] , 
        \wAIn101[1] , \wAIn101[0] }), .BIn({\wBIn101[31] , \wBIn101[30] , 
        \wBIn101[29] , \wBIn101[28] , \wBIn101[27] , \wBIn101[26] , 
        \wBIn101[25] , \wBIn101[24] , \wBIn101[23] , \wBIn101[22] , 
        \wBIn101[21] , \wBIn101[20] , \wBIn101[19] , \wBIn101[18] , 
        \wBIn101[17] , \wBIn101[16] , \wBIn101[15] , \wBIn101[14] , 
        \wBIn101[13] , \wBIn101[12] , \wBIn101[11] , \wBIn101[10] , 
        \wBIn101[9] , \wBIn101[8] , \wBIn101[7] , \wBIn101[6] , \wBIn101[5] , 
        \wBIn101[4] , \wBIn101[3] , \wBIn101[2] , \wBIn101[1] , \wBIn101[0] }), 
        .HiOut({\wBMid100[31] , \wBMid100[30] , \wBMid100[29] , \wBMid100[28] , 
        \wBMid100[27] , \wBMid100[26] , \wBMid100[25] , \wBMid100[24] , 
        \wBMid100[23] , \wBMid100[22] , \wBMid100[21] , \wBMid100[20] , 
        \wBMid100[19] , \wBMid100[18] , \wBMid100[17] , \wBMid100[16] , 
        \wBMid100[15] , \wBMid100[14] , \wBMid100[13] , \wBMid100[12] , 
        \wBMid100[11] , \wBMid100[10] , \wBMid100[9] , \wBMid100[8] , 
        \wBMid100[7] , \wBMid100[6] , \wBMid100[5] , \wBMid100[4] , 
        \wBMid100[3] , \wBMid100[2] , \wBMid100[1] , \wBMid100[0] }), .LoOut({
        \wAMid101[31] , \wAMid101[30] , \wAMid101[29] , \wAMid101[28] , 
        \wAMid101[27] , \wAMid101[26] , \wAMid101[25] , \wAMid101[24] , 
        \wAMid101[23] , \wAMid101[22] , \wAMid101[21] , \wAMid101[20] , 
        \wAMid101[19] , \wAMid101[18] , \wAMid101[17] , \wAMid101[16] , 
        \wAMid101[15] , \wAMid101[14] , \wAMid101[13] , \wAMid101[12] , 
        \wAMid101[11] , \wAMid101[10] , \wAMid101[9] , \wAMid101[8] , 
        \wAMid101[7] , \wAMid101[6] , \wAMid101[5] , \wAMid101[4] , 
        \wAMid101[3] , \wAMid101[2] , \wAMid101[1] , \wAMid101[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid41[31] , \wAMid41[30] , \wAMid41[29] , \wAMid41[28] , 
        \wAMid41[27] , \wAMid41[26] , \wAMid41[25] , \wAMid41[24] , 
        \wAMid41[23] , \wAMid41[22] , \wAMid41[21] , \wAMid41[20] , 
        \wAMid41[19] , \wAMid41[18] , \wAMid41[17] , \wAMid41[16] , 
        \wAMid41[15] , \wAMid41[14] , \wAMid41[13] , \wAMid41[12] , 
        \wAMid41[11] , \wAMid41[10] , \wAMid41[9] , \wAMid41[8] , \wAMid41[7] , 
        \wAMid41[6] , \wAMid41[5] , \wAMid41[4] , \wAMid41[3] , \wAMid41[2] , 
        \wAMid41[1] , \wAMid41[0] }), .BIn({\wBMid41[31] , \wBMid41[30] , 
        \wBMid41[29] , \wBMid41[28] , \wBMid41[27] , \wBMid41[26] , 
        \wBMid41[25] , \wBMid41[24] , \wBMid41[23] , \wBMid41[22] , 
        \wBMid41[21] , \wBMid41[20] , \wBMid41[19] , \wBMid41[18] , 
        \wBMid41[17] , \wBMid41[16] , \wBMid41[15] , \wBMid41[14] , 
        \wBMid41[13] , \wBMid41[12] , \wBMid41[11] , \wBMid41[10] , 
        \wBMid41[9] , \wBMid41[8] , \wBMid41[7] , \wBMid41[6] , \wBMid41[5] , 
        \wBMid41[4] , \wBMid41[3] , \wBMid41[2] , \wBMid41[1] , \wBMid41[0] }), 
        .HiOut({\wRegInB41[31] , \wRegInB41[30] , \wRegInB41[29] , 
        \wRegInB41[28] , \wRegInB41[27] , \wRegInB41[26] , \wRegInB41[25] , 
        \wRegInB41[24] , \wRegInB41[23] , \wRegInB41[22] , \wRegInB41[21] , 
        \wRegInB41[20] , \wRegInB41[19] , \wRegInB41[18] , \wRegInB41[17] , 
        \wRegInB41[16] , \wRegInB41[15] , \wRegInB41[14] , \wRegInB41[13] , 
        \wRegInB41[12] , \wRegInB41[11] , \wRegInB41[10] , \wRegInB41[9] , 
        \wRegInB41[8] , \wRegInB41[7] , \wRegInB41[6] , \wRegInB41[5] , 
        \wRegInB41[4] , \wRegInB41[3] , \wRegInB41[2] , \wRegInB41[1] , 
        \wRegInB41[0] }), .LoOut({\wRegInA42[31] , \wRegInA42[30] , 
        \wRegInA42[29] , \wRegInA42[28] , \wRegInA42[27] , \wRegInA42[26] , 
        \wRegInA42[25] , \wRegInA42[24] , \wRegInA42[23] , \wRegInA42[22] , 
        \wRegInA42[21] , \wRegInA42[20] , \wRegInA42[19] , \wRegInA42[18] , 
        \wRegInA42[17] , \wRegInA42[16] , \wRegInA42[15] , \wRegInA42[14] , 
        \wRegInA42[13] , \wRegInA42[12] , \wRegInA42[11] , \wRegInA42[10] , 
        \wRegInA42[9] , \wRegInA42[8] , \wRegInA42[7] , \wRegInA42[6] , 
        \wRegInA42[5] , \wRegInA42[4] , \wRegInA42[3] , \wRegInA42[2] , 
        \wRegInA42[1] , \wRegInA42[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_24 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink25[31] , \ScanLink25[30] , \ScanLink25[29] , 
        \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , \ScanLink25[25] , 
        \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , \ScanLink25[21] , 
        \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , \ScanLink25[17] , 
        \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , \ScanLink25[13] , 
        \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , \ScanLink25[9] , 
        \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , \ScanLink25[5] , 
        \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , \ScanLink25[1] , 
        \ScanLink25[0] }), .ScanOut({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB115[31] , \wRegInB115[30] , 
        \wRegInB115[29] , \wRegInB115[28] , \wRegInB115[27] , \wRegInB115[26] , 
        \wRegInB115[25] , \wRegInB115[24] , \wRegInB115[23] , \wRegInB115[22] , 
        \wRegInB115[21] , \wRegInB115[20] , \wRegInB115[19] , \wRegInB115[18] , 
        \wRegInB115[17] , \wRegInB115[16] , \wRegInB115[15] , \wRegInB115[14] , 
        \wRegInB115[13] , \wRegInB115[12] , \wRegInB115[11] , \wRegInB115[10] , 
        \wRegInB115[9] , \wRegInB115[8] , \wRegInB115[7] , \wRegInB115[6] , 
        \wRegInB115[5] , \wRegInB115[4] , \wRegInB115[3] , \wRegInB115[2] , 
        \wRegInB115[1] , \wRegInB115[0] }), .Out({\wBIn115[31] , \wBIn115[30] , 
        \wBIn115[29] , \wBIn115[28] , \wBIn115[27] , \wBIn115[26] , 
        \wBIn115[25] , \wBIn115[24] , \wBIn115[23] , \wBIn115[22] , 
        \wBIn115[21] , \wBIn115[20] , \wBIn115[19] , \wBIn115[18] , 
        \wBIn115[17] , \wBIn115[16] , \wBIn115[15] , \wBIn115[14] , 
        \wBIn115[13] , \wBIn115[12] , \wBIn115[11] , \wBIn115[10] , 
        \wBIn115[9] , \wBIn115[8] , \wBIn115[7] , \wBIn115[6] , \wBIn115[5] , 
        \wBIn115[4] , \wBIn115[3] , \wBIn115[2] , \wBIn115[1] , \wBIn115[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_174 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink175[31] , \ScanLink175[30] , \ScanLink175[29] , 
        \ScanLink175[28] , \ScanLink175[27] , \ScanLink175[26] , 
        \ScanLink175[25] , \ScanLink175[24] , \ScanLink175[23] , 
        \ScanLink175[22] , \ScanLink175[21] , \ScanLink175[20] , 
        \ScanLink175[19] , \ScanLink175[18] , \ScanLink175[17] , 
        \ScanLink175[16] , \ScanLink175[15] , \ScanLink175[14] , 
        \ScanLink175[13] , \ScanLink175[12] , \ScanLink175[11] , 
        \ScanLink175[10] , \ScanLink175[9] , \ScanLink175[8] , 
        \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , \ScanLink175[4] , 
        \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , \ScanLink175[0] 
        }), .ScanOut({\ScanLink174[31] , \ScanLink174[30] , \ScanLink174[29] , 
        \ScanLink174[28] , \ScanLink174[27] , \ScanLink174[26] , 
        \ScanLink174[25] , \ScanLink174[24] , \ScanLink174[23] , 
        \ScanLink174[22] , \ScanLink174[21] , \ScanLink174[20] , 
        \ScanLink174[19] , \ScanLink174[18] , \ScanLink174[17] , 
        \ScanLink174[16] , \ScanLink174[15] , \ScanLink174[14] , 
        \ScanLink174[13] , \ScanLink174[12] , \ScanLink174[11] , 
        \ScanLink174[10] , \ScanLink174[9] , \ScanLink174[8] , 
        \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , \ScanLink174[4] , 
        \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , \ScanLink174[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB40[31] , \wRegInB40[30] , \wRegInB40[29] , 
        \wRegInB40[28] , \wRegInB40[27] , \wRegInB40[26] , \wRegInB40[25] , 
        \wRegInB40[24] , \wRegInB40[23] , \wRegInB40[22] , \wRegInB40[21] , 
        \wRegInB40[20] , \wRegInB40[19] , \wRegInB40[18] , \wRegInB40[17] , 
        \wRegInB40[16] , \wRegInB40[15] , \wRegInB40[14] , \wRegInB40[13] , 
        \wRegInB40[12] , \wRegInB40[11] , \wRegInB40[10] , \wRegInB40[9] , 
        \wRegInB40[8] , \wRegInB40[7] , \wRegInB40[6] , \wRegInB40[5] , 
        \wRegInB40[4] , \wRegInB40[3] , \wRegInB40[2] , \wRegInB40[1] , 
        \wRegInB40[0] }), .Out({\wBIn40[31] , \wBIn40[30] , \wBIn40[29] , 
        \wBIn40[28] , \wBIn40[27] , \wBIn40[26] , \wBIn40[25] , \wBIn40[24] , 
        \wBIn40[23] , \wBIn40[22] , \wBIn40[21] , \wBIn40[20] , \wBIn40[19] , 
        \wBIn40[18] , \wBIn40[17] , \wBIn40[16] , \wBIn40[15] , \wBIn40[14] , 
        \wBIn40[13] , \wBIn40[12] , \wBIn40[11] , \wBIn40[10] , \wBIn40[9] , 
        \wBIn40[8] , \wBIn40[7] , \wBIn40[6] , \wBIn40[5] , \wBIn40[4] , 
        \wBIn40[3] , \wBIn40[2] , \wBIn40[1] , \wBIn40[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid110[31] , \wAMid110[30] , \wAMid110[29] , \wAMid110[28] , 
        \wAMid110[27] , \wAMid110[26] , \wAMid110[25] , \wAMid110[24] , 
        \wAMid110[23] , \wAMid110[22] , \wAMid110[21] , \wAMid110[20] , 
        \wAMid110[19] , \wAMid110[18] , \wAMid110[17] , \wAMid110[16] , 
        \wAMid110[15] , \wAMid110[14] , \wAMid110[13] , \wAMid110[12] , 
        \wAMid110[11] , \wAMid110[10] , \wAMid110[9] , \wAMid110[8] , 
        \wAMid110[7] , \wAMid110[6] , \wAMid110[5] , \wAMid110[4] , 
        \wAMid110[3] , \wAMid110[2] , \wAMid110[1] , \wAMid110[0] }), .BIn({
        \wBMid110[31] , \wBMid110[30] , \wBMid110[29] , \wBMid110[28] , 
        \wBMid110[27] , \wBMid110[26] , \wBMid110[25] , \wBMid110[24] , 
        \wBMid110[23] , \wBMid110[22] , \wBMid110[21] , \wBMid110[20] , 
        \wBMid110[19] , \wBMid110[18] , \wBMid110[17] , \wBMid110[16] , 
        \wBMid110[15] , \wBMid110[14] , \wBMid110[13] , \wBMid110[12] , 
        \wBMid110[11] , \wBMid110[10] , \wBMid110[9] , \wBMid110[8] , 
        \wBMid110[7] , \wBMid110[6] , \wBMid110[5] , \wBMid110[4] , 
        \wBMid110[3] , \wBMid110[2] , \wBMid110[1] , \wBMid110[0] }), .HiOut({
        \wRegInB110[31] , \wRegInB110[30] , \wRegInB110[29] , \wRegInB110[28] , 
        \wRegInB110[27] , \wRegInB110[26] , \wRegInB110[25] , \wRegInB110[24] , 
        \wRegInB110[23] , \wRegInB110[22] , \wRegInB110[21] , \wRegInB110[20] , 
        \wRegInB110[19] , \wRegInB110[18] , \wRegInB110[17] , \wRegInB110[16] , 
        \wRegInB110[15] , \wRegInB110[14] , \wRegInB110[13] , \wRegInB110[12] , 
        \wRegInB110[11] , \wRegInB110[10] , \wRegInB110[9] , \wRegInB110[8] , 
        \wRegInB110[7] , \wRegInB110[6] , \wRegInB110[5] , \wRegInB110[4] , 
        \wRegInB110[3] , \wRegInB110[2] , \wRegInB110[1] , \wRegInB110[0] }), 
        .LoOut({\wRegInA111[31] , \wRegInA111[30] , \wRegInA111[29] , 
        \wRegInA111[28] , \wRegInA111[27] , \wRegInA111[26] , \wRegInA111[25] , 
        \wRegInA111[24] , \wRegInA111[23] , \wRegInA111[22] , \wRegInA111[21] , 
        \wRegInA111[20] , \wRegInA111[19] , \wRegInA111[18] , \wRegInA111[17] , 
        \wRegInA111[16] , \wRegInA111[15] , \wRegInA111[14] , \wRegInA111[13] , 
        \wRegInA111[12] , \wRegInA111[11] , \wRegInA111[10] , \wRegInA111[9] , 
        \wRegInA111[8] , \wRegInA111[7] , \wRegInA111[6] , \wRegInA111[5] , 
        \wRegInA111[4] , \wRegInA111[3] , \wRegInA111[2] , \wRegInA111[1] , 
        \wRegInA111[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_244 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink245[31] , \ScanLink245[30] , \ScanLink245[29] , 
        \ScanLink245[28] , \ScanLink245[27] , \ScanLink245[26] , 
        \ScanLink245[25] , \ScanLink245[24] , \ScanLink245[23] , 
        \ScanLink245[22] , \ScanLink245[21] , \ScanLink245[20] , 
        \ScanLink245[19] , \ScanLink245[18] , \ScanLink245[17] , 
        \ScanLink245[16] , \ScanLink245[15] , \ScanLink245[14] , 
        \ScanLink245[13] , \ScanLink245[12] , \ScanLink245[11] , 
        \ScanLink245[10] , \ScanLink245[9] , \ScanLink245[8] , 
        \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , \ScanLink245[4] , 
        \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , \ScanLink245[0] 
        }), .ScanOut({\ScanLink244[31] , \ScanLink244[30] , \ScanLink244[29] , 
        \ScanLink244[28] , \ScanLink244[27] , \ScanLink244[26] , 
        \ScanLink244[25] , \ScanLink244[24] , \ScanLink244[23] , 
        \ScanLink244[22] , \ScanLink244[21] , \ScanLink244[20] , 
        \ScanLink244[19] , \ScanLink244[18] , \ScanLink244[17] , 
        \ScanLink244[16] , \ScanLink244[15] , \ScanLink244[14] , 
        \ScanLink244[13] , \ScanLink244[12] , \ScanLink244[11] , 
        \ScanLink244[10] , \ScanLink244[9] , \ScanLink244[8] , 
        \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , \ScanLink244[4] , 
        \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , \ScanLink244[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB5[31] , \wRegInB5[30] , \wRegInB5[29] , \wRegInB5[28] , 
        \wRegInB5[27] , \wRegInB5[26] , \wRegInB5[25] , \wRegInB5[24] , 
        \wRegInB5[23] , \wRegInB5[22] , \wRegInB5[21] , \wRegInB5[20] , 
        \wRegInB5[19] , \wRegInB5[18] , \wRegInB5[17] , \wRegInB5[16] , 
        \wRegInB5[15] , \wRegInB5[14] , \wRegInB5[13] , \wRegInB5[12] , 
        \wRegInB5[11] , \wRegInB5[10] , \wRegInB5[9] , \wRegInB5[8] , 
        \wRegInB5[7] , \wRegInB5[6] , \wRegInB5[5] , \wRegInB5[4] , 
        \wRegInB5[3] , \wRegInB5[2] , \wRegInB5[1] , \wRegInB5[0] }), .Out({
        \wBIn5[31] , \wBIn5[30] , \wBIn5[29] , \wBIn5[28] , \wBIn5[27] , 
        \wBIn5[26] , \wBIn5[25] , \wBIn5[24] , \wBIn5[23] , \wBIn5[22] , 
        \wBIn5[21] , \wBIn5[20] , \wBIn5[19] , \wBIn5[18] , \wBIn5[17] , 
        \wBIn5[16] , \wBIn5[15] , \wBIn5[14] , \wBIn5[13] , \wBIn5[12] , 
        \wBIn5[11] , \wBIn5[10] , \wBIn5[9] , \wBIn5[8] , \wBIn5[7] , 
        \wBIn5[6] , \wBIn5[5] , \wBIn5[4] , \wBIn5[3] , \wBIn5[2] , \wBIn5[1] , 
        \wBIn5[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_148 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink149[31] , \ScanLink149[30] , \ScanLink149[29] , 
        \ScanLink149[28] , \ScanLink149[27] , \ScanLink149[26] , 
        \ScanLink149[25] , \ScanLink149[24] , \ScanLink149[23] , 
        \ScanLink149[22] , \ScanLink149[21] , \ScanLink149[20] , 
        \ScanLink149[19] , \ScanLink149[18] , \ScanLink149[17] , 
        \ScanLink149[16] , \ScanLink149[15] , \ScanLink149[14] , 
        \ScanLink149[13] , \ScanLink149[12] , \ScanLink149[11] , 
        \ScanLink149[10] , \ScanLink149[9] , \ScanLink149[8] , 
        \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , \ScanLink149[4] , 
        \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , \ScanLink149[0] 
        }), .ScanOut({\ScanLink148[31] , \ScanLink148[30] , \ScanLink148[29] , 
        \ScanLink148[28] , \ScanLink148[27] , \ScanLink148[26] , 
        \ScanLink148[25] , \ScanLink148[24] , \ScanLink148[23] , 
        \ScanLink148[22] , \ScanLink148[21] , \ScanLink148[20] , 
        \ScanLink148[19] , \ScanLink148[18] , \ScanLink148[17] , 
        \ScanLink148[16] , \ScanLink148[15] , \ScanLink148[14] , 
        \ScanLink148[13] , \ScanLink148[12] , \ScanLink148[11] , 
        \ScanLink148[10] , \ScanLink148[9] , \ScanLink148[8] , 
        \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , \ScanLink148[4] , 
        \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , \ScanLink148[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB53[31] , \wRegInB53[30] , \wRegInB53[29] , 
        \wRegInB53[28] , \wRegInB53[27] , \wRegInB53[26] , \wRegInB53[25] , 
        \wRegInB53[24] , \wRegInB53[23] , \wRegInB53[22] , \wRegInB53[21] , 
        \wRegInB53[20] , \wRegInB53[19] , \wRegInB53[18] , \wRegInB53[17] , 
        \wRegInB53[16] , \wRegInB53[15] , \wRegInB53[14] , \wRegInB53[13] , 
        \wRegInB53[12] , \wRegInB53[11] , \wRegInB53[10] , \wRegInB53[9] , 
        \wRegInB53[8] , \wRegInB53[7] , \wRegInB53[6] , \wRegInB53[5] , 
        \wRegInB53[4] , \wRegInB53[3] , \wRegInB53[2] , \wRegInB53[1] , 
        \wRegInB53[0] }), .Out({\wBIn53[31] , \wBIn53[30] , \wBIn53[29] , 
        \wBIn53[28] , \wBIn53[27] , \wBIn53[26] , \wBIn53[25] , \wBIn53[24] , 
        \wBIn53[23] , \wBIn53[22] , \wBIn53[21] , \wBIn53[20] , \wBIn53[19] , 
        \wBIn53[18] , \wBIn53[17] , \wBIn53[16] , \wBIn53[15] , \wBIn53[14] , 
        \wBIn53[13] , \wBIn53[12] , \wBIn53[11] , \wBIn53[10] , \wBIn53[9] , 
        \wBIn53[8] , \wBIn53[7] , \wBIn53[6] , \wBIn53[5] , \wBIn53[4] , 
        \wBIn53[3] , \wBIn53[2] , \wBIn53[1] , \wBIn53[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_93 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink94[31] , \ScanLink94[30] , \ScanLink94[29] , 
        \ScanLink94[28] , \ScanLink94[27] , \ScanLink94[26] , \ScanLink94[25] , 
        \ScanLink94[24] , \ScanLink94[23] , \ScanLink94[22] , \ScanLink94[21] , 
        \ScanLink94[20] , \ScanLink94[19] , \ScanLink94[18] , \ScanLink94[17] , 
        \ScanLink94[16] , \ScanLink94[15] , \ScanLink94[14] , \ScanLink94[13] , 
        \ScanLink94[12] , \ScanLink94[11] , \ScanLink94[10] , \ScanLink94[9] , 
        \ScanLink94[8] , \ScanLink94[7] , \ScanLink94[6] , \ScanLink94[5] , 
        \ScanLink94[4] , \ScanLink94[3] , \ScanLink94[2] , \ScanLink94[1] , 
        \ScanLink94[0] }), .ScanOut({\ScanLink93[31] , \ScanLink93[30] , 
        \ScanLink93[29] , \ScanLink93[28] , \ScanLink93[27] , \ScanLink93[26] , 
        \ScanLink93[25] , \ScanLink93[24] , \ScanLink93[23] , \ScanLink93[22] , 
        \ScanLink93[21] , \ScanLink93[20] , \ScanLink93[19] , \ScanLink93[18] , 
        \ScanLink93[17] , \ScanLink93[16] , \ScanLink93[15] , \ScanLink93[14] , 
        \ScanLink93[13] , \ScanLink93[12] , \ScanLink93[11] , \ScanLink93[10] , 
        \ScanLink93[9] , \ScanLink93[8] , \ScanLink93[7] , \ScanLink93[6] , 
        \ScanLink93[5] , \ScanLink93[4] , \ScanLink93[3] , \ScanLink93[2] , 
        \ScanLink93[1] , \ScanLink93[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA81[31] , \wRegInA81[30] , 
        \wRegInA81[29] , \wRegInA81[28] , \wRegInA81[27] , \wRegInA81[26] , 
        \wRegInA81[25] , \wRegInA81[24] , \wRegInA81[23] , \wRegInA81[22] , 
        \wRegInA81[21] , \wRegInA81[20] , \wRegInA81[19] , \wRegInA81[18] , 
        \wRegInA81[17] , \wRegInA81[16] , \wRegInA81[15] , \wRegInA81[14] , 
        \wRegInA81[13] , \wRegInA81[12] , \wRegInA81[11] , \wRegInA81[10] , 
        \wRegInA81[9] , \wRegInA81[8] , \wRegInA81[7] , \wRegInA81[6] , 
        \wRegInA81[5] , \wRegInA81[4] , \wRegInA81[3] , \wRegInA81[2] , 
        \wRegInA81[1] , \wRegInA81[0] }), .Out({\wAIn81[31] , \wAIn81[30] , 
        \wAIn81[29] , \wAIn81[28] , \wAIn81[27] , \wAIn81[26] , \wAIn81[25] , 
        \wAIn81[24] , \wAIn81[23] , \wAIn81[22] , \wAIn81[21] , \wAIn81[20] , 
        \wAIn81[19] , \wAIn81[18] , \wAIn81[17] , \wAIn81[16] , \wAIn81[15] , 
        \wAIn81[14] , \wAIn81[13] , \wAIn81[12] , \wAIn81[11] , \wAIn81[10] , 
        \wAIn81[9] , \wAIn81[8] , \wAIn81[7] , \wAIn81[6] , \wAIn81[5] , 
        \wAIn81[4] , \wAIn81[3] , \wAIn81[2] , \wAIn81[1] , \wAIn81[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_18 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink19[31] , \ScanLink19[30] , \ScanLink19[29] , 
        \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , \ScanLink19[25] , 
        \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , \ScanLink19[21] , 
        \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , \ScanLink19[17] , 
        \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , \ScanLink19[13] , 
        \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , \ScanLink19[9] , 
        \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , \ScanLink19[5] , 
        \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , \ScanLink19[1] , 
        \ScanLink19[0] }), .ScanOut({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB118[31] , \wRegInB118[30] , 
        \wRegInB118[29] , \wRegInB118[28] , \wRegInB118[27] , \wRegInB118[26] , 
        \wRegInB118[25] , \wRegInB118[24] , \wRegInB118[23] , \wRegInB118[22] , 
        \wRegInB118[21] , \wRegInB118[20] , \wRegInB118[19] , \wRegInB118[18] , 
        \wRegInB118[17] , \wRegInB118[16] , \wRegInB118[15] , \wRegInB118[14] , 
        \wRegInB118[13] , \wRegInB118[12] , \wRegInB118[11] , \wRegInB118[10] , 
        \wRegInB118[9] , \wRegInB118[8] , \wRegInB118[7] , \wRegInB118[6] , 
        \wRegInB118[5] , \wRegInB118[4] , \wRegInB118[3] , \wRegInB118[2] , 
        \wRegInB118[1] , \wRegInB118[0] }), .Out({\wBIn118[31] , \wBIn118[30] , 
        \wBIn118[29] , \wBIn118[28] , \wBIn118[27] , \wBIn118[26] , 
        \wBIn118[25] , \wBIn118[24] , \wBIn118[23] , \wBIn118[22] , 
        \wBIn118[21] , \wBIn118[20] , \wBIn118[19] , \wBIn118[18] , 
        \wBIn118[17] , \wBIn118[16] , \wBIn118[15] , \wBIn118[14] , 
        \wBIn118[13] , \wBIn118[12] , \wBIn118[11] , \wBIn118[10] , 
        \wBIn118[9] , \wBIn118[8] , \wBIn118[7] , \wBIn118[6] , \wBIn118[5] , 
        \wBIn118[4] , \wBIn118[3] , \wBIn118[2] , \wBIn118[1] , \wBIn118[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn16[31] , \wAIn16[30] , \wAIn16[29] , \wAIn16[28] , \wAIn16[27] , 
        \wAIn16[26] , \wAIn16[25] , \wAIn16[24] , \wAIn16[23] , \wAIn16[22] , 
        \wAIn16[21] , \wAIn16[20] , \wAIn16[19] , \wAIn16[18] , \wAIn16[17] , 
        \wAIn16[16] , \wAIn16[15] , \wAIn16[14] , \wAIn16[13] , \wAIn16[12] , 
        \wAIn16[11] , \wAIn16[10] , \wAIn16[9] , \wAIn16[8] , \wAIn16[7] , 
        \wAIn16[6] , \wAIn16[5] , \wAIn16[4] , \wAIn16[3] , \wAIn16[2] , 
        \wAIn16[1] , \wAIn16[0] }), .BIn({\wBIn16[31] , \wBIn16[30] , 
        \wBIn16[29] , \wBIn16[28] , \wBIn16[27] , \wBIn16[26] , \wBIn16[25] , 
        \wBIn16[24] , \wBIn16[23] , \wBIn16[22] , \wBIn16[21] , \wBIn16[20] , 
        \wBIn16[19] , \wBIn16[18] , \wBIn16[17] , \wBIn16[16] , \wBIn16[15] , 
        \wBIn16[14] , \wBIn16[13] , \wBIn16[12] , \wBIn16[11] , \wBIn16[10] , 
        \wBIn16[9] , \wBIn16[8] , \wBIn16[7] , \wBIn16[6] , \wBIn16[5] , 
        \wBIn16[4] , \wBIn16[3] , \wBIn16[2] , \wBIn16[1] , \wBIn16[0] }), 
        .HiOut({\wBMid15[31] , \wBMid15[30] , \wBMid15[29] , \wBMid15[28] , 
        \wBMid15[27] , \wBMid15[26] , \wBMid15[25] , \wBMid15[24] , 
        \wBMid15[23] , \wBMid15[22] , \wBMid15[21] , \wBMid15[20] , 
        \wBMid15[19] , \wBMid15[18] , \wBMid15[17] , \wBMid15[16] , 
        \wBMid15[15] , \wBMid15[14] , \wBMid15[13] , \wBMid15[12] , 
        \wBMid15[11] , \wBMid15[10] , \wBMid15[9] , \wBMid15[8] , \wBMid15[7] , 
        \wBMid15[6] , \wBMid15[5] , \wBMid15[4] , \wBMid15[3] , \wBMid15[2] , 
        \wBMid15[1] , \wBMid15[0] }), .LoOut({\wAMid16[31] , \wAMid16[30] , 
        \wAMid16[29] , \wAMid16[28] , \wAMid16[27] , \wAMid16[26] , 
        \wAMid16[25] , \wAMid16[24] , \wAMid16[23] , \wAMid16[22] , 
        \wAMid16[21] , \wAMid16[20] , \wAMid16[19] , \wAMid16[18] , 
        \wAMid16[17] , \wAMid16[16] , \wAMid16[15] , \wAMid16[14] , 
        \wAMid16[13] , \wAMid16[12] , \wAMid16[11] , \wAMid16[10] , 
        \wAMid16[9] , \wAMid16[8] , \wAMid16[7] , \wAMid16[6] , \wAMid16[5] , 
        \wAMid16[4] , \wAMid16[3] , \wAMid16[2] , \wAMid16[1] , \wAMid16[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn23[31] , \wAIn23[30] , \wAIn23[29] , \wAIn23[28] , \wAIn23[27] , 
        \wAIn23[26] , \wAIn23[25] , \wAIn23[24] , \wAIn23[23] , \wAIn23[22] , 
        \wAIn23[21] , \wAIn23[20] , \wAIn23[19] , \wAIn23[18] , \wAIn23[17] , 
        \wAIn23[16] , \wAIn23[15] , \wAIn23[14] , \wAIn23[13] , \wAIn23[12] , 
        \wAIn23[11] , \wAIn23[10] , \wAIn23[9] , \wAIn23[8] , \wAIn23[7] , 
        \wAIn23[6] , \wAIn23[5] , \wAIn23[4] , \wAIn23[3] , \wAIn23[2] , 
        \wAIn23[1] , \wAIn23[0] }), .BIn({\wBIn23[31] , \wBIn23[30] , 
        \wBIn23[29] , \wBIn23[28] , \wBIn23[27] , \wBIn23[26] , \wBIn23[25] , 
        \wBIn23[24] , \wBIn23[23] , \wBIn23[22] , \wBIn23[21] , \wBIn23[20] , 
        \wBIn23[19] , \wBIn23[18] , \wBIn23[17] , \wBIn23[16] , \wBIn23[15] , 
        \wBIn23[14] , \wBIn23[13] , \wBIn23[12] , \wBIn23[11] , \wBIn23[10] , 
        \wBIn23[9] , \wBIn23[8] , \wBIn23[7] , \wBIn23[6] , \wBIn23[5] , 
        \wBIn23[4] , \wBIn23[3] , \wBIn23[2] , \wBIn23[1] , \wBIn23[0] }), 
        .HiOut({\wBMid22[31] , \wBMid22[30] , \wBMid22[29] , \wBMid22[28] , 
        \wBMid22[27] , \wBMid22[26] , \wBMid22[25] , \wBMid22[24] , 
        \wBMid22[23] , \wBMid22[22] , \wBMid22[21] , \wBMid22[20] , 
        \wBMid22[19] , \wBMid22[18] , \wBMid22[17] , \wBMid22[16] , 
        \wBMid22[15] , \wBMid22[14] , \wBMid22[13] , \wBMid22[12] , 
        \wBMid22[11] , \wBMid22[10] , \wBMid22[9] , \wBMid22[8] , \wBMid22[7] , 
        \wBMid22[6] , \wBMid22[5] , \wBMid22[4] , \wBMid22[3] , \wBMid22[2] , 
        \wBMid22[1] , \wBMid22[0] }), .LoOut({\wAMid23[31] , \wAMid23[30] , 
        \wAMid23[29] , \wAMid23[28] , \wAMid23[27] , \wAMid23[26] , 
        \wAMid23[25] , \wAMid23[24] , \wAMid23[23] , \wAMid23[22] , 
        \wAMid23[21] , \wAMid23[20] , \wAMid23[19] , \wAMid23[18] , 
        \wAMid23[17] , \wAMid23[16] , \wAMid23[15] , \wAMid23[14] , 
        \wAMid23[13] , \wAMid23[12] , \wAMid23[11] , \wAMid23[10] , 
        \wAMid23[9] , \wAMid23[8] , \wAMid23[7] , \wAMid23[6] , \wAMid23[5] , 
        \wAMid23[4] , \wAMid23[3] , \wAMid23[2] , \wAMid23[1] , \wAMid23[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid13[31] , \wAMid13[30] , \wAMid13[29] , \wAMid13[28] , 
        \wAMid13[27] , \wAMid13[26] , \wAMid13[25] , \wAMid13[24] , 
        \wAMid13[23] , \wAMid13[22] , \wAMid13[21] , \wAMid13[20] , 
        \wAMid13[19] , \wAMid13[18] , \wAMid13[17] , \wAMid13[16] , 
        \wAMid13[15] , \wAMid13[14] , \wAMid13[13] , \wAMid13[12] , 
        \wAMid13[11] , \wAMid13[10] , \wAMid13[9] , \wAMid13[8] , \wAMid13[7] , 
        \wAMid13[6] , \wAMid13[5] , \wAMid13[4] , \wAMid13[3] , \wAMid13[2] , 
        \wAMid13[1] , \wAMid13[0] }), .BIn({\wBMid13[31] , \wBMid13[30] , 
        \wBMid13[29] , \wBMid13[28] , \wBMid13[27] , \wBMid13[26] , 
        \wBMid13[25] , \wBMid13[24] , \wBMid13[23] , \wBMid13[22] , 
        \wBMid13[21] , \wBMid13[20] , \wBMid13[19] , \wBMid13[18] , 
        \wBMid13[17] , \wBMid13[16] , \wBMid13[15] , \wBMid13[14] , 
        \wBMid13[13] , \wBMid13[12] , \wBMid13[11] , \wBMid13[10] , 
        \wBMid13[9] , \wBMid13[8] , \wBMid13[7] , \wBMid13[6] , \wBMid13[5] , 
        \wBMid13[4] , \wBMid13[3] , \wBMid13[2] , \wBMid13[1] , \wBMid13[0] }), 
        .HiOut({\wRegInB13[31] , \wRegInB13[30] , \wRegInB13[29] , 
        \wRegInB13[28] , \wRegInB13[27] , \wRegInB13[26] , \wRegInB13[25] , 
        \wRegInB13[24] , \wRegInB13[23] , \wRegInB13[22] , \wRegInB13[21] , 
        \wRegInB13[20] , \wRegInB13[19] , \wRegInB13[18] , \wRegInB13[17] , 
        \wRegInB13[16] , \wRegInB13[15] , \wRegInB13[14] , \wRegInB13[13] , 
        \wRegInB13[12] , \wRegInB13[11] , \wRegInB13[10] , \wRegInB13[9] , 
        \wRegInB13[8] , \wRegInB13[7] , \wRegInB13[6] , \wRegInB13[5] , 
        \wRegInB13[4] , \wRegInB13[3] , \wRegInB13[2] , \wRegInB13[1] , 
        \wRegInB13[0] }), .LoOut({\wRegInA14[31] , \wRegInA14[30] , 
        \wRegInA14[29] , \wRegInA14[28] , \wRegInA14[27] , \wRegInA14[26] , 
        \wRegInA14[25] , \wRegInA14[24] , \wRegInA14[23] , \wRegInA14[22] , 
        \wRegInA14[21] , \wRegInA14[20] , \wRegInA14[19] , \wRegInA14[18] , 
        \wRegInA14[17] , \wRegInA14[16] , \wRegInA14[15] , \wRegInA14[14] , 
        \wRegInA14[13] , \wRegInA14[12] , \wRegInA14[11] , \wRegInA14[10] , 
        \wRegInA14[9] , \wRegInA14[8] , \wRegInA14[7] , \wRegInA14[6] , 
        \wRegInA14[5] , \wRegInA14[4] , \wRegInA14[3] , \wRegInA14[2] , 
        \wRegInA14[1] , \wRegInA14[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid98[31] , \wAMid98[30] , \wAMid98[29] , \wAMid98[28] , 
        \wAMid98[27] , \wAMid98[26] , \wAMid98[25] , \wAMid98[24] , 
        \wAMid98[23] , \wAMid98[22] , \wAMid98[21] , \wAMid98[20] , 
        \wAMid98[19] , \wAMid98[18] , \wAMid98[17] , \wAMid98[16] , 
        \wAMid98[15] , \wAMid98[14] , \wAMid98[13] , \wAMid98[12] , 
        \wAMid98[11] , \wAMid98[10] , \wAMid98[9] , \wAMid98[8] , \wAMid98[7] , 
        \wAMid98[6] , \wAMid98[5] , \wAMid98[4] , \wAMid98[3] , \wAMid98[2] , 
        \wAMid98[1] , \wAMid98[0] }), .BIn({\wBMid98[31] , \wBMid98[30] , 
        \wBMid98[29] , \wBMid98[28] , \wBMid98[27] , \wBMid98[26] , 
        \wBMid98[25] , \wBMid98[24] , \wBMid98[23] , \wBMid98[22] , 
        \wBMid98[21] , \wBMid98[20] , \wBMid98[19] , \wBMid98[18] , 
        \wBMid98[17] , \wBMid98[16] , \wBMid98[15] , \wBMid98[14] , 
        \wBMid98[13] , \wBMid98[12] , \wBMid98[11] , \wBMid98[10] , 
        \wBMid98[9] , \wBMid98[8] , \wBMid98[7] , \wBMid98[6] , \wBMid98[5] , 
        \wBMid98[4] , \wBMid98[3] , \wBMid98[2] , \wBMid98[1] , \wBMid98[0] }), 
        .HiOut({\wRegInB98[31] , \wRegInB98[30] , \wRegInB98[29] , 
        \wRegInB98[28] , \wRegInB98[27] , \wRegInB98[26] , \wRegInB98[25] , 
        \wRegInB98[24] , \wRegInB98[23] , \wRegInB98[22] , \wRegInB98[21] , 
        \wRegInB98[20] , \wRegInB98[19] , \wRegInB98[18] , \wRegInB98[17] , 
        \wRegInB98[16] , \wRegInB98[15] , \wRegInB98[14] , \wRegInB98[13] , 
        \wRegInB98[12] , \wRegInB98[11] , \wRegInB98[10] , \wRegInB98[9] , 
        \wRegInB98[8] , \wRegInB98[7] , \wRegInB98[6] , \wRegInB98[5] , 
        \wRegInB98[4] , \wRegInB98[3] , \wRegInB98[2] , \wRegInB98[1] , 
        \wRegInB98[0] }), .LoOut({\wRegInA99[31] , \wRegInA99[30] , 
        \wRegInA99[29] , \wRegInA99[28] , \wRegInA99[27] , \wRegInA99[26] , 
        \wRegInA99[25] , \wRegInA99[24] , \wRegInA99[23] , \wRegInA99[22] , 
        \wRegInA99[21] , \wRegInA99[20] , \wRegInA99[19] , \wRegInA99[18] , 
        \wRegInA99[17] , \wRegInA99[16] , \wRegInA99[15] , \wRegInA99[14] , 
        \wRegInA99[13] , \wRegInA99[12] , \wRegInA99[11] , \wRegInA99[10] , 
        \wRegInA99[9] , \wRegInA99[8] , \wRegInA99[7] , \wRegInA99[6] , 
        \wRegInA99[5] , \wRegInA99[4] , \wRegInA99[3] , \wRegInA99[2] , 
        \wRegInA99[1] , \wRegInA99[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_126 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink127[31] , \ScanLink127[30] , \ScanLink127[29] , 
        \ScanLink127[28] , \ScanLink127[27] , \ScanLink127[26] , 
        \ScanLink127[25] , \ScanLink127[24] , \ScanLink127[23] , 
        \ScanLink127[22] , \ScanLink127[21] , \ScanLink127[20] , 
        \ScanLink127[19] , \ScanLink127[18] , \ScanLink127[17] , 
        \ScanLink127[16] , \ScanLink127[15] , \ScanLink127[14] , 
        \ScanLink127[13] , \ScanLink127[12] , \ScanLink127[11] , 
        \ScanLink127[10] , \ScanLink127[9] , \ScanLink127[8] , 
        \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , \ScanLink127[4] , 
        \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , \ScanLink127[0] 
        }), .ScanOut({\ScanLink126[31] , \ScanLink126[30] , \ScanLink126[29] , 
        \ScanLink126[28] , \ScanLink126[27] , \ScanLink126[26] , 
        \ScanLink126[25] , \ScanLink126[24] , \ScanLink126[23] , 
        \ScanLink126[22] , \ScanLink126[21] , \ScanLink126[20] , 
        \ScanLink126[19] , \ScanLink126[18] , \ScanLink126[17] , 
        \ScanLink126[16] , \ScanLink126[15] , \ScanLink126[14] , 
        \ScanLink126[13] , \ScanLink126[12] , \ScanLink126[11] , 
        \ScanLink126[10] , \ScanLink126[9] , \ScanLink126[8] , 
        \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , \ScanLink126[4] , 
        \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , \ScanLink126[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB64[31] , \wRegInB64[30] , \wRegInB64[29] , 
        \wRegInB64[28] , \wRegInB64[27] , \wRegInB64[26] , \wRegInB64[25] , 
        \wRegInB64[24] , \wRegInB64[23] , \wRegInB64[22] , \wRegInB64[21] , 
        \wRegInB64[20] , \wRegInB64[19] , \wRegInB64[18] , \wRegInB64[17] , 
        \wRegInB64[16] , \wRegInB64[15] , \wRegInB64[14] , \wRegInB64[13] , 
        \wRegInB64[12] , \wRegInB64[11] , \wRegInB64[10] , \wRegInB64[9] , 
        \wRegInB64[8] , \wRegInB64[7] , \wRegInB64[6] , \wRegInB64[5] , 
        \wRegInB64[4] , \wRegInB64[3] , \wRegInB64[2] , \wRegInB64[1] , 
        \wRegInB64[0] }), .Out({\wBIn64[31] , \wBIn64[30] , \wBIn64[29] , 
        \wBIn64[28] , \wBIn64[27] , \wBIn64[26] , \wBIn64[25] , \wBIn64[24] , 
        \wBIn64[23] , \wBIn64[22] , \wBIn64[21] , \wBIn64[20] , \wBIn64[19] , 
        \wBIn64[18] , \wBIn64[17] , \wBIn64[16] , \wBIn64[15] , \wBIn64[14] , 
        \wBIn64[13] , \wBIn64[12] , \wBIn64[11] , \wBIn64[10] , \wBIn64[9] , 
        \wBIn64[8] , \wBIn64[7] , \wBIn64[6] , \wBIn64[5] , \wBIn64[4] , 
        \wBIn64[3] , \wBIn64[2] , \wBIn64[1] , \wBIn64[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_76 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink77[31] , \ScanLink77[30] , \ScanLink77[29] , 
        \ScanLink77[28] , \ScanLink77[27] , \ScanLink77[26] , \ScanLink77[25] , 
        \ScanLink77[24] , \ScanLink77[23] , \ScanLink77[22] , \ScanLink77[21] , 
        \ScanLink77[20] , \ScanLink77[19] , \ScanLink77[18] , \ScanLink77[17] , 
        \ScanLink77[16] , \ScanLink77[15] , \ScanLink77[14] , \ScanLink77[13] , 
        \ScanLink77[12] , \ScanLink77[11] , \ScanLink77[10] , \ScanLink77[9] , 
        \ScanLink77[8] , \ScanLink77[7] , \ScanLink77[6] , \ScanLink77[5] , 
        \ScanLink77[4] , \ScanLink77[3] , \ScanLink77[2] , \ScanLink77[1] , 
        \ScanLink77[0] }), .ScanOut({\ScanLink76[31] , \ScanLink76[30] , 
        \ScanLink76[29] , \ScanLink76[28] , \ScanLink76[27] , \ScanLink76[26] , 
        \ScanLink76[25] , \ScanLink76[24] , \ScanLink76[23] , \ScanLink76[22] , 
        \ScanLink76[21] , \ScanLink76[20] , \ScanLink76[19] , \ScanLink76[18] , 
        \ScanLink76[17] , \ScanLink76[16] , \ScanLink76[15] , \ScanLink76[14] , 
        \ScanLink76[13] , \ScanLink76[12] , \ScanLink76[11] , \ScanLink76[10] , 
        \ScanLink76[9] , \ScanLink76[8] , \ScanLink76[7] , \ScanLink76[6] , 
        \ScanLink76[5] , \ScanLink76[4] , \ScanLink76[3] , \ScanLink76[2] , 
        \ScanLink76[1] , \ScanLink76[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB89[31] , \wRegInB89[30] , 
        \wRegInB89[29] , \wRegInB89[28] , \wRegInB89[27] , \wRegInB89[26] , 
        \wRegInB89[25] , \wRegInB89[24] , \wRegInB89[23] , \wRegInB89[22] , 
        \wRegInB89[21] , \wRegInB89[20] , \wRegInB89[19] , \wRegInB89[18] , 
        \wRegInB89[17] , \wRegInB89[16] , \wRegInB89[15] , \wRegInB89[14] , 
        \wRegInB89[13] , \wRegInB89[12] , \wRegInB89[11] , \wRegInB89[10] , 
        \wRegInB89[9] , \wRegInB89[8] , \wRegInB89[7] , \wRegInB89[6] , 
        \wRegInB89[5] , \wRegInB89[4] , \wRegInB89[3] , \wRegInB89[2] , 
        \wRegInB89[1] , \wRegInB89[0] }), .Out({\wBIn89[31] , \wBIn89[30] , 
        \wBIn89[29] , \wBIn89[28] , \wBIn89[27] , \wBIn89[26] , \wBIn89[25] , 
        \wBIn89[24] , \wBIn89[23] , \wBIn89[22] , \wBIn89[21] , \wBIn89[20] , 
        \wBIn89[19] , \wBIn89[18] , \wBIn89[17] , \wBIn89[16] , \wBIn89[15] , 
        \wBIn89[14] , \wBIn89[13] , \wBIn89[12] , \wBIn89[11] , \wBIn89[10] , 
        \wBIn89[9] , \wBIn89[8] , \wBIn89[7] , \wBIn89[6] , \wBIn89[5] , 
        \wBIn89[4] , \wBIn89[3] , \wBIn89[2] , \wBIn89[1] , \wBIn89[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn31[31] , \wAIn31[30] , \wAIn31[29] , \wAIn31[28] , \wAIn31[27] , 
        \wAIn31[26] , \wAIn31[25] , \wAIn31[24] , \wAIn31[23] , \wAIn31[22] , 
        \wAIn31[21] , \wAIn31[20] , \wAIn31[19] , \wAIn31[18] , \wAIn31[17] , 
        \wAIn31[16] , \wAIn31[15] , \wAIn31[14] , \wAIn31[13] , \wAIn31[12] , 
        \wAIn31[11] , \wAIn31[10] , \wAIn31[9] , \wAIn31[8] , \wAIn31[7] , 
        \wAIn31[6] , \wAIn31[5] , \wAIn31[4] , \wAIn31[3] , \wAIn31[2] , 
        \wAIn31[1] , \wAIn31[0] }), .BIn({\wBIn31[31] , \wBIn31[30] , 
        \wBIn31[29] , \wBIn31[28] , \wBIn31[27] , \wBIn31[26] , \wBIn31[25] , 
        \wBIn31[24] , \wBIn31[23] , \wBIn31[22] , \wBIn31[21] , \wBIn31[20] , 
        \wBIn31[19] , \wBIn31[18] , \wBIn31[17] , \wBIn31[16] , \wBIn31[15] , 
        \wBIn31[14] , \wBIn31[13] , \wBIn31[12] , \wBIn31[11] , \wBIn31[10] , 
        \wBIn31[9] , \wBIn31[8] , \wBIn31[7] , \wBIn31[6] , \wBIn31[5] , 
        \wBIn31[4] , \wBIn31[3] , \wBIn31[2] , \wBIn31[1] , \wBIn31[0] }), 
        .HiOut({\wBMid30[31] , \wBMid30[30] , \wBMid30[29] , \wBMid30[28] , 
        \wBMid30[27] , \wBMid30[26] , \wBMid30[25] , \wBMid30[24] , 
        \wBMid30[23] , \wBMid30[22] , \wBMid30[21] , \wBMid30[20] , 
        \wBMid30[19] , \wBMid30[18] , \wBMid30[17] , \wBMid30[16] , 
        \wBMid30[15] , \wBMid30[14] , \wBMid30[13] , \wBMid30[12] , 
        \wBMid30[11] , \wBMid30[10] , \wBMid30[9] , \wBMid30[8] , \wBMid30[7] , 
        \wBMid30[6] , \wBMid30[5] , \wBMid30[4] , \wBMid30[3] , \wBMid30[2] , 
        \wBMid30[1] , \wBMid30[0] }), .LoOut({\wAMid31[31] , \wAMid31[30] , 
        \wAMid31[29] , \wAMid31[28] , \wAMid31[27] , \wAMid31[26] , 
        \wAMid31[25] , \wAMid31[24] , \wAMid31[23] , \wAMid31[22] , 
        \wAMid31[21] , \wAMid31[20] , \wAMid31[19] , \wAMid31[18] , 
        \wAMid31[17] , \wAMid31[16] , \wAMid31[15] , \wAMid31[14] , 
        \wAMid31[13] , \wAMid31[12] , \wAMid31[11] , \wAMid31[10] , 
        \wAMid31[9] , \wAMid31[8] , \wAMid31[7] , \wAMid31[6] , \wAMid31[5] , 
        \wAMid31[4] , \wAMid31[3] , \wAMid31[2] , \wAMid31[1] , \wAMid31[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid34[31] , \wAMid34[30] , \wAMid34[29] , \wAMid34[28] , 
        \wAMid34[27] , \wAMid34[26] , \wAMid34[25] , \wAMid34[24] , 
        \wAMid34[23] , \wAMid34[22] , \wAMid34[21] , \wAMid34[20] , 
        \wAMid34[19] , \wAMid34[18] , \wAMid34[17] , \wAMid34[16] , 
        \wAMid34[15] , \wAMid34[14] , \wAMid34[13] , \wAMid34[12] , 
        \wAMid34[11] , \wAMid34[10] , \wAMid34[9] , \wAMid34[8] , \wAMid34[7] , 
        \wAMid34[6] , \wAMid34[5] , \wAMid34[4] , \wAMid34[3] , \wAMid34[2] , 
        \wAMid34[1] , \wAMid34[0] }), .BIn({\wBMid34[31] , \wBMid34[30] , 
        \wBMid34[29] , \wBMid34[28] , \wBMid34[27] , \wBMid34[26] , 
        \wBMid34[25] , \wBMid34[24] , \wBMid34[23] , \wBMid34[22] , 
        \wBMid34[21] , \wBMid34[20] , \wBMid34[19] , \wBMid34[18] , 
        \wBMid34[17] , \wBMid34[16] , \wBMid34[15] , \wBMid34[14] , 
        \wBMid34[13] , \wBMid34[12] , \wBMid34[11] , \wBMid34[10] , 
        \wBMid34[9] , \wBMid34[8] , \wBMid34[7] , \wBMid34[6] , \wBMid34[5] , 
        \wBMid34[4] , \wBMid34[3] , \wBMid34[2] , \wBMid34[1] , \wBMid34[0] }), 
        .HiOut({\wRegInB34[31] , \wRegInB34[30] , \wRegInB34[29] , 
        \wRegInB34[28] , \wRegInB34[27] , \wRegInB34[26] , \wRegInB34[25] , 
        \wRegInB34[24] , \wRegInB34[23] , \wRegInB34[22] , \wRegInB34[21] , 
        \wRegInB34[20] , \wRegInB34[19] , \wRegInB34[18] , \wRegInB34[17] , 
        \wRegInB34[16] , \wRegInB34[15] , \wRegInB34[14] , \wRegInB34[13] , 
        \wRegInB34[12] , \wRegInB34[11] , \wRegInB34[10] , \wRegInB34[9] , 
        \wRegInB34[8] , \wRegInB34[7] , \wRegInB34[6] , \wRegInB34[5] , 
        \wRegInB34[4] , \wRegInB34[3] , \wRegInB34[2] , \wRegInB34[1] , 
        \wRegInB34[0] }), .LoOut({\wRegInA35[31] , \wRegInA35[30] , 
        \wRegInA35[29] , \wRegInA35[28] , \wRegInA35[27] , \wRegInA35[26] , 
        \wRegInA35[25] , \wRegInA35[24] , \wRegInA35[23] , \wRegInA35[22] , 
        \wRegInA35[21] , \wRegInA35[20] , \wRegInA35[19] , \wRegInA35[18] , 
        \wRegInA35[17] , \wRegInA35[16] , \wRegInA35[15] , \wRegInA35[14] , 
        \wRegInA35[13] , \wRegInA35[12] , \wRegInA35[11] , \wRegInA35[10] , 
        \wRegInA35[9] , \wRegInA35[8] , \wRegInA35[7] , \wRegInA35[6] , 
        \wRegInA35[5] , \wRegInA35[4] , \wRegInA35[3] , \wRegInA35[2] , 
        \wRegInA35[1] , \wRegInA35[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_231 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink232[31] , \ScanLink232[30] , \ScanLink232[29] , 
        \ScanLink232[28] , \ScanLink232[27] , \ScanLink232[26] , 
        \ScanLink232[25] , \ScanLink232[24] , \ScanLink232[23] , 
        \ScanLink232[22] , \ScanLink232[21] , \ScanLink232[20] , 
        \ScanLink232[19] , \ScanLink232[18] , \ScanLink232[17] , 
        \ScanLink232[16] , \ScanLink232[15] , \ScanLink232[14] , 
        \ScanLink232[13] , \ScanLink232[12] , \ScanLink232[11] , 
        \ScanLink232[10] , \ScanLink232[9] , \ScanLink232[8] , 
        \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , \ScanLink232[4] , 
        \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , \ScanLink232[0] 
        }), .ScanOut({\ScanLink231[31] , \ScanLink231[30] , \ScanLink231[29] , 
        \ScanLink231[28] , \ScanLink231[27] , \ScanLink231[26] , 
        \ScanLink231[25] , \ScanLink231[24] , \ScanLink231[23] , 
        \ScanLink231[22] , \ScanLink231[21] , \ScanLink231[20] , 
        \ScanLink231[19] , \ScanLink231[18] , \ScanLink231[17] , 
        \ScanLink231[16] , \ScanLink231[15] , \ScanLink231[14] , 
        \ScanLink231[13] , \ScanLink231[12] , \ScanLink231[11] , 
        \ScanLink231[10] , \ScanLink231[9] , \ScanLink231[8] , 
        \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , \ScanLink231[4] , 
        \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , \ScanLink231[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA12[31] , \wRegInA12[30] , \wRegInA12[29] , 
        \wRegInA12[28] , \wRegInA12[27] , \wRegInA12[26] , \wRegInA12[25] , 
        \wRegInA12[24] , \wRegInA12[23] , \wRegInA12[22] , \wRegInA12[21] , 
        \wRegInA12[20] , \wRegInA12[19] , \wRegInA12[18] , \wRegInA12[17] , 
        \wRegInA12[16] , \wRegInA12[15] , \wRegInA12[14] , \wRegInA12[13] , 
        \wRegInA12[12] , \wRegInA12[11] , \wRegInA12[10] , \wRegInA12[9] , 
        \wRegInA12[8] , \wRegInA12[7] , \wRegInA12[6] , \wRegInA12[5] , 
        \wRegInA12[4] , \wRegInA12[3] , \wRegInA12[2] , \wRegInA12[1] , 
        \wRegInA12[0] }), .Out({\wAIn12[31] , \wAIn12[30] , \wAIn12[29] , 
        \wAIn12[28] , \wAIn12[27] , \wAIn12[26] , \wAIn12[25] , \wAIn12[24] , 
        \wAIn12[23] , \wAIn12[22] , \wAIn12[21] , \wAIn12[20] , \wAIn12[19] , 
        \wAIn12[18] , \wAIn12[17] , \wAIn12[16] , \wAIn12[15] , \wAIn12[14] , 
        \wAIn12[13] , \wAIn12[12] , \wAIn12[11] , \wAIn12[10] , \wAIn12[9] , 
        \wAIn12[8] , \wAIn12[7] , \wAIn12[6] , \wAIn12[5] , \wAIn12[4] , 
        \wAIn12[3] , \wAIn12[2] , \wAIn12[1] , \wAIn12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_216 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink217[31] , \ScanLink217[30] , \ScanLink217[29] , 
        \ScanLink217[28] , \ScanLink217[27] , \ScanLink217[26] , 
        \ScanLink217[25] , \ScanLink217[24] , \ScanLink217[23] , 
        \ScanLink217[22] , \ScanLink217[21] , \ScanLink217[20] , 
        \ScanLink217[19] , \ScanLink217[18] , \ScanLink217[17] , 
        \ScanLink217[16] , \ScanLink217[15] , \ScanLink217[14] , 
        \ScanLink217[13] , \ScanLink217[12] , \ScanLink217[11] , 
        \ScanLink217[10] , \ScanLink217[9] , \ScanLink217[8] , 
        \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , \ScanLink217[4] , 
        \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , \ScanLink217[0] 
        }), .ScanOut({\ScanLink216[31] , \ScanLink216[30] , \ScanLink216[29] , 
        \ScanLink216[28] , \ScanLink216[27] , \ScanLink216[26] , 
        \ScanLink216[25] , \ScanLink216[24] , \ScanLink216[23] , 
        \ScanLink216[22] , \ScanLink216[21] , \ScanLink216[20] , 
        \ScanLink216[19] , \ScanLink216[18] , \ScanLink216[17] , 
        \ScanLink216[16] , \ScanLink216[15] , \ScanLink216[14] , 
        \ScanLink216[13] , \ScanLink216[12] , \ScanLink216[11] , 
        \ScanLink216[10] , \ScanLink216[9] , \ScanLink216[8] , 
        \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , \ScanLink216[4] , 
        \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , \ScanLink216[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB19[31] , \wRegInB19[30] , \wRegInB19[29] , 
        \wRegInB19[28] , \wRegInB19[27] , \wRegInB19[26] , \wRegInB19[25] , 
        \wRegInB19[24] , \wRegInB19[23] , \wRegInB19[22] , \wRegInB19[21] , 
        \wRegInB19[20] , \wRegInB19[19] , \wRegInB19[18] , \wRegInB19[17] , 
        \wRegInB19[16] , \wRegInB19[15] , \wRegInB19[14] , \wRegInB19[13] , 
        \wRegInB19[12] , \wRegInB19[11] , \wRegInB19[10] , \wRegInB19[9] , 
        \wRegInB19[8] , \wRegInB19[7] , \wRegInB19[6] , \wRegInB19[5] , 
        \wRegInB19[4] , \wRegInB19[3] , \wRegInB19[2] , \wRegInB19[1] , 
        \wRegInB19[0] }), .Out({\wBIn19[31] , \wBIn19[30] , \wBIn19[29] , 
        \wBIn19[28] , \wBIn19[27] , \wBIn19[26] , \wBIn19[25] , \wBIn19[24] , 
        \wBIn19[23] , \wBIn19[22] , \wBIn19[21] , \wBIn19[20] , \wBIn19[19] , 
        \wBIn19[18] , \wBIn19[17] , \wBIn19[16] , \wBIn19[15] , \wBIn19[14] , 
        \wBIn19[13] , \wBIn19[12] , \wBIn19[11] , \wBIn19[10] , \wBIn19[9] , 
        \wBIn19[8] , \wBIn19[7] , \wBIn19[6] , \wBIn19[5] , \wBIn19[4] , 
        \wBIn19[3] , \wBIn19[2] , \wBIn19[1] , \wBIn19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_51 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink52[31] , \ScanLink52[30] , \ScanLink52[29] , 
        \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , \ScanLink52[25] , 
        \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , \ScanLink52[21] , 
        \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , \ScanLink52[17] , 
        \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , \ScanLink52[13] , 
        \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , \ScanLink52[9] , 
        \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , \ScanLink52[5] , 
        \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , \ScanLink52[1] , 
        \ScanLink52[0] }), .ScanOut({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA102[31] , \wRegInA102[30] , 
        \wRegInA102[29] , \wRegInA102[28] , \wRegInA102[27] , \wRegInA102[26] , 
        \wRegInA102[25] , \wRegInA102[24] , \wRegInA102[23] , \wRegInA102[22] , 
        \wRegInA102[21] , \wRegInA102[20] , \wRegInA102[19] , \wRegInA102[18] , 
        \wRegInA102[17] , \wRegInA102[16] , \wRegInA102[15] , \wRegInA102[14] , 
        \wRegInA102[13] , \wRegInA102[12] , \wRegInA102[11] , \wRegInA102[10] , 
        \wRegInA102[9] , \wRegInA102[8] , \wRegInA102[7] , \wRegInA102[6] , 
        \wRegInA102[5] , \wRegInA102[4] , \wRegInA102[3] , \wRegInA102[2] , 
        \wRegInA102[1] , \wRegInA102[0] }), .Out({\wAIn102[31] , \wAIn102[30] , 
        \wAIn102[29] , \wAIn102[28] , \wAIn102[27] , \wAIn102[26] , 
        \wAIn102[25] , \wAIn102[24] , \wAIn102[23] , \wAIn102[22] , 
        \wAIn102[21] , \wAIn102[20] , \wAIn102[19] , \wAIn102[18] , 
        \wAIn102[17] , \wAIn102[16] , \wAIn102[15] , \wAIn102[14] , 
        \wAIn102[13] , \wAIn102[12] , \wAIn102[11] , \wAIn102[10] , 
        \wAIn102[9] , \wAIn102[8] , \wAIn102[7] , \wAIn102[6] , \wAIn102[5] , 
        \wAIn102[4] , \wAIn102[3] , \wAIn102[2] , \wAIn102[1] , \wAIn102[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_134 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink135[31] , \ScanLink135[30] , \ScanLink135[29] , 
        \ScanLink135[28] , \ScanLink135[27] , \ScanLink135[26] , 
        \ScanLink135[25] , \ScanLink135[24] , \ScanLink135[23] , 
        \ScanLink135[22] , \ScanLink135[21] , \ScanLink135[20] , 
        \ScanLink135[19] , \ScanLink135[18] , \ScanLink135[17] , 
        \ScanLink135[16] , \ScanLink135[15] , \ScanLink135[14] , 
        \ScanLink135[13] , \ScanLink135[12] , \ScanLink135[11] , 
        \ScanLink135[10] , \ScanLink135[9] , \ScanLink135[8] , 
        \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , \ScanLink135[4] , 
        \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , \ScanLink135[0] 
        }), .ScanOut({\ScanLink134[31] , \ScanLink134[30] , \ScanLink134[29] , 
        \ScanLink134[28] , \ScanLink134[27] , \ScanLink134[26] , 
        \ScanLink134[25] , \ScanLink134[24] , \ScanLink134[23] , 
        \ScanLink134[22] , \ScanLink134[21] , \ScanLink134[20] , 
        \ScanLink134[19] , \ScanLink134[18] , \ScanLink134[17] , 
        \ScanLink134[16] , \ScanLink134[15] , \ScanLink134[14] , 
        \ScanLink134[13] , \ScanLink134[12] , \ScanLink134[11] , 
        \ScanLink134[10] , \ScanLink134[9] , \ScanLink134[8] , 
        \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , \ScanLink134[4] , 
        \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , \ScanLink134[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB60[31] , \wRegInB60[30] , \wRegInB60[29] , 
        \wRegInB60[28] , \wRegInB60[27] , \wRegInB60[26] , \wRegInB60[25] , 
        \wRegInB60[24] , \wRegInB60[23] , \wRegInB60[22] , \wRegInB60[21] , 
        \wRegInB60[20] , \wRegInB60[19] , \wRegInB60[18] , \wRegInB60[17] , 
        \wRegInB60[16] , \wRegInB60[15] , \wRegInB60[14] , \wRegInB60[13] , 
        \wRegInB60[12] , \wRegInB60[11] , \wRegInB60[10] , \wRegInB60[9] , 
        \wRegInB60[8] , \wRegInB60[7] , \wRegInB60[6] , \wRegInB60[5] , 
        \wRegInB60[4] , \wRegInB60[3] , \wRegInB60[2] , \wRegInB60[1] , 
        \wRegInB60[0] }), .Out({\wBIn60[31] , \wBIn60[30] , \wBIn60[29] , 
        \wBIn60[28] , \wBIn60[27] , \wBIn60[26] , \wBIn60[25] , \wBIn60[24] , 
        \wBIn60[23] , \wBIn60[22] , \wBIn60[21] , \wBIn60[20] , \wBIn60[19] , 
        \wBIn60[18] , \wBIn60[17] , \wBIn60[16] , \wBIn60[15] , \wBIn60[14] , 
        \wBIn60[13] , \wBIn60[12] , \wBIn60[11] , \wBIn60[10] , \wBIn60[9] , 
        \wBIn60[8] , \wBIn60[7] , \wBIn60[6] , \wBIn60[5] , \wBIn60[4] , 
        \wBIn60[3] , \wBIn60[2] , \wBIn60[1] , \wBIn60[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_101 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink102[31] , \ScanLink102[30] , \ScanLink102[29] , 
        \ScanLink102[28] , \ScanLink102[27] , \ScanLink102[26] , 
        \ScanLink102[25] , \ScanLink102[24] , \ScanLink102[23] , 
        \ScanLink102[22] , \ScanLink102[21] , \ScanLink102[20] , 
        \ScanLink102[19] , \ScanLink102[18] , \ScanLink102[17] , 
        \ScanLink102[16] , \ScanLink102[15] , \ScanLink102[14] , 
        \ScanLink102[13] , \ScanLink102[12] , \ScanLink102[11] , 
        \ScanLink102[10] , \ScanLink102[9] , \ScanLink102[8] , 
        \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , \ScanLink102[4] , 
        \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , \ScanLink102[0] 
        }), .ScanOut({\ScanLink101[31] , \ScanLink101[30] , \ScanLink101[29] , 
        \ScanLink101[28] , \ScanLink101[27] , \ScanLink101[26] , 
        \ScanLink101[25] , \ScanLink101[24] , \ScanLink101[23] , 
        \ScanLink101[22] , \ScanLink101[21] , \ScanLink101[20] , 
        \ScanLink101[19] , \ScanLink101[18] , \ScanLink101[17] , 
        \ScanLink101[16] , \ScanLink101[15] , \ScanLink101[14] , 
        \ScanLink101[13] , \ScanLink101[12] , \ScanLink101[11] , 
        \ScanLink101[10] , \ScanLink101[9] , \ScanLink101[8] , 
        \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , \ScanLink101[4] , 
        \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , \ScanLink101[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA77[31] , \wRegInA77[30] , \wRegInA77[29] , 
        \wRegInA77[28] , \wRegInA77[27] , \wRegInA77[26] , \wRegInA77[25] , 
        \wRegInA77[24] , \wRegInA77[23] , \wRegInA77[22] , \wRegInA77[21] , 
        \wRegInA77[20] , \wRegInA77[19] , \wRegInA77[18] , \wRegInA77[17] , 
        \wRegInA77[16] , \wRegInA77[15] , \wRegInA77[14] , \wRegInA77[13] , 
        \wRegInA77[12] , \wRegInA77[11] , \wRegInA77[10] , \wRegInA77[9] , 
        \wRegInA77[8] , \wRegInA77[7] , \wRegInA77[6] , \wRegInA77[5] , 
        \wRegInA77[4] , \wRegInA77[3] , \wRegInA77[2] , \wRegInA77[1] , 
        \wRegInA77[0] }), .Out({\wAIn77[31] , \wAIn77[30] , \wAIn77[29] , 
        \wAIn77[28] , \wAIn77[27] , \wAIn77[26] , \wAIn77[25] , \wAIn77[24] , 
        \wAIn77[23] , \wAIn77[22] , \wAIn77[21] , \wAIn77[20] , \wAIn77[19] , 
        \wAIn77[18] , \wAIn77[17] , \wAIn77[16] , \wAIn77[15] , \wAIn77[14] , 
        \wAIn77[13] , \wAIn77[12] , \wAIn77[11] , \wAIn77[10] , \wAIn77[9] , 
        \wAIn77[8] , \wAIn77[7] , \wAIn77[6] , \wAIn77[5] , \wAIn77[4] , 
        \wAIn77[3] , \wAIn77[2] , \wAIn77[1] , \wAIn77[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_64 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink65[31] , \ScanLink65[30] , \ScanLink65[29] , 
        \ScanLink65[28] , \ScanLink65[27] , \ScanLink65[26] , \ScanLink65[25] , 
        \ScanLink65[24] , \ScanLink65[23] , \ScanLink65[22] , \ScanLink65[21] , 
        \ScanLink65[20] , \ScanLink65[19] , \ScanLink65[18] , \ScanLink65[17] , 
        \ScanLink65[16] , \ScanLink65[15] , \ScanLink65[14] , \ScanLink65[13] , 
        \ScanLink65[12] , \ScanLink65[11] , \ScanLink65[10] , \ScanLink65[9] , 
        \ScanLink65[8] , \ScanLink65[7] , \ScanLink65[6] , \ScanLink65[5] , 
        \ScanLink65[4] , \ScanLink65[3] , \ScanLink65[2] , \ScanLink65[1] , 
        \ScanLink65[0] }), .ScanOut({\ScanLink64[31] , \ScanLink64[30] , 
        \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , 
        \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , 
        \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , 
        \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , 
        \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , 
        \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , 
        \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , 
        \ScanLink64[1] , \ScanLink64[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB95[31] , \wRegInB95[30] , 
        \wRegInB95[29] , \wRegInB95[28] , \wRegInB95[27] , \wRegInB95[26] , 
        \wRegInB95[25] , \wRegInB95[24] , \wRegInB95[23] , \wRegInB95[22] , 
        \wRegInB95[21] , \wRegInB95[20] , \wRegInB95[19] , \wRegInB95[18] , 
        \wRegInB95[17] , \wRegInB95[16] , \wRegInB95[15] , \wRegInB95[14] , 
        \wRegInB95[13] , \wRegInB95[12] , \wRegInB95[11] , \wRegInB95[10] , 
        \wRegInB95[9] , \wRegInB95[8] , \wRegInB95[7] , \wRegInB95[6] , 
        \wRegInB95[5] , \wRegInB95[4] , \wRegInB95[3] , \wRegInB95[2] , 
        \wRegInB95[1] , \wRegInB95[0] }), .Out({\wBIn95[31] , \wBIn95[30] , 
        \wBIn95[29] , \wBIn95[28] , \wBIn95[27] , \wBIn95[26] , \wBIn95[25] , 
        \wBIn95[24] , \wBIn95[23] , \wBIn95[22] , \wBIn95[21] , \wBIn95[20] , 
        \wBIn95[19] , \wBIn95[18] , \wBIn95[17] , \wBIn95[16] , \wBIn95[15] , 
        \wBIn95[14] , \wBIn95[13] , \wBIn95[12] , \wBIn95[11] , \wBIn95[10] , 
        \wBIn95[9] , \wBIn95[8] , \wBIn95[7] , \wBIn95[6] , \wBIn95[5] , 
        \wBIn95[4] , \wBIn95[3] , \wBIn95[2] , \wBIn95[1] , \wBIn95[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid26[31] , \wAMid26[30] , \wAMid26[29] , \wAMid26[28] , 
        \wAMid26[27] , \wAMid26[26] , \wAMid26[25] , \wAMid26[24] , 
        \wAMid26[23] , \wAMid26[22] , \wAMid26[21] , \wAMid26[20] , 
        \wAMid26[19] , \wAMid26[18] , \wAMid26[17] , \wAMid26[16] , 
        \wAMid26[15] , \wAMid26[14] , \wAMid26[13] , \wAMid26[12] , 
        \wAMid26[11] , \wAMid26[10] , \wAMid26[9] , \wAMid26[8] , \wAMid26[7] , 
        \wAMid26[6] , \wAMid26[5] , \wAMid26[4] , \wAMid26[3] , \wAMid26[2] , 
        \wAMid26[1] , \wAMid26[0] }), .BIn({\wBMid26[31] , \wBMid26[30] , 
        \wBMid26[29] , \wBMid26[28] , \wBMid26[27] , \wBMid26[26] , 
        \wBMid26[25] , \wBMid26[24] , \wBMid26[23] , \wBMid26[22] , 
        \wBMid26[21] , \wBMid26[20] , \wBMid26[19] , \wBMid26[18] , 
        \wBMid26[17] , \wBMid26[16] , \wBMid26[15] , \wBMid26[14] , 
        \wBMid26[13] , \wBMid26[12] , \wBMid26[11] , \wBMid26[10] , 
        \wBMid26[9] , \wBMid26[8] , \wBMid26[7] , \wBMid26[6] , \wBMid26[5] , 
        \wBMid26[4] , \wBMid26[3] , \wBMid26[2] , \wBMid26[1] , \wBMid26[0] }), 
        .HiOut({\wRegInB26[31] , \wRegInB26[30] , \wRegInB26[29] , 
        \wRegInB26[28] , \wRegInB26[27] , \wRegInB26[26] , \wRegInB26[25] , 
        \wRegInB26[24] , \wRegInB26[23] , \wRegInB26[22] , \wRegInB26[21] , 
        \wRegInB26[20] , \wRegInB26[19] , \wRegInB26[18] , \wRegInB26[17] , 
        \wRegInB26[16] , \wRegInB26[15] , \wRegInB26[14] , \wRegInB26[13] , 
        \wRegInB26[12] , \wRegInB26[11] , \wRegInB26[10] , \wRegInB26[9] , 
        \wRegInB26[8] , \wRegInB26[7] , \wRegInB26[6] , \wRegInB26[5] , 
        \wRegInB26[4] , \wRegInB26[3] , \wRegInB26[2] , \wRegInB26[1] , 
        \wRegInB26[0] }), .LoOut({\wRegInA27[31] , \wRegInA27[30] , 
        \wRegInA27[29] , \wRegInA27[28] , \wRegInA27[27] , \wRegInA27[26] , 
        \wRegInA27[25] , \wRegInA27[24] , \wRegInA27[23] , \wRegInA27[22] , 
        \wRegInA27[21] , \wRegInA27[20] , \wRegInA27[19] , \wRegInA27[18] , 
        \wRegInA27[17] , \wRegInA27[16] , \wRegInA27[15] , \wRegInA27[14] , 
        \wRegInA27[13] , \wRegInA27[12] , \wRegInA27[11] , \wRegInA27[10] , 
        \wRegInA27[9] , \wRegInA27[8] , \wRegInA27[7] , \wRegInA27[6] , 
        \wRegInA27[5] , \wRegInA27[4] , \wRegInA27[3] , \wRegInA27[2] , 
        \wRegInA27[1] , \wRegInA27[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_223 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink224[31] , \ScanLink224[30] , \ScanLink224[29] , 
        \ScanLink224[28] , \ScanLink224[27] , \ScanLink224[26] , 
        \ScanLink224[25] , \ScanLink224[24] , \ScanLink224[23] , 
        \ScanLink224[22] , \ScanLink224[21] , \ScanLink224[20] , 
        \ScanLink224[19] , \ScanLink224[18] , \ScanLink224[17] , 
        \ScanLink224[16] , \ScanLink224[15] , \ScanLink224[14] , 
        \ScanLink224[13] , \ScanLink224[12] , \ScanLink224[11] , 
        \ScanLink224[10] , \ScanLink224[9] , \ScanLink224[8] , 
        \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , \ScanLink224[4] , 
        \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , \ScanLink224[0] 
        }), .ScanOut({\ScanLink223[31] , \ScanLink223[30] , \ScanLink223[29] , 
        \ScanLink223[28] , \ScanLink223[27] , \ScanLink223[26] , 
        \ScanLink223[25] , \ScanLink223[24] , \ScanLink223[23] , 
        \ScanLink223[22] , \ScanLink223[21] , \ScanLink223[20] , 
        \ScanLink223[19] , \ScanLink223[18] , \ScanLink223[17] , 
        \ScanLink223[16] , \ScanLink223[15] , \ScanLink223[14] , 
        \ScanLink223[13] , \ScanLink223[12] , \ScanLink223[11] , 
        \ScanLink223[10] , \ScanLink223[9] , \ScanLink223[8] , 
        \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , \ScanLink223[4] , 
        \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , \ScanLink223[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA16[31] , \wRegInA16[30] , \wRegInA16[29] , 
        \wRegInA16[28] , \wRegInA16[27] , \wRegInA16[26] , \wRegInA16[25] , 
        \wRegInA16[24] , \wRegInA16[23] , \wRegInA16[22] , \wRegInA16[21] , 
        \wRegInA16[20] , \wRegInA16[19] , \wRegInA16[18] , \wRegInA16[17] , 
        \wRegInA16[16] , \wRegInA16[15] , \wRegInA16[14] , \wRegInA16[13] , 
        \wRegInA16[12] , \wRegInA16[11] , \wRegInA16[10] , \wRegInA16[9] , 
        \wRegInA16[8] , \wRegInA16[7] , \wRegInA16[6] , \wRegInA16[5] , 
        \wRegInA16[4] , \wRegInA16[3] , \wRegInA16[2] , \wRegInA16[1] , 
        \wRegInA16[0] }), .Out({\wAIn16[31] , \wAIn16[30] , \wAIn16[29] , 
        \wAIn16[28] , \wAIn16[27] , \wAIn16[26] , \wAIn16[25] , \wAIn16[24] , 
        \wAIn16[23] , \wAIn16[22] , \wAIn16[21] , \wAIn16[20] , \wAIn16[19] , 
        \wAIn16[18] , \wAIn16[17] , \wAIn16[16] , \wAIn16[15] , \wAIn16[14] , 
        \wAIn16[13] , \wAIn16[12] , \wAIn16[11] , \wAIn16[10] , \wAIn16[9] , 
        \wAIn16[8] , \wAIn16[7] , \wAIn16[6] , \wAIn16[5] , \wAIn16[4] , 
        \wAIn16[3] , \wAIn16[2] , \wAIn16[1] , \wAIn16[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_204 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink205[31] , \ScanLink205[30] , \ScanLink205[29] , 
        \ScanLink205[28] , \ScanLink205[27] , \ScanLink205[26] , 
        \ScanLink205[25] , \ScanLink205[24] , \ScanLink205[23] , 
        \ScanLink205[22] , \ScanLink205[21] , \ScanLink205[20] , 
        \ScanLink205[19] , \ScanLink205[18] , \ScanLink205[17] , 
        \ScanLink205[16] , \ScanLink205[15] , \ScanLink205[14] , 
        \ScanLink205[13] , \ScanLink205[12] , \ScanLink205[11] , 
        \ScanLink205[10] , \ScanLink205[9] , \ScanLink205[8] , 
        \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , \ScanLink205[4] , 
        \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , \ScanLink205[0] 
        }), .ScanOut({\ScanLink204[31] , \ScanLink204[30] , \ScanLink204[29] , 
        \ScanLink204[28] , \ScanLink204[27] , \ScanLink204[26] , 
        \ScanLink204[25] , \ScanLink204[24] , \ScanLink204[23] , 
        \ScanLink204[22] , \ScanLink204[21] , \ScanLink204[20] , 
        \ScanLink204[19] , \ScanLink204[18] , \ScanLink204[17] , 
        \ScanLink204[16] , \ScanLink204[15] , \ScanLink204[14] , 
        \ScanLink204[13] , \ScanLink204[12] , \ScanLink204[11] , 
        \ScanLink204[10] , \ScanLink204[9] , \ScanLink204[8] , 
        \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , \ScanLink204[4] , 
        \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , \ScanLink204[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB25[31] , \wRegInB25[30] , \wRegInB25[29] , 
        \wRegInB25[28] , \wRegInB25[27] , \wRegInB25[26] , \wRegInB25[25] , 
        \wRegInB25[24] , \wRegInB25[23] , \wRegInB25[22] , \wRegInB25[21] , 
        \wRegInB25[20] , \wRegInB25[19] , \wRegInB25[18] , \wRegInB25[17] , 
        \wRegInB25[16] , \wRegInB25[15] , \wRegInB25[14] , \wRegInB25[13] , 
        \wRegInB25[12] , \wRegInB25[11] , \wRegInB25[10] , \wRegInB25[9] , 
        \wRegInB25[8] , \wRegInB25[7] , \wRegInB25[6] , \wRegInB25[5] , 
        \wRegInB25[4] , \wRegInB25[3] , \wRegInB25[2] , \wRegInB25[1] , 
        \wRegInB25[0] }), .Out({\wBIn25[31] , \wBIn25[30] , \wBIn25[29] , 
        \wBIn25[28] , \wBIn25[27] , \wBIn25[26] , \wBIn25[25] , \wBIn25[24] , 
        \wBIn25[23] , \wBIn25[22] , \wBIn25[21] , \wBIn25[20] , \wBIn25[19] , 
        \wBIn25[18] , \wBIn25[17] , \wBIn25[16] , \wBIn25[15] , \wBIn25[14] , 
        \wBIn25[13] , \wBIn25[12] , \wBIn25[11] , \wBIn25[10] , \wBIn25[9] , 
        \wBIn25[8] , \wBIn25[7] , \wBIn25[6] , \wBIn25[5] , \wBIn25[4] , 
        \wBIn25[3] , \wBIn25[2] , \wBIn25[1] , \wBIn25[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_0 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB127[31] , \wRegInB127[30] , 
        \wRegInB127[29] , \wRegInB127[28] , \wRegInB127[27] , \wRegInB127[26] , 
        \wRegInB127[25] , \wRegInB127[24] , \wRegInB127[23] , \wRegInB127[22] , 
        \wRegInB127[21] , \wRegInB127[20] , \wRegInB127[19] , \wRegInB127[18] , 
        \wRegInB127[17] , \wRegInB127[16] , \wRegInB127[15] , \wRegInB127[14] , 
        \wRegInB127[13] , \wRegInB127[12] , \wRegInB127[11] , \wRegInB127[10] , 
        \wRegInB127[9] , \wRegInB127[8] , \wRegInB127[7] , \wRegInB127[6] , 
        \wRegInB127[5] , \wRegInB127[4] , \wRegInB127[3] , \wRegInB127[2] , 
        \wRegInB127[1] , \wRegInB127[0] }), .Out({\wBIn127[31] , \wBIn127[30] , 
        \wBIn127[29] , \wBIn127[28] , \wBIn127[27] , \wBIn127[26] , 
        \wBIn127[25] , \wBIn127[24] , \wBIn127[23] , \wBIn127[22] , 
        \wBIn127[21] , \wBIn127[20] , \wBIn127[19] , \wBIn127[18] , 
        \wBIn127[17] , \wBIn127[16] , \wBIn127[15] , \wBIn127[14] , 
        \wBIn127[13] , \wBIn127[12] , \wBIn127[11] , \wBIn127[10] , 
        \wBIn127[9] , \wBIn127[8] , \wBIn127[7] , \wBIn127[6] , \wBIn127[5] , 
        \wBIn127[4] , \wBIn127[3] , \wBIn127[2] , \wBIn127[1] , \wBIn127[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_113 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink114[31] , \ScanLink114[30] , \ScanLink114[29] , 
        \ScanLink114[28] , \ScanLink114[27] , \ScanLink114[26] , 
        \ScanLink114[25] , \ScanLink114[24] , \ScanLink114[23] , 
        \ScanLink114[22] , \ScanLink114[21] , \ScanLink114[20] , 
        \ScanLink114[19] , \ScanLink114[18] , \ScanLink114[17] , 
        \ScanLink114[16] , \ScanLink114[15] , \ScanLink114[14] , 
        \ScanLink114[13] , \ScanLink114[12] , \ScanLink114[11] , 
        \ScanLink114[10] , \ScanLink114[9] , \ScanLink114[8] , 
        \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , \ScanLink114[4] , 
        \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , \ScanLink114[0] 
        }), .ScanOut({\ScanLink113[31] , \ScanLink113[30] , \ScanLink113[29] , 
        \ScanLink113[28] , \ScanLink113[27] , \ScanLink113[26] , 
        \ScanLink113[25] , \ScanLink113[24] , \ScanLink113[23] , 
        \ScanLink113[22] , \ScanLink113[21] , \ScanLink113[20] , 
        \ScanLink113[19] , \ScanLink113[18] , \ScanLink113[17] , 
        \ScanLink113[16] , \ScanLink113[15] , \ScanLink113[14] , 
        \ScanLink113[13] , \ScanLink113[12] , \ScanLink113[11] , 
        \ScanLink113[10] , \ScanLink113[9] , \ScanLink113[8] , 
        \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , \ScanLink113[4] , 
        \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , \ScanLink113[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA71[31] , \wRegInA71[30] , \wRegInA71[29] , 
        \wRegInA71[28] , \wRegInA71[27] , \wRegInA71[26] , \wRegInA71[25] , 
        \wRegInA71[24] , \wRegInA71[23] , \wRegInA71[22] , \wRegInA71[21] , 
        \wRegInA71[20] , \wRegInA71[19] , \wRegInA71[18] , \wRegInA71[17] , 
        \wRegInA71[16] , \wRegInA71[15] , \wRegInA71[14] , \wRegInA71[13] , 
        \wRegInA71[12] , \wRegInA71[11] , \wRegInA71[10] , \wRegInA71[9] , 
        \wRegInA71[8] , \wRegInA71[7] , \wRegInA71[6] , \wRegInA71[5] , 
        \wRegInA71[4] , \wRegInA71[3] , \wRegInA71[2] , \wRegInA71[1] , 
        \wRegInA71[0] }), .Out({\wAIn71[31] , \wAIn71[30] , \wAIn71[29] , 
        \wAIn71[28] , \wAIn71[27] , \wAIn71[26] , \wAIn71[25] , \wAIn71[24] , 
        \wAIn71[23] , \wAIn71[22] , \wAIn71[21] , \wAIn71[20] , \wAIn71[19] , 
        \wAIn71[18] , \wAIn71[17] , \wAIn71[16] , \wAIn71[15] , \wAIn71[14] , 
        \wAIn71[13] , \wAIn71[12] , \wAIn71[11] , \wAIn71[10] , \wAIn71[9] , 
        \wAIn71[8] , \wAIn71[7] , \wAIn71[6] , \wAIn71[5] , \wAIn71[4] , 
        \wAIn71[3] , \wAIn71[2] , \wAIn71[1] , \wAIn71[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_43 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink44[31] , \ScanLink44[30] , \ScanLink44[29] , 
        \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , \ScanLink44[25] , 
        \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , \ScanLink44[21] , 
        \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , \ScanLink44[17] , 
        \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , \ScanLink44[13] , 
        \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , \ScanLink44[9] , 
        \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , \ScanLink44[5] , 
        \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , \ScanLink44[1] , 
        \ScanLink44[0] }), .ScanOut({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA106[31] , \wRegInA106[30] , 
        \wRegInA106[29] , \wRegInA106[28] , \wRegInA106[27] , \wRegInA106[26] , 
        \wRegInA106[25] , \wRegInA106[24] , \wRegInA106[23] , \wRegInA106[22] , 
        \wRegInA106[21] , \wRegInA106[20] , \wRegInA106[19] , \wRegInA106[18] , 
        \wRegInA106[17] , \wRegInA106[16] , \wRegInA106[15] , \wRegInA106[14] , 
        \wRegInA106[13] , \wRegInA106[12] , \wRegInA106[11] , \wRegInA106[10] , 
        \wRegInA106[9] , \wRegInA106[8] , \wRegInA106[7] , \wRegInA106[6] , 
        \wRegInA106[5] , \wRegInA106[4] , \wRegInA106[3] , \wRegInA106[2] , 
        \wRegInA106[1] , \wRegInA106[0] }), .Out({\wAIn106[31] , \wAIn106[30] , 
        \wAIn106[29] , \wAIn106[28] , \wAIn106[27] , \wAIn106[26] , 
        \wAIn106[25] , \wAIn106[24] , \wAIn106[23] , \wAIn106[22] , 
        \wAIn106[21] , \wAIn106[20] , \wAIn106[19] , \wAIn106[18] , 
        \wAIn106[17] , \wAIn106[16] , \wAIn106[15] , \wAIn106[14] , 
        \wAIn106[13] , \wAIn106[12] , \wAIn106[11] , \wAIn106[10] , 
        \wAIn106[9] , \wAIn106[8] , \wAIn106[7] , \wAIn106[6] , \wAIn106[5] , 
        \wAIn106[4] , \wAIn106[3] , \wAIn106[2] , \wAIn106[1] , \wAIn106[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn44[31] , \wAIn44[30] , \wAIn44[29] , \wAIn44[28] , \wAIn44[27] , 
        \wAIn44[26] , \wAIn44[25] , \wAIn44[24] , \wAIn44[23] , \wAIn44[22] , 
        \wAIn44[21] , \wAIn44[20] , \wAIn44[19] , \wAIn44[18] , \wAIn44[17] , 
        \wAIn44[16] , \wAIn44[15] , \wAIn44[14] , \wAIn44[13] , \wAIn44[12] , 
        \wAIn44[11] , \wAIn44[10] , \wAIn44[9] , \wAIn44[8] , \wAIn44[7] , 
        \wAIn44[6] , \wAIn44[5] , \wAIn44[4] , \wAIn44[3] , \wAIn44[2] , 
        \wAIn44[1] , \wAIn44[0] }), .BIn({\wBIn44[31] , \wBIn44[30] , 
        \wBIn44[29] , \wBIn44[28] , \wBIn44[27] , \wBIn44[26] , \wBIn44[25] , 
        \wBIn44[24] , \wBIn44[23] , \wBIn44[22] , \wBIn44[21] , \wBIn44[20] , 
        \wBIn44[19] , \wBIn44[18] , \wBIn44[17] , \wBIn44[16] , \wBIn44[15] , 
        \wBIn44[14] , \wBIn44[13] , \wBIn44[12] , \wBIn44[11] , \wBIn44[10] , 
        \wBIn44[9] , \wBIn44[8] , \wBIn44[7] , \wBIn44[6] , \wBIn44[5] , 
        \wBIn44[4] , \wBIn44[3] , \wBIn44[2] , \wBIn44[1] , \wBIn44[0] }), 
        .HiOut({\wBMid43[31] , \wBMid43[30] , \wBMid43[29] , \wBMid43[28] , 
        \wBMid43[27] , \wBMid43[26] , \wBMid43[25] , \wBMid43[24] , 
        \wBMid43[23] , \wBMid43[22] , \wBMid43[21] , \wBMid43[20] , 
        \wBMid43[19] , \wBMid43[18] , \wBMid43[17] , \wBMid43[16] , 
        \wBMid43[15] , \wBMid43[14] , \wBMid43[13] , \wBMid43[12] , 
        \wBMid43[11] , \wBMid43[10] , \wBMid43[9] , \wBMid43[8] , \wBMid43[7] , 
        \wBMid43[6] , \wBMid43[5] , \wBMid43[4] , \wBMid43[3] , \wBMid43[2] , 
        \wBMid43[1] , \wBMid43[0] }), .LoOut({\wAMid44[31] , \wAMid44[30] , 
        \wAMid44[29] , \wAMid44[28] , \wAMid44[27] , \wAMid44[26] , 
        \wAMid44[25] , \wAMid44[24] , \wAMid44[23] , \wAMid44[22] , 
        \wAMid44[21] , \wAMid44[20] , \wAMid44[19] , \wAMid44[18] , 
        \wAMid44[17] , \wAMid44[16] , \wAMid44[15] , \wAMid44[14] , 
        \wAMid44[13] , \wAMid44[12] , \wAMid44[11] , \wAMid44[10] , 
        \wAMid44[9] , \wAMid44[8] , \wAMid44[7] , \wAMid44[6] , \wAMid44[5] , 
        \wAMid44[4] , \wAMid44[3] , \wAMid44[2] , \wAMid44[1] , \wAMid44[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn78[31] , \wAIn78[30] , \wAIn78[29] , \wAIn78[28] , \wAIn78[27] , 
        \wAIn78[26] , \wAIn78[25] , \wAIn78[24] , \wAIn78[23] , \wAIn78[22] , 
        \wAIn78[21] , \wAIn78[20] , \wAIn78[19] , \wAIn78[18] , \wAIn78[17] , 
        \wAIn78[16] , \wAIn78[15] , \wAIn78[14] , \wAIn78[13] , \wAIn78[12] , 
        \wAIn78[11] , \wAIn78[10] , \wAIn78[9] , \wAIn78[8] , \wAIn78[7] , 
        \wAIn78[6] , \wAIn78[5] , \wAIn78[4] , \wAIn78[3] , \wAIn78[2] , 
        \wAIn78[1] , \wAIn78[0] }), .BIn({\wBIn78[31] , \wBIn78[30] , 
        \wBIn78[29] , \wBIn78[28] , \wBIn78[27] , \wBIn78[26] , \wBIn78[25] , 
        \wBIn78[24] , \wBIn78[23] , \wBIn78[22] , \wBIn78[21] , \wBIn78[20] , 
        \wBIn78[19] , \wBIn78[18] , \wBIn78[17] , \wBIn78[16] , \wBIn78[15] , 
        \wBIn78[14] , \wBIn78[13] , \wBIn78[12] , \wBIn78[11] , \wBIn78[10] , 
        \wBIn78[9] , \wBIn78[8] , \wBIn78[7] , \wBIn78[6] , \wBIn78[5] , 
        \wBIn78[4] , \wBIn78[3] , \wBIn78[2] , \wBIn78[1] , \wBIn78[0] }), 
        .HiOut({\wBMid77[31] , \wBMid77[30] , \wBMid77[29] , \wBMid77[28] , 
        \wBMid77[27] , \wBMid77[26] , \wBMid77[25] , \wBMid77[24] , 
        \wBMid77[23] , \wBMid77[22] , \wBMid77[21] , \wBMid77[20] , 
        \wBMid77[19] , \wBMid77[18] , \wBMid77[17] , \wBMid77[16] , 
        \wBMid77[15] , \wBMid77[14] , \wBMid77[13] , \wBMid77[12] , 
        \wBMid77[11] , \wBMid77[10] , \wBMid77[9] , \wBMid77[8] , \wBMid77[7] , 
        \wBMid77[6] , \wBMid77[5] , \wBMid77[4] , \wBMid77[3] , \wBMid77[2] , 
        \wBMid77[1] , \wBMid77[0] }), .LoOut({\wAMid78[31] , \wAMid78[30] , 
        \wAMid78[29] , \wAMid78[28] , \wAMid78[27] , \wAMid78[26] , 
        \wAMid78[25] , \wAMid78[24] , \wAMid78[23] , \wAMid78[22] , 
        \wAMid78[21] , \wAMid78[20] , \wAMid78[19] , \wAMid78[18] , 
        \wAMid78[17] , \wAMid78[16] , \wAMid78[15] , \wAMid78[14] , 
        \wAMid78[13] , \wAMid78[12] , \wAMid78[11] , \wAMid78[10] , 
        \wAMid78[9] , \wAMid78[8] , \wAMid78[7] , \wAMid78[6] , \wAMid78[5] , 
        \wAMid78[4] , \wAMid78[3] , \wAMid78[2] , \wAMid78[1] , \wAMid78[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn108[31] , \wAIn108[30] , \wAIn108[29] , \wAIn108[28] , 
        \wAIn108[27] , \wAIn108[26] , \wAIn108[25] , \wAIn108[24] , 
        \wAIn108[23] , \wAIn108[22] , \wAIn108[21] , \wAIn108[20] , 
        \wAIn108[19] , \wAIn108[18] , \wAIn108[17] , \wAIn108[16] , 
        \wAIn108[15] , \wAIn108[14] , \wAIn108[13] , \wAIn108[12] , 
        \wAIn108[11] , \wAIn108[10] , \wAIn108[9] , \wAIn108[8] , \wAIn108[7] , 
        \wAIn108[6] , \wAIn108[5] , \wAIn108[4] , \wAIn108[3] , \wAIn108[2] , 
        \wAIn108[1] , \wAIn108[0] }), .BIn({\wBIn108[31] , \wBIn108[30] , 
        \wBIn108[29] , \wBIn108[28] , \wBIn108[27] , \wBIn108[26] , 
        \wBIn108[25] , \wBIn108[24] , \wBIn108[23] , \wBIn108[22] , 
        \wBIn108[21] , \wBIn108[20] , \wBIn108[19] , \wBIn108[18] , 
        \wBIn108[17] , \wBIn108[16] , \wBIn108[15] , \wBIn108[14] , 
        \wBIn108[13] , \wBIn108[12] , \wBIn108[11] , \wBIn108[10] , 
        \wBIn108[9] , \wBIn108[8] , \wBIn108[7] , \wBIn108[6] , \wBIn108[5] , 
        \wBIn108[4] , \wBIn108[3] , \wBIn108[2] , \wBIn108[1] , \wBIn108[0] }), 
        .HiOut({\wBMid107[31] , \wBMid107[30] , \wBMid107[29] , \wBMid107[28] , 
        \wBMid107[27] , \wBMid107[26] , \wBMid107[25] , \wBMid107[24] , 
        \wBMid107[23] , \wBMid107[22] , \wBMid107[21] , \wBMid107[20] , 
        \wBMid107[19] , \wBMid107[18] , \wBMid107[17] , \wBMid107[16] , 
        \wBMid107[15] , \wBMid107[14] , \wBMid107[13] , \wBMid107[12] , 
        \wBMid107[11] , \wBMid107[10] , \wBMid107[9] , \wBMid107[8] , 
        \wBMid107[7] , \wBMid107[6] , \wBMid107[5] , \wBMid107[4] , 
        \wBMid107[3] , \wBMid107[2] , \wBMid107[1] , \wBMid107[0] }), .LoOut({
        \wAMid108[31] , \wAMid108[30] , \wAMid108[29] , \wAMid108[28] , 
        \wAMid108[27] , \wAMid108[26] , \wAMid108[25] , \wAMid108[24] , 
        \wAMid108[23] , \wAMid108[22] , \wAMid108[21] , \wAMid108[20] , 
        \wAMid108[19] , \wAMid108[18] , \wAMid108[17] , \wAMid108[16] , 
        \wAMid108[15] , \wAMid108[14] , \wAMid108[13] , \wAMid108[12] , 
        \wAMid108[11] , \wAMid108[10] , \wAMid108[9] , \wAMid108[8] , 
        \wAMid108[7] , \wAMid108[6] , \wAMid108[5] , \wAMid108[4] , 
        \wAMid108[3] , \wAMid108[2] , \wAMid108[1] , \wAMid108[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid102[31] , \wAMid102[30] , \wAMid102[29] , \wAMid102[28] , 
        \wAMid102[27] , \wAMid102[26] , \wAMid102[25] , \wAMid102[24] , 
        \wAMid102[23] , \wAMid102[22] , \wAMid102[21] , \wAMid102[20] , 
        \wAMid102[19] , \wAMid102[18] , \wAMid102[17] , \wAMid102[16] , 
        \wAMid102[15] , \wAMid102[14] , \wAMid102[13] , \wAMid102[12] , 
        \wAMid102[11] , \wAMid102[10] , \wAMid102[9] , \wAMid102[8] , 
        \wAMid102[7] , \wAMid102[6] , \wAMid102[5] , \wAMid102[4] , 
        \wAMid102[3] , \wAMid102[2] , \wAMid102[1] , \wAMid102[0] }), .BIn({
        \wBMid102[31] , \wBMid102[30] , \wBMid102[29] , \wBMid102[28] , 
        \wBMid102[27] , \wBMid102[26] , \wBMid102[25] , \wBMid102[24] , 
        \wBMid102[23] , \wBMid102[22] , \wBMid102[21] , \wBMid102[20] , 
        \wBMid102[19] , \wBMid102[18] , \wBMid102[17] , \wBMid102[16] , 
        \wBMid102[15] , \wBMid102[14] , \wBMid102[13] , \wBMid102[12] , 
        \wBMid102[11] , \wBMid102[10] , \wBMid102[9] , \wBMid102[8] , 
        \wBMid102[7] , \wBMid102[6] , \wBMid102[5] , \wBMid102[4] , 
        \wBMid102[3] , \wBMid102[2] , \wBMid102[1] , \wBMid102[0] }), .HiOut({
        \wRegInB102[31] , \wRegInB102[30] , \wRegInB102[29] , \wRegInB102[28] , 
        \wRegInB102[27] , \wRegInB102[26] , \wRegInB102[25] , \wRegInB102[24] , 
        \wRegInB102[23] , \wRegInB102[22] , \wRegInB102[21] , \wRegInB102[20] , 
        \wRegInB102[19] , \wRegInB102[18] , \wRegInB102[17] , \wRegInB102[16] , 
        \wRegInB102[15] , \wRegInB102[14] , \wRegInB102[13] , \wRegInB102[12] , 
        \wRegInB102[11] , \wRegInB102[10] , \wRegInB102[9] , \wRegInB102[8] , 
        \wRegInB102[7] , \wRegInB102[6] , \wRegInB102[5] , \wRegInB102[4] , 
        \wRegInB102[3] , \wRegInB102[2] , \wRegInB102[1] , \wRegInB102[0] }), 
        .LoOut({\wRegInA103[31] , \wRegInA103[30] , \wRegInA103[29] , 
        \wRegInA103[28] , \wRegInA103[27] , \wRegInA103[26] , \wRegInA103[25] , 
        \wRegInA103[24] , \wRegInA103[23] , \wRegInA103[22] , \wRegInA103[21] , 
        \wRegInA103[20] , \wRegInA103[19] , \wRegInA103[18] , \wRegInA103[17] , 
        \wRegInA103[16] , \wRegInA103[15] , \wRegInA103[14] , \wRegInA103[13] , 
        \wRegInA103[12] , \wRegInA103[11] , \wRegInA103[10] , \wRegInA103[9] , 
        \wRegInA103[8] , \wRegInA103[7] , \wRegInA103[6] , \wRegInA103[5] , 
        \wRegInA103[4] , \wRegInA103[3] , \wRegInA103[2] , \wRegInA103[1] , 
        \wRegInA103[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid125[31] , \wAMid125[30] , \wAMid125[29] , \wAMid125[28] , 
        \wAMid125[27] , \wAMid125[26] , \wAMid125[25] , \wAMid125[24] , 
        \wAMid125[23] , \wAMid125[22] , \wAMid125[21] , \wAMid125[20] , 
        \wAMid125[19] , \wAMid125[18] , \wAMid125[17] , \wAMid125[16] , 
        \wAMid125[15] , \wAMid125[14] , \wAMid125[13] , \wAMid125[12] , 
        \wAMid125[11] , \wAMid125[10] , \wAMid125[9] , \wAMid125[8] , 
        \wAMid125[7] , \wAMid125[6] , \wAMid125[5] , \wAMid125[4] , 
        \wAMid125[3] , \wAMid125[2] , \wAMid125[1] , \wAMid125[0] }), .BIn({
        \wBMid125[31] , \wBMid125[30] , \wBMid125[29] , \wBMid125[28] , 
        \wBMid125[27] , \wBMid125[26] , \wBMid125[25] , \wBMid125[24] , 
        \wBMid125[23] , \wBMid125[22] , \wBMid125[21] , \wBMid125[20] , 
        \wBMid125[19] , \wBMid125[18] , \wBMid125[17] , \wBMid125[16] , 
        \wBMid125[15] , \wBMid125[14] , \wBMid125[13] , \wBMid125[12] , 
        \wBMid125[11] , \wBMid125[10] , \wBMid125[9] , \wBMid125[8] , 
        \wBMid125[7] , \wBMid125[6] , \wBMid125[5] , \wBMid125[4] , 
        \wBMid125[3] , \wBMid125[2] , \wBMid125[1] , \wBMid125[0] }), .HiOut({
        \wRegInB125[31] , \wRegInB125[30] , \wRegInB125[29] , \wRegInB125[28] , 
        \wRegInB125[27] , \wRegInB125[26] , \wRegInB125[25] , \wRegInB125[24] , 
        \wRegInB125[23] , \wRegInB125[22] , \wRegInB125[21] , \wRegInB125[20] , 
        \wRegInB125[19] , \wRegInB125[18] , \wRegInB125[17] , \wRegInB125[16] , 
        \wRegInB125[15] , \wRegInB125[14] , \wRegInB125[13] , \wRegInB125[12] , 
        \wRegInB125[11] , \wRegInB125[10] , \wRegInB125[9] , \wRegInB125[8] , 
        \wRegInB125[7] , \wRegInB125[6] , \wRegInB125[5] , \wRegInB125[4] , 
        \wRegInB125[3] , \wRegInB125[2] , \wRegInB125[1] , \wRegInB125[0] }), 
        .LoOut({\wRegInA126[31] , \wRegInA126[30] , \wRegInA126[29] , 
        \wRegInA126[28] , \wRegInA126[27] , \wRegInA126[26] , \wRegInA126[25] , 
        \wRegInA126[24] , \wRegInA126[23] , \wRegInA126[22] , \wRegInA126[21] , 
        \wRegInA126[20] , \wRegInA126[19] , \wRegInA126[18] , \wRegInA126[17] , 
        \wRegInA126[16] , \wRegInA126[15] , \wRegInA126[14] , \wRegInA126[13] , 
        \wRegInA126[12] , \wRegInA126[11] , \wRegInA126[10] , \wRegInA126[9] , 
        \wRegInA126[8] , \wRegInA126[7] , \wRegInA126[6] , \wRegInA126[5] , 
        \wRegInA126[4] , \wRegInA126[3] , \wRegInA126[2] , \wRegInA126[1] , 
        \wRegInA126[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_198 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink199[31] , \ScanLink199[30] , \ScanLink199[29] , 
        \ScanLink199[28] , \ScanLink199[27] , \ScanLink199[26] , 
        \ScanLink199[25] , \ScanLink199[24] , \ScanLink199[23] , 
        \ScanLink199[22] , \ScanLink199[21] , \ScanLink199[20] , 
        \ScanLink199[19] , \ScanLink199[18] , \ScanLink199[17] , 
        \ScanLink199[16] , \ScanLink199[15] , \ScanLink199[14] , 
        \ScanLink199[13] , \ScanLink199[12] , \ScanLink199[11] , 
        \ScanLink199[10] , \ScanLink199[9] , \ScanLink199[8] , 
        \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , \ScanLink199[4] , 
        \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , \ScanLink199[0] 
        }), .ScanOut({\ScanLink198[31] , \ScanLink198[30] , \ScanLink198[29] , 
        \ScanLink198[28] , \ScanLink198[27] , \ScanLink198[26] , 
        \ScanLink198[25] , \ScanLink198[24] , \ScanLink198[23] , 
        \ScanLink198[22] , \ScanLink198[21] , \ScanLink198[20] , 
        \ScanLink198[19] , \ScanLink198[18] , \ScanLink198[17] , 
        \ScanLink198[16] , \ScanLink198[15] , \ScanLink198[14] , 
        \ScanLink198[13] , \ScanLink198[12] , \ScanLink198[11] , 
        \ScanLink198[10] , \ScanLink198[9] , \ScanLink198[8] , 
        \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , \ScanLink198[4] , 
        \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , \ScanLink198[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB28[31] , \wRegInB28[30] , \wRegInB28[29] , 
        \wRegInB28[28] , \wRegInB28[27] , \wRegInB28[26] , \wRegInB28[25] , 
        \wRegInB28[24] , \wRegInB28[23] , \wRegInB28[22] , \wRegInB28[21] , 
        \wRegInB28[20] , \wRegInB28[19] , \wRegInB28[18] , \wRegInB28[17] , 
        \wRegInB28[16] , \wRegInB28[15] , \wRegInB28[14] , \wRegInB28[13] , 
        \wRegInB28[12] , \wRegInB28[11] , \wRegInB28[10] , \wRegInB28[9] , 
        \wRegInB28[8] , \wRegInB28[7] , \wRegInB28[6] , \wRegInB28[5] , 
        \wRegInB28[4] , \wRegInB28[3] , \wRegInB28[2] , \wRegInB28[1] , 
        \wRegInB28[0] }), .Out({\wBIn28[31] , \wBIn28[30] , \wBIn28[29] , 
        \wBIn28[28] , \wBIn28[27] , \wBIn28[26] , \wBIn28[25] , \wBIn28[24] , 
        \wBIn28[23] , \wBIn28[22] , \wBIn28[21] , \wBIn28[20] , \wBIn28[19] , 
        \wBIn28[18] , \wBIn28[17] , \wBIn28[16] , \wBIn28[15] , \wBIn28[14] , 
        \wBIn28[13] , \wBIn28[12] , \wBIn28[11] , \wBIn28[10] , \wBIn28[9] , 
        \wBIn28[8] , \wBIn28[7] , \wBIn28[6] , \wBIn28[5] , \wBIn28[4] , 
        \wBIn28[3] , \wBIn28[2] , \wBIn28[1] , \wBIn28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_81 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink82[31] , \ScanLink82[30] , \ScanLink82[29] , 
        \ScanLink82[28] , \ScanLink82[27] , \ScanLink82[26] , \ScanLink82[25] , 
        \ScanLink82[24] , \ScanLink82[23] , \ScanLink82[22] , \ScanLink82[21] , 
        \ScanLink82[20] , \ScanLink82[19] , \ScanLink82[18] , \ScanLink82[17] , 
        \ScanLink82[16] , \ScanLink82[15] , \ScanLink82[14] , \ScanLink82[13] , 
        \ScanLink82[12] , \ScanLink82[11] , \ScanLink82[10] , \ScanLink82[9] , 
        \ScanLink82[8] , \ScanLink82[7] , \ScanLink82[6] , \ScanLink82[5] , 
        \ScanLink82[4] , \ScanLink82[3] , \ScanLink82[2] , \ScanLink82[1] , 
        \ScanLink82[0] }), .ScanOut({\ScanLink81[31] , \ScanLink81[30] , 
        \ScanLink81[29] , \ScanLink81[28] , \ScanLink81[27] , \ScanLink81[26] , 
        \ScanLink81[25] , \ScanLink81[24] , \ScanLink81[23] , \ScanLink81[22] , 
        \ScanLink81[21] , \ScanLink81[20] , \ScanLink81[19] , \ScanLink81[18] , 
        \ScanLink81[17] , \ScanLink81[16] , \ScanLink81[15] , \ScanLink81[14] , 
        \ScanLink81[13] , \ScanLink81[12] , \ScanLink81[11] , \ScanLink81[10] , 
        \ScanLink81[9] , \ScanLink81[8] , \ScanLink81[7] , \ScanLink81[6] , 
        \ScanLink81[5] , \ScanLink81[4] , \ScanLink81[3] , \ScanLink81[2] , 
        \ScanLink81[1] , \ScanLink81[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA87[31] , \wRegInA87[30] , 
        \wRegInA87[29] , \wRegInA87[28] , \wRegInA87[27] , \wRegInA87[26] , 
        \wRegInA87[25] , \wRegInA87[24] , \wRegInA87[23] , \wRegInA87[22] , 
        \wRegInA87[21] , \wRegInA87[20] , \wRegInA87[19] , \wRegInA87[18] , 
        \wRegInA87[17] , \wRegInA87[16] , \wRegInA87[15] , \wRegInA87[14] , 
        \wRegInA87[13] , \wRegInA87[12] , \wRegInA87[11] , \wRegInA87[10] , 
        \wRegInA87[9] , \wRegInA87[8] , \wRegInA87[7] , \wRegInA87[6] , 
        \wRegInA87[5] , \wRegInA87[4] , \wRegInA87[3] , \wRegInA87[2] , 
        \wRegInA87[1] , \wRegInA87[0] }), .Out({\wAIn87[31] , \wAIn87[30] , 
        \wAIn87[29] , \wAIn87[28] , \wAIn87[27] , \wAIn87[26] , \wAIn87[25] , 
        \wAIn87[24] , \wAIn87[23] , \wAIn87[22] , \wAIn87[21] , \wAIn87[20] , 
        \wAIn87[19] , \wAIn87[18] , \wAIn87[17] , \wAIn87[16] , \wAIn87[15] , 
        \wAIn87[14] , \wAIn87[13] , \wAIn87[12] , \wAIn87[11] , \wAIn87[10] , 
        \wAIn87[9] , \wAIn87[8] , \wAIn87[7] , \wAIn87[6] , \wAIn87[5] , 
        \wAIn87[4] , \wAIn87[3] , \wAIn87[2] , \wAIn87[1] , \wAIn87[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid48[31] , \wAMid48[30] , \wAMid48[29] , \wAMid48[28] , 
        \wAMid48[27] , \wAMid48[26] , \wAMid48[25] , \wAMid48[24] , 
        \wAMid48[23] , \wAMid48[22] , \wAMid48[21] , \wAMid48[20] , 
        \wAMid48[19] , \wAMid48[18] , \wAMid48[17] , \wAMid48[16] , 
        \wAMid48[15] , \wAMid48[14] , \wAMid48[13] , \wAMid48[12] , 
        \wAMid48[11] , \wAMid48[10] , \wAMid48[9] , \wAMid48[8] , \wAMid48[7] , 
        \wAMid48[6] , \wAMid48[5] , \wAMid48[4] , \wAMid48[3] , \wAMid48[2] , 
        \wAMid48[1] , \wAMid48[0] }), .BIn({\wBMid48[31] , \wBMid48[30] , 
        \wBMid48[29] , \wBMid48[28] , \wBMid48[27] , \wBMid48[26] , 
        \wBMid48[25] , \wBMid48[24] , \wBMid48[23] , \wBMid48[22] , 
        \wBMid48[21] , \wBMid48[20] , \wBMid48[19] , \wBMid48[18] , 
        \wBMid48[17] , \wBMid48[16] , \wBMid48[15] , \wBMid48[14] , 
        \wBMid48[13] , \wBMid48[12] , \wBMid48[11] , \wBMid48[10] , 
        \wBMid48[9] , \wBMid48[8] , \wBMid48[7] , \wBMid48[6] , \wBMid48[5] , 
        \wBMid48[4] , \wBMid48[3] , \wBMid48[2] , \wBMid48[1] , \wBMid48[0] }), 
        .HiOut({\wRegInB48[31] , \wRegInB48[30] , \wRegInB48[29] , 
        \wRegInB48[28] , \wRegInB48[27] , \wRegInB48[26] , \wRegInB48[25] , 
        \wRegInB48[24] , \wRegInB48[23] , \wRegInB48[22] , \wRegInB48[21] , 
        \wRegInB48[20] , \wRegInB48[19] , \wRegInB48[18] , \wRegInB48[17] , 
        \wRegInB48[16] , \wRegInB48[15] , \wRegInB48[14] , \wRegInB48[13] , 
        \wRegInB48[12] , \wRegInB48[11] , \wRegInB48[10] , \wRegInB48[9] , 
        \wRegInB48[8] , \wRegInB48[7] , \wRegInB48[6] , \wRegInB48[5] , 
        \wRegInB48[4] , \wRegInB48[3] , \wRegInB48[2] , \wRegInB48[1] , 
        \wRegInB48[0] }), .LoOut({\wRegInA49[31] , \wRegInA49[30] , 
        \wRegInA49[29] , \wRegInA49[28] , \wRegInA49[27] , \wRegInA49[26] , 
        \wRegInA49[25] , \wRegInA49[24] , \wRegInA49[23] , \wRegInA49[22] , 
        \wRegInA49[21] , \wRegInA49[20] , \wRegInA49[19] , \wRegInA49[18] , 
        \wRegInA49[17] , \wRegInA49[16] , \wRegInA49[15] , \wRegInA49[14] , 
        \wRegInA49[13] , \wRegInA49[12] , \wRegInA49[11] , \wRegInA49[10] , 
        \wRegInA49[9] , \wRegInA49[8] , \wRegInA49[7] , \wRegInA49[6] , 
        \wRegInA49[5] , \wRegInA49[4] , \wRegInA49[3] , \wRegInA49[2] , 
        \wRegInA49[1] , \wRegInA49[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn63[31] , \wAIn63[30] , \wAIn63[29] , \wAIn63[28] , \wAIn63[27] , 
        \wAIn63[26] , \wAIn63[25] , \wAIn63[24] , \wAIn63[23] , \wAIn63[22] , 
        \wAIn63[21] , \wAIn63[20] , \wAIn63[19] , \wAIn63[18] , \wAIn63[17] , 
        \wAIn63[16] , \wAIn63[15] , \wAIn63[14] , \wAIn63[13] , \wAIn63[12] , 
        \wAIn63[11] , \wAIn63[10] , \wAIn63[9] , \wAIn63[8] , \wAIn63[7] , 
        \wAIn63[6] , \wAIn63[5] , \wAIn63[4] , \wAIn63[3] , \wAIn63[2] , 
        \wAIn63[1] , \wAIn63[0] }), .BIn({\wBIn63[31] , \wBIn63[30] , 
        \wBIn63[29] , \wBIn63[28] , \wBIn63[27] , \wBIn63[26] , \wBIn63[25] , 
        \wBIn63[24] , \wBIn63[23] , \wBIn63[22] , \wBIn63[21] , \wBIn63[20] , 
        \wBIn63[19] , \wBIn63[18] , \wBIn63[17] , \wBIn63[16] , \wBIn63[15] , 
        \wBIn63[14] , \wBIn63[13] , \wBIn63[12] , \wBIn63[11] , \wBIn63[10] , 
        \wBIn63[9] , \wBIn63[8] , \wBIn63[7] , \wBIn63[6] , \wBIn63[5] , 
        \wBIn63[4] , \wBIn63[3] , \wBIn63[2] , \wBIn63[1] , \wBIn63[0] }), 
        .HiOut({\wBMid62[31] , \wBMid62[30] , \wBMid62[29] , \wBMid62[28] , 
        \wBMid62[27] , \wBMid62[26] , \wBMid62[25] , \wBMid62[24] , 
        \wBMid62[23] , \wBMid62[22] , \wBMid62[21] , \wBMid62[20] , 
        \wBMid62[19] , \wBMid62[18] , \wBMid62[17] , \wBMid62[16] , 
        \wBMid62[15] , \wBMid62[14] , \wBMid62[13] , \wBMid62[12] , 
        \wBMid62[11] , \wBMid62[10] , \wBMid62[9] , \wBMid62[8] , \wBMid62[7] , 
        \wBMid62[6] , \wBMid62[5] , \wBMid62[4] , \wBMid62[3] , \wBMid62[2] , 
        \wBMid62[1] , \wBMid62[0] }), .LoOut({\wAMid63[31] , \wAMid63[30] , 
        \wAMid63[29] , \wAMid63[28] , \wAMid63[27] , \wAMid63[26] , 
        \wAMid63[25] , \wAMid63[24] , \wAMid63[23] , \wAMid63[22] , 
        \wAMid63[21] , \wAMid63[20] , \wAMid63[19] , \wAMid63[18] , 
        \wAMid63[17] , \wAMid63[16] , \wAMid63[15] , \wAMid63[14] , 
        \wAMid63[13] , \wAMid63[12] , \wAMid63[11] , \wAMid63[10] , 
        \wAMid63[9] , \wAMid63[8] , \wAMid63[7] , \wAMid63[6] , \wAMid63[5] , 
        \wAMid63[4] , \wAMid63[3] , \wAMid63[2] , \wAMid63[1] , \wAMid63[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid74[31] , \wAMid74[30] , \wAMid74[29] , \wAMid74[28] , 
        \wAMid74[27] , \wAMid74[26] , \wAMid74[25] , \wAMid74[24] , 
        \wAMid74[23] , \wAMid74[22] , \wAMid74[21] , \wAMid74[20] , 
        \wAMid74[19] , \wAMid74[18] , \wAMid74[17] , \wAMid74[16] , 
        \wAMid74[15] , \wAMid74[14] , \wAMid74[13] , \wAMid74[12] , 
        \wAMid74[11] , \wAMid74[10] , \wAMid74[9] , \wAMid74[8] , \wAMid74[7] , 
        \wAMid74[6] , \wAMid74[5] , \wAMid74[4] , \wAMid74[3] , \wAMid74[2] , 
        \wAMid74[1] , \wAMid74[0] }), .BIn({\wBMid74[31] , \wBMid74[30] , 
        \wBMid74[29] , \wBMid74[28] , \wBMid74[27] , \wBMid74[26] , 
        \wBMid74[25] , \wBMid74[24] , \wBMid74[23] , \wBMid74[22] , 
        \wBMid74[21] , \wBMid74[20] , \wBMid74[19] , \wBMid74[18] , 
        \wBMid74[17] , \wBMid74[16] , \wBMid74[15] , \wBMid74[14] , 
        \wBMid74[13] , \wBMid74[12] , \wBMid74[11] , \wBMid74[10] , 
        \wBMid74[9] , \wBMid74[8] , \wBMid74[7] , \wBMid74[6] , \wBMid74[5] , 
        \wBMid74[4] , \wBMid74[3] , \wBMid74[2] , \wBMid74[1] , \wBMid74[0] }), 
        .HiOut({\wRegInB74[31] , \wRegInB74[30] , \wRegInB74[29] , 
        \wRegInB74[28] , \wRegInB74[27] , \wRegInB74[26] , \wRegInB74[25] , 
        \wRegInB74[24] , \wRegInB74[23] , \wRegInB74[22] , \wRegInB74[21] , 
        \wRegInB74[20] , \wRegInB74[19] , \wRegInB74[18] , \wRegInB74[17] , 
        \wRegInB74[16] , \wRegInB74[15] , \wRegInB74[14] , \wRegInB74[13] , 
        \wRegInB74[12] , \wRegInB74[11] , \wRegInB74[10] , \wRegInB74[9] , 
        \wRegInB74[8] , \wRegInB74[7] , \wRegInB74[6] , \wRegInB74[5] , 
        \wRegInB74[4] , \wRegInB74[3] , \wRegInB74[2] , \wRegInB74[1] , 
        \wRegInB74[0] }), .LoOut({\wRegInA75[31] , \wRegInA75[30] , 
        \wRegInA75[29] , \wRegInA75[28] , \wRegInA75[27] , \wRegInA75[26] , 
        \wRegInA75[25] , \wRegInA75[24] , \wRegInA75[23] , \wRegInA75[22] , 
        \wRegInA75[21] , \wRegInA75[20] , \wRegInA75[19] , \wRegInA75[18] , 
        \wRegInA75[17] , \wRegInA75[16] , \wRegInA75[15] , \wRegInA75[14] , 
        \wRegInA75[13] , \wRegInA75[12] , \wRegInA75[11] , \wRegInA75[10] , 
        \wRegInA75[9] , \wRegInA75[8] , \wRegInA75[7] , \wRegInA75[6] , 
        \wRegInA75[5] , \wRegInA75[4] , \wRegInA75[3] , \wRegInA75[2] , 
        \wRegInA75[1] , \wRegInA75[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_141 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink142[31] , \ScanLink142[30] , \ScanLink142[29] , 
        \ScanLink142[28] , \ScanLink142[27] , \ScanLink142[26] , 
        \ScanLink142[25] , \ScanLink142[24] , \ScanLink142[23] , 
        \ScanLink142[22] , \ScanLink142[21] , \ScanLink142[20] , 
        \ScanLink142[19] , \ScanLink142[18] , \ScanLink142[17] , 
        \ScanLink142[16] , \ScanLink142[15] , \ScanLink142[14] , 
        \ScanLink142[13] , \ScanLink142[12] , \ScanLink142[11] , 
        \ScanLink142[10] , \ScanLink142[9] , \ScanLink142[8] , 
        \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , \ScanLink142[4] , 
        \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , \ScanLink142[0] 
        }), .ScanOut({\ScanLink141[31] , \ScanLink141[30] , \ScanLink141[29] , 
        \ScanLink141[28] , \ScanLink141[27] , \ScanLink141[26] , 
        \ScanLink141[25] , \ScanLink141[24] , \ScanLink141[23] , 
        \ScanLink141[22] , \ScanLink141[21] , \ScanLink141[20] , 
        \ScanLink141[19] , \ScanLink141[18] , \ScanLink141[17] , 
        \ScanLink141[16] , \ScanLink141[15] , \ScanLink141[14] , 
        \ScanLink141[13] , \ScanLink141[12] , \ScanLink141[11] , 
        \ScanLink141[10] , \ScanLink141[9] , \ScanLink141[8] , 
        \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , \ScanLink141[4] , 
        \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , \ScanLink141[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA57[31] , \wRegInA57[30] , \wRegInA57[29] , 
        \wRegInA57[28] , \wRegInA57[27] , \wRegInA57[26] , \wRegInA57[25] , 
        \wRegInA57[24] , \wRegInA57[23] , \wRegInA57[22] , \wRegInA57[21] , 
        \wRegInA57[20] , \wRegInA57[19] , \wRegInA57[18] , \wRegInA57[17] , 
        \wRegInA57[16] , \wRegInA57[15] , \wRegInA57[14] , \wRegInA57[13] , 
        \wRegInA57[12] , \wRegInA57[11] , \wRegInA57[10] , \wRegInA57[9] , 
        \wRegInA57[8] , \wRegInA57[7] , \wRegInA57[6] , \wRegInA57[5] , 
        \wRegInA57[4] , \wRegInA57[3] , \wRegInA57[2] , \wRegInA57[1] , 
        \wRegInA57[0] }), .Out({\wAIn57[31] , \wAIn57[30] , \wAIn57[29] , 
        \wAIn57[28] , \wAIn57[27] , \wAIn57[26] , \wAIn57[25] , \wAIn57[24] , 
        \wAIn57[23] , \wAIn57[22] , \wAIn57[21] , \wAIn57[20] , \wAIn57[19] , 
        \wAIn57[18] , \wAIn57[17] , \wAIn57[16] , \wAIn57[15] , \wAIn57[14] , 
        \wAIn57[13] , \wAIn57[12] , \wAIn57[11] , \wAIn57[10] , \wAIn57[9] , 
        \wAIn57[8] , \wAIn57[7] , \wAIn57[6] , \wAIn57[5] , \wAIn57[4] , 
        \wAIn57[3] , \wAIn57[2] , \wAIn57[1] , \wAIn57[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_11 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[31] , \ScanLink12[30] , \ScanLink12[29] , 
        \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , \ScanLink12[25] , 
        \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , \ScanLink12[21] , 
        \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , \ScanLink12[17] , 
        \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , \ScanLink12[13] , 
        \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , \ScanLink12[9] , 
        \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA122[31] , \wRegInA122[30] , 
        \wRegInA122[29] , \wRegInA122[28] , \wRegInA122[27] , \wRegInA122[26] , 
        \wRegInA122[25] , \wRegInA122[24] , \wRegInA122[23] , \wRegInA122[22] , 
        \wRegInA122[21] , \wRegInA122[20] , \wRegInA122[19] , \wRegInA122[18] , 
        \wRegInA122[17] , \wRegInA122[16] , \wRegInA122[15] , \wRegInA122[14] , 
        \wRegInA122[13] , \wRegInA122[12] , \wRegInA122[11] , \wRegInA122[10] , 
        \wRegInA122[9] , \wRegInA122[8] , \wRegInA122[7] , \wRegInA122[6] , 
        \wRegInA122[5] , \wRegInA122[4] , \wRegInA122[3] , \wRegInA122[2] , 
        \wRegInA122[1] , \wRegInA122[0] }), .Out({\wAIn122[31] , \wAIn122[30] , 
        \wAIn122[29] , \wAIn122[28] , \wAIn122[27] , \wAIn122[26] , 
        \wAIn122[25] , \wAIn122[24] , \wAIn122[23] , \wAIn122[22] , 
        \wAIn122[21] , \wAIn122[20] , \wAIn122[19] , \wAIn122[18] , 
        \wAIn122[17] , \wAIn122[16] , \wAIn122[15] , \wAIn122[14] , 
        \wAIn122[13] , \wAIn122[12] , \wAIn122[11] , \wAIn122[10] , 
        \wAIn122[9] , \wAIn122[8] , \wAIn122[7] , \wAIn122[6] , \wAIn122[5] , 
        \wAIn122[4] , \wAIn122[3] , \wAIn122[2] , \wAIn122[1] , \wAIn122[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn86[31] , \wAIn86[30] , \wAIn86[29] , \wAIn86[28] , \wAIn86[27] , 
        \wAIn86[26] , \wAIn86[25] , \wAIn86[24] , \wAIn86[23] , \wAIn86[22] , 
        \wAIn86[21] , \wAIn86[20] , \wAIn86[19] , \wAIn86[18] , \wAIn86[17] , 
        \wAIn86[16] , \wAIn86[15] , \wAIn86[14] , \wAIn86[13] , \wAIn86[12] , 
        \wAIn86[11] , \wAIn86[10] , \wAIn86[9] , \wAIn86[8] , \wAIn86[7] , 
        \wAIn86[6] , \wAIn86[5] , \wAIn86[4] , \wAIn86[3] , \wAIn86[2] , 
        \wAIn86[1] , \wAIn86[0] }), .BIn({\wBIn86[31] , \wBIn86[30] , 
        \wBIn86[29] , \wBIn86[28] , \wBIn86[27] , \wBIn86[26] , \wBIn86[25] , 
        \wBIn86[24] , \wBIn86[23] , \wBIn86[22] , \wBIn86[21] , \wBIn86[20] , 
        \wBIn86[19] , \wBIn86[18] , \wBIn86[17] , \wBIn86[16] , \wBIn86[15] , 
        \wBIn86[14] , \wBIn86[13] , \wBIn86[12] , \wBIn86[11] , \wBIn86[10] , 
        \wBIn86[9] , \wBIn86[8] , \wBIn86[7] , \wBIn86[6] , \wBIn86[5] , 
        \wBIn86[4] , \wBIn86[3] , \wBIn86[2] , \wBIn86[1] , \wBIn86[0] }), 
        .HiOut({\wBMid85[31] , \wBMid85[30] , \wBMid85[29] , \wBMid85[28] , 
        \wBMid85[27] , \wBMid85[26] , \wBMid85[25] , \wBMid85[24] , 
        \wBMid85[23] , \wBMid85[22] , \wBMid85[21] , \wBMid85[20] , 
        \wBMid85[19] , \wBMid85[18] , \wBMid85[17] , \wBMid85[16] , 
        \wBMid85[15] , \wBMid85[14] , \wBMid85[13] , \wBMid85[12] , 
        \wBMid85[11] , \wBMid85[10] , \wBMid85[9] , \wBMid85[8] , \wBMid85[7] , 
        \wBMid85[6] , \wBMid85[5] , \wBMid85[4] , \wBMid85[3] , \wBMid85[2] , 
        \wBMid85[1] , \wBMid85[0] }), .LoOut({\wAMid86[31] , \wAMid86[30] , 
        \wAMid86[29] , \wAMid86[28] , \wAMid86[27] , \wAMid86[26] , 
        \wAMid86[25] , \wAMid86[24] , \wAMid86[23] , \wAMid86[22] , 
        \wAMid86[21] , \wAMid86[20] , \wAMid86[19] , \wAMid86[18] , 
        \wAMid86[17] , \wAMid86[16] , \wAMid86[15] , \wAMid86[14] , 
        \wAMid86[13] , \wAMid86[12] , \wAMid86[11] , \wAMid86[10] , 
        \wAMid86[9] , \wAMid86[8] , \wAMid86[7] , \wAMid86[6] , \wAMid86[5] , 
        \wAMid86[4] , \wAMid86[3] , \wAMid86[2] , \wAMid86[1] , \wAMid86[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn113[31] , \wAIn113[30] , \wAIn113[29] , \wAIn113[28] , 
        \wAIn113[27] , \wAIn113[26] , \wAIn113[25] , \wAIn113[24] , 
        \wAIn113[23] , \wAIn113[22] , \wAIn113[21] , \wAIn113[20] , 
        \wAIn113[19] , \wAIn113[18] , \wAIn113[17] , \wAIn113[16] , 
        \wAIn113[15] , \wAIn113[14] , \wAIn113[13] , \wAIn113[12] , 
        \wAIn113[11] , \wAIn113[10] , \wAIn113[9] , \wAIn113[8] , \wAIn113[7] , 
        \wAIn113[6] , \wAIn113[5] , \wAIn113[4] , \wAIn113[3] , \wAIn113[2] , 
        \wAIn113[1] , \wAIn113[0] }), .BIn({\wBIn113[31] , \wBIn113[30] , 
        \wBIn113[29] , \wBIn113[28] , \wBIn113[27] , \wBIn113[26] , 
        \wBIn113[25] , \wBIn113[24] , \wBIn113[23] , \wBIn113[22] , 
        \wBIn113[21] , \wBIn113[20] , \wBIn113[19] , \wBIn113[18] , 
        \wBIn113[17] , \wBIn113[16] , \wBIn113[15] , \wBIn113[14] , 
        \wBIn113[13] , \wBIn113[12] , \wBIn113[11] , \wBIn113[10] , 
        \wBIn113[9] , \wBIn113[8] , \wBIn113[7] , \wBIn113[6] , \wBIn113[5] , 
        \wBIn113[4] , \wBIn113[3] , \wBIn113[2] , \wBIn113[1] , \wBIn113[0] }), 
        .HiOut({\wBMid112[31] , \wBMid112[30] , \wBMid112[29] , \wBMid112[28] , 
        \wBMid112[27] , \wBMid112[26] , \wBMid112[25] , \wBMid112[24] , 
        \wBMid112[23] , \wBMid112[22] , \wBMid112[21] , \wBMid112[20] , 
        \wBMid112[19] , \wBMid112[18] , \wBMid112[17] , \wBMid112[16] , 
        \wBMid112[15] , \wBMid112[14] , \wBMid112[13] , \wBMid112[12] , 
        \wBMid112[11] , \wBMid112[10] , \wBMid112[9] , \wBMid112[8] , 
        \wBMid112[7] , \wBMid112[6] , \wBMid112[5] , \wBMid112[4] , 
        \wBMid112[3] , \wBMid112[2] , \wBMid112[1] , \wBMid112[0] }), .LoOut({
        \wAMid113[31] , \wAMid113[30] , \wAMid113[29] , \wAMid113[28] , 
        \wAMid113[27] , \wAMid113[26] , \wAMid113[25] , \wAMid113[24] , 
        \wAMid113[23] , \wAMid113[22] , \wAMid113[21] , \wAMid113[20] , 
        \wAMid113[19] , \wAMid113[18] , \wAMid113[17] , \wAMid113[16] , 
        \wAMid113[15] , \wAMid113[14] , \wAMid113[13] , \wAMid113[12] , 
        \wAMid113[11] , \wAMid113[10] , \wAMid113[9] , \wAMid113[8] , 
        \wAMid113[7] , \wAMid113[6] , \wAMid113[5] , \wAMid113[4] , 
        \wAMid113[3] , \wAMid113[2] , \wAMid113[1] , \wAMid113[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid53[31] , \wAMid53[30] , \wAMid53[29] , \wAMid53[28] , 
        \wAMid53[27] , \wAMid53[26] , \wAMid53[25] , \wAMid53[24] , 
        \wAMid53[23] , \wAMid53[22] , \wAMid53[21] , \wAMid53[20] , 
        \wAMid53[19] , \wAMid53[18] , \wAMid53[17] , \wAMid53[16] , 
        \wAMid53[15] , \wAMid53[14] , \wAMid53[13] , \wAMid53[12] , 
        \wAMid53[11] , \wAMid53[10] , \wAMid53[9] , \wAMid53[8] , \wAMid53[7] , 
        \wAMid53[6] , \wAMid53[5] , \wAMid53[4] , \wAMid53[3] , \wAMid53[2] , 
        \wAMid53[1] , \wAMid53[0] }), .BIn({\wBMid53[31] , \wBMid53[30] , 
        \wBMid53[29] , \wBMid53[28] , \wBMid53[27] , \wBMid53[26] , 
        \wBMid53[25] , \wBMid53[24] , \wBMid53[23] , \wBMid53[22] , 
        \wBMid53[21] , \wBMid53[20] , \wBMid53[19] , \wBMid53[18] , 
        \wBMid53[17] , \wBMid53[16] , \wBMid53[15] , \wBMid53[14] , 
        \wBMid53[13] , \wBMid53[12] , \wBMid53[11] , \wBMid53[10] , 
        \wBMid53[9] , \wBMid53[8] , \wBMid53[7] , \wBMid53[6] , \wBMid53[5] , 
        \wBMid53[4] , \wBMid53[3] , \wBMid53[2] , \wBMid53[1] , \wBMid53[0] }), 
        .HiOut({\wRegInB53[31] , \wRegInB53[30] , \wRegInB53[29] , 
        \wRegInB53[28] , \wRegInB53[27] , \wRegInB53[26] , \wRegInB53[25] , 
        \wRegInB53[24] , \wRegInB53[23] , \wRegInB53[22] , \wRegInB53[21] , 
        \wRegInB53[20] , \wRegInB53[19] , \wRegInB53[18] , \wRegInB53[17] , 
        \wRegInB53[16] , \wRegInB53[15] , \wRegInB53[14] , \wRegInB53[13] , 
        \wRegInB53[12] , \wRegInB53[11] , \wRegInB53[10] , \wRegInB53[9] , 
        \wRegInB53[8] , \wRegInB53[7] , \wRegInB53[6] , \wRegInB53[5] , 
        \wRegInB53[4] , \wRegInB53[3] , \wRegInB53[2] , \wRegInB53[1] , 
        \wRegInB53[0] }), .LoOut({\wRegInA54[31] , \wRegInA54[30] , 
        \wRegInA54[29] , \wRegInA54[28] , \wRegInA54[27] , \wRegInA54[26] , 
        \wRegInA54[25] , \wRegInA54[24] , \wRegInA54[23] , \wRegInA54[22] , 
        \wRegInA54[21] , \wRegInA54[20] , \wRegInA54[19] , \wRegInA54[18] , 
        \wRegInA54[17] , \wRegInA54[16] , \wRegInA54[15] , \wRegInA54[14] , 
        \wRegInA54[13] , \wRegInA54[12] , \wRegInA54[11] , \wRegInA54[10] , 
        \wRegInA54[9] , \wRegInA54[8] , \wRegInA54[7] , \wRegInA54[6] , 
        \wRegInA54[5] , \wRegInA54[4] , \wRegInA54[3] , \wRegInA54[2] , 
        \wRegInA54[1] , \wRegInA54[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_166 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink167[31] , \ScanLink167[30] , \ScanLink167[29] , 
        \ScanLink167[28] , \ScanLink167[27] , \ScanLink167[26] , 
        \ScanLink167[25] , \ScanLink167[24] , \ScanLink167[23] , 
        \ScanLink167[22] , \ScanLink167[21] , \ScanLink167[20] , 
        \ScanLink167[19] , \ScanLink167[18] , \ScanLink167[17] , 
        \ScanLink167[16] , \ScanLink167[15] , \ScanLink167[14] , 
        \ScanLink167[13] , \ScanLink167[12] , \ScanLink167[11] , 
        \ScanLink167[10] , \ScanLink167[9] , \ScanLink167[8] , 
        \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , \ScanLink167[4] , 
        \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , \ScanLink167[0] 
        }), .ScanOut({\ScanLink166[31] , \ScanLink166[30] , \ScanLink166[29] , 
        \ScanLink166[28] , \ScanLink166[27] , \ScanLink166[26] , 
        \ScanLink166[25] , \ScanLink166[24] , \ScanLink166[23] , 
        \ScanLink166[22] , \ScanLink166[21] , \ScanLink166[20] , 
        \ScanLink166[19] , \ScanLink166[18] , \ScanLink166[17] , 
        \ScanLink166[16] , \ScanLink166[15] , \ScanLink166[14] , 
        \ScanLink166[13] , \ScanLink166[12] , \ScanLink166[11] , 
        \ScanLink166[10] , \ScanLink166[9] , \ScanLink166[8] , 
        \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , \ScanLink166[4] , 
        \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , \ScanLink166[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB44[31] , \wRegInB44[30] , \wRegInB44[29] , 
        \wRegInB44[28] , \wRegInB44[27] , \wRegInB44[26] , \wRegInB44[25] , 
        \wRegInB44[24] , \wRegInB44[23] , \wRegInB44[22] , \wRegInB44[21] , 
        \wRegInB44[20] , \wRegInB44[19] , \wRegInB44[18] , \wRegInB44[17] , 
        \wRegInB44[16] , \wRegInB44[15] , \wRegInB44[14] , \wRegInB44[13] , 
        \wRegInB44[12] , \wRegInB44[11] , \wRegInB44[10] , \wRegInB44[9] , 
        \wRegInB44[8] , \wRegInB44[7] , \wRegInB44[6] , \wRegInB44[5] , 
        \wRegInB44[4] , \wRegInB44[3] , \wRegInB44[2] , \wRegInB44[1] , 
        \wRegInB44[0] }), .Out({\wBIn44[31] , \wBIn44[30] , \wBIn44[29] , 
        \wBIn44[28] , \wBIn44[27] , \wBIn44[26] , \wBIn44[25] , \wBIn44[24] , 
        \wBIn44[23] , \wBIn44[22] , \wBIn44[21] , \wBIn44[20] , \wBIn44[19] , 
        \wBIn44[18] , \wBIn44[17] , \wBIn44[16] , \wBIn44[15] , \wBIn44[14] , 
        \wBIn44[13] , \wBIn44[12] , \wBIn44[11] , \wBIn44[10] , \wBIn44[9] , 
        \wBIn44[8] , \wBIn44[7] , \wBIn44[6] , \wBIn44[5] , \wBIn44[4] , 
        \wBIn44[3] , \wBIn44[2] , \wBIn44[1] , \wBIn44[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_36 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink37[31] , \ScanLink37[30] , \ScanLink37[29] , 
        \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , \ScanLink37[25] , 
        \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , \ScanLink37[21] , 
        \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , \ScanLink37[17] , 
        \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , \ScanLink37[13] , 
        \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , \ScanLink37[9] , 
        \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , \ScanLink37[5] , 
        \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , \ScanLink37[1] , 
        \ScanLink37[0] }), .ScanOut({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB109[31] , \wRegInB109[30] , 
        \wRegInB109[29] , \wRegInB109[28] , \wRegInB109[27] , \wRegInB109[26] , 
        \wRegInB109[25] , \wRegInB109[24] , \wRegInB109[23] , \wRegInB109[22] , 
        \wRegInB109[21] , \wRegInB109[20] , \wRegInB109[19] , \wRegInB109[18] , 
        \wRegInB109[17] , \wRegInB109[16] , \wRegInB109[15] , \wRegInB109[14] , 
        \wRegInB109[13] , \wRegInB109[12] , \wRegInB109[11] , \wRegInB109[10] , 
        \wRegInB109[9] , \wRegInB109[8] , \wRegInB109[7] , \wRegInB109[6] , 
        \wRegInB109[5] , \wRegInB109[4] , \wRegInB109[3] , \wRegInB109[2] , 
        \wRegInB109[1] , \wRegInB109[0] }), .Out({\wBIn109[31] , \wBIn109[30] , 
        \wBIn109[29] , \wBIn109[28] , \wBIn109[27] , \wBIn109[26] , 
        \wBIn109[25] , \wBIn109[24] , \wBIn109[23] , \wBIn109[22] , 
        \wBIn109[21] , \wBIn109[20] , \wBIn109[19] , \wBIn109[18] , 
        \wBIn109[17] , \wBIn109[16] , \wBIn109[15] , \wBIn109[14] , 
        \wBIn109[13] , \wBIn109[12] , \wBIn109[11] , \wBIn109[10] , 
        \wBIn109[9] , \wBIn109[8] , \wBIn109[7] , \wBIn109[6] , \wBIn109[5] , 
        \wBIn109[4] , \wBIn109[3] , \wBIn109[2] , \wBIn109[1] , \wBIn109[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid119[31] , \wAMid119[30] , \wAMid119[29] , \wAMid119[28] , 
        \wAMid119[27] , \wAMid119[26] , \wAMid119[25] , \wAMid119[24] , 
        \wAMid119[23] , \wAMid119[22] , \wAMid119[21] , \wAMid119[20] , 
        \wAMid119[19] , \wAMid119[18] , \wAMid119[17] , \wAMid119[16] , 
        \wAMid119[15] , \wAMid119[14] , \wAMid119[13] , \wAMid119[12] , 
        \wAMid119[11] , \wAMid119[10] , \wAMid119[9] , \wAMid119[8] , 
        \wAMid119[7] , \wAMid119[6] , \wAMid119[5] , \wAMid119[4] , 
        \wAMid119[3] , \wAMid119[2] , \wAMid119[1] , \wAMid119[0] }), .BIn({
        \wBMid119[31] , \wBMid119[30] , \wBMid119[29] , \wBMid119[28] , 
        \wBMid119[27] , \wBMid119[26] , \wBMid119[25] , \wBMid119[24] , 
        \wBMid119[23] , \wBMid119[22] , \wBMid119[21] , \wBMid119[20] , 
        \wBMid119[19] , \wBMid119[18] , \wBMid119[17] , \wBMid119[16] , 
        \wBMid119[15] , \wBMid119[14] , \wBMid119[13] , \wBMid119[12] , 
        \wBMid119[11] , \wBMid119[10] , \wBMid119[9] , \wBMid119[8] , 
        \wBMid119[7] , \wBMid119[6] , \wBMid119[5] , \wBMid119[4] , 
        \wBMid119[3] , \wBMid119[2] , \wBMid119[1] , \wBMid119[0] }), .HiOut({
        \wRegInB119[31] , \wRegInB119[30] , \wRegInB119[29] , \wRegInB119[28] , 
        \wRegInB119[27] , \wRegInB119[26] , \wRegInB119[25] , \wRegInB119[24] , 
        \wRegInB119[23] , \wRegInB119[22] , \wRegInB119[21] , \wRegInB119[20] , 
        \wRegInB119[19] , \wRegInB119[18] , \wRegInB119[17] , \wRegInB119[16] , 
        \wRegInB119[15] , \wRegInB119[14] , \wRegInB119[13] , \wRegInB119[12] , 
        \wRegInB119[11] , \wRegInB119[10] , \wRegInB119[9] , \wRegInB119[8] , 
        \wRegInB119[7] , \wRegInB119[6] , \wRegInB119[5] , \wRegInB119[4] , 
        \wRegInB119[3] , \wRegInB119[2] , \wRegInB119[1] , \wRegInB119[0] }), 
        .LoOut({\wRegInA120[31] , \wRegInA120[30] , \wRegInA120[29] , 
        \wRegInA120[28] , \wRegInA120[27] , \wRegInA120[26] , \wRegInA120[25] , 
        \wRegInA120[24] , \wRegInA120[23] , \wRegInA120[22] , \wRegInA120[21] , 
        \wRegInA120[20] , \wRegInA120[19] , \wRegInA120[18] , \wRegInA120[17] , 
        \wRegInA120[16] , \wRegInA120[15] , \wRegInA120[14] , \wRegInA120[13] , 
        \wRegInA120[12] , \wRegInA120[11] , \wRegInA120[10] , \wRegInA120[9] , 
        \wRegInA120[8] , \wRegInA120[7] , \wRegInA120[6] , \wRegInA120[5] , 
        \wRegInA120[4] , \wRegInA120[3] , \wRegInA120[2] , \wRegInA120[1] , 
        \wRegInA120[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_183 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink184[31] , \ScanLink184[30] , \ScanLink184[29] , 
        \ScanLink184[28] , \ScanLink184[27] , \ScanLink184[26] , 
        \ScanLink184[25] , \ScanLink184[24] , \ScanLink184[23] , 
        \ScanLink184[22] , \ScanLink184[21] , \ScanLink184[20] , 
        \ScanLink184[19] , \ScanLink184[18] , \ScanLink184[17] , 
        \ScanLink184[16] , \ScanLink184[15] , \ScanLink184[14] , 
        \ScanLink184[13] , \ScanLink184[12] , \ScanLink184[11] , 
        \ScanLink184[10] , \ScanLink184[9] , \ScanLink184[8] , 
        \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , \ScanLink184[4] , 
        \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , \ScanLink184[0] 
        }), .ScanOut({\ScanLink183[31] , \ScanLink183[30] , \ScanLink183[29] , 
        \ScanLink183[28] , \ScanLink183[27] , \ScanLink183[26] , 
        \ScanLink183[25] , \ScanLink183[24] , \ScanLink183[23] , 
        \ScanLink183[22] , \ScanLink183[21] , \ScanLink183[20] , 
        \ScanLink183[19] , \ScanLink183[18] , \ScanLink183[17] , 
        \ScanLink183[16] , \ScanLink183[15] , \ScanLink183[14] , 
        \ScanLink183[13] , \ScanLink183[12] , \ScanLink183[11] , 
        \ScanLink183[10] , \ScanLink183[9] , \ScanLink183[8] , 
        \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , \ScanLink183[4] , 
        \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , \ScanLink183[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA36[31] , \wRegInA36[30] , \wRegInA36[29] , 
        \wRegInA36[28] , \wRegInA36[27] , \wRegInA36[26] , \wRegInA36[25] , 
        \wRegInA36[24] , \wRegInA36[23] , \wRegInA36[22] , \wRegInA36[21] , 
        \wRegInA36[20] , \wRegInA36[19] , \wRegInA36[18] , \wRegInA36[17] , 
        \wRegInA36[16] , \wRegInA36[15] , \wRegInA36[14] , \wRegInA36[13] , 
        \wRegInA36[12] , \wRegInA36[11] , \wRegInA36[10] , \wRegInA36[9] , 
        \wRegInA36[8] , \wRegInA36[7] , \wRegInA36[6] , \wRegInA36[5] , 
        \wRegInA36[4] , \wRegInA36[3] , \wRegInA36[2] , \wRegInA36[1] , 
        \wRegInA36[0] }), .Out({\wAIn36[31] , \wAIn36[30] , \wAIn36[29] , 
        \wAIn36[28] , \wAIn36[27] , \wAIn36[26] , \wAIn36[25] , \wAIn36[24] , 
        \wAIn36[23] , \wAIn36[22] , \wAIn36[21] , \wAIn36[20] , \wAIn36[19] , 
        \wAIn36[18] , \wAIn36[17] , \wAIn36[16] , \wAIn36[15] , \wAIn36[14] , 
        \wAIn36[13] , \wAIn36[12] , \wAIn36[11] , \wAIn36[10] , \wAIn36[9] , 
        \wAIn36[8] , \wAIn36[7] , \wAIn36[6] , \wAIn36[5] , \wAIn36[4] , 
        \wAIn36[3] , \wAIn36[2] , \wAIn36[1] , \wAIn36[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid91[31] , \wAMid91[30] , \wAMid91[29] , \wAMid91[28] , 
        \wAMid91[27] , \wAMid91[26] , \wAMid91[25] , \wAMid91[24] , 
        \wAMid91[23] , \wAMid91[22] , \wAMid91[21] , \wAMid91[20] , 
        \wAMid91[19] , \wAMid91[18] , \wAMid91[17] , \wAMid91[16] , 
        \wAMid91[15] , \wAMid91[14] , \wAMid91[13] , \wAMid91[12] , 
        \wAMid91[11] , \wAMid91[10] , \wAMid91[9] , \wAMid91[8] , \wAMid91[7] , 
        \wAMid91[6] , \wAMid91[5] , \wAMid91[4] , \wAMid91[3] , \wAMid91[2] , 
        \wAMid91[1] , \wAMid91[0] }), .BIn({\wBMid91[31] , \wBMid91[30] , 
        \wBMid91[29] , \wBMid91[28] , \wBMid91[27] , \wBMid91[26] , 
        \wBMid91[25] , \wBMid91[24] , \wBMid91[23] , \wBMid91[22] , 
        \wBMid91[21] , \wBMid91[20] , \wBMid91[19] , \wBMid91[18] , 
        \wBMid91[17] , \wBMid91[16] , \wBMid91[15] , \wBMid91[14] , 
        \wBMid91[13] , \wBMid91[12] , \wBMid91[11] , \wBMid91[10] , 
        \wBMid91[9] , \wBMid91[8] , \wBMid91[7] , \wBMid91[6] , \wBMid91[5] , 
        \wBMid91[4] , \wBMid91[3] , \wBMid91[2] , \wBMid91[1] , \wBMid91[0] }), 
        .HiOut({\wRegInB91[31] , \wRegInB91[30] , \wRegInB91[29] , 
        \wRegInB91[28] , \wRegInB91[27] , \wRegInB91[26] , \wRegInB91[25] , 
        \wRegInB91[24] , \wRegInB91[23] , \wRegInB91[22] , \wRegInB91[21] , 
        \wRegInB91[20] , \wRegInB91[19] , \wRegInB91[18] , \wRegInB91[17] , 
        \wRegInB91[16] , \wRegInB91[15] , \wRegInB91[14] , \wRegInB91[13] , 
        \wRegInB91[12] , \wRegInB91[11] , \wRegInB91[10] , \wRegInB91[9] , 
        \wRegInB91[8] , \wRegInB91[7] , \wRegInB91[6] , \wRegInB91[5] , 
        \wRegInB91[4] , \wRegInB91[3] , \wRegInB91[2] , \wRegInB91[1] , 
        \wRegInB91[0] }), .LoOut({\wRegInA92[31] , \wRegInA92[30] , 
        \wRegInA92[29] , \wRegInA92[28] , \wRegInA92[27] , \wRegInA92[26] , 
        \wRegInA92[25] , \wRegInA92[24] , \wRegInA92[23] , \wRegInA92[22] , 
        \wRegInA92[21] , \wRegInA92[20] , \wRegInA92[19] , \wRegInA92[18] , 
        \wRegInA92[17] , \wRegInA92[16] , \wRegInA92[15] , \wRegInA92[14] , 
        \wRegInA92[13] , \wRegInA92[12] , \wRegInA92[11] , \wRegInA92[10] , 
        \wRegInA92[9] , \wRegInA92[8] , \wRegInA92[7] , \wRegInA92[6] , 
        \wRegInA92[5] , \wRegInA92[4] , \wRegInA92[3] , \wRegInA92[2] , 
        \wRegInA92[1] , \wRegInA92[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn1[31] , 
        \wAIn1[30] , \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , \wAIn1[26] , 
        \wAIn1[25] , \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , \wAIn1[21] , 
        \wAIn1[20] , \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , \wAIn1[16] , 
        \wAIn1[15] , \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , \wAIn1[11] , 
        \wAIn1[10] , \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , \wAIn1[6] , 
        \wAIn1[5] , \wAIn1[4] , \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , \wAIn1[0] 
        }), .BIn({\wBIn1[31] , \wBIn1[30] , \wBIn1[29] , \wBIn1[28] , 
        \wBIn1[27] , \wBIn1[26] , \wBIn1[25] , \wBIn1[24] , \wBIn1[23] , 
        \wBIn1[22] , \wBIn1[21] , \wBIn1[20] , \wBIn1[19] , \wBIn1[18] , 
        \wBIn1[17] , \wBIn1[16] , \wBIn1[15] , \wBIn1[14] , \wBIn1[13] , 
        \wBIn1[12] , \wBIn1[11] , \wBIn1[10] , \wBIn1[9] , \wBIn1[8] , 
        \wBIn1[7] , \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , \wBIn1[3] , \wBIn1[2] , 
        \wBIn1[1] , \wBIn1[0] }), .HiOut({\wBMid0[31] , \wBMid0[30] , 
        \wBMid0[29] , \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , 
        \wBMid0[24] , \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , 
        \wBMid0[19] , \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , 
        \wBMid0[14] , \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , 
        \wBMid0[9] , \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , 
        \wBMid0[4] , \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), 
        .LoOut({\wAMid1[31] , \wAMid1[30] , \wAMid1[29] , \wAMid1[28] , 
        \wAMid1[27] , \wAMid1[26] , \wAMid1[25] , \wAMid1[24] , \wAMid1[23] , 
        \wAMid1[22] , \wAMid1[21] , \wAMid1[20] , \wAMid1[19] , \wAMid1[18] , 
        \wAMid1[17] , \wAMid1[16] , \wAMid1[15] , \wAMid1[14] , \wAMid1[13] , 
        \wAMid1[12] , \wAMid1[11] , \wAMid1[10] , \wAMid1[9] , \wAMid1[8] , 
        \wAMid1[7] , \wAMid1[6] , \wAMid1[5] , \wAMid1[4] , \wAMid1[3] , 
        \wAMid1[2] , \wAMid1[1] , \wAMid1[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn8[31] , 
        \wAIn8[30] , \wAIn8[29] , \wAIn8[28] , \wAIn8[27] , \wAIn8[26] , 
        \wAIn8[25] , \wAIn8[24] , \wAIn8[23] , \wAIn8[22] , \wAIn8[21] , 
        \wAIn8[20] , \wAIn8[19] , \wAIn8[18] , \wAIn8[17] , \wAIn8[16] , 
        \wAIn8[15] , \wAIn8[14] , \wAIn8[13] , \wAIn8[12] , \wAIn8[11] , 
        \wAIn8[10] , \wAIn8[9] , \wAIn8[8] , \wAIn8[7] , \wAIn8[6] , 
        \wAIn8[5] , \wAIn8[4] , \wAIn8[3] , \wAIn8[2] , \wAIn8[1] , \wAIn8[0] 
        }), .BIn({\wBIn8[31] , \wBIn8[30] , \wBIn8[29] , \wBIn8[28] , 
        \wBIn8[27] , \wBIn8[26] , \wBIn8[25] , \wBIn8[24] , \wBIn8[23] , 
        \wBIn8[22] , \wBIn8[21] , \wBIn8[20] , \wBIn8[19] , \wBIn8[18] , 
        \wBIn8[17] , \wBIn8[16] , \wBIn8[15] , \wBIn8[14] , \wBIn8[13] , 
        \wBIn8[12] , \wBIn8[11] , \wBIn8[10] , \wBIn8[9] , \wBIn8[8] , 
        \wBIn8[7] , \wBIn8[6] , \wBIn8[5] , \wBIn8[4] , \wBIn8[3] , \wBIn8[2] , 
        \wBIn8[1] , \wBIn8[0] }), .HiOut({\wBMid7[31] , \wBMid7[30] , 
        \wBMid7[29] , \wBMid7[28] , \wBMid7[27] , \wBMid7[26] , \wBMid7[25] , 
        \wBMid7[24] , \wBMid7[23] , \wBMid7[22] , \wBMid7[21] , \wBMid7[20] , 
        \wBMid7[19] , \wBMid7[18] , \wBMid7[17] , \wBMid7[16] , \wBMid7[15] , 
        \wBMid7[14] , \wBMid7[13] , \wBMid7[12] , \wBMid7[11] , \wBMid7[10] , 
        \wBMid7[9] , \wBMid7[8] , \wBMid7[7] , \wBMid7[6] , \wBMid7[5] , 
        \wBMid7[4] , \wBMid7[3] , \wBMid7[2] , \wBMid7[1] , \wBMid7[0] }), 
        .LoOut({\wAMid8[31] , \wAMid8[30] , \wAMid8[29] , \wAMid8[28] , 
        \wAMid8[27] , \wAMid8[26] , \wAMid8[25] , \wAMid8[24] , \wAMid8[23] , 
        \wAMid8[22] , \wAMid8[21] , \wAMid8[20] , \wAMid8[19] , \wAMid8[18] , 
        \wAMid8[17] , \wAMid8[16] , \wAMid8[15] , \wAMid8[14] , \wAMid8[13] , 
        \wAMid8[12] , \wAMid8[11] , \wAMid8[10] , \wAMid8[9] , \wAMid8[8] , 
        \wAMid8[7] , \wAMid8[6] , \wAMid8[5] , \wAMid8[4] , \wAMid8[3] , 
        \wAMid8[2] , \wAMid8[1] , \wAMid8[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid99[31] , \wAMid99[30] , \wAMid99[29] , \wAMid99[28] , 
        \wAMid99[27] , \wAMid99[26] , \wAMid99[25] , \wAMid99[24] , 
        \wAMid99[23] , \wAMid99[22] , \wAMid99[21] , \wAMid99[20] , 
        \wAMid99[19] , \wAMid99[18] , \wAMid99[17] , \wAMid99[16] , 
        \wAMid99[15] , \wAMid99[14] , \wAMid99[13] , \wAMid99[12] , 
        \wAMid99[11] , \wAMid99[10] , \wAMid99[9] , \wAMid99[8] , \wAMid99[7] , 
        \wAMid99[6] , \wAMid99[5] , \wAMid99[4] , \wAMid99[3] , \wAMid99[2] , 
        \wAMid99[1] , \wAMid99[0] }), .BIn({\wBMid99[31] , \wBMid99[30] , 
        \wBMid99[29] , \wBMid99[28] , \wBMid99[27] , \wBMid99[26] , 
        \wBMid99[25] , \wBMid99[24] , \wBMid99[23] , \wBMid99[22] , 
        \wBMid99[21] , \wBMid99[20] , \wBMid99[19] , \wBMid99[18] , 
        \wBMid99[17] , \wBMid99[16] , \wBMid99[15] , \wBMid99[14] , 
        \wBMid99[13] , \wBMid99[12] , \wBMid99[11] , \wBMid99[10] , 
        \wBMid99[9] , \wBMid99[8] , \wBMid99[7] , \wBMid99[6] , \wBMid99[5] , 
        \wBMid99[4] , \wBMid99[3] , \wBMid99[2] , \wBMid99[1] , \wBMid99[0] }), 
        .HiOut({\wRegInB99[31] , \wRegInB99[30] , \wRegInB99[29] , 
        \wRegInB99[28] , \wRegInB99[27] , \wRegInB99[26] , \wRegInB99[25] , 
        \wRegInB99[24] , \wRegInB99[23] , \wRegInB99[22] , \wRegInB99[21] , 
        \wRegInB99[20] , \wRegInB99[19] , \wRegInB99[18] , \wRegInB99[17] , 
        \wRegInB99[16] , \wRegInB99[15] , \wRegInB99[14] , \wRegInB99[13] , 
        \wRegInB99[12] , \wRegInB99[11] , \wRegInB99[10] , \wRegInB99[9] , 
        \wRegInB99[8] , \wRegInB99[7] , \wRegInB99[6] , \wRegInB99[5] , 
        \wRegInB99[4] , \wRegInB99[3] , \wRegInB99[2] , \wRegInB99[1] , 
        \wRegInB99[0] }), .LoOut({\wRegInA100[31] , \wRegInA100[30] , 
        \wRegInA100[29] , \wRegInA100[28] , \wRegInA100[27] , \wRegInA100[26] , 
        \wRegInA100[25] , \wRegInA100[24] , \wRegInA100[23] , \wRegInA100[22] , 
        \wRegInA100[21] , \wRegInA100[20] , \wRegInA100[19] , \wRegInA100[18] , 
        \wRegInA100[17] , \wRegInA100[16] , \wRegInA100[15] , \wRegInA100[14] , 
        \wRegInA100[13] , \wRegInA100[12] , \wRegInA100[11] , \wRegInA100[10] , 
        \wRegInA100[9] , \wRegInA100[8] , \wRegInA100[7] , \wRegInA100[6] , 
        \wRegInA100[5] , \wRegInA100[4] , \wRegInA100[3] , \wRegInA100[2] , 
        \wRegInA100[1] , \wRegInA100[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_238 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink239[31] , \ScanLink239[30] , \ScanLink239[29] , 
        \ScanLink239[28] , \ScanLink239[27] , \ScanLink239[26] , 
        \ScanLink239[25] , \ScanLink239[24] , \ScanLink239[23] , 
        \ScanLink239[22] , \ScanLink239[21] , \ScanLink239[20] , 
        \ScanLink239[19] , \ScanLink239[18] , \ScanLink239[17] , 
        \ScanLink239[16] , \ScanLink239[15] , \ScanLink239[14] , 
        \ScanLink239[13] , \ScanLink239[12] , \ScanLink239[11] , 
        \ScanLink239[10] , \ScanLink239[9] , \ScanLink239[8] , 
        \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , \ScanLink239[4] , 
        \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , \ScanLink239[0] 
        }), .ScanOut({\ScanLink238[31] , \ScanLink238[30] , \ScanLink238[29] , 
        \ScanLink238[28] , \ScanLink238[27] , \ScanLink238[26] , 
        \ScanLink238[25] , \ScanLink238[24] , \ScanLink238[23] , 
        \ScanLink238[22] , \ScanLink238[21] , \ScanLink238[20] , 
        \ScanLink238[19] , \ScanLink238[18] , \ScanLink238[17] , 
        \ScanLink238[16] , \ScanLink238[15] , \ScanLink238[14] , 
        \ScanLink238[13] , \ScanLink238[12] , \ScanLink238[11] , 
        \ScanLink238[10] , \ScanLink238[9] , \ScanLink238[8] , 
        \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , \ScanLink238[4] , 
        \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , \ScanLink238[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB8[31] , \wRegInB8[30] , \wRegInB8[29] , \wRegInB8[28] , 
        \wRegInB8[27] , \wRegInB8[26] , \wRegInB8[25] , \wRegInB8[24] , 
        \wRegInB8[23] , \wRegInB8[22] , \wRegInB8[21] , \wRegInB8[20] , 
        \wRegInB8[19] , \wRegInB8[18] , \wRegInB8[17] , \wRegInB8[16] , 
        \wRegInB8[15] , \wRegInB8[14] , \wRegInB8[13] , \wRegInB8[12] , 
        \wRegInB8[11] , \wRegInB8[10] , \wRegInB8[9] , \wRegInB8[8] , 
        \wRegInB8[7] , \wRegInB8[6] , \wRegInB8[5] , \wRegInB8[4] , 
        \wRegInB8[3] , \wRegInB8[2] , \wRegInB8[1] , \wRegInB8[0] }), .Out({
        \wBIn8[31] , \wBIn8[30] , \wBIn8[29] , \wBIn8[28] , \wBIn8[27] , 
        \wBIn8[26] , \wBIn8[25] , \wBIn8[24] , \wBIn8[23] , \wBIn8[22] , 
        \wBIn8[21] , \wBIn8[20] , \wBIn8[19] , \wBIn8[18] , \wBIn8[17] , 
        \wBIn8[16] , \wBIn8[15] , \wBIn8[14] , \wBIn8[13] , \wBIn8[12] , 
        \wBIn8[11] , \wBIn8[10] , \wBIn8[9] , \wBIn8[8] , \wBIn8[7] , 
        \wBIn8[6] , \wBIn8[5] , \wBIn8[4] , \wBIn8[3] , \wBIn8[2] , \wBIn8[1] , 
        \wBIn8[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_108 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink109[31] , \ScanLink109[30] , \ScanLink109[29] , 
        \ScanLink109[28] , \ScanLink109[27] , \ScanLink109[26] , 
        \ScanLink109[25] , \ScanLink109[24] , \ScanLink109[23] , 
        \ScanLink109[22] , \ScanLink109[21] , \ScanLink109[20] , 
        \ScanLink109[19] , \ScanLink109[18] , \ScanLink109[17] , 
        \ScanLink109[16] , \ScanLink109[15] , \ScanLink109[14] , 
        \ScanLink109[13] , \ScanLink109[12] , \ScanLink109[11] , 
        \ScanLink109[10] , \ScanLink109[9] , \ScanLink109[8] , 
        \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , \ScanLink109[4] , 
        \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , \ScanLink109[0] 
        }), .ScanOut({\ScanLink108[31] , \ScanLink108[30] , \ScanLink108[29] , 
        \ScanLink108[28] , \ScanLink108[27] , \ScanLink108[26] , 
        \ScanLink108[25] , \ScanLink108[24] , \ScanLink108[23] , 
        \ScanLink108[22] , \ScanLink108[21] , \ScanLink108[20] , 
        \ScanLink108[19] , \ScanLink108[18] , \ScanLink108[17] , 
        \ScanLink108[16] , \ScanLink108[15] , \ScanLink108[14] , 
        \ScanLink108[13] , \ScanLink108[12] , \ScanLink108[11] , 
        \ScanLink108[10] , \ScanLink108[9] , \ScanLink108[8] , 
        \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , \ScanLink108[4] , 
        \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , \ScanLink108[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB73[31] , \wRegInB73[30] , \wRegInB73[29] , 
        \wRegInB73[28] , \wRegInB73[27] , \wRegInB73[26] , \wRegInB73[25] , 
        \wRegInB73[24] , \wRegInB73[23] , \wRegInB73[22] , \wRegInB73[21] , 
        \wRegInB73[20] , \wRegInB73[19] , \wRegInB73[18] , \wRegInB73[17] , 
        \wRegInB73[16] , \wRegInB73[15] , \wRegInB73[14] , \wRegInB73[13] , 
        \wRegInB73[12] , \wRegInB73[11] , \wRegInB73[10] , \wRegInB73[9] , 
        \wRegInB73[8] , \wRegInB73[7] , \wRegInB73[6] , \wRegInB73[5] , 
        \wRegInB73[4] , \wRegInB73[3] , \wRegInB73[2] , \wRegInB73[1] , 
        \wRegInB73[0] }), .Out({\wBIn73[31] , \wBIn73[30] , \wBIn73[29] , 
        \wBIn73[28] , \wBIn73[27] , \wBIn73[26] , \wBIn73[25] , \wBIn73[24] , 
        \wBIn73[23] , \wBIn73[22] , \wBIn73[21] , \wBIn73[20] , \wBIn73[19] , 
        \wBIn73[18] , \wBIn73[17] , \wBIn73[16] , \wBIn73[15] , \wBIn73[14] , 
        \wBIn73[13] , \wBIn73[12] , \wBIn73[11] , \wBIn73[10] , \wBIn73[9] , 
        \wBIn73[8] , \wBIn73[7] , \wBIn73[6] , \wBIn73[5] , \wBIn73[4] , 
        \wBIn73[3] , \wBIn73[2] , \wBIn73[1] , \wBIn73[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_58 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink59[31] , \ScanLink59[30] , \ScanLink59[29] , 
        \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , \ScanLink59[25] , 
        \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , \ScanLink59[21] , 
        \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , \ScanLink59[17] , 
        \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , \ScanLink59[13] , 
        \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , \ScanLink59[9] , 
        \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , \ScanLink59[5] , 
        \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , \ScanLink59[1] , 
        \ScanLink59[0] }), .ScanOut({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB98[31] , \wRegInB98[30] , 
        \wRegInB98[29] , \wRegInB98[28] , \wRegInB98[27] , \wRegInB98[26] , 
        \wRegInB98[25] , \wRegInB98[24] , \wRegInB98[23] , \wRegInB98[22] , 
        \wRegInB98[21] , \wRegInB98[20] , \wRegInB98[19] , \wRegInB98[18] , 
        \wRegInB98[17] , \wRegInB98[16] , \wRegInB98[15] , \wRegInB98[14] , 
        \wRegInB98[13] , \wRegInB98[12] , \wRegInB98[11] , \wRegInB98[10] , 
        \wRegInB98[9] , \wRegInB98[8] , \wRegInB98[7] , \wRegInB98[6] , 
        \wRegInB98[5] , \wRegInB98[4] , \wRegInB98[3] , \wRegInB98[2] , 
        \wRegInB98[1] , \wRegInB98[0] }), .Out({\wBIn98[31] , \wBIn98[30] , 
        \wBIn98[29] , \wBIn98[28] , \wBIn98[27] , \wBIn98[26] , \wBIn98[25] , 
        \wBIn98[24] , \wBIn98[23] , \wBIn98[22] , \wBIn98[21] , \wBIn98[20] , 
        \wBIn98[19] , \wBIn98[18] , \wBIn98[17] , \wBIn98[16] , \wBIn98[15] , 
        \wBIn98[14] , \wBIn98[13] , \wBIn98[12] , \wBIn98[11] , \wBIn98[10] , 
        \wBIn98[9] , \wBIn98[8] , \wBIn98[7] , \wBIn98[6] , \wBIn98[5] , 
        \wBIn98[4] , \wBIn98[3] , \wBIn98[2] , \wBIn98[1] , \wBIn98[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn22[31] , \wAIn22[30] , \wAIn22[29] , \wAIn22[28] , \wAIn22[27] , 
        \wAIn22[26] , \wAIn22[25] , \wAIn22[24] , \wAIn22[23] , \wAIn22[22] , 
        \wAIn22[21] , \wAIn22[20] , \wAIn22[19] , \wAIn22[18] , \wAIn22[17] , 
        \wAIn22[16] , \wAIn22[15] , \wAIn22[14] , \wAIn22[13] , \wAIn22[12] , 
        \wAIn22[11] , \wAIn22[10] , \wAIn22[9] , \wAIn22[8] , \wAIn22[7] , 
        \wAIn22[6] , \wAIn22[5] , \wAIn22[4] , \wAIn22[3] , \wAIn22[2] , 
        \wAIn22[1] , \wAIn22[0] }), .BIn({\wBIn22[31] , \wBIn22[30] , 
        \wBIn22[29] , \wBIn22[28] , \wBIn22[27] , \wBIn22[26] , \wBIn22[25] , 
        \wBIn22[24] , \wBIn22[23] , \wBIn22[22] , \wBIn22[21] , \wBIn22[20] , 
        \wBIn22[19] , \wBIn22[18] , \wBIn22[17] , \wBIn22[16] , \wBIn22[15] , 
        \wBIn22[14] , \wBIn22[13] , \wBIn22[12] , \wBIn22[11] , \wBIn22[10] , 
        \wBIn22[9] , \wBIn22[8] , \wBIn22[7] , \wBIn22[6] , \wBIn22[5] , 
        \wBIn22[4] , \wBIn22[3] , \wBIn22[2] , \wBIn22[1] , \wBIn22[0] }), 
        .HiOut({\wBMid21[31] , \wBMid21[30] , \wBMid21[29] , \wBMid21[28] , 
        \wBMid21[27] , \wBMid21[26] , \wBMid21[25] , \wBMid21[24] , 
        \wBMid21[23] , \wBMid21[22] , \wBMid21[21] , \wBMid21[20] , 
        \wBMid21[19] , \wBMid21[18] , \wBMid21[17] , \wBMid21[16] , 
        \wBMid21[15] , \wBMid21[14] , \wBMid21[13] , \wBMid21[12] , 
        \wBMid21[11] , \wBMid21[10] , \wBMid21[9] , \wBMid21[8] , \wBMid21[7] , 
        \wBMid21[6] , \wBMid21[5] , \wBMid21[4] , \wBMid21[3] , \wBMid21[2] , 
        \wBMid21[1] , \wBMid21[0] }), .LoOut({\wAMid22[31] , \wAMid22[30] , 
        \wAMid22[29] , \wAMid22[28] , \wAMid22[27] , \wAMid22[26] , 
        \wAMid22[25] , \wAMid22[24] , \wAMid22[23] , \wAMid22[22] , 
        \wAMid22[21] , \wAMid22[20] , \wAMid22[19] , \wAMid22[18] , 
        \wAMid22[17] , \wAMid22[16] , \wAMid22[15] , \wAMid22[14] , 
        \wAMid22[13] , \wAMid22[12] , \wAMid22[11] , \wAMid22[10] , 
        \wAMid22[9] , \wAMid22[8] , \wAMid22[7] , \wAMid22[6] , \wAMid22[5] , 
        \wAMid22[4] , \wAMid22[3] , \wAMid22[2] , \wAMid22[1] , \wAMid22[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn39[31] , \wAIn39[30] , \wAIn39[29] , \wAIn39[28] , \wAIn39[27] , 
        \wAIn39[26] , \wAIn39[25] , \wAIn39[24] , \wAIn39[23] , \wAIn39[22] , 
        \wAIn39[21] , \wAIn39[20] , \wAIn39[19] , \wAIn39[18] , \wAIn39[17] , 
        \wAIn39[16] , \wAIn39[15] , \wAIn39[14] , \wAIn39[13] , \wAIn39[12] , 
        \wAIn39[11] , \wAIn39[10] , \wAIn39[9] , \wAIn39[8] , \wAIn39[7] , 
        \wAIn39[6] , \wAIn39[5] , \wAIn39[4] , \wAIn39[3] , \wAIn39[2] , 
        \wAIn39[1] , \wAIn39[0] }), .BIn({\wBIn39[31] , \wBIn39[30] , 
        \wBIn39[29] , \wBIn39[28] , \wBIn39[27] , \wBIn39[26] , \wBIn39[25] , 
        \wBIn39[24] , \wBIn39[23] , \wBIn39[22] , \wBIn39[21] , \wBIn39[20] , 
        \wBIn39[19] , \wBIn39[18] , \wBIn39[17] , \wBIn39[16] , \wBIn39[15] , 
        \wBIn39[14] , \wBIn39[13] , \wBIn39[12] , \wBIn39[11] , \wBIn39[10] , 
        \wBIn39[9] , \wBIn39[8] , \wBIn39[7] , \wBIn39[6] , \wBIn39[5] , 
        \wBIn39[4] , \wBIn39[3] , \wBIn39[2] , \wBIn39[1] , \wBIn39[0] }), 
        .HiOut({\wBMid38[31] , \wBMid38[30] , \wBMid38[29] , \wBMid38[28] , 
        \wBMid38[27] , \wBMid38[26] , \wBMid38[25] , \wBMid38[24] , 
        \wBMid38[23] , \wBMid38[22] , \wBMid38[21] , \wBMid38[20] , 
        \wBMid38[19] , \wBMid38[18] , \wBMid38[17] , \wBMid38[16] , 
        \wBMid38[15] , \wBMid38[14] , \wBMid38[13] , \wBMid38[12] , 
        \wBMid38[11] , \wBMid38[10] , \wBMid38[9] , \wBMid38[8] , \wBMid38[7] , 
        \wBMid38[6] , \wBMid38[5] , \wBMid38[4] , \wBMid38[3] , \wBMid38[2] , 
        \wBMid38[1] , \wBMid38[0] }), .LoOut({\wAMid39[31] , \wAMid39[30] , 
        \wAMid39[29] , \wAMid39[28] , \wAMid39[27] , \wAMid39[26] , 
        \wAMid39[25] , \wAMid39[24] , \wAMid39[23] , \wAMid39[22] , 
        \wAMid39[21] , \wAMid39[20] , \wAMid39[19] , \wAMid39[18] , 
        \wAMid39[17] , \wAMid39[16] , \wAMid39[15] , \wAMid39[14] , 
        \wAMid39[13] , \wAMid39[12] , \wAMid39[11] , \wAMid39[10] , 
        \wAMid39[9] , \wAMid39[8] , \wAMid39[7] , \wAMid39[6] , \wAMid39[5] , 
        \wAMid39[4] , \wAMid39[3] , \wAMid39[2] , \wAMid39[1] , \wAMid39[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn57[31] , \wAIn57[30] , \wAIn57[29] , \wAIn57[28] , \wAIn57[27] , 
        \wAIn57[26] , \wAIn57[25] , \wAIn57[24] , \wAIn57[23] , \wAIn57[22] , 
        \wAIn57[21] , \wAIn57[20] , \wAIn57[19] , \wAIn57[18] , \wAIn57[17] , 
        \wAIn57[16] , \wAIn57[15] , \wAIn57[14] , \wAIn57[13] , \wAIn57[12] , 
        \wAIn57[11] , \wAIn57[10] , \wAIn57[9] , \wAIn57[8] , \wAIn57[7] , 
        \wAIn57[6] , \wAIn57[5] , \wAIn57[4] , \wAIn57[3] , \wAIn57[2] , 
        \wAIn57[1] , \wAIn57[0] }), .BIn({\wBIn57[31] , \wBIn57[30] , 
        \wBIn57[29] , \wBIn57[28] , \wBIn57[27] , \wBIn57[26] , \wBIn57[25] , 
        \wBIn57[24] , \wBIn57[23] , \wBIn57[22] , \wBIn57[21] , \wBIn57[20] , 
        \wBIn57[19] , \wBIn57[18] , \wBIn57[17] , \wBIn57[16] , \wBIn57[15] , 
        \wBIn57[14] , \wBIn57[13] , \wBIn57[12] , \wBIn57[11] , \wBIn57[10] , 
        \wBIn57[9] , \wBIn57[8] , \wBIn57[7] , \wBIn57[6] , \wBIn57[5] , 
        \wBIn57[4] , \wBIn57[3] , \wBIn57[2] , \wBIn57[1] , \wBIn57[0] }), 
        .HiOut({\wBMid56[31] , \wBMid56[30] , \wBMid56[29] , \wBMid56[28] , 
        \wBMid56[27] , \wBMid56[26] , \wBMid56[25] , \wBMid56[24] , 
        \wBMid56[23] , \wBMid56[22] , \wBMid56[21] , \wBMid56[20] , 
        \wBMid56[19] , \wBMid56[18] , \wBMid56[17] , \wBMid56[16] , 
        \wBMid56[15] , \wBMid56[14] , \wBMid56[13] , \wBMid56[12] , 
        \wBMid56[11] , \wBMid56[10] , \wBMid56[9] , \wBMid56[8] , \wBMid56[7] , 
        \wBMid56[6] , \wBMid56[5] , \wBMid56[4] , \wBMid56[3] , \wBMid56[2] , 
        \wBMid56[1] , \wBMid56[0] }), .LoOut({\wAMid57[31] , \wAMid57[30] , 
        \wAMid57[29] , \wAMid57[28] , \wAMid57[27] , \wAMid57[26] , 
        \wAMid57[25] , \wAMid57[24] , \wAMid57[23] , \wAMid57[22] , 
        \wAMid57[21] , \wAMid57[20] , \wAMid57[19] , \wAMid57[18] , 
        \wAMid57[17] , \wAMid57[16] , \wAMid57[15] , \wAMid57[14] , 
        \wAMid57[13] , \wAMid57[12] , \wAMid57[11] , \wAMid57[10] , 
        \wAMid57[9] , \wAMid57[8] , \wAMid57[7] , \wAMid57[6] , \wAMid57[5] , 
        \wAMid57[4] , \wAMid57[3] , \wAMid57[2] , \wAMid57[1] , \wAMid57[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn127[31] , \wAIn127[30] , \wAIn127[29] , \wAIn127[28] , 
        \wAIn127[27] , \wAIn127[26] , \wAIn127[25] , \wAIn127[24] , 
        \wAIn127[23] , \wAIn127[22] , \wAIn127[21] , \wAIn127[20] , 
        \wAIn127[19] , \wAIn127[18] , \wAIn127[17] , \wAIn127[16] , 
        \wAIn127[15] , \wAIn127[14] , \wAIn127[13] , \wAIn127[12] , 
        \wAIn127[11] , \wAIn127[10] , \wAIn127[9] , \wAIn127[8] , \wAIn127[7] , 
        \wAIn127[6] , \wAIn127[5] , \wAIn127[4] , \wAIn127[3] , \wAIn127[2] , 
        \wAIn127[1] , \wAIn127[0] }), .BIn({\wBIn127[31] , \wBIn127[30] , 
        \wBIn127[29] , \wBIn127[28] , \wBIn127[27] , \wBIn127[26] , 
        \wBIn127[25] , \wBIn127[24] , \wBIn127[23] , \wBIn127[22] , 
        \wBIn127[21] , \wBIn127[20] , \wBIn127[19] , \wBIn127[18] , 
        \wBIn127[17] , \wBIn127[16] , \wBIn127[15] , \wBIn127[14] , 
        \wBIn127[13] , \wBIn127[12] , \wBIn127[11] , \wBIn127[10] , 
        \wBIn127[9] , \wBIn127[8] , \wBIn127[7] , \wBIn127[6] , \wBIn127[5] , 
        \wBIn127[4] , \wBIn127[3] , \wBIn127[2] , \wBIn127[1] , \wBIn127[0] }), 
        .HiOut({\wBMid126[31] , \wBMid126[30] , \wBMid126[29] , \wBMid126[28] , 
        \wBMid126[27] , \wBMid126[26] , \wBMid126[25] , \wBMid126[24] , 
        \wBMid126[23] , \wBMid126[22] , \wBMid126[21] , \wBMid126[20] , 
        \wBMid126[19] , \wBMid126[18] , \wBMid126[17] , \wBMid126[16] , 
        \wBMid126[15] , \wBMid126[14] , \wBMid126[13] , \wBMid126[12] , 
        \wBMid126[11] , \wBMid126[10] , \wBMid126[9] , \wBMid126[8] , 
        \wBMid126[7] , \wBMid126[6] , \wBMid126[5] , \wBMid126[4] , 
        \wBMid126[3] , \wBMid126[2] , \wBMid126[1] , \wBMid126[0] }), .LoOut({
        \wRegInB127[31] , \wRegInB127[30] , \wRegInB127[29] , \wRegInB127[28] , 
        \wRegInB127[27] , \wRegInB127[26] , \wRegInB127[25] , \wRegInB127[24] , 
        \wRegInB127[23] , \wRegInB127[22] , \wRegInB127[21] , \wRegInB127[20] , 
        \wRegInB127[19] , \wRegInB127[18] , \wRegInB127[17] , \wRegInB127[16] , 
        \wRegInB127[15] , \wRegInB127[14] , \wRegInB127[13] , \wRegInB127[12] , 
        \wRegInB127[11] , \wRegInB127[10] , \wRegInB127[9] , \wRegInB127[8] , 
        \wRegInB127[7] , \wRegInB127[6] , \wRegInB127[5] , \wRegInB127[4] , 
        \wRegInB127[3] , \wRegInB127[2] , \wRegInB127[1] , \wRegInB127[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid12[31] , \wAMid12[30] , \wAMid12[29] , \wAMid12[28] , 
        \wAMid12[27] , \wAMid12[26] , \wAMid12[25] , \wAMid12[24] , 
        \wAMid12[23] , \wAMid12[22] , \wAMid12[21] , \wAMid12[20] , 
        \wAMid12[19] , \wAMid12[18] , \wAMid12[17] , \wAMid12[16] , 
        \wAMid12[15] , \wAMid12[14] , \wAMid12[13] , \wAMid12[12] , 
        \wAMid12[11] , \wAMid12[10] , \wAMid12[9] , \wAMid12[8] , \wAMid12[7] , 
        \wAMid12[6] , \wAMid12[5] , \wAMid12[4] , \wAMid12[3] , \wAMid12[2] , 
        \wAMid12[1] , \wAMid12[0] }), .BIn({\wBMid12[31] , \wBMid12[30] , 
        \wBMid12[29] , \wBMid12[28] , \wBMid12[27] , \wBMid12[26] , 
        \wBMid12[25] , \wBMid12[24] , \wBMid12[23] , \wBMid12[22] , 
        \wBMid12[21] , \wBMid12[20] , \wBMid12[19] , \wBMid12[18] , 
        \wBMid12[17] , \wBMid12[16] , \wBMid12[15] , \wBMid12[14] , 
        \wBMid12[13] , \wBMid12[12] , \wBMid12[11] , \wBMid12[10] , 
        \wBMid12[9] , \wBMid12[8] , \wBMid12[7] , \wBMid12[6] , \wBMid12[5] , 
        \wBMid12[4] , \wBMid12[3] , \wBMid12[2] , \wBMid12[1] , \wBMid12[0] }), 
        .HiOut({\wRegInB12[31] , \wRegInB12[30] , \wRegInB12[29] , 
        \wRegInB12[28] , \wRegInB12[27] , \wRegInB12[26] , \wRegInB12[25] , 
        \wRegInB12[24] , \wRegInB12[23] , \wRegInB12[22] , \wRegInB12[21] , 
        \wRegInB12[20] , \wRegInB12[19] , \wRegInB12[18] , \wRegInB12[17] , 
        \wRegInB12[16] , \wRegInB12[15] , \wRegInB12[14] , \wRegInB12[13] , 
        \wRegInB12[12] , \wRegInB12[11] , \wRegInB12[10] , \wRegInB12[9] , 
        \wRegInB12[8] , \wRegInB12[7] , \wRegInB12[6] , \wRegInB12[5] , 
        \wRegInB12[4] , \wRegInB12[3] , \wRegInB12[2] , \wRegInB12[1] , 
        \wRegInB12[0] }), .LoOut({\wRegInA13[31] , \wRegInA13[30] , 
        \wRegInA13[29] , \wRegInA13[28] , \wRegInA13[27] , \wRegInA13[26] , 
        \wRegInA13[25] , \wRegInA13[24] , \wRegInA13[23] , \wRegInA13[22] , 
        \wRegInA13[21] , \wRegInA13[20] , \wRegInA13[19] , \wRegInA13[18] , 
        \wRegInA13[17] , \wRegInA13[16] , \wRegInA13[15] , \wRegInA13[14] , 
        \wRegInA13[13] , \wRegInA13[12] , \wRegInA13[11] , \wRegInA13[10] , 
        \wRegInA13[9] , \wRegInA13[8] , \wRegInA13[7] , \wRegInA13[6] , 
        \wRegInA13[5] , \wRegInA13[4] , \wRegInA13[3] , \wRegInA13[2] , 
        \wRegInA13[1] , \wRegInA13[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid35[31] , \wAMid35[30] , \wAMid35[29] , \wAMid35[28] , 
        \wAMid35[27] , \wAMid35[26] , \wAMid35[25] , \wAMid35[24] , 
        \wAMid35[23] , \wAMid35[22] , \wAMid35[21] , \wAMid35[20] , 
        \wAMid35[19] , \wAMid35[18] , \wAMid35[17] , \wAMid35[16] , 
        \wAMid35[15] , \wAMid35[14] , \wAMid35[13] , \wAMid35[12] , 
        \wAMid35[11] , \wAMid35[10] , \wAMid35[9] , \wAMid35[8] , \wAMid35[7] , 
        \wAMid35[6] , \wAMid35[5] , \wAMid35[4] , \wAMid35[3] , \wAMid35[2] , 
        \wAMid35[1] , \wAMid35[0] }), .BIn({\wBMid35[31] , \wBMid35[30] , 
        \wBMid35[29] , \wBMid35[28] , \wBMid35[27] , \wBMid35[26] , 
        \wBMid35[25] , \wBMid35[24] , \wBMid35[23] , \wBMid35[22] , 
        \wBMid35[21] , \wBMid35[20] , \wBMid35[19] , \wBMid35[18] , 
        \wBMid35[17] , \wBMid35[16] , \wBMid35[15] , \wBMid35[14] , 
        \wBMid35[13] , \wBMid35[12] , \wBMid35[11] , \wBMid35[10] , 
        \wBMid35[9] , \wBMid35[8] , \wBMid35[7] , \wBMid35[6] , \wBMid35[5] , 
        \wBMid35[4] , \wBMid35[3] , \wBMid35[2] , \wBMid35[1] , \wBMid35[0] }), 
        .HiOut({\wRegInB35[31] , \wRegInB35[30] , \wRegInB35[29] , 
        \wRegInB35[28] , \wRegInB35[27] , \wRegInB35[26] , \wRegInB35[25] , 
        \wRegInB35[24] , \wRegInB35[23] , \wRegInB35[22] , \wRegInB35[21] , 
        \wRegInB35[20] , \wRegInB35[19] , \wRegInB35[18] , \wRegInB35[17] , 
        \wRegInB35[16] , \wRegInB35[15] , \wRegInB35[14] , \wRegInB35[13] , 
        \wRegInB35[12] , \wRegInB35[11] , \wRegInB35[10] , \wRegInB35[9] , 
        \wRegInB35[8] , \wRegInB35[7] , \wRegInB35[6] , \wRegInB35[5] , 
        \wRegInB35[4] , \wRegInB35[3] , \wRegInB35[2] , \wRegInB35[1] , 
        \wRegInB35[0] }), .LoOut({\wRegInA36[31] , \wRegInA36[30] , 
        \wRegInA36[29] , \wRegInA36[28] , \wRegInA36[27] , \wRegInA36[26] , 
        \wRegInA36[25] , \wRegInA36[24] , \wRegInA36[23] , \wRegInA36[22] , 
        \wRegInA36[21] , \wRegInA36[20] , \wRegInA36[19] , \wRegInA36[18] , 
        \wRegInA36[17] , \wRegInA36[16] , \wRegInA36[15] , \wRegInA36[14] , 
        \wRegInA36[13] , \wRegInA36[12] , \wRegInA36[11] , \wRegInA36[10] , 
        \wRegInA36[9] , \wRegInA36[8] , \wRegInA36[7] , \wRegInA36[6] , 
        \wRegInA36[5] , \wRegInA36[4] , \wRegInA36[3] , \wRegInA36[2] , 
        \wRegInA36[1] , \wRegInA36[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_230 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink231[31] , \ScanLink231[30] , \ScanLink231[29] , 
        \ScanLink231[28] , \ScanLink231[27] , \ScanLink231[26] , 
        \ScanLink231[25] , \ScanLink231[24] , \ScanLink231[23] , 
        \ScanLink231[22] , \ScanLink231[21] , \ScanLink231[20] , 
        \ScanLink231[19] , \ScanLink231[18] , \ScanLink231[17] , 
        \ScanLink231[16] , \ScanLink231[15] , \ScanLink231[14] , 
        \ScanLink231[13] , \ScanLink231[12] , \ScanLink231[11] , 
        \ScanLink231[10] , \ScanLink231[9] , \ScanLink231[8] , 
        \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , \ScanLink231[4] , 
        \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , \ScanLink231[0] 
        }), .ScanOut({\ScanLink230[31] , \ScanLink230[30] , \ScanLink230[29] , 
        \ScanLink230[28] , \ScanLink230[27] , \ScanLink230[26] , 
        \ScanLink230[25] , \ScanLink230[24] , \ScanLink230[23] , 
        \ScanLink230[22] , \ScanLink230[21] , \ScanLink230[20] , 
        \ScanLink230[19] , \ScanLink230[18] , \ScanLink230[17] , 
        \ScanLink230[16] , \ScanLink230[15] , \ScanLink230[14] , 
        \ScanLink230[13] , \ScanLink230[12] , \ScanLink230[11] , 
        \ScanLink230[10] , \ScanLink230[9] , \ScanLink230[8] , 
        \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , \ScanLink230[4] , 
        \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , \ScanLink230[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB12[31] , \wRegInB12[30] , \wRegInB12[29] , 
        \wRegInB12[28] , \wRegInB12[27] , \wRegInB12[26] , \wRegInB12[25] , 
        \wRegInB12[24] , \wRegInB12[23] , \wRegInB12[22] , \wRegInB12[21] , 
        \wRegInB12[20] , \wRegInB12[19] , \wRegInB12[18] , \wRegInB12[17] , 
        \wRegInB12[16] , \wRegInB12[15] , \wRegInB12[14] , \wRegInB12[13] , 
        \wRegInB12[12] , \wRegInB12[11] , \wRegInB12[10] , \wRegInB12[9] , 
        \wRegInB12[8] , \wRegInB12[7] , \wRegInB12[6] , \wRegInB12[5] , 
        \wRegInB12[4] , \wRegInB12[3] , \wRegInB12[2] , \wRegInB12[1] , 
        \wRegInB12[0] }), .Out({\wBIn12[31] , \wBIn12[30] , \wBIn12[29] , 
        \wBIn12[28] , \wBIn12[27] , \wBIn12[26] , \wBIn12[25] , \wBIn12[24] , 
        \wBIn12[23] , \wBIn12[22] , \wBIn12[21] , \wBIn12[20] , \wBIn12[19] , 
        \wBIn12[18] , \wBIn12[17] , \wBIn12[16] , \wBIn12[15] , \wBIn12[14] , 
        \wBIn12[13] , \wBIn12[12] , \wBIn12[11] , \wBIn12[10] , \wBIn12[9] , 
        \wBIn12[8] , \wBIn12[7] , \wBIn12[6] , \wBIn12[5] , \wBIn12[4] , 
        \wBIn12[3] , \wBIn12[2] , \wBIn12[1] , \wBIn12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_217 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink218[31] , \ScanLink218[30] , \ScanLink218[29] , 
        \ScanLink218[28] , \ScanLink218[27] , \ScanLink218[26] , 
        \ScanLink218[25] , \ScanLink218[24] , \ScanLink218[23] , 
        \ScanLink218[22] , \ScanLink218[21] , \ScanLink218[20] , 
        \ScanLink218[19] , \ScanLink218[18] , \ScanLink218[17] , 
        \ScanLink218[16] , \ScanLink218[15] , \ScanLink218[14] , 
        \ScanLink218[13] , \ScanLink218[12] , \ScanLink218[11] , 
        \ScanLink218[10] , \ScanLink218[9] , \ScanLink218[8] , 
        \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , \ScanLink218[4] , 
        \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , \ScanLink218[0] 
        }), .ScanOut({\ScanLink217[31] , \ScanLink217[30] , \ScanLink217[29] , 
        \ScanLink217[28] , \ScanLink217[27] , \ScanLink217[26] , 
        \ScanLink217[25] , \ScanLink217[24] , \ScanLink217[23] , 
        \ScanLink217[22] , \ScanLink217[21] , \ScanLink217[20] , 
        \ScanLink217[19] , \ScanLink217[18] , \ScanLink217[17] , 
        \ScanLink217[16] , \ScanLink217[15] , \ScanLink217[14] , 
        \ScanLink217[13] , \ScanLink217[12] , \ScanLink217[11] , 
        \ScanLink217[10] , \ScanLink217[9] , \ScanLink217[8] , 
        \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , \ScanLink217[4] , 
        \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , \ScanLink217[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA19[31] , \wRegInA19[30] , \wRegInA19[29] , 
        \wRegInA19[28] , \wRegInA19[27] , \wRegInA19[26] , \wRegInA19[25] , 
        \wRegInA19[24] , \wRegInA19[23] , \wRegInA19[22] , \wRegInA19[21] , 
        \wRegInA19[20] , \wRegInA19[19] , \wRegInA19[18] , \wRegInA19[17] , 
        \wRegInA19[16] , \wRegInA19[15] , \wRegInA19[14] , \wRegInA19[13] , 
        \wRegInA19[12] , \wRegInA19[11] , \wRegInA19[10] , \wRegInA19[9] , 
        \wRegInA19[8] , \wRegInA19[7] , \wRegInA19[6] , \wRegInA19[5] , 
        \wRegInA19[4] , \wRegInA19[3] , \wRegInA19[2] , \wRegInA19[1] , 
        \wRegInA19[0] }), .Out({\wAIn19[31] , \wAIn19[30] , \wAIn19[29] , 
        \wAIn19[28] , \wAIn19[27] , \wAIn19[26] , \wAIn19[25] , \wAIn19[24] , 
        \wAIn19[23] , \wAIn19[22] , \wAIn19[21] , \wAIn19[20] , \wAIn19[19] , 
        \wAIn19[18] , \wAIn19[17] , \wAIn19[16] , \wAIn19[15] , \wAIn19[14] , 
        \wAIn19[13] , \wAIn19[12] , \wAIn19[11] , \wAIn19[10] , \wAIn19[9] , 
        \wAIn19[8] , \wAIn19[7] , \wAIn19[6] , \wAIn19[5] , \wAIn19[4] , 
        \wAIn19[3] , \wAIn19[2] , \wAIn19[1] , \wAIn19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_127 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink128[31] , \ScanLink128[30] , \ScanLink128[29] , 
        \ScanLink128[28] , \ScanLink128[27] , \ScanLink128[26] , 
        \ScanLink128[25] , \ScanLink128[24] , \ScanLink128[23] , 
        \ScanLink128[22] , \ScanLink128[21] , \ScanLink128[20] , 
        \ScanLink128[19] , \ScanLink128[18] , \ScanLink128[17] , 
        \ScanLink128[16] , \ScanLink128[15] , \ScanLink128[14] , 
        \ScanLink128[13] , \ScanLink128[12] , \ScanLink128[11] , 
        \ScanLink128[10] , \ScanLink128[9] , \ScanLink128[8] , 
        \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , \ScanLink128[4] , 
        \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , \ScanLink128[0] 
        }), .ScanOut({\ScanLink127[31] , \ScanLink127[30] , \ScanLink127[29] , 
        \ScanLink127[28] , \ScanLink127[27] , \ScanLink127[26] , 
        \ScanLink127[25] , \ScanLink127[24] , \ScanLink127[23] , 
        \ScanLink127[22] , \ScanLink127[21] , \ScanLink127[20] , 
        \ScanLink127[19] , \ScanLink127[18] , \ScanLink127[17] , 
        \ScanLink127[16] , \ScanLink127[15] , \ScanLink127[14] , 
        \ScanLink127[13] , \ScanLink127[12] , \ScanLink127[11] , 
        \ScanLink127[10] , \ScanLink127[9] , \ScanLink127[8] , 
        \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , \ScanLink127[4] , 
        \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , \ScanLink127[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA64[31] , \wRegInA64[30] , \wRegInA64[29] , 
        \wRegInA64[28] , \wRegInA64[27] , \wRegInA64[26] , \wRegInA64[25] , 
        \wRegInA64[24] , \wRegInA64[23] , \wRegInA64[22] , \wRegInA64[21] , 
        \wRegInA64[20] , \wRegInA64[19] , \wRegInA64[18] , \wRegInA64[17] , 
        \wRegInA64[16] , \wRegInA64[15] , \wRegInA64[14] , \wRegInA64[13] , 
        \wRegInA64[12] , \wRegInA64[11] , \wRegInA64[10] , \wRegInA64[9] , 
        \wRegInA64[8] , \wRegInA64[7] , \wRegInA64[6] , \wRegInA64[5] , 
        \wRegInA64[4] , \wRegInA64[3] , \wRegInA64[2] , \wRegInA64[1] , 
        \wRegInA64[0] }), .Out({\wAIn64[31] , \wAIn64[30] , \wAIn64[29] , 
        \wAIn64[28] , \wAIn64[27] , \wAIn64[26] , \wAIn64[25] , \wAIn64[24] , 
        \wAIn64[23] , \wAIn64[22] , \wAIn64[21] , \wAIn64[20] , \wAIn64[19] , 
        \wAIn64[18] , \wAIn64[17] , \wAIn64[16] , \wAIn64[15] , \wAIn64[14] , 
        \wAIn64[13] , \wAIn64[12] , \wAIn64[11] , \wAIn64[10] , \wAIn64[9] , 
        \wAIn64[8] , \wAIn64[7] , \wAIn64[6] , \wAIn64[5] , \wAIn64[4] , 
        \wAIn64[3] , \wAIn64[2] , \wAIn64[1] , \wAIn64[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_77 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink78[31] , \ScanLink78[30] , \ScanLink78[29] , 
        \ScanLink78[28] , \ScanLink78[27] , \ScanLink78[26] , \ScanLink78[25] , 
        \ScanLink78[24] , \ScanLink78[23] , \ScanLink78[22] , \ScanLink78[21] , 
        \ScanLink78[20] , \ScanLink78[19] , \ScanLink78[18] , \ScanLink78[17] , 
        \ScanLink78[16] , \ScanLink78[15] , \ScanLink78[14] , \ScanLink78[13] , 
        \ScanLink78[12] , \ScanLink78[11] , \ScanLink78[10] , \ScanLink78[9] , 
        \ScanLink78[8] , \ScanLink78[7] , \ScanLink78[6] , \ScanLink78[5] , 
        \ScanLink78[4] , \ScanLink78[3] , \ScanLink78[2] , \ScanLink78[1] , 
        \ScanLink78[0] }), .ScanOut({\ScanLink77[31] , \ScanLink77[30] , 
        \ScanLink77[29] , \ScanLink77[28] , \ScanLink77[27] , \ScanLink77[26] , 
        \ScanLink77[25] , \ScanLink77[24] , \ScanLink77[23] , \ScanLink77[22] , 
        \ScanLink77[21] , \ScanLink77[20] , \ScanLink77[19] , \ScanLink77[18] , 
        \ScanLink77[17] , \ScanLink77[16] , \ScanLink77[15] , \ScanLink77[14] , 
        \ScanLink77[13] , \ScanLink77[12] , \ScanLink77[11] , \ScanLink77[10] , 
        \ScanLink77[9] , \ScanLink77[8] , \ScanLink77[7] , \ScanLink77[6] , 
        \ScanLink77[5] , \ScanLink77[4] , \ScanLink77[3] , \ScanLink77[2] , 
        \ScanLink77[1] , \ScanLink77[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA89[31] , \wRegInA89[30] , 
        \wRegInA89[29] , \wRegInA89[28] , \wRegInA89[27] , \wRegInA89[26] , 
        \wRegInA89[25] , \wRegInA89[24] , \wRegInA89[23] , \wRegInA89[22] , 
        \wRegInA89[21] , \wRegInA89[20] , \wRegInA89[19] , \wRegInA89[18] , 
        \wRegInA89[17] , \wRegInA89[16] , \wRegInA89[15] , \wRegInA89[14] , 
        \wRegInA89[13] , \wRegInA89[12] , \wRegInA89[11] , \wRegInA89[10] , 
        \wRegInA89[9] , \wRegInA89[8] , \wRegInA89[7] , \wRegInA89[6] , 
        \wRegInA89[5] , \wRegInA89[4] , \wRegInA89[3] , \wRegInA89[2] , 
        \wRegInA89[1] , \wRegInA89[0] }), .Out({\wAIn89[31] , \wAIn89[30] , 
        \wAIn89[29] , \wAIn89[28] , \wAIn89[27] , \wAIn89[26] , \wAIn89[25] , 
        \wAIn89[24] , \wAIn89[23] , \wAIn89[22] , \wAIn89[21] , \wAIn89[20] , 
        \wAIn89[19] , \wAIn89[18] , \wAIn89[17] , \wAIn89[16] , \wAIn89[15] , 
        \wAIn89[14] , \wAIn89[13] , \wAIn89[12] , \wAIn89[11] , \wAIn89[10] , 
        \wAIn89[9] , \wAIn89[8] , \wAIn89[7] , \wAIn89[6] , \wAIn89[5] , 
        \wAIn89[4] , \wAIn89[3] , \wAIn89[2] , \wAIn89[1] , \wAIn89[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_50 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink51[31] , \ScanLink51[30] , \ScanLink51[29] , 
        \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , \ScanLink51[25] , 
        \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , \ScanLink51[21] , 
        \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , \ScanLink51[17] , 
        \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , \ScanLink51[13] , 
        \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , \ScanLink51[9] , 
        \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , \ScanLink51[5] , 
        \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , \ScanLink51[1] , 
        \ScanLink51[0] }), .ScanOut({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB102[31] , \wRegInB102[30] , 
        \wRegInB102[29] , \wRegInB102[28] , \wRegInB102[27] , \wRegInB102[26] , 
        \wRegInB102[25] , \wRegInB102[24] , \wRegInB102[23] , \wRegInB102[22] , 
        \wRegInB102[21] , \wRegInB102[20] , \wRegInB102[19] , \wRegInB102[18] , 
        \wRegInB102[17] , \wRegInB102[16] , \wRegInB102[15] , \wRegInB102[14] , 
        \wRegInB102[13] , \wRegInB102[12] , \wRegInB102[11] , \wRegInB102[10] , 
        \wRegInB102[9] , \wRegInB102[8] , \wRegInB102[7] , \wRegInB102[6] , 
        \wRegInB102[5] , \wRegInB102[4] , \wRegInB102[3] , \wRegInB102[2] , 
        \wRegInB102[1] , \wRegInB102[0] }), .Out({\wBIn102[31] , \wBIn102[30] , 
        \wBIn102[29] , \wBIn102[28] , \wBIn102[27] , \wBIn102[26] , 
        \wBIn102[25] , \wBIn102[24] , \wBIn102[23] , \wBIn102[22] , 
        \wBIn102[21] , \wBIn102[20] , \wBIn102[19] , \wBIn102[18] , 
        \wBIn102[17] , \wBIn102[16] , \wBIn102[15] , \wBIn102[14] , 
        \wBIn102[13] , \wBIn102[12] , \wBIn102[11] , \wBIn102[10] , 
        \wBIn102[9] , \wBIn102[8] , \wBIn102[7] , \wBIn102[6] , \wBIn102[5] , 
        \wBIn102[4] , \wBIn102[3] , \wBIn102[2] , \wBIn102[1] , \wBIn102[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid111[31] , \wAMid111[30] , \wAMid111[29] , \wAMid111[28] , 
        \wAMid111[27] , \wAMid111[26] , \wAMid111[25] , \wAMid111[24] , 
        \wAMid111[23] , \wAMid111[22] , \wAMid111[21] , \wAMid111[20] , 
        \wAMid111[19] , \wAMid111[18] , \wAMid111[17] , \wAMid111[16] , 
        \wAMid111[15] , \wAMid111[14] , \wAMid111[13] , \wAMid111[12] , 
        \wAMid111[11] , \wAMid111[10] , \wAMid111[9] , \wAMid111[8] , 
        \wAMid111[7] , \wAMid111[6] , \wAMid111[5] , \wAMid111[4] , 
        \wAMid111[3] , \wAMid111[2] , \wAMid111[1] , \wAMid111[0] }), .BIn({
        \wBMid111[31] , \wBMid111[30] , \wBMid111[29] , \wBMid111[28] , 
        \wBMid111[27] , \wBMid111[26] , \wBMid111[25] , \wBMid111[24] , 
        \wBMid111[23] , \wBMid111[22] , \wBMid111[21] , \wBMid111[20] , 
        \wBMid111[19] , \wBMid111[18] , \wBMid111[17] , \wBMid111[16] , 
        \wBMid111[15] , \wBMid111[14] , \wBMid111[13] , \wBMid111[12] , 
        \wBMid111[11] , \wBMid111[10] , \wBMid111[9] , \wBMid111[8] , 
        \wBMid111[7] , \wBMid111[6] , \wBMid111[5] , \wBMid111[4] , 
        \wBMid111[3] , \wBMid111[2] , \wBMid111[1] , \wBMid111[0] }), .HiOut({
        \wRegInB111[31] , \wRegInB111[30] , \wRegInB111[29] , \wRegInB111[28] , 
        \wRegInB111[27] , \wRegInB111[26] , \wRegInB111[25] , \wRegInB111[24] , 
        \wRegInB111[23] , \wRegInB111[22] , \wRegInB111[21] , \wRegInB111[20] , 
        \wRegInB111[19] , \wRegInB111[18] , \wRegInB111[17] , \wRegInB111[16] , 
        \wRegInB111[15] , \wRegInB111[14] , \wRegInB111[13] , \wRegInB111[12] , 
        \wRegInB111[11] , \wRegInB111[10] , \wRegInB111[9] , \wRegInB111[8] , 
        \wRegInB111[7] , \wRegInB111[6] , \wRegInB111[5] , \wRegInB111[4] , 
        \wRegInB111[3] , \wRegInB111[2] , \wRegInB111[1] , \wRegInB111[0] }), 
        .LoOut({\wRegInA112[31] , \wRegInA112[30] , \wRegInA112[29] , 
        \wRegInA112[28] , \wRegInA112[27] , \wRegInA112[26] , \wRegInA112[25] , 
        \wRegInA112[24] , \wRegInA112[23] , \wRegInA112[22] , \wRegInA112[21] , 
        \wRegInA112[20] , \wRegInA112[19] , \wRegInA112[18] , \wRegInA112[17] , 
        \wRegInA112[16] , \wRegInA112[15] , \wRegInA112[14] , \wRegInA112[13] , 
        \wRegInA112[12] , \wRegInA112[11] , \wRegInA112[10] , \wRegInA112[9] , 
        \wRegInA112[8] , \wRegInA112[7] , \wRegInA112[6] , \wRegInA112[5] , 
        \wRegInA112[4] , \wRegInA112[3] , \wRegInA112[2] , \wRegInA112[1] , 
        \wRegInA112[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_149 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink150[31] , \ScanLink150[30] , \ScanLink150[29] , 
        \ScanLink150[28] , \ScanLink150[27] , \ScanLink150[26] , 
        \ScanLink150[25] , \ScanLink150[24] , \ScanLink150[23] , 
        \ScanLink150[22] , \ScanLink150[21] , \ScanLink150[20] , 
        \ScanLink150[19] , \ScanLink150[18] , \ScanLink150[17] , 
        \ScanLink150[16] , \ScanLink150[15] , \ScanLink150[14] , 
        \ScanLink150[13] , \ScanLink150[12] , \ScanLink150[11] , 
        \ScanLink150[10] , \ScanLink150[9] , \ScanLink150[8] , 
        \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , \ScanLink150[4] , 
        \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , \ScanLink150[0] 
        }), .ScanOut({\ScanLink149[31] , \ScanLink149[30] , \ScanLink149[29] , 
        \ScanLink149[28] , \ScanLink149[27] , \ScanLink149[26] , 
        \ScanLink149[25] , \ScanLink149[24] , \ScanLink149[23] , 
        \ScanLink149[22] , \ScanLink149[21] , \ScanLink149[20] , 
        \ScanLink149[19] , \ScanLink149[18] , \ScanLink149[17] , 
        \ScanLink149[16] , \ScanLink149[15] , \ScanLink149[14] , 
        \ScanLink149[13] , \ScanLink149[12] , \ScanLink149[11] , 
        \ScanLink149[10] , \ScanLink149[9] , \ScanLink149[8] , 
        \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , \ScanLink149[4] , 
        \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , \ScanLink149[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA53[31] , \wRegInA53[30] , \wRegInA53[29] , 
        \wRegInA53[28] , \wRegInA53[27] , \wRegInA53[26] , \wRegInA53[25] , 
        \wRegInA53[24] , \wRegInA53[23] , \wRegInA53[22] , \wRegInA53[21] , 
        \wRegInA53[20] , \wRegInA53[19] , \wRegInA53[18] , \wRegInA53[17] , 
        \wRegInA53[16] , \wRegInA53[15] , \wRegInA53[14] , \wRegInA53[13] , 
        \wRegInA53[12] , \wRegInA53[11] , \wRegInA53[10] , \wRegInA53[9] , 
        \wRegInA53[8] , \wRegInA53[7] , \wRegInA53[6] , \wRegInA53[5] , 
        \wRegInA53[4] , \wRegInA53[3] , \wRegInA53[2] , \wRegInA53[1] , 
        \wRegInA53[0] }), .Out({\wAIn53[31] , \wAIn53[30] , \wAIn53[29] , 
        \wAIn53[28] , \wAIn53[27] , \wAIn53[26] , \wAIn53[25] , \wAIn53[24] , 
        \wAIn53[23] , \wAIn53[22] , \wAIn53[21] , \wAIn53[20] , \wAIn53[19] , 
        \wAIn53[18] , \wAIn53[17] , \wAIn53[16] , \wAIn53[15] , \wAIn53[14] , 
        \wAIn53[13] , \wAIn53[12] , \wAIn53[11] , \wAIn53[10] , \wAIn53[9] , 
        \wAIn53[8] , \wAIn53[7] , \wAIn53[6] , \wAIn53[5] , \wAIn53[4] , 
        \wAIn53[3] , \wAIn53[2] , \wAIn53[1] , \wAIn53[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_100 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink101[31] , \ScanLink101[30] , \ScanLink101[29] , 
        \ScanLink101[28] , \ScanLink101[27] , \ScanLink101[26] , 
        \ScanLink101[25] , \ScanLink101[24] , \ScanLink101[23] , 
        \ScanLink101[22] , \ScanLink101[21] , \ScanLink101[20] , 
        \ScanLink101[19] , \ScanLink101[18] , \ScanLink101[17] , 
        \ScanLink101[16] , \ScanLink101[15] , \ScanLink101[14] , 
        \ScanLink101[13] , \ScanLink101[12] , \ScanLink101[11] , 
        \ScanLink101[10] , \ScanLink101[9] , \ScanLink101[8] , 
        \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , \ScanLink101[4] , 
        \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , \ScanLink101[0] 
        }), .ScanOut({\ScanLink100[31] , \ScanLink100[30] , \ScanLink100[29] , 
        \ScanLink100[28] , \ScanLink100[27] , \ScanLink100[26] , 
        \ScanLink100[25] , \ScanLink100[24] , \ScanLink100[23] , 
        \ScanLink100[22] , \ScanLink100[21] , \ScanLink100[20] , 
        \ScanLink100[19] , \ScanLink100[18] , \ScanLink100[17] , 
        \ScanLink100[16] , \ScanLink100[15] , \ScanLink100[14] , 
        \ScanLink100[13] , \ScanLink100[12] , \ScanLink100[11] , 
        \ScanLink100[10] , \ScanLink100[9] , \ScanLink100[8] , 
        \ScanLink100[7] , \ScanLink100[6] , \ScanLink100[5] , \ScanLink100[4] , 
        \ScanLink100[3] , \ScanLink100[2] , \ScanLink100[1] , \ScanLink100[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB77[31] , \wRegInB77[30] , \wRegInB77[29] , 
        \wRegInB77[28] , \wRegInB77[27] , \wRegInB77[26] , \wRegInB77[25] , 
        \wRegInB77[24] , \wRegInB77[23] , \wRegInB77[22] , \wRegInB77[21] , 
        \wRegInB77[20] , \wRegInB77[19] , \wRegInB77[18] , \wRegInB77[17] , 
        \wRegInB77[16] , \wRegInB77[15] , \wRegInB77[14] , \wRegInB77[13] , 
        \wRegInB77[12] , \wRegInB77[11] , \wRegInB77[10] , \wRegInB77[9] , 
        \wRegInB77[8] , \wRegInB77[7] , \wRegInB77[6] , \wRegInB77[5] , 
        \wRegInB77[4] , \wRegInB77[3] , \wRegInB77[2] , \wRegInB77[1] , 
        \wRegInB77[0] }), .Out({\wBIn77[31] , \wBIn77[30] , \wBIn77[29] , 
        \wBIn77[28] , \wBIn77[27] , \wBIn77[26] , \wBIn77[25] , \wBIn77[24] , 
        \wBIn77[23] , \wBIn77[22] , \wBIn77[21] , \wBIn77[20] , \wBIn77[19] , 
        \wBIn77[18] , \wBIn77[17] , \wBIn77[16] , \wBIn77[15] , \wBIn77[14] , 
        \wBIn77[13] , \wBIn77[12] , \wBIn77[11] , \wBIn77[10] , \wBIn77[9] , 
        \wBIn77[8] , \wBIn77[7] , \wBIn77[6] , \wBIn77[5] , \wBIn77[4] , 
        \wBIn77[3] , \wBIn77[2] , \wBIn77[1] , \wBIn77[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_92 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink93[31] , \ScanLink93[30] , \ScanLink93[29] , 
        \ScanLink93[28] , \ScanLink93[27] , \ScanLink93[26] , \ScanLink93[25] , 
        \ScanLink93[24] , \ScanLink93[23] , \ScanLink93[22] , \ScanLink93[21] , 
        \ScanLink93[20] , \ScanLink93[19] , \ScanLink93[18] , \ScanLink93[17] , 
        \ScanLink93[16] , \ScanLink93[15] , \ScanLink93[14] , \ScanLink93[13] , 
        \ScanLink93[12] , \ScanLink93[11] , \ScanLink93[10] , \ScanLink93[9] , 
        \ScanLink93[8] , \ScanLink93[7] , \ScanLink93[6] , \ScanLink93[5] , 
        \ScanLink93[4] , \ScanLink93[3] , \ScanLink93[2] , \ScanLink93[1] , 
        \ScanLink93[0] }), .ScanOut({\ScanLink92[31] , \ScanLink92[30] , 
        \ScanLink92[29] , \ScanLink92[28] , \ScanLink92[27] , \ScanLink92[26] , 
        \ScanLink92[25] , \ScanLink92[24] , \ScanLink92[23] , \ScanLink92[22] , 
        \ScanLink92[21] , \ScanLink92[20] , \ScanLink92[19] , \ScanLink92[18] , 
        \ScanLink92[17] , \ScanLink92[16] , \ScanLink92[15] , \ScanLink92[14] , 
        \ScanLink92[13] , \ScanLink92[12] , \ScanLink92[11] , \ScanLink92[10] , 
        \ScanLink92[9] , \ScanLink92[8] , \ScanLink92[7] , \ScanLink92[6] , 
        \ScanLink92[5] , \ScanLink92[4] , \ScanLink92[3] , \ScanLink92[2] , 
        \ScanLink92[1] , \ScanLink92[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB81[31] , \wRegInB81[30] , 
        \wRegInB81[29] , \wRegInB81[28] , \wRegInB81[27] , \wRegInB81[26] , 
        \wRegInB81[25] , \wRegInB81[24] , \wRegInB81[23] , \wRegInB81[22] , 
        \wRegInB81[21] , \wRegInB81[20] , \wRegInB81[19] , \wRegInB81[18] , 
        \wRegInB81[17] , \wRegInB81[16] , \wRegInB81[15] , \wRegInB81[14] , 
        \wRegInB81[13] , \wRegInB81[12] , \wRegInB81[11] , \wRegInB81[10] , 
        \wRegInB81[9] , \wRegInB81[8] , \wRegInB81[7] , \wRegInB81[6] , 
        \wRegInB81[5] , \wRegInB81[4] , \wRegInB81[3] , \wRegInB81[2] , 
        \wRegInB81[1] , \wRegInB81[0] }), .Out({\wBIn81[31] , \wBIn81[30] , 
        \wBIn81[29] , \wBIn81[28] , \wBIn81[27] , \wBIn81[26] , \wBIn81[25] , 
        \wBIn81[24] , \wBIn81[23] , \wBIn81[22] , \wBIn81[21] , \wBIn81[20] , 
        \wBIn81[19] , \wBIn81[18] , \wBIn81[17] , \wBIn81[16] , \wBIn81[15] , 
        \wBIn81[14] , \wBIn81[13] , \wBIn81[12] , \wBIn81[11] , \wBIn81[10] , 
        \wBIn81[9] , \wBIn81[8] , \wBIn81[7] , \wBIn81[6] , \wBIn81[5] , 
        \wBIn81[4] , \wBIn81[3] , \wBIn81[2] , \wBIn81[1] , \wBIn81[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_19 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink20[31] , \ScanLink20[30] , \ScanLink20[29] , 
        \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , \ScanLink20[25] , 
        \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , \ScanLink20[21] , 
        \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , \ScanLink20[17] , 
        \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , \ScanLink20[13] , 
        \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , \ScanLink20[9] , 
        \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , \ScanLink20[5] , 
        \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , \ScanLink20[1] , 
        \ScanLink20[0] }), .ScanOut({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA118[31] , \wRegInA118[30] , 
        \wRegInA118[29] , \wRegInA118[28] , \wRegInA118[27] , \wRegInA118[26] , 
        \wRegInA118[25] , \wRegInA118[24] , \wRegInA118[23] , \wRegInA118[22] , 
        \wRegInA118[21] , \wRegInA118[20] , \wRegInA118[19] , \wRegInA118[18] , 
        \wRegInA118[17] , \wRegInA118[16] , \wRegInA118[15] , \wRegInA118[14] , 
        \wRegInA118[13] , \wRegInA118[12] , \wRegInA118[11] , \wRegInA118[10] , 
        \wRegInA118[9] , \wRegInA118[8] , \wRegInA118[7] , \wRegInA118[6] , 
        \wRegInA118[5] , \wRegInA118[4] , \wRegInA118[3] , \wRegInA118[2] , 
        \wRegInA118[1] , \wRegInA118[0] }), .Out({\wAIn118[31] , \wAIn118[30] , 
        \wAIn118[29] , \wAIn118[28] , \wAIn118[27] , \wAIn118[26] , 
        \wAIn118[25] , \wAIn118[24] , \wAIn118[23] , \wAIn118[22] , 
        \wAIn118[21] , \wAIn118[20] , \wAIn118[19] , \wAIn118[18] , 
        \wAIn118[17] , \wAIn118[16] , \wAIn118[15] , \wAIn118[14] , 
        \wAIn118[13] , \wAIn118[12] , \wAIn118[11] , \wAIn118[10] , 
        \wAIn118[9] , \wAIn118[8] , \wAIn118[7] , \wAIn118[6] , \wAIn118[5] , 
        \wAIn118[4] , \wAIn118[3] , \wAIn118[2] , \wAIn118[1] , \wAIn118[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_89 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink90[31] , \ScanLink90[30] , \ScanLink90[29] , 
        \ScanLink90[28] , \ScanLink90[27] , \ScanLink90[26] , \ScanLink90[25] , 
        \ScanLink90[24] , \ScanLink90[23] , \ScanLink90[22] , \ScanLink90[21] , 
        \ScanLink90[20] , \ScanLink90[19] , \ScanLink90[18] , \ScanLink90[17] , 
        \ScanLink90[16] , \ScanLink90[15] , \ScanLink90[14] , \ScanLink90[13] , 
        \ScanLink90[12] , \ScanLink90[11] , \ScanLink90[10] , \ScanLink90[9] , 
        \ScanLink90[8] , \ScanLink90[7] , \ScanLink90[6] , \ScanLink90[5] , 
        \ScanLink90[4] , \ScanLink90[3] , \ScanLink90[2] , \ScanLink90[1] , 
        \ScanLink90[0] }), .ScanOut({\ScanLink89[31] , \ScanLink89[30] , 
        \ScanLink89[29] , \ScanLink89[28] , \ScanLink89[27] , \ScanLink89[26] , 
        \ScanLink89[25] , \ScanLink89[24] , \ScanLink89[23] , \ScanLink89[22] , 
        \ScanLink89[21] , \ScanLink89[20] , \ScanLink89[19] , \ScanLink89[18] , 
        \ScanLink89[17] , \ScanLink89[16] , \ScanLink89[15] , \ScanLink89[14] , 
        \ScanLink89[13] , \ScanLink89[12] , \ScanLink89[11] , \ScanLink89[10] , 
        \ScanLink89[9] , \ScanLink89[8] , \ScanLink89[7] , \ScanLink89[6] , 
        \ScanLink89[5] , \ScanLink89[4] , \ScanLink89[3] , \ScanLink89[2] , 
        \ScanLink89[1] , \ScanLink89[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA83[31] , \wRegInA83[30] , 
        \wRegInA83[29] , \wRegInA83[28] , \wRegInA83[27] , \wRegInA83[26] , 
        \wRegInA83[25] , \wRegInA83[24] , \wRegInA83[23] , \wRegInA83[22] , 
        \wRegInA83[21] , \wRegInA83[20] , \wRegInA83[19] , \wRegInA83[18] , 
        \wRegInA83[17] , \wRegInA83[16] , \wRegInA83[15] , \wRegInA83[14] , 
        \wRegInA83[13] , \wRegInA83[12] , \wRegInA83[11] , \wRegInA83[10] , 
        \wRegInA83[9] , \wRegInA83[8] , \wRegInA83[7] , \wRegInA83[6] , 
        \wRegInA83[5] , \wRegInA83[4] , \wRegInA83[3] , \wRegInA83[2] , 
        \wRegInA83[1] , \wRegInA83[0] }), .Out({\wAIn83[31] , \wAIn83[30] , 
        \wAIn83[29] , \wAIn83[28] , \wAIn83[27] , \wAIn83[26] , \wAIn83[25] , 
        \wAIn83[24] , \wAIn83[23] , \wAIn83[22] , \wAIn83[21] , \wAIn83[20] , 
        \wAIn83[19] , \wAIn83[18] , \wAIn83[17] , \wAIn83[16] , \wAIn83[15] , 
        \wAIn83[14] , \wAIn83[13] , \wAIn83[12] , \wAIn83[11] , \wAIn83[10] , 
        \wAIn83[9] , \wAIn83[8] , \wAIn83[7] , \wAIn83[6] , \wAIn83[5] , 
        \wAIn83[4] , \wAIn83[3] , \wAIn83[2] , \wAIn83[1] , \wAIn83[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid67[31] , \wAMid67[30] , \wAMid67[29] , \wAMid67[28] , 
        \wAMid67[27] , \wAMid67[26] , \wAMid67[25] , \wAMid67[24] , 
        \wAMid67[23] , \wAMid67[22] , \wAMid67[21] , \wAMid67[20] , 
        \wAMid67[19] , \wAMid67[18] , \wAMid67[17] , \wAMid67[16] , 
        \wAMid67[15] , \wAMid67[14] , \wAMid67[13] , \wAMid67[12] , 
        \wAMid67[11] , \wAMid67[10] , \wAMid67[9] , \wAMid67[8] , \wAMid67[7] , 
        \wAMid67[6] , \wAMid67[5] , \wAMid67[4] , \wAMid67[3] , \wAMid67[2] , 
        \wAMid67[1] , \wAMid67[0] }), .BIn({\wBMid67[31] , \wBMid67[30] , 
        \wBMid67[29] , \wBMid67[28] , \wBMid67[27] , \wBMid67[26] , 
        \wBMid67[25] , \wBMid67[24] , \wBMid67[23] , \wBMid67[22] , 
        \wBMid67[21] , \wBMid67[20] , \wBMid67[19] , \wBMid67[18] , 
        \wBMid67[17] , \wBMid67[16] , \wBMid67[15] , \wBMid67[14] , 
        \wBMid67[13] , \wBMid67[12] , \wBMid67[11] , \wBMid67[10] , 
        \wBMid67[9] , \wBMid67[8] , \wBMid67[7] , \wBMid67[6] , \wBMid67[5] , 
        \wBMid67[4] , \wBMid67[3] , \wBMid67[2] , \wBMid67[1] , \wBMid67[0] }), 
        .HiOut({\wRegInB67[31] , \wRegInB67[30] , \wRegInB67[29] , 
        \wRegInB67[28] , \wRegInB67[27] , \wRegInB67[26] , \wRegInB67[25] , 
        \wRegInB67[24] , \wRegInB67[23] , \wRegInB67[22] , \wRegInB67[21] , 
        \wRegInB67[20] , \wRegInB67[19] , \wRegInB67[18] , \wRegInB67[17] , 
        \wRegInB67[16] , \wRegInB67[15] , \wRegInB67[14] , \wRegInB67[13] , 
        \wRegInB67[12] , \wRegInB67[11] , \wRegInB67[10] , \wRegInB67[9] , 
        \wRegInB67[8] , \wRegInB67[7] , \wRegInB67[6] , \wRegInB67[5] , 
        \wRegInB67[4] , \wRegInB67[3] , \wRegInB67[2] , \wRegInB67[1] , 
        \wRegInB67[0] }), .LoOut({\wRegInA68[31] , \wRegInA68[30] , 
        \wRegInA68[29] , \wRegInA68[28] , \wRegInA68[27] , \wRegInA68[26] , 
        \wRegInA68[25] , \wRegInA68[24] , \wRegInA68[23] , \wRegInA68[22] , 
        \wRegInA68[21] , \wRegInA68[20] , \wRegInA68[19] , \wRegInA68[18] , 
        \wRegInA68[17] , \wRegInA68[16] , \wRegInA68[15] , \wRegInA68[14] , 
        \wRegInA68[13] , \wRegInA68[12] , \wRegInA68[11] , \wRegInA68[10] , 
        \wRegInA68[9] , \wRegInA68[8] , \wRegInA68[7] , \wRegInA68[6] , 
        \wRegInA68[5] , \wRegInA68[4] , \wRegInA68[3] , \wRegInA68[2] , 
        \wRegInA68[1] , \wRegInA68[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_152 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink153[31] , \ScanLink153[30] , \ScanLink153[29] , 
        \ScanLink153[28] , \ScanLink153[27] , \ScanLink153[26] , 
        \ScanLink153[25] , \ScanLink153[24] , \ScanLink153[23] , 
        \ScanLink153[22] , \ScanLink153[21] , \ScanLink153[20] , 
        \ScanLink153[19] , \ScanLink153[18] , \ScanLink153[17] , 
        \ScanLink153[16] , \ScanLink153[15] , \ScanLink153[14] , 
        \ScanLink153[13] , \ScanLink153[12] , \ScanLink153[11] , 
        \ScanLink153[10] , \ScanLink153[9] , \ScanLink153[8] , 
        \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , \ScanLink153[4] , 
        \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , \ScanLink153[0] 
        }), .ScanOut({\ScanLink152[31] , \ScanLink152[30] , \ScanLink152[29] , 
        \ScanLink152[28] , \ScanLink152[27] , \ScanLink152[26] , 
        \ScanLink152[25] , \ScanLink152[24] , \ScanLink152[23] , 
        \ScanLink152[22] , \ScanLink152[21] , \ScanLink152[20] , 
        \ScanLink152[19] , \ScanLink152[18] , \ScanLink152[17] , 
        \ScanLink152[16] , \ScanLink152[15] , \ScanLink152[14] , 
        \ScanLink152[13] , \ScanLink152[12] , \ScanLink152[11] , 
        \ScanLink152[10] , \ScanLink152[9] , \ScanLink152[8] , 
        \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , \ScanLink152[4] , 
        \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , \ScanLink152[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB51[31] , \wRegInB51[30] , \wRegInB51[29] , 
        \wRegInB51[28] , \wRegInB51[27] , \wRegInB51[26] , \wRegInB51[25] , 
        \wRegInB51[24] , \wRegInB51[23] , \wRegInB51[22] , \wRegInB51[21] , 
        \wRegInB51[20] , \wRegInB51[19] , \wRegInB51[18] , \wRegInB51[17] , 
        \wRegInB51[16] , \wRegInB51[15] , \wRegInB51[14] , \wRegInB51[13] , 
        \wRegInB51[12] , \wRegInB51[11] , \wRegInB51[10] , \wRegInB51[9] , 
        \wRegInB51[8] , \wRegInB51[7] , \wRegInB51[6] , \wRegInB51[5] , 
        \wRegInB51[4] , \wRegInB51[3] , \wRegInB51[2] , \wRegInB51[1] , 
        \wRegInB51[0] }), .Out({\wBIn51[31] , \wBIn51[30] , \wBIn51[29] , 
        \wBIn51[28] , \wBIn51[27] , \wBIn51[26] , \wBIn51[25] , \wBIn51[24] , 
        \wBIn51[23] , \wBIn51[22] , \wBIn51[21] , \wBIn51[20] , \wBIn51[19] , 
        \wBIn51[18] , \wBIn51[17] , \wBIn51[16] , \wBIn51[15] , \wBIn51[14] , 
        \wBIn51[13] , \wBIn51[12] , \wBIn51[11] , \wBIn51[10] , \wBIn51[9] , 
        \wBIn51[8] , \wBIn51[7] , \wBIn51[6] , \wBIn51[5] , \wBIn51[4] , 
        \wBIn51[3] , \wBIn51[2] , \wBIn51[1] , \wBIn51[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn70[31] , \wAIn70[30] , \wAIn70[29] , \wAIn70[28] , \wAIn70[27] , 
        \wAIn70[26] , \wAIn70[25] , \wAIn70[24] , \wAIn70[23] , \wAIn70[22] , 
        \wAIn70[21] , \wAIn70[20] , \wAIn70[19] , \wAIn70[18] , \wAIn70[17] , 
        \wAIn70[16] , \wAIn70[15] , \wAIn70[14] , \wAIn70[13] , \wAIn70[12] , 
        \wAIn70[11] , \wAIn70[10] , \wAIn70[9] , \wAIn70[8] , \wAIn70[7] , 
        \wAIn70[6] , \wAIn70[5] , \wAIn70[4] , \wAIn70[3] , \wAIn70[2] , 
        \wAIn70[1] , \wAIn70[0] }), .BIn({\wBIn70[31] , \wBIn70[30] , 
        \wBIn70[29] , \wBIn70[28] , \wBIn70[27] , \wBIn70[26] , \wBIn70[25] , 
        \wBIn70[24] , \wBIn70[23] , \wBIn70[22] , \wBIn70[21] , \wBIn70[20] , 
        \wBIn70[19] , \wBIn70[18] , \wBIn70[17] , \wBIn70[16] , \wBIn70[15] , 
        \wBIn70[14] , \wBIn70[13] , \wBIn70[12] , \wBIn70[11] , \wBIn70[10] , 
        \wBIn70[9] , \wBIn70[8] , \wBIn70[7] , \wBIn70[6] , \wBIn70[5] , 
        \wBIn70[4] , \wBIn70[3] , \wBIn70[2] , \wBIn70[1] , \wBIn70[0] }), 
        .HiOut({\wBMid69[31] , \wBMid69[30] , \wBMid69[29] , \wBMid69[28] , 
        \wBMid69[27] , \wBMid69[26] , \wBMid69[25] , \wBMid69[24] , 
        \wBMid69[23] , \wBMid69[22] , \wBMid69[21] , \wBMid69[20] , 
        \wBMid69[19] , \wBMid69[18] , \wBMid69[17] , \wBMid69[16] , 
        \wBMid69[15] , \wBMid69[14] , \wBMid69[13] , \wBMid69[12] , 
        \wBMid69[11] , \wBMid69[10] , \wBMid69[9] , \wBMid69[8] , \wBMid69[7] , 
        \wBMid69[6] , \wBMid69[5] , \wBMid69[4] , \wBMid69[3] , \wBMid69[2] , 
        \wBMid69[1] , \wBMid69[0] }), .LoOut({\wAMid70[31] , \wAMid70[30] , 
        \wAMid70[29] , \wAMid70[28] , \wAMid70[27] , \wAMid70[26] , 
        \wAMid70[25] , \wAMid70[24] , \wAMid70[23] , \wAMid70[22] , 
        \wAMid70[21] , \wAMid70[20] , \wAMid70[19] , \wAMid70[18] , 
        \wAMid70[17] , \wAMid70[16] , \wAMid70[15] , \wAMid70[14] , 
        \wAMid70[13] , \wAMid70[12] , \wAMid70[11] , \wAMid70[10] , 
        \wAMid70[9] , \wAMid70[8] , \wAMid70[7] , \wAMid70[6] , \wAMid70[5] , 
        \wAMid70[4] , \wAMid70[3] , \wAMid70[2] , \wAMid70[1] , \wAMid70[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid40[31] , \wAMid40[30] , \wAMid40[29] , \wAMid40[28] , 
        \wAMid40[27] , \wAMid40[26] , \wAMid40[25] , \wAMid40[24] , 
        \wAMid40[23] , \wAMid40[22] , \wAMid40[21] , \wAMid40[20] , 
        \wAMid40[19] , \wAMid40[18] , \wAMid40[17] , \wAMid40[16] , 
        \wAMid40[15] , \wAMid40[14] , \wAMid40[13] , \wAMid40[12] , 
        \wAMid40[11] , \wAMid40[10] , \wAMid40[9] , \wAMid40[8] , \wAMid40[7] , 
        \wAMid40[6] , \wAMid40[5] , \wAMid40[4] , \wAMid40[3] , \wAMid40[2] , 
        \wAMid40[1] , \wAMid40[0] }), .BIn({\wBMid40[31] , \wBMid40[30] , 
        \wBMid40[29] , \wBMid40[28] , \wBMid40[27] , \wBMid40[26] , 
        \wBMid40[25] , \wBMid40[24] , \wBMid40[23] , \wBMid40[22] , 
        \wBMid40[21] , \wBMid40[20] , \wBMid40[19] , \wBMid40[18] , 
        \wBMid40[17] , \wBMid40[16] , \wBMid40[15] , \wBMid40[14] , 
        \wBMid40[13] , \wBMid40[12] , \wBMid40[11] , \wBMid40[10] , 
        \wBMid40[9] , \wBMid40[8] , \wBMid40[7] , \wBMid40[6] , \wBMid40[5] , 
        \wBMid40[4] , \wBMid40[3] , \wBMid40[2] , \wBMid40[1] , \wBMid40[0] }), 
        .HiOut({\wRegInB40[31] , \wRegInB40[30] , \wRegInB40[29] , 
        \wRegInB40[28] , \wRegInB40[27] , \wRegInB40[26] , \wRegInB40[25] , 
        \wRegInB40[24] , \wRegInB40[23] , \wRegInB40[22] , \wRegInB40[21] , 
        \wRegInB40[20] , \wRegInB40[19] , \wRegInB40[18] , \wRegInB40[17] , 
        \wRegInB40[16] , \wRegInB40[15] , \wRegInB40[14] , \wRegInB40[13] , 
        \wRegInB40[12] , \wRegInB40[11] , \wRegInB40[10] , \wRegInB40[9] , 
        \wRegInB40[8] , \wRegInB40[7] , \wRegInB40[6] , \wRegInB40[5] , 
        \wRegInB40[4] , \wRegInB40[3] , \wRegInB40[2] , \wRegInB40[1] , 
        \wRegInB40[0] }), .LoOut({\wRegInA41[31] , \wRegInA41[30] , 
        \wRegInA41[29] , \wRegInA41[28] , \wRegInA41[27] , \wRegInA41[26] , 
        \wRegInA41[25] , \wRegInA41[24] , \wRegInA41[23] , \wRegInA41[22] , 
        \wRegInA41[21] , \wRegInA41[20] , \wRegInA41[19] , \wRegInA41[18] , 
        \wRegInA41[17] , \wRegInA41[16] , \wRegInA41[15] , \wRegInA41[14] , 
        \wRegInA41[13] , \wRegInA41[12] , \wRegInA41[11] , \wRegInA41[10] , 
        \wRegInA41[9] , \wRegInA41[8] , \wRegInA41[7] , \wRegInA41[6] , 
        \wRegInA41[5] , \wRegInA41[4] , \wRegInA41[3] , \wRegInA41[2] , 
        \wRegInA41[1] , \wRegInA41[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_25 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink26[31] , \ScanLink26[30] , \ScanLink26[29] , 
        \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , \ScanLink26[25] , 
        \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , \ScanLink26[21] , 
        \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , \ScanLink26[17] , 
        \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , \ScanLink26[13] , 
        \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , \ScanLink26[9] , 
        \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , \ScanLink26[5] , 
        \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , \ScanLink26[1] , 
        \ScanLink26[0] }), .ScanOut({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA115[31] , \wRegInA115[30] , 
        \wRegInA115[29] , \wRegInA115[28] , \wRegInA115[27] , \wRegInA115[26] , 
        \wRegInA115[25] , \wRegInA115[24] , \wRegInA115[23] , \wRegInA115[22] , 
        \wRegInA115[21] , \wRegInA115[20] , \wRegInA115[19] , \wRegInA115[18] , 
        \wRegInA115[17] , \wRegInA115[16] , \wRegInA115[15] , \wRegInA115[14] , 
        \wRegInA115[13] , \wRegInA115[12] , \wRegInA115[11] , \wRegInA115[10] , 
        \wRegInA115[9] , \wRegInA115[8] , \wRegInA115[7] , \wRegInA115[6] , 
        \wRegInA115[5] , \wRegInA115[4] , \wRegInA115[3] , \wRegInA115[2] , 
        \wRegInA115[1] , \wRegInA115[0] }), .Out({\wAIn115[31] , \wAIn115[30] , 
        \wAIn115[29] , \wAIn115[28] , \wAIn115[27] , \wAIn115[26] , 
        \wAIn115[25] , \wAIn115[24] , \wAIn115[23] , \wAIn115[22] , 
        \wAIn115[21] , \wAIn115[20] , \wAIn115[19] , \wAIn115[18] , 
        \wAIn115[17] , \wAIn115[16] , \wAIn115[15] , \wAIn115[14] , 
        \wAIn115[13] , \wAIn115[12] , \wAIn115[11] , \wAIn115[10] , 
        \wAIn115[9] , \wAIn115[8] , \wAIn115[7] , \wAIn115[6] , \wAIn115[5] , 
        \wAIn115[4] , \wAIn115[3] , \wAIn115[2] , \wAIn115[1] , \wAIn115[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_175 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink176[31] , \ScanLink176[30] , \ScanLink176[29] , 
        \ScanLink176[28] , \ScanLink176[27] , \ScanLink176[26] , 
        \ScanLink176[25] , \ScanLink176[24] , \ScanLink176[23] , 
        \ScanLink176[22] , \ScanLink176[21] , \ScanLink176[20] , 
        \ScanLink176[19] , \ScanLink176[18] , \ScanLink176[17] , 
        \ScanLink176[16] , \ScanLink176[15] , \ScanLink176[14] , 
        \ScanLink176[13] , \ScanLink176[12] , \ScanLink176[11] , 
        \ScanLink176[10] , \ScanLink176[9] , \ScanLink176[8] , 
        \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , \ScanLink176[4] , 
        \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , \ScanLink176[0] 
        }), .ScanOut({\ScanLink175[31] , \ScanLink175[30] , \ScanLink175[29] , 
        \ScanLink175[28] , \ScanLink175[27] , \ScanLink175[26] , 
        \ScanLink175[25] , \ScanLink175[24] , \ScanLink175[23] , 
        \ScanLink175[22] , \ScanLink175[21] , \ScanLink175[20] , 
        \ScanLink175[19] , \ScanLink175[18] , \ScanLink175[17] , 
        \ScanLink175[16] , \ScanLink175[15] , \ScanLink175[14] , 
        \ScanLink175[13] , \ScanLink175[12] , \ScanLink175[11] , 
        \ScanLink175[10] , \ScanLink175[9] , \ScanLink175[8] , 
        \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , \ScanLink175[4] , 
        \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , \ScanLink175[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA40[31] , \wRegInA40[30] , \wRegInA40[29] , 
        \wRegInA40[28] , \wRegInA40[27] , \wRegInA40[26] , \wRegInA40[25] , 
        \wRegInA40[24] , \wRegInA40[23] , \wRegInA40[22] , \wRegInA40[21] , 
        \wRegInA40[20] , \wRegInA40[19] , \wRegInA40[18] , \wRegInA40[17] , 
        \wRegInA40[16] , \wRegInA40[15] , \wRegInA40[14] , \wRegInA40[13] , 
        \wRegInA40[12] , \wRegInA40[11] , \wRegInA40[10] , \wRegInA40[9] , 
        \wRegInA40[8] , \wRegInA40[7] , \wRegInA40[6] , \wRegInA40[5] , 
        \wRegInA40[4] , \wRegInA40[3] , \wRegInA40[2] , \wRegInA40[1] , 
        \wRegInA40[0] }), .Out({\wAIn40[31] , \wAIn40[30] , \wAIn40[29] , 
        \wAIn40[28] , \wAIn40[27] , \wAIn40[26] , \wAIn40[25] , \wAIn40[24] , 
        \wAIn40[23] , \wAIn40[22] , \wAIn40[21] , \wAIn40[20] , \wAIn40[19] , 
        \wAIn40[18] , \wAIn40[17] , \wAIn40[16] , \wAIn40[15] , \wAIn40[14] , 
        \wAIn40[13] , \wAIn40[12] , \wAIn40[11] , \wAIn40[10] , \wAIn40[9] , 
        \wAIn40[8] , \wAIn40[7] , \wAIn40[6] , \wAIn40[5] , \wAIn40[4] , 
        \wAIn40[3] , \wAIn40[2] , \wAIn40[1] , \wAIn40[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn100[31] , \wAIn100[30] , \wAIn100[29] , \wAIn100[28] , 
        \wAIn100[27] , \wAIn100[26] , \wAIn100[25] , \wAIn100[24] , 
        \wAIn100[23] , \wAIn100[22] , \wAIn100[21] , \wAIn100[20] , 
        \wAIn100[19] , \wAIn100[18] , \wAIn100[17] , \wAIn100[16] , 
        \wAIn100[15] , \wAIn100[14] , \wAIn100[13] , \wAIn100[12] , 
        \wAIn100[11] , \wAIn100[10] , \wAIn100[9] , \wAIn100[8] , \wAIn100[7] , 
        \wAIn100[6] , \wAIn100[5] , \wAIn100[4] , \wAIn100[3] , \wAIn100[2] , 
        \wAIn100[1] , \wAIn100[0] }), .BIn({\wBIn100[31] , \wBIn100[30] , 
        \wBIn100[29] , \wBIn100[28] , \wBIn100[27] , \wBIn100[26] , 
        \wBIn100[25] , \wBIn100[24] , \wBIn100[23] , \wBIn100[22] , 
        \wBIn100[21] , \wBIn100[20] , \wBIn100[19] , \wBIn100[18] , 
        \wBIn100[17] , \wBIn100[16] , \wBIn100[15] , \wBIn100[14] , 
        \wBIn100[13] , \wBIn100[12] , \wBIn100[11] , \wBIn100[10] , 
        \wBIn100[9] , \wBIn100[8] , \wBIn100[7] , \wBIn100[6] , \wBIn100[5] , 
        \wBIn100[4] , \wBIn100[3] , \wBIn100[2] , \wBIn100[1] , \wBIn100[0] }), 
        .HiOut({\wBMid99[31] , \wBMid99[30] , \wBMid99[29] , \wBMid99[28] , 
        \wBMid99[27] , \wBMid99[26] , \wBMid99[25] , \wBMid99[24] , 
        \wBMid99[23] , \wBMid99[22] , \wBMid99[21] , \wBMid99[20] , 
        \wBMid99[19] , \wBMid99[18] , \wBMid99[17] , \wBMid99[16] , 
        \wBMid99[15] , \wBMid99[14] , \wBMid99[13] , \wBMid99[12] , 
        \wBMid99[11] , \wBMid99[10] , \wBMid99[9] , \wBMid99[8] , \wBMid99[7] , 
        \wBMid99[6] , \wBMid99[5] , \wBMid99[4] , \wBMid99[3] , \wBMid99[2] , 
        \wBMid99[1] , \wBMid99[0] }), .LoOut({\wAMid100[31] , \wAMid100[30] , 
        \wAMid100[29] , \wAMid100[28] , \wAMid100[27] , \wAMid100[26] , 
        \wAMid100[25] , \wAMid100[24] , \wAMid100[23] , \wAMid100[22] , 
        \wAMid100[21] , \wAMid100[20] , \wAMid100[19] , \wAMid100[18] , 
        \wAMid100[17] , \wAMid100[16] , \wAMid100[15] , \wAMid100[14] , 
        \wAMid100[13] , \wAMid100[12] , \wAMid100[11] , \wAMid100[10] , 
        \wAMid100[9] , \wAMid100[8] , \wAMid100[7] , \wAMid100[6] , 
        \wAMid100[5] , \wAMid100[4] , \wAMid100[3] , \wAMid100[2] , 
        \wAMid100[1] , \wAMid100[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_245 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink246[31] , \ScanLink246[30] , \ScanLink246[29] , 
        \ScanLink246[28] , \ScanLink246[27] , \ScanLink246[26] , 
        \ScanLink246[25] , \ScanLink246[24] , \ScanLink246[23] , 
        \ScanLink246[22] , \ScanLink246[21] , \ScanLink246[20] , 
        \ScanLink246[19] , \ScanLink246[18] , \ScanLink246[17] , 
        \ScanLink246[16] , \ScanLink246[15] , \ScanLink246[14] , 
        \ScanLink246[13] , \ScanLink246[12] , \ScanLink246[11] , 
        \ScanLink246[10] , \ScanLink246[9] , \ScanLink246[8] , 
        \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , \ScanLink246[4] , 
        \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , \ScanLink246[0] 
        }), .ScanOut({\ScanLink245[31] , \ScanLink245[30] , \ScanLink245[29] , 
        \ScanLink245[28] , \ScanLink245[27] , \ScanLink245[26] , 
        \ScanLink245[25] , \ScanLink245[24] , \ScanLink245[23] , 
        \ScanLink245[22] , \ScanLink245[21] , \ScanLink245[20] , 
        \ScanLink245[19] , \ScanLink245[18] , \ScanLink245[17] , 
        \ScanLink245[16] , \ScanLink245[15] , \ScanLink245[14] , 
        \ScanLink245[13] , \ScanLink245[12] , \ScanLink245[11] , 
        \ScanLink245[10] , \ScanLink245[9] , \ScanLink245[8] , 
        \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , \ScanLink245[4] , 
        \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , \ScanLink245[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA5[31] , \wRegInA5[30] , \wRegInA5[29] , \wRegInA5[28] , 
        \wRegInA5[27] , \wRegInA5[26] , \wRegInA5[25] , \wRegInA5[24] , 
        \wRegInA5[23] , \wRegInA5[22] , \wRegInA5[21] , \wRegInA5[20] , 
        \wRegInA5[19] , \wRegInA5[18] , \wRegInA5[17] , \wRegInA5[16] , 
        \wRegInA5[15] , \wRegInA5[14] , \wRegInA5[13] , \wRegInA5[12] , 
        \wRegInA5[11] , \wRegInA5[10] , \wRegInA5[9] , \wRegInA5[8] , 
        \wRegInA5[7] , \wRegInA5[6] , \wRegInA5[5] , \wRegInA5[4] , 
        \wRegInA5[3] , \wRegInA5[2] , \wRegInA5[1] , \wRegInA5[0] }), .Out({
        \wAIn5[31] , \wAIn5[30] , \wAIn5[29] , \wAIn5[28] , \wAIn5[27] , 
        \wAIn5[26] , \wAIn5[25] , \wAIn5[24] , \wAIn5[23] , \wAIn5[22] , 
        \wAIn5[21] , \wAIn5[20] , \wAIn5[19] , \wAIn5[18] , \wAIn5[17] , 
        \wAIn5[16] , \wAIn5[15] , \wAIn5[14] , \wAIn5[13] , \wAIn5[12] , 
        \wAIn5[11] , \wAIn5[10] , \wAIn5[9] , \wAIn5[8] , \wAIn5[7] , 
        \wAIn5[6] , \wAIn5[5] , \wAIn5[4] , \wAIn5[3] , \wAIn5[2] , \wAIn5[1] , 
        \wAIn5[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_8 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[31] , \ScanLink9[30] , \ScanLink9[29] , 
        \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , \ScanLink9[25] , 
        \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , \ScanLink9[21] , 
        \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , \ScanLink9[17] , 
        \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , \ScanLink9[13] , 
        \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , \ScanLink9[9] , 
        \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB123[31] , \wRegInB123[30] , 
        \wRegInB123[29] , \wRegInB123[28] , \wRegInB123[27] , \wRegInB123[26] , 
        \wRegInB123[25] , \wRegInB123[24] , \wRegInB123[23] , \wRegInB123[22] , 
        \wRegInB123[21] , \wRegInB123[20] , \wRegInB123[19] , \wRegInB123[18] , 
        \wRegInB123[17] , \wRegInB123[16] , \wRegInB123[15] , \wRegInB123[14] , 
        \wRegInB123[13] , \wRegInB123[12] , \wRegInB123[11] , \wRegInB123[10] , 
        \wRegInB123[9] , \wRegInB123[8] , \wRegInB123[7] , \wRegInB123[6] , 
        \wRegInB123[5] , \wRegInB123[4] , \wRegInB123[3] , \wRegInB123[2] , 
        \wRegInB123[1] , \wRegInB123[0] }), .Out({\wBIn123[31] , \wBIn123[30] , 
        \wBIn123[29] , \wBIn123[28] , \wBIn123[27] , \wBIn123[26] , 
        \wBIn123[25] , \wBIn123[24] , \wBIn123[23] , \wBIn123[22] , 
        \wBIn123[21] , \wBIn123[20] , \wBIn123[19] , \wBIn123[18] , 
        \wBIn123[17] , \wBIn123[16] , \wBIn123[15] , \wBIn123[14] , 
        \wBIn123[13] , \wBIn123[12] , \wBIn123[11] , \wBIn123[10] , 
        \wBIn123[9] , \wBIn123[8] , \wBIn123[7] , \wBIn123[6] , \wBIn123[5] , 
        \wBIn123[4] , \wBIn123[3] , \wBIn123[2] , \wBIn123[1] , \wBIn123[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn87[31] , \wAIn87[30] , \wAIn87[29] , \wAIn87[28] , \wAIn87[27] , 
        \wAIn87[26] , \wAIn87[25] , \wAIn87[24] , \wAIn87[23] , \wAIn87[22] , 
        \wAIn87[21] , \wAIn87[20] , \wAIn87[19] , \wAIn87[18] , \wAIn87[17] , 
        \wAIn87[16] , \wAIn87[15] , \wAIn87[14] , \wAIn87[13] , \wAIn87[12] , 
        \wAIn87[11] , \wAIn87[10] , \wAIn87[9] , \wAIn87[8] , \wAIn87[7] , 
        \wAIn87[6] , \wAIn87[5] , \wAIn87[4] , \wAIn87[3] , \wAIn87[2] , 
        \wAIn87[1] , \wAIn87[0] }), .BIn({\wBIn87[31] , \wBIn87[30] , 
        \wBIn87[29] , \wBIn87[28] , \wBIn87[27] , \wBIn87[26] , \wBIn87[25] , 
        \wBIn87[24] , \wBIn87[23] , \wBIn87[22] , \wBIn87[21] , \wBIn87[20] , 
        \wBIn87[19] , \wBIn87[18] , \wBIn87[17] , \wBIn87[16] , \wBIn87[15] , 
        \wBIn87[14] , \wBIn87[13] , \wBIn87[12] , \wBIn87[11] , \wBIn87[10] , 
        \wBIn87[9] , \wBIn87[8] , \wBIn87[7] , \wBIn87[6] , \wBIn87[5] , 
        \wBIn87[4] , \wBIn87[3] , \wBIn87[2] , \wBIn87[1] , \wBIn87[0] }), 
        .HiOut({\wBMid86[31] , \wBMid86[30] , \wBMid86[29] , \wBMid86[28] , 
        \wBMid86[27] , \wBMid86[26] , \wBMid86[25] , \wBMid86[24] , 
        \wBMid86[23] , \wBMid86[22] , \wBMid86[21] , \wBMid86[20] , 
        \wBMid86[19] , \wBMid86[18] , \wBMid86[17] , \wBMid86[16] , 
        \wBMid86[15] , \wBMid86[14] , \wBMid86[13] , \wBMid86[12] , 
        \wBMid86[11] , \wBMid86[10] , \wBMid86[9] , \wBMid86[8] , \wBMid86[7] , 
        \wBMid86[6] , \wBMid86[5] , \wBMid86[4] , \wBMid86[3] , \wBMid86[2] , 
        \wBMid86[1] , \wBMid86[0] }), .LoOut({\wAMid87[31] , \wAMid87[30] , 
        \wAMid87[29] , \wAMid87[28] , \wAMid87[27] , \wAMid87[26] , 
        \wAMid87[25] , \wAMid87[24] , \wAMid87[23] , \wAMid87[22] , 
        \wAMid87[21] , \wAMid87[20] , \wAMid87[19] , \wAMid87[18] , 
        \wAMid87[17] , \wAMid87[16] , \wAMid87[15] , \wAMid87[14] , 
        \wAMid87[13] , \wAMid87[12] , \wAMid87[11] , \wAMid87[10] , 
        \wAMid87[9] , \wAMid87[8] , \wAMid87[7] , \wAMid87[6] , \wAMid87[5] , 
        \wAMid87[4] , \wAMid87[3] , \wAMid87[2] , \wAMid87[1] , \wAMid87[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn95[31] , \wAIn95[30] , \wAIn95[29] , \wAIn95[28] , \wAIn95[27] , 
        \wAIn95[26] , \wAIn95[25] , \wAIn95[24] , \wAIn95[23] , \wAIn95[22] , 
        \wAIn95[21] , \wAIn95[20] , \wAIn95[19] , \wAIn95[18] , \wAIn95[17] , 
        \wAIn95[16] , \wAIn95[15] , \wAIn95[14] , \wAIn95[13] , \wAIn95[12] , 
        \wAIn95[11] , \wAIn95[10] , \wAIn95[9] , \wAIn95[8] , \wAIn95[7] , 
        \wAIn95[6] , \wAIn95[5] , \wAIn95[4] , \wAIn95[3] , \wAIn95[2] , 
        \wAIn95[1] , \wAIn95[0] }), .BIn({\wBIn95[31] , \wBIn95[30] , 
        \wBIn95[29] , \wBIn95[28] , \wBIn95[27] , \wBIn95[26] , \wBIn95[25] , 
        \wBIn95[24] , \wBIn95[23] , \wBIn95[22] , \wBIn95[21] , \wBIn95[20] , 
        \wBIn95[19] , \wBIn95[18] , \wBIn95[17] , \wBIn95[16] , \wBIn95[15] , 
        \wBIn95[14] , \wBIn95[13] , \wBIn95[12] , \wBIn95[11] , \wBIn95[10] , 
        \wBIn95[9] , \wBIn95[8] , \wBIn95[7] , \wBIn95[6] , \wBIn95[5] , 
        \wBIn95[4] , \wBIn95[3] , \wBIn95[2] , \wBIn95[1] , \wBIn95[0] }), 
        .HiOut({\wBMid94[31] , \wBMid94[30] , \wBMid94[29] , \wBMid94[28] , 
        \wBMid94[27] , \wBMid94[26] , \wBMid94[25] , \wBMid94[24] , 
        \wBMid94[23] , \wBMid94[22] , \wBMid94[21] , \wBMid94[20] , 
        \wBMid94[19] , \wBMid94[18] , \wBMid94[17] , \wBMid94[16] , 
        \wBMid94[15] , \wBMid94[14] , \wBMid94[13] , \wBMid94[12] , 
        \wBMid94[11] , \wBMid94[10] , \wBMid94[9] , \wBMid94[8] , \wBMid94[7] , 
        \wBMid94[6] , \wBMid94[5] , \wBMid94[4] , \wBMid94[3] , \wBMid94[2] , 
        \wBMid94[1] , \wBMid94[0] }), .LoOut({\wAMid95[31] , \wAMid95[30] , 
        \wAMid95[29] , \wAMid95[28] , \wAMid95[27] , \wAMid95[26] , 
        \wAMid95[25] , \wAMid95[24] , \wAMid95[23] , \wAMid95[22] , 
        \wAMid95[21] , \wAMid95[20] , \wAMid95[19] , \wAMid95[18] , 
        \wAMid95[17] , \wAMid95[16] , \wAMid95[15] , \wAMid95[14] , 
        \wAMid95[13] , \wAMid95[12] , \wAMid95[11] , \wAMid95[10] , 
        \wAMid95[9] , \wAMid95[8] , \wAMid95[7] , \wAMid95[6] , \wAMid95[5] , 
        \wAMid95[4] , \wAMid95[3] , \wAMid95[2] , \wAMid95[1] , \wAMid95[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid4[31] , 
        \wAMid4[30] , \wAMid4[29] , \wAMid4[28] , \wAMid4[27] , \wAMid4[26] , 
        \wAMid4[25] , \wAMid4[24] , \wAMid4[23] , \wAMid4[22] , \wAMid4[21] , 
        \wAMid4[20] , \wAMid4[19] , \wAMid4[18] , \wAMid4[17] , \wAMid4[16] , 
        \wAMid4[15] , \wAMid4[14] , \wAMid4[13] , \wAMid4[12] , \wAMid4[11] , 
        \wAMid4[10] , \wAMid4[9] , \wAMid4[8] , \wAMid4[7] , \wAMid4[6] , 
        \wAMid4[5] , \wAMid4[4] , \wAMid4[3] , \wAMid4[2] , \wAMid4[1] , 
        \wAMid4[0] }), .BIn({\wBMid4[31] , \wBMid4[30] , \wBMid4[29] , 
        \wBMid4[28] , \wBMid4[27] , \wBMid4[26] , \wBMid4[25] , \wBMid4[24] , 
        \wBMid4[23] , \wBMid4[22] , \wBMid4[21] , \wBMid4[20] , \wBMid4[19] , 
        \wBMid4[18] , \wBMid4[17] , \wBMid4[16] , \wBMid4[15] , \wBMid4[14] , 
        \wBMid4[13] , \wBMid4[12] , \wBMid4[11] , \wBMid4[10] , \wBMid4[9] , 
        \wBMid4[8] , \wBMid4[7] , \wBMid4[6] , \wBMid4[5] , \wBMid4[4] , 
        \wBMid4[3] , \wBMid4[2] , \wBMid4[1] , \wBMid4[0] }), .HiOut({
        \wRegInB4[31] , \wRegInB4[30] , \wRegInB4[29] , \wRegInB4[28] , 
        \wRegInB4[27] , \wRegInB4[26] , \wRegInB4[25] , \wRegInB4[24] , 
        \wRegInB4[23] , \wRegInB4[22] , \wRegInB4[21] , \wRegInB4[20] , 
        \wRegInB4[19] , \wRegInB4[18] , \wRegInB4[17] , \wRegInB4[16] , 
        \wRegInB4[15] , \wRegInB4[14] , \wRegInB4[13] , \wRegInB4[12] , 
        \wRegInB4[11] , \wRegInB4[10] , \wRegInB4[9] , \wRegInB4[8] , 
        \wRegInB4[7] , \wRegInB4[6] , \wRegInB4[5] , \wRegInB4[4] , 
        \wRegInB4[3] , \wRegInB4[2] , \wRegInB4[1] , \wRegInB4[0] }), .LoOut({
        \wRegInA5[31] , \wRegInA5[30] , \wRegInA5[29] , \wRegInA5[28] , 
        \wRegInA5[27] , \wRegInA5[26] , \wRegInA5[25] , \wRegInA5[24] , 
        \wRegInA5[23] , \wRegInA5[22] , \wRegInA5[21] , \wRegInA5[20] , 
        \wRegInA5[19] , \wRegInA5[18] , \wRegInA5[17] , \wRegInA5[16] , 
        \wRegInA5[15] , \wRegInA5[14] , \wRegInA5[13] , \wRegInA5[12] , 
        \wRegInA5[11] , \wRegInA5[10] , \wRegInA5[9] , \wRegInA5[8] , 
        \wRegInA5[7] , \wRegInA5[6] , \wRegInA5[5] , \wRegInA5[4] , 
        \wRegInA5[3] , \wRegInA5[2] , \wRegInA5[1] , \wRegInA5[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_190 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink191[31] , \ScanLink191[30] , \ScanLink191[29] , 
        \ScanLink191[28] , \ScanLink191[27] , \ScanLink191[26] , 
        \ScanLink191[25] , \ScanLink191[24] , \ScanLink191[23] , 
        \ScanLink191[22] , \ScanLink191[21] , \ScanLink191[20] , 
        \ScanLink191[19] , \ScanLink191[18] , \ScanLink191[17] , 
        \ScanLink191[16] , \ScanLink191[15] , \ScanLink191[14] , 
        \ScanLink191[13] , \ScanLink191[12] , \ScanLink191[11] , 
        \ScanLink191[10] , \ScanLink191[9] , \ScanLink191[8] , 
        \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , \ScanLink191[4] , 
        \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , \ScanLink191[0] 
        }), .ScanOut({\ScanLink190[31] , \ScanLink190[30] , \ScanLink190[29] , 
        \ScanLink190[28] , \ScanLink190[27] , \ScanLink190[26] , 
        \ScanLink190[25] , \ScanLink190[24] , \ScanLink190[23] , 
        \ScanLink190[22] , \ScanLink190[21] , \ScanLink190[20] , 
        \ScanLink190[19] , \ScanLink190[18] , \ScanLink190[17] , 
        \ScanLink190[16] , \ScanLink190[15] , \ScanLink190[14] , 
        \ScanLink190[13] , \ScanLink190[12] , \ScanLink190[11] , 
        \ScanLink190[10] , \ScanLink190[9] , \ScanLink190[8] , 
        \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , \ScanLink190[4] , 
        \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , \ScanLink190[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB32[31] , \wRegInB32[30] , \wRegInB32[29] , 
        \wRegInB32[28] , \wRegInB32[27] , \wRegInB32[26] , \wRegInB32[25] , 
        \wRegInB32[24] , \wRegInB32[23] , \wRegInB32[22] , \wRegInB32[21] , 
        \wRegInB32[20] , \wRegInB32[19] , \wRegInB32[18] , \wRegInB32[17] , 
        \wRegInB32[16] , \wRegInB32[15] , \wRegInB32[14] , \wRegInB32[13] , 
        \wRegInB32[12] , \wRegInB32[11] , \wRegInB32[10] , \wRegInB32[9] , 
        \wRegInB32[8] , \wRegInB32[7] , \wRegInB32[6] , \wRegInB32[5] , 
        \wRegInB32[4] , \wRegInB32[3] , \wRegInB32[2] , \wRegInB32[1] , 
        \wRegInB32[0] }), .Out({\wBIn32[31] , \wBIn32[30] , \wBIn32[29] , 
        \wBIn32[28] , \wBIn32[27] , \wBIn32[26] , \wBIn32[25] , \wBIn32[24] , 
        \wBIn32[23] , \wBIn32[22] , \wBIn32[21] , \wBIn32[20] , \wBIn32[19] , 
        \wBIn32[18] , \wBIn32[17] , \wBIn32[16] , \wBIn32[15] , \wBIn32[14] , 
        \wBIn32[13] , \wBIn32[12] , \wBIn32[11] , \wBIn32[10] , \wBIn32[9] , 
        \wBIn32[8] , \wBIn32[7] , \wBIn32[6] , \wBIn32[5] , \wBIn32[4] , 
        \wBIn32[3] , \wBIn32[2] , \wBIn32[1] , \wBIn32[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid82[31] , \wAMid82[30] , \wAMid82[29] , \wAMid82[28] , 
        \wAMid82[27] , \wAMid82[26] , \wAMid82[25] , \wAMid82[24] , 
        \wAMid82[23] , \wAMid82[22] , \wAMid82[21] , \wAMid82[20] , 
        \wAMid82[19] , \wAMid82[18] , \wAMid82[17] , \wAMid82[16] , 
        \wAMid82[15] , \wAMid82[14] , \wAMid82[13] , \wAMid82[12] , 
        \wAMid82[11] , \wAMid82[10] , \wAMid82[9] , \wAMid82[8] , \wAMid82[7] , 
        \wAMid82[6] , \wAMid82[5] , \wAMid82[4] , \wAMid82[3] , \wAMid82[2] , 
        \wAMid82[1] , \wAMid82[0] }), .BIn({\wBMid82[31] , \wBMid82[30] , 
        \wBMid82[29] , \wBMid82[28] , \wBMid82[27] , \wBMid82[26] , 
        \wBMid82[25] , \wBMid82[24] , \wBMid82[23] , \wBMid82[22] , 
        \wBMid82[21] , \wBMid82[20] , \wBMid82[19] , \wBMid82[18] , 
        \wBMid82[17] , \wBMid82[16] , \wBMid82[15] , \wBMid82[14] , 
        \wBMid82[13] , \wBMid82[12] , \wBMid82[11] , \wBMid82[10] , 
        \wBMid82[9] , \wBMid82[8] , \wBMid82[7] , \wBMid82[6] , \wBMid82[5] , 
        \wBMid82[4] , \wBMid82[3] , \wBMid82[2] , \wBMid82[1] , \wBMid82[0] }), 
        .HiOut({\wRegInB82[31] , \wRegInB82[30] , \wRegInB82[29] , 
        \wRegInB82[28] , \wRegInB82[27] , \wRegInB82[26] , \wRegInB82[25] , 
        \wRegInB82[24] , \wRegInB82[23] , \wRegInB82[22] , \wRegInB82[21] , 
        \wRegInB82[20] , \wRegInB82[19] , \wRegInB82[18] , \wRegInB82[17] , 
        \wRegInB82[16] , \wRegInB82[15] , \wRegInB82[14] , \wRegInB82[13] , 
        \wRegInB82[12] , \wRegInB82[11] , \wRegInB82[10] , \wRegInB82[9] , 
        \wRegInB82[8] , \wRegInB82[7] , \wRegInB82[6] , \wRegInB82[5] , 
        \wRegInB82[4] , \wRegInB82[3] , \wRegInB82[2] , \wRegInB82[1] , 
        \wRegInB82[0] }), .LoOut({\wRegInA83[31] , \wRegInA83[30] , 
        \wRegInA83[29] , \wRegInA83[28] , \wRegInA83[27] , \wRegInA83[26] , 
        \wRegInA83[25] , \wRegInA83[24] , \wRegInA83[23] , \wRegInA83[22] , 
        \wRegInA83[21] , \wRegInA83[20] , \wRegInA83[19] , \wRegInA83[18] , 
        \wRegInA83[17] , \wRegInA83[16] , \wRegInA83[15] , \wRegInA83[14] , 
        \wRegInA83[13] , \wRegInA83[12] , \wRegInA83[11] , \wRegInA83[10] , 
        \wRegInA83[9] , \wRegInA83[8] , \wRegInA83[7] , \wRegInA83[6] , 
        \wRegInA83[5] , \wRegInA83[4] , \wRegInA83[3] , \wRegInA83[2] , 
        \wRegInA83[1] , \wRegInA83[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_182 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink183[31] , \ScanLink183[30] , \ScanLink183[29] , 
        \ScanLink183[28] , \ScanLink183[27] , \ScanLink183[26] , 
        \ScanLink183[25] , \ScanLink183[24] , \ScanLink183[23] , 
        \ScanLink183[22] , \ScanLink183[21] , \ScanLink183[20] , 
        \ScanLink183[19] , \ScanLink183[18] , \ScanLink183[17] , 
        \ScanLink183[16] , \ScanLink183[15] , \ScanLink183[14] , 
        \ScanLink183[13] , \ScanLink183[12] , \ScanLink183[11] , 
        \ScanLink183[10] , \ScanLink183[9] , \ScanLink183[8] , 
        \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , \ScanLink183[4] , 
        \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , \ScanLink183[0] 
        }), .ScanOut({\ScanLink182[31] , \ScanLink182[30] , \ScanLink182[29] , 
        \ScanLink182[28] , \ScanLink182[27] , \ScanLink182[26] , 
        \ScanLink182[25] , \ScanLink182[24] , \ScanLink182[23] , 
        \ScanLink182[22] , \ScanLink182[21] , \ScanLink182[20] , 
        \ScanLink182[19] , \ScanLink182[18] , \ScanLink182[17] , 
        \ScanLink182[16] , \ScanLink182[15] , \ScanLink182[14] , 
        \ScanLink182[13] , \ScanLink182[12] , \ScanLink182[11] , 
        \ScanLink182[10] , \ScanLink182[9] , \ScanLink182[8] , 
        \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , \ScanLink182[4] , 
        \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , \ScanLink182[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB36[31] , \wRegInB36[30] , \wRegInB36[29] , 
        \wRegInB36[28] , \wRegInB36[27] , \wRegInB36[26] , \wRegInB36[25] , 
        \wRegInB36[24] , \wRegInB36[23] , \wRegInB36[22] , \wRegInB36[21] , 
        \wRegInB36[20] , \wRegInB36[19] , \wRegInB36[18] , \wRegInB36[17] , 
        \wRegInB36[16] , \wRegInB36[15] , \wRegInB36[14] , \wRegInB36[13] , 
        \wRegInB36[12] , \wRegInB36[11] , \wRegInB36[10] , \wRegInB36[9] , 
        \wRegInB36[8] , \wRegInB36[7] , \wRegInB36[6] , \wRegInB36[5] , 
        \wRegInB36[4] , \wRegInB36[3] , \wRegInB36[2] , \wRegInB36[1] , 
        \wRegInB36[0] }), .Out({\wBIn36[31] , \wBIn36[30] , \wBIn36[29] , 
        \wBIn36[28] , \wBIn36[27] , \wBIn36[26] , \wBIn36[25] , \wBIn36[24] , 
        \wBIn36[23] , \wBIn36[22] , \wBIn36[21] , \wBIn36[20] , \wBIn36[19] , 
        \wBIn36[18] , \wBIn36[17] , \wBIn36[16] , \wBIn36[15] , \wBIn36[14] , 
        \wBIn36[13] , \wBIn36[12] , \wBIn36[11] , \wBIn36[10] , \wBIn36[9] , 
        \wBIn36[8] , \wBIn36[7] , \wBIn36[6] , \wBIn36[5] , \wBIn36[4] , 
        \wBIn36[3] , \wBIn36[2] , \wBIn36[1] , \wBIn36[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn6[31] , 
        \wAIn6[30] , \wAIn6[29] , \wAIn6[28] , \wAIn6[27] , \wAIn6[26] , 
        \wAIn6[25] , \wAIn6[24] , \wAIn6[23] , \wAIn6[22] , \wAIn6[21] , 
        \wAIn6[20] , \wAIn6[19] , \wAIn6[18] , \wAIn6[17] , \wAIn6[16] , 
        \wAIn6[15] , \wAIn6[14] , \wAIn6[13] , \wAIn6[12] , \wAIn6[11] , 
        \wAIn6[10] , \wAIn6[9] , \wAIn6[8] , \wAIn6[7] , \wAIn6[6] , 
        \wAIn6[5] , \wAIn6[4] , \wAIn6[3] , \wAIn6[2] , \wAIn6[1] , \wAIn6[0] 
        }), .BIn({\wBIn6[31] , \wBIn6[30] , \wBIn6[29] , \wBIn6[28] , 
        \wBIn6[27] , \wBIn6[26] , \wBIn6[25] , \wBIn6[24] , \wBIn6[23] , 
        \wBIn6[22] , \wBIn6[21] , \wBIn6[20] , \wBIn6[19] , \wBIn6[18] , 
        \wBIn6[17] , \wBIn6[16] , \wBIn6[15] , \wBIn6[14] , \wBIn6[13] , 
        \wBIn6[12] , \wBIn6[11] , \wBIn6[10] , \wBIn6[9] , \wBIn6[8] , 
        \wBIn6[7] , \wBIn6[6] , \wBIn6[5] , \wBIn6[4] , \wBIn6[3] , \wBIn6[2] , 
        \wBIn6[1] , \wBIn6[0] }), .HiOut({\wBMid5[31] , \wBMid5[30] , 
        \wBMid5[29] , \wBMid5[28] , \wBMid5[27] , \wBMid5[26] , \wBMid5[25] , 
        \wBMid5[24] , \wBMid5[23] , \wBMid5[22] , \wBMid5[21] , \wBMid5[20] , 
        \wBMid5[19] , \wBMid5[18] , \wBMid5[17] , \wBMid5[16] , \wBMid5[15] , 
        \wBMid5[14] , \wBMid5[13] , \wBMid5[12] , \wBMid5[11] , \wBMid5[10] , 
        \wBMid5[9] , \wBMid5[8] , \wBMid5[7] , \wBMid5[6] , \wBMid5[5] , 
        \wBMid5[4] , \wBMid5[3] , \wBMid5[2] , \wBMid5[1] , \wBMid5[0] }), 
        .LoOut({\wAMid6[31] , \wAMid6[30] , \wAMid6[29] , \wAMid6[28] , 
        \wAMid6[27] , \wAMid6[26] , \wAMid6[25] , \wAMid6[24] , \wAMid6[23] , 
        \wAMid6[22] , \wAMid6[21] , \wAMid6[20] , \wAMid6[19] , \wAMid6[18] , 
        \wAMid6[17] , \wAMid6[16] , \wAMid6[15] , \wAMid6[14] , \wAMid6[13] , 
        \wAMid6[12] , \wAMid6[11] , \wAMid6[10] , \wAMid6[9] , \wAMid6[8] , 
        \wAMid6[7] , \wAMid6[6] , \wAMid6[5] , \wAMid6[4] , \wAMid6[3] , 
        \wAMid6[2] , \wAMid6[1] , \wAMid6[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn10[31] , \wAIn10[30] , \wAIn10[29] , \wAIn10[28] , \wAIn10[27] , 
        \wAIn10[26] , \wAIn10[25] , \wAIn10[24] , \wAIn10[23] , \wAIn10[22] , 
        \wAIn10[21] , \wAIn10[20] , \wAIn10[19] , \wAIn10[18] , \wAIn10[17] , 
        \wAIn10[16] , \wAIn10[15] , \wAIn10[14] , \wAIn10[13] , \wAIn10[12] , 
        \wAIn10[11] , \wAIn10[10] , \wAIn10[9] , \wAIn10[8] , \wAIn10[7] , 
        \wAIn10[6] , \wAIn10[5] , \wAIn10[4] , \wAIn10[3] , \wAIn10[2] , 
        \wAIn10[1] , \wAIn10[0] }), .BIn({\wBIn10[31] , \wBIn10[30] , 
        \wBIn10[29] , \wBIn10[28] , \wBIn10[27] , \wBIn10[26] , \wBIn10[25] , 
        \wBIn10[24] , \wBIn10[23] , \wBIn10[22] , \wBIn10[21] , \wBIn10[20] , 
        \wBIn10[19] , \wBIn10[18] , \wBIn10[17] , \wBIn10[16] , \wBIn10[15] , 
        \wBIn10[14] , \wBIn10[13] , \wBIn10[12] , \wBIn10[11] , \wBIn10[10] , 
        \wBIn10[9] , \wBIn10[8] , \wBIn10[7] , \wBIn10[6] , \wBIn10[5] , 
        \wBIn10[4] , \wBIn10[3] , \wBIn10[2] , \wBIn10[1] , \wBIn10[0] }), 
        .HiOut({\wBMid9[31] , \wBMid9[30] , \wBMid9[29] , \wBMid9[28] , 
        \wBMid9[27] , \wBMid9[26] , \wBMid9[25] , \wBMid9[24] , \wBMid9[23] , 
        \wBMid9[22] , \wBMid9[21] , \wBMid9[20] , \wBMid9[19] , \wBMid9[18] , 
        \wBMid9[17] , \wBMid9[16] , \wBMid9[15] , \wBMid9[14] , \wBMid9[13] , 
        \wBMid9[12] , \wBMid9[11] , \wBMid9[10] , \wBMid9[9] , \wBMid9[8] , 
        \wBMid9[7] , \wBMid9[6] , \wBMid9[5] , \wBMid9[4] , \wBMid9[3] , 
        \wBMid9[2] , \wBMid9[1] , \wBMid9[0] }), .LoOut({\wAMid10[31] , 
        \wAMid10[30] , \wAMid10[29] , \wAMid10[28] , \wAMid10[27] , 
        \wAMid10[26] , \wAMid10[25] , \wAMid10[24] , \wAMid10[23] , 
        \wAMid10[22] , \wAMid10[21] , \wAMid10[20] , \wAMid10[19] , 
        \wAMid10[18] , \wAMid10[17] , \wAMid10[16] , \wAMid10[15] , 
        \wAMid10[14] , \wAMid10[13] , \wAMid10[12] , \wAMid10[11] , 
        \wAMid10[10] , \wAMid10[9] , \wAMid10[8] , \wAMid10[7] , \wAMid10[6] , 
        \wAMid10[5] , \wAMid10[4] , \wAMid10[3] , \wAMid10[2] , \wAMid10[1] , 
        \wAMid10[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn17[31] , \wAIn17[30] , \wAIn17[29] , \wAIn17[28] , \wAIn17[27] , 
        \wAIn17[26] , \wAIn17[25] , \wAIn17[24] , \wAIn17[23] , \wAIn17[22] , 
        \wAIn17[21] , \wAIn17[20] , \wAIn17[19] , \wAIn17[18] , \wAIn17[17] , 
        \wAIn17[16] , \wAIn17[15] , \wAIn17[14] , \wAIn17[13] , \wAIn17[12] , 
        \wAIn17[11] , \wAIn17[10] , \wAIn17[9] , \wAIn17[8] , \wAIn17[7] , 
        \wAIn17[6] , \wAIn17[5] , \wAIn17[4] , \wAIn17[3] , \wAIn17[2] , 
        \wAIn17[1] , \wAIn17[0] }), .BIn({\wBIn17[31] , \wBIn17[30] , 
        \wBIn17[29] , \wBIn17[28] , \wBIn17[27] , \wBIn17[26] , \wBIn17[25] , 
        \wBIn17[24] , \wBIn17[23] , \wBIn17[22] , \wBIn17[21] , \wBIn17[20] , 
        \wBIn17[19] , \wBIn17[18] , \wBIn17[17] , \wBIn17[16] , \wBIn17[15] , 
        \wBIn17[14] , \wBIn17[13] , \wBIn17[12] , \wBIn17[11] , \wBIn17[10] , 
        \wBIn17[9] , \wBIn17[8] , \wBIn17[7] , \wBIn17[6] , \wBIn17[5] , 
        \wBIn17[4] , \wBIn17[3] , \wBIn17[2] , \wBIn17[1] , \wBIn17[0] }), 
        .HiOut({\wBMid16[31] , \wBMid16[30] , \wBMid16[29] , \wBMid16[28] , 
        \wBMid16[27] , \wBMid16[26] , \wBMid16[25] , \wBMid16[24] , 
        \wBMid16[23] , \wBMid16[22] , \wBMid16[21] , \wBMid16[20] , 
        \wBMid16[19] , \wBMid16[18] , \wBMid16[17] , \wBMid16[16] , 
        \wBMid16[15] , \wBMid16[14] , \wBMid16[13] , \wBMid16[12] , 
        \wBMid16[11] , \wBMid16[10] , \wBMid16[9] , \wBMid16[8] , \wBMid16[7] , 
        \wBMid16[6] , \wBMid16[5] , \wBMid16[4] , \wBMid16[3] , \wBMid16[2] , 
        \wBMid16[1] , \wBMid16[0] }), .LoOut({\wAMid17[31] , \wAMid17[30] , 
        \wAMid17[29] , \wAMid17[28] , \wAMid17[27] , \wAMid17[26] , 
        \wAMid17[25] , \wAMid17[24] , \wAMid17[23] , \wAMid17[22] , 
        \wAMid17[21] , \wAMid17[20] , \wAMid17[19] , \wAMid17[18] , 
        \wAMid17[17] , \wAMid17[16] , \wAMid17[15] , \wAMid17[14] , 
        \wAMid17[13] , \wAMid17[12] , \wAMid17[11] , \wAMid17[10] , 
        \wAMid17[9] , \wAMid17[8] , \wAMid17[7] , \wAMid17[6] , \wAMid17[5] , 
        \wAMid17[4] , \wAMid17[3] , \wAMid17[2] , \wAMid17[1] , \wAMid17[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn30[31] , \wAIn30[30] , \wAIn30[29] , \wAIn30[28] , \wAIn30[27] , 
        \wAIn30[26] , \wAIn30[25] , \wAIn30[24] , \wAIn30[23] , \wAIn30[22] , 
        \wAIn30[21] , \wAIn30[20] , \wAIn30[19] , \wAIn30[18] , \wAIn30[17] , 
        \wAIn30[16] , \wAIn30[15] , \wAIn30[14] , \wAIn30[13] , \wAIn30[12] , 
        \wAIn30[11] , \wAIn30[10] , \wAIn30[9] , \wAIn30[8] , \wAIn30[7] , 
        \wAIn30[6] , \wAIn30[5] , \wAIn30[4] , \wAIn30[3] , \wAIn30[2] , 
        \wAIn30[1] , \wAIn30[0] }), .BIn({\wBIn30[31] , \wBIn30[30] , 
        \wBIn30[29] , \wBIn30[28] , \wBIn30[27] , \wBIn30[26] , \wBIn30[25] , 
        \wBIn30[24] , \wBIn30[23] , \wBIn30[22] , \wBIn30[21] , \wBIn30[20] , 
        \wBIn30[19] , \wBIn30[18] , \wBIn30[17] , \wBIn30[16] , \wBIn30[15] , 
        \wBIn30[14] , \wBIn30[13] , \wBIn30[12] , \wBIn30[11] , \wBIn30[10] , 
        \wBIn30[9] , \wBIn30[8] , \wBIn30[7] , \wBIn30[6] , \wBIn30[5] , 
        \wBIn30[4] , \wBIn30[3] , \wBIn30[2] , \wBIn30[1] , \wBIn30[0] }), 
        .HiOut({\wBMid29[31] , \wBMid29[30] , \wBMid29[29] , \wBMid29[28] , 
        \wBMid29[27] , \wBMid29[26] , \wBMid29[25] , \wBMid29[24] , 
        \wBMid29[23] , \wBMid29[22] , \wBMid29[21] , \wBMid29[20] , 
        \wBMid29[19] , \wBMid29[18] , \wBMid29[17] , \wBMid29[16] , 
        \wBMid29[15] , \wBMid29[14] , \wBMid29[13] , \wBMid29[12] , 
        \wBMid29[11] , \wBMid29[10] , \wBMid29[9] , \wBMid29[8] , \wBMid29[7] , 
        \wBMid29[6] , \wBMid29[5] , \wBMid29[4] , \wBMid29[3] , \wBMid29[2] , 
        \wBMid29[1] , \wBMid29[0] }), .LoOut({\wAMid30[31] , \wAMid30[30] , 
        \wAMid30[29] , \wAMid30[28] , \wAMid30[27] , \wAMid30[26] , 
        \wAMid30[25] , \wAMid30[24] , \wAMid30[23] , \wAMid30[22] , 
        \wAMid30[21] , \wAMid30[20] , \wAMid30[19] , \wAMid30[18] , 
        \wAMid30[17] , \wAMid30[16] , \wAMid30[15] , \wAMid30[14] , 
        \wAMid30[13] , \wAMid30[12] , \wAMid30[11] , \wAMid30[10] , 
        \wAMid30[9] , \wAMid30[8] , \wAMid30[7] , \wAMid30[6] , \wAMid30[5] , 
        \wAMid30[4] , \wAMid30[3] , \wAMid30[2] , \wAMid30[1] , \wAMid30[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn45[31] , \wAIn45[30] , \wAIn45[29] , \wAIn45[28] , \wAIn45[27] , 
        \wAIn45[26] , \wAIn45[25] , \wAIn45[24] , \wAIn45[23] , \wAIn45[22] , 
        \wAIn45[21] , \wAIn45[20] , \wAIn45[19] , \wAIn45[18] , \wAIn45[17] , 
        \wAIn45[16] , \wAIn45[15] , \wAIn45[14] , \wAIn45[13] , \wAIn45[12] , 
        \wAIn45[11] , \wAIn45[10] , \wAIn45[9] , \wAIn45[8] , \wAIn45[7] , 
        \wAIn45[6] , \wAIn45[5] , \wAIn45[4] , \wAIn45[3] , \wAIn45[2] , 
        \wAIn45[1] , \wAIn45[0] }), .BIn({\wBIn45[31] , \wBIn45[30] , 
        \wBIn45[29] , \wBIn45[28] , \wBIn45[27] , \wBIn45[26] , \wBIn45[25] , 
        \wBIn45[24] , \wBIn45[23] , \wBIn45[22] , \wBIn45[21] , \wBIn45[20] , 
        \wBIn45[19] , \wBIn45[18] , \wBIn45[17] , \wBIn45[16] , \wBIn45[15] , 
        \wBIn45[14] , \wBIn45[13] , \wBIn45[12] , \wBIn45[11] , \wBIn45[10] , 
        \wBIn45[9] , \wBIn45[8] , \wBIn45[7] , \wBIn45[6] , \wBIn45[5] , 
        \wBIn45[4] , \wBIn45[3] , \wBIn45[2] , \wBIn45[1] , \wBIn45[0] }), 
        .HiOut({\wBMid44[31] , \wBMid44[30] , \wBMid44[29] , \wBMid44[28] , 
        \wBMid44[27] , \wBMid44[26] , \wBMid44[25] , \wBMid44[24] , 
        \wBMid44[23] , \wBMid44[22] , \wBMid44[21] , \wBMid44[20] , 
        \wBMid44[19] , \wBMid44[18] , \wBMid44[17] , \wBMid44[16] , 
        \wBMid44[15] , \wBMid44[14] , \wBMid44[13] , \wBMid44[12] , 
        \wBMid44[11] , \wBMid44[10] , \wBMid44[9] , \wBMid44[8] , \wBMid44[7] , 
        \wBMid44[6] , \wBMid44[5] , \wBMid44[4] , \wBMid44[3] , \wBMid44[2] , 
        \wBMid44[1] , \wBMid44[0] }), .LoOut({\wAMid45[31] , \wAMid45[30] , 
        \wAMid45[29] , \wAMid45[28] , \wAMid45[27] , \wAMid45[26] , 
        \wAMid45[25] , \wAMid45[24] , \wAMid45[23] , \wAMid45[22] , 
        \wAMid45[21] , \wAMid45[20] , \wAMid45[19] , \wAMid45[18] , 
        \wAMid45[17] , \wAMid45[16] , \wAMid45[15] , \wAMid45[14] , 
        \wAMid45[13] , \wAMid45[12] , \wAMid45[11] , \wAMid45[10] , 
        \wAMid45[9] , \wAMid45[8] , \wAMid45[7] , \wAMid45[6] , \wAMid45[5] , 
        \wAMid45[4] , \wAMid45[3] , \wAMid45[2] , \wAMid45[1] , \wAMid45[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid75[31] , \wAMid75[30] , \wAMid75[29] , \wAMid75[28] , 
        \wAMid75[27] , \wAMid75[26] , \wAMid75[25] , \wAMid75[24] , 
        \wAMid75[23] , \wAMid75[22] , \wAMid75[21] , \wAMid75[20] , 
        \wAMid75[19] , \wAMid75[18] , \wAMid75[17] , \wAMid75[16] , 
        \wAMid75[15] , \wAMid75[14] , \wAMid75[13] , \wAMid75[12] , 
        \wAMid75[11] , \wAMid75[10] , \wAMid75[9] , \wAMid75[8] , \wAMid75[7] , 
        \wAMid75[6] , \wAMid75[5] , \wAMid75[4] , \wAMid75[3] , \wAMid75[2] , 
        \wAMid75[1] , \wAMid75[0] }), .BIn({\wBMid75[31] , \wBMid75[30] , 
        \wBMid75[29] , \wBMid75[28] , \wBMid75[27] , \wBMid75[26] , 
        \wBMid75[25] , \wBMid75[24] , \wBMid75[23] , \wBMid75[22] , 
        \wBMid75[21] , \wBMid75[20] , \wBMid75[19] , \wBMid75[18] , 
        \wBMid75[17] , \wBMid75[16] , \wBMid75[15] , \wBMid75[14] , 
        \wBMid75[13] , \wBMid75[12] , \wBMid75[11] , \wBMid75[10] , 
        \wBMid75[9] , \wBMid75[8] , \wBMid75[7] , \wBMid75[6] , \wBMid75[5] , 
        \wBMid75[4] , \wBMid75[3] , \wBMid75[2] , \wBMid75[1] , \wBMid75[0] }), 
        .HiOut({\wRegInB75[31] , \wRegInB75[30] , \wRegInB75[29] , 
        \wRegInB75[28] , \wRegInB75[27] , \wRegInB75[26] , \wRegInB75[25] , 
        \wRegInB75[24] , \wRegInB75[23] , \wRegInB75[22] , \wRegInB75[21] , 
        \wRegInB75[20] , \wRegInB75[19] , \wRegInB75[18] , \wRegInB75[17] , 
        \wRegInB75[16] , \wRegInB75[15] , \wRegInB75[14] , \wRegInB75[13] , 
        \wRegInB75[12] , \wRegInB75[11] , \wRegInB75[10] , \wRegInB75[9] , 
        \wRegInB75[8] , \wRegInB75[7] , \wRegInB75[6] , \wRegInB75[5] , 
        \wRegInB75[4] , \wRegInB75[3] , \wRegInB75[2] , \wRegInB75[1] , 
        \wRegInB75[0] }), .LoOut({\wRegInA76[31] , \wRegInA76[30] , 
        \wRegInA76[29] , \wRegInA76[28] , \wRegInA76[27] , \wRegInA76[26] , 
        \wRegInA76[25] , \wRegInA76[24] , \wRegInA76[23] , \wRegInA76[22] , 
        \wRegInA76[21] , \wRegInA76[20] , \wRegInA76[19] , \wRegInA76[18] , 
        \wRegInA76[17] , \wRegInA76[16] , \wRegInA76[15] , \wRegInA76[14] , 
        \wRegInA76[13] , \wRegInA76[12] , \wRegInA76[11] , \wRegInA76[10] , 
        \wRegInA76[9] , \wRegInA76[8] , \wRegInA76[7] , \wRegInA76[6] , 
        \wRegInA76[5] , \wRegInA76[4] , \wRegInA76[3] , \wRegInA76[2] , 
        \wRegInA76[1] , \wRegInA76[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid90[31] , \wAMid90[30] , \wAMid90[29] , \wAMid90[28] , 
        \wAMid90[27] , \wAMid90[26] , \wAMid90[25] , \wAMid90[24] , 
        \wAMid90[23] , \wAMid90[22] , \wAMid90[21] , \wAMid90[20] , 
        \wAMid90[19] , \wAMid90[18] , \wAMid90[17] , \wAMid90[16] , 
        \wAMid90[15] , \wAMid90[14] , \wAMid90[13] , \wAMid90[12] , 
        \wAMid90[11] , \wAMid90[10] , \wAMid90[9] , \wAMid90[8] , \wAMid90[7] , 
        \wAMid90[6] , \wAMid90[5] , \wAMid90[4] , \wAMid90[3] , \wAMid90[2] , 
        \wAMid90[1] , \wAMid90[0] }), .BIn({\wBMid90[31] , \wBMid90[30] , 
        \wBMid90[29] , \wBMid90[28] , \wBMid90[27] , \wBMid90[26] , 
        \wBMid90[25] , \wBMid90[24] , \wBMid90[23] , \wBMid90[22] , 
        \wBMid90[21] , \wBMid90[20] , \wBMid90[19] , \wBMid90[18] , 
        \wBMid90[17] , \wBMid90[16] , \wBMid90[15] , \wBMid90[14] , 
        \wBMid90[13] , \wBMid90[12] , \wBMid90[11] , \wBMid90[10] , 
        \wBMid90[9] , \wBMid90[8] , \wBMid90[7] , \wBMid90[6] , \wBMid90[5] , 
        \wBMid90[4] , \wBMid90[3] , \wBMid90[2] , \wBMid90[1] , \wBMid90[0] }), 
        .HiOut({\wRegInB90[31] , \wRegInB90[30] , \wRegInB90[29] , 
        \wRegInB90[28] , \wRegInB90[27] , \wRegInB90[26] , \wRegInB90[25] , 
        \wRegInB90[24] , \wRegInB90[23] , \wRegInB90[22] , \wRegInB90[21] , 
        \wRegInB90[20] , \wRegInB90[19] , \wRegInB90[18] , \wRegInB90[17] , 
        \wRegInB90[16] , \wRegInB90[15] , \wRegInB90[14] , \wRegInB90[13] , 
        \wRegInB90[12] , \wRegInB90[11] , \wRegInB90[10] , \wRegInB90[9] , 
        \wRegInB90[8] , \wRegInB90[7] , \wRegInB90[6] , \wRegInB90[5] , 
        \wRegInB90[4] , \wRegInB90[3] , \wRegInB90[2] , \wRegInB90[1] , 
        \wRegInB90[0] }), .LoOut({\wRegInA91[31] , \wRegInA91[30] , 
        \wRegInA91[29] , \wRegInA91[28] , \wRegInA91[27] , \wRegInA91[26] , 
        \wRegInA91[25] , \wRegInA91[24] , \wRegInA91[23] , \wRegInA91[22] , 
        \wRegInA91[21] , \wRegInA91[20] , \wRegInA91[19] , \wRegInA91[18] , 
        \wRegInA91[17] , \wRegInA91[16] , \wRegInA91[15] , \wRegInA91[14] , 
        \wRegInA91[13] , \wRegInA91[12] , \wRegInA91[11] , \wRegInA91[10] , 
        \wRegInA91[9] , \wRegInA91[8] , \wRegInA91[7] , \wRegInA91[6] , 
        \wRegInA91[5] , \wRegInA91[4] , \wRegInA91[3] , \wRegInA91[2] , 
        \wRegInA91[1] , \wRegInA91[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_239 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink240[31] , \ScanLink240[30] , \ScanLink240[29] , 
        \ScanLink240[28] , \ScanLink240[27] , \ScanLink240[26] , 
        \ScanLink240[25] , \ScanLink240[24] , \ScanLink240[23] , 
        \ScanLink240[22] , \ScanLink240[21] , \ScanLink240[20] , 
        \ScanLink240[19] , \ScanLink240[18] , \ScanLink240[17] , 
        \ScanLink240[16] , \ScanLink240[15] , \ScanLink240[14] , 
        \ScanLink240[13] , \ScanLink240[12] , \ScanLink240[11] , 
        \ScanLink240[10] , \ScanLink240[9] , \ScanLink240[8] , 
        \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , \ScanLink240[4] , 
        \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , \ScanLink240[0] 
        }), .ScanOut({\ScanLink239[31] , \ScanLink239[30] , \ScanLink239[29] , 
        \ScanLink239[28] , \ScanLink239[27] , \ScanLink239[26] , 
        \ScanLink239[25] , \ScanLink239[24] , \ScanLink239[23] , 
        \ScanLink239[22] , \ScanLink239[21] , \ScanLink239[20] , 
        \ScanLink239[19] , \ScanLink239[18] , \ScanLink239[17] , 
        \ScanLink239[16] , \ScanLink239[15] , \ScanLink239[14] , 
        \ScanLink239[13] , \ScanLink239[12] , \ScanLink239[11] , 
        \ScanLink239[10] , \ScanLink239[9] , \ScanLink239[8] , 
        \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , \ScanLink239[4] , 
        \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , \ScanLink239[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA8[31] , \wRegInA8[30] , \wRegInA8[29] , \wRegInA8[28] , 
        \wRegInA8[27] , \wRegInA8[26] , \wRegInA8[25] , \wRegInA8[24] , 
        \wRegInA8[23] , \wRegInA8[22] , \wRegInA8[21] , \wRegInA8[20] , 
        \wRegInA8[19] , \wRegInA8[18] , \wRegInA8[17] , \wRegInA8[16] , 
        \wRegInA8[15] , \wRegInA8[14] , \wRegInA8[13] , \wRegInA8[12] , 
        \wRegInA8[11] , \wRegInA8[10] , \wRegInA8[9] , \wRegInA8[8] , 
        \wRegInA8[7] , \wRegInA8[6] , \wRegInA8[5] , \wRegInA8[4] , 
        \wRegInA8[3] , \wRegInA8[2] , \wRegInA8[1] , \wRegInA8[0] }), .Out({
        \wAIn8[31] , \wAIn8[30] , \wAIn8[29] , \wAIn8[28] , \wAIn8[27] , 
        \wAIn8[26] , \wAIn8[25] , \wAIn8[24] , \wAIn8[23] , \wAIn8[22] , 
        \wAIn8[21] , \wAIn8[20] , \wAIn8[19] , \wAIn8[18] , \wAIn8[17] , 
        \wAIn8[16] , \wAIn8[15] , \wAIn8[14] , \wAIn8[13] , \wAIn8[12] , 
        \wAIn8[11] , \wAIn8[10] , \wAIn8[9] , \wAIn8[8] , \wAIn8[7] , 
        \wAIn8[6] , \wAIn8[5] , \wAIn8[4] , \wAIn8[3] , \wAIn8[2] , \wAIn8[1] , 
        \wAIn8[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_109 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink110[31] , \ScanLink110[30] , \ScanLink110[29] , 
        \ScanLink110[28] , \ScanLink110[27] , \ScanLink110[26] , 
        \ScanLink110[25] , \ScanLink110[24] , \ScanLink110[23] , 
        \ScanLink110[22] , \ScanLink110[21] , \ScanLink110[20] , 
        \ScanLink110[19] , \ScanLink110[18] , \ScanLink110[17] , 
        \ScanLink110[16] , \ScanLink110[15] , \ScanLink110[14] , 
        \ScanLink110[13] , \ScanLink110[12] , \ScanLink110[11] , 
        \ScanLink110[10] , \ScanLink110[9] , \ScanLink110[8] , 
        \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , \ScanLink110[4] , 
        \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , \ScanLink110[0] 
        }), .ScanOut({\ScanLink109[31] , \ScanLink109[30] , \ScanLink109[29] , 
        \ScanLink109[28] , \ScanLink109[27] , \ScanLink109[26] , 
        \ScanLink109[25] , \ScanLink109[24] , \ScanLink109[23] , 
        \ScanLink109[22] , \ScanLink109[21] , \ScanLink109[20] , 
        \ScanLink109[19] , \ScanLink109[18] , \ScanLink109[17] , 
        \ScanLink109[16] , \ScanLink109[15] , \ScanLink109[14] , 
        \ScanLink109[13] , \ScanLink109[12] , \ScanLink109[11] , 
        \ScanLink109[10] , \ScanLink109[9] , \ScanLink109[8] , 
        \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , \ScanLink109[4] , 
        \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , \ScanLink109[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA73[31] , \wRegInA73[30] , \wRegInA73[29] , 
        \wRegInA73[28] , \wRegInA73[27] , \wRegInA73[26] , \wRegInA73[25] , 
        \wRegInA73[24] , \wRegInA73[23] , \wRegInA73[22] , \wRegInA73[21] , 
        \wRegInA73[20] , \wRegInA73[19] , \wRegInA73[18] , \wRegInA73[17] , 
        \wRegInA73[16] , \wRegInA73[15] , \wRegInA73[14] , \wRegInA73[13] , 
        \wRegInA73[12] , \wRegInA73[11] , \wRegInA73[10] , \wRegInA73[9] , 
        \wRegInA73[8] , \wRegInA73[7] , \wRegInA73[6] , \wRegInA73[5] , 
        \wRegInA73[4] , \wRegInA73[3] , \wRegInA73[2] , \wRegInA73[1] , 
        \wRegInA73[0] }), .Out({\wAIn73[31] , \wAIn73[30] , \wAIn73[29] , 
        \wAIn73[28] , \wAIn73[27] , \wAIn73[26] , \wAIn73[25] , \wAIn73[24] , 
        \wAIn73[23] , \wAIn73[22] , \wAIn73[21] , \wAIn73[20] , \wAIn73[19] , 
        \wAIn73[18] , \wAIn73[17] , \wAIn73[16] , \wAIn73[15] , \wAIn73[14] , 
        \wAIn73[13] , \wAIn73[12] , \wAIn73[11] , \wAIn73[10] , \wAIn73[9] , 
        \wAIn73[8] , \wAIn73[7] , \wAIn73[6] , \wAIn73[5] , \wAIn73[4] , 
        \wAIn73[3] , \wAIn73[2] , \wAIn73[1] , \wAIn73[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_59 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink60[31] , \ScanLink60[30] , \ScanLink60[29] , 
        \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , \ScanLink60[25] , 
        \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , \ScanLink60[21] , 
        \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , \ScanLink60[17] , 
        \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , \ScanLink60[13] , 
        \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , \ScanLink60[9] , 
        \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , \ScanLink60[5] , 
        \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , \ScanLink60[1] , 
        \ScanLink60[0] }), .ScanOut({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA98[31] , \wRegInA98[30] , 
        \wRegInA98[29] , \wRegInA98[28] , \wRegInA98[27] , \wRegInA98[26] , 
        \wRegInA98[25] , \wRegInA98[24] , \wRegInA98[23] , \wRegInA98[22] , 
        \wRegInA98[21] , \wRegInA98[20] , \wRegInA98[19] , \wRegInA98[18] , 
        \wRegInA98[17] , \wRegInA98[16] , \wRegInA98[15] , \wRegInA98[14] , 
        \wRegInA98[13] , \wRegInA98[12] , \wRegInA98[11] , \wRegInA98[10] , 
        \wRegInA98[9] , \wRegInA98[8] , \wRegInA98[7] , \wRegInA98[6] , 
        \wRegInA98[5] , \wRegInA98[4] , \wRegInA98[3] , \wRegInA98[2] , 
        \wRegInA98[1] , \wRegInA98[0] }), .Out({\wAIn98[31] , \wAIn98[30] , 
        \wAIn98[29] , \wAIn98[28] , \wAIn98[27] , \wAIn98[26] , \wAIn98[25] , 
        \wAIn98[24] , \wAIn98[23] , \wAIn98[22] , \wAIn98[21] , \wAIn98[20] , 
        \wAIn98[19] , \wAIn98[18] , \wAIn98[17] , \wAIn98[16] , \wAIn98[15] , 
        \wAIn98[14] , \wAIn98[13] , \wAIn98[12] , \wAIn98[11] , \wAIn98[10] , 
        \wAIn98[9] , \wAIn98[8] , \wAIn98[7] , \wAIn98[6] , \wAIn98[5] , 
        \wAIn98[4] , \wAIn98[3] , \wAIn98[2] , \wAIn98[1] , \wAIn98[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_140 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink141[31] , \ScanLink141[30] , \ScanLink141[29] , 
        \ScanLink141[28] , \ScanLink141[27] , \ScanLink141[26] , 
        \ScanLink141[25] , \ScanLink141[24] , \ScanLink141[23] , 
        \ScanLink141[22] , \ScanLink141[21] , \ScanLink141[20] , 
        \ScanLink141[19] , \ScanLink141[18] , \ScanLink141[17] , 
        \ScanLink141[16] , \ScanLink141[15] , \ScanLink141[14] , 
        \ScanLink141[13] , \ScanLink141[12] , \ScanLink141[11] , 
        \ScanLink141[10] , \ScanLink141[9] , \ScanLink141[8] , 
        \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , \ScanLink141[4] , 
        \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , \ScanLink141[0] 
        }), .ScanOut({\ScanLink140[31] , \ScanLink140[30] , \ScanLink140[29] , 
        \ScanLink140[28] , \ScanLink140[27] , \ScanLink140[26] , 
        \ScanLink140[25] , \ScanLink140[24] , \ScanLink140[23] , 
        \ScanLink140[22] , \ScanLink140[21] , \ScanLink140[20] , 
        \ScanLink140[19] , \ScanLink140[18] , \ScanLink140[17] , 
        \ScanLink140[16] , \ScanLink140[15] , \ScanLink140[14] , 
        \ScanLink140[13] , \ScanLink140[12] , \ScanLink140[11] , 
        \ScanLink140[10] , \ScanLink140[9] , \ScanLink140[8] , 
        \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , \ScanLink140[4] , 
        \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , \ScanLink140[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB57[31] , \wRegInB57[30] , \wRegInB57[29] , 
        \wRegInB57[28] , \wRegInB57[27] , \wRegInB57[26] , \wRegInB57[25] , 
        \wRegInB57[24] , \wRegInB57[23] , \wRegInB57[22] , \wRegInB57[21] , 
        \wRegInB57[20] , \wRegInB57[19] , \wRegInB57[18] , \wRegInB57[17] , 
        \wRegInB57[16] , \wRegInB57[15] , \wRegInB57[14] , \wRegInB57[13] , 
        \wRegInB57[12] , \wRegInB57[11] , \wRegInB57[10] , \wRegInB57[9] , 
        \wRegInB57[8] , \wRegInB57[7] , \wRegInB57[6] , \wRegInB57[5] , 
        \wRegInB57[4] , \wRegInB57[3] , \wRegInB57[2] , \wRegInB57[1] , 
        \wRegInB57[0] }), .Out({\wBIn57[31] , \wBIn57[30] , \wBIn57[29] , 
        \wBIn57[28] , \wBIn57[27] , \wBIn57[26] , \wBIn57[25] , \wBIn57[24] , 
        \wBIn57[23] , \wBIn57[22] , \wBIn57[21] , \wBIn57[20] , \wBIn57[19] , 
        \wBIn57[18] , \wBIn57[17] , \wBIn57[16] , \wBIn57[15] , \wBIn57[14] , 
        \wBIn57[13] , \wBIn57[12] , \wBIn57[11] , \wBIn57[10] , \wBIn57[9] , 
        \wBIn57[8] , \wBIn57[7] , \wBIn57[6] , \wBIn57[5] , \wBIn57[4] , 
        \wBIn57[3] , \wBIn57[2] , \wBIn57[1] , \wBIn57[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_10 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[31] , \ScanLink11[30] , \ScanLink11[29] , 
        \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , \ScanLink11[25] , 
        \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , \ScanLink11[21] , 
        \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , \ScanLink11[17] , 
        \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , \ScanLink11[13] , 
        \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , \ScanLink11[9] , 
        \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB122[31] , \wRegInB122[30] , 
        \wRegInB122[29] , \wRegInB122[28] , \wRegInB122[27] , \wRegInB122[26] , 
        \wRegInB122[25] , \wRegInB122[24] , \wRegInB122[23] , \wRegInB122[22] , 
        \wRegInB122[21] , \wRegInB122[20] , \wRegInB122[19] , \wRegInB122[18] , 
        \wRegInB122[17] , \wRegInB122[16] , \wRegInB122[15] , \wRegInB122[14] , 
        \wRegInB122[13] , \wRegInB122[12] , \wRegInB122[11] , \wRegInB122[10] , 
        \wRegInB122[9] , \wRegInB122[8] , \wRegInB122[7] , \wRegInB122[6] , 
        \wRegInB122[5] , \wRegInB122[4] , \wRegInB122[3] , \wRegInB122[2] , 
        \wRegInB122[1] , \wRegInB122[0] }), .Out({\wBIn122[31] , \wBIn122[30] , 
        \wBIn122[29] , \wBIn122[28] , \wBIn122[27] , \wBIn122[26] , 
        \wBIn122[25] , \wBIn122[24] , \wBIn122[23] , \wBIn122[22] , 
        \wBIn122[21] , \wBIn122[20] , \wBIn122[19] , \wBIn122[18] , 
        \wBIn122[17] , \wBIn122[16] , \wBIn122[15] , \wBIn122[14] , 
        \wBIn122[13] , \wBIn122[12] , \wBIn122[11] , \wBIn122[10] , 
        \wBIn122[9] , \wBIn122[8] , \wBIn122[7] , \wBIn122[6] , \wBIn122[5] , 
        \wBIn122[4] , \wBIn122[3] , \wBIn122[2] , \wBIn122[1] , \wBIn122[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn62[31] , \wAIn62[30] , \wAIn62[29] , \wAIn62[28] , \wAIn62[27] , 
        \wAIn62[26] , \wAIn62[25] , \wAIn62[24] , \wAIn62[23] , \wAIn62[22] , 
        \wAIn62[21] , \wAIn62[20] , \wAIn62[19] , \wAIn62[18] , \wAIn62[17] , 
        \wAIn62[16] , \wAIn62[15] , \wAIn62[14] , \wAIn62[13] , \wAIn62[12] , 
        \wAIn62[11] , \wAIn62[10] , \wAIn62[9] , \wAIn62[8] , \wAIn62[7] , 
        \wAIn62[6] , \wAIn62[5] , \wAIn62[4] , \wAIn62[3] , \wAIn62[2] , 
        \wAIn62[1] , \wAIn62[0] }), .BIn({\wBIn62[31] , \wBIn62[30] , 
        \wBIn62[29] , \wBIn62[28] , \wBIn62[27] , \wBIn62[26] , \wBIn62[25] , 
        \wBIn62[24] , \wBIn62[23] , \wBIn62[22] , \wBIn62[21] , \wBIn62[20] , 
        \wBIn62[19] , \wBIn62[18] , \wBIn62[17] , \wBIn62[16] , \wBIn62[15] , 
        \wBIn62[14] , \wBIn62[13] , \wBIn62[12] , \wBIn62[11] , \wBIn62[10] , 
        \wBIn62[9] , \wBIn62[8] , \wBIn62[7] , \wBIn62[6] , \wBIn62[5] , 
        \wBIn62[4] , \wBIn62[3] , \wBIn62[2] , \wBIn62[1] , \wBIn62[0] }), 
        .HiOut({\wBMid61[31] , \wBMid61[30] , \wBMid61[29] , \wBMid61[28] , 
        \wBMid61[27] , \wBMid61[26] , \wBMid61[25] , \wBMid61[24] , 
        \wBMid61[23] , \wBMid61[22] , \wBMid61[21] , \wBMid61[20] , 
        \wBMid61[19] , \wBMid61[18] , \wBMid61[17] , \wBMid61[16] , 
        \wBMid61[15] , \wBMid61[14] , \wBMid61[13] , \wBMid61[12] , 
        \wBMid61[11] , \wBMid61[10] , \wBMid61[9] , \wBMid61[8] , \wBMid61[7] , 
        \wBMid61[6] , \wBMid61[5] , \wBMid61[4] , \wBMid61[3] , \wBMid61[2] , 
        \wBMid61[1] , \wBMid61[0] }), .LoOut({\wAMid62[31] , \wAMid62[30] , 
        \wAMid62[29] , \wAMid62[28] , \wAMid62[27] , \wAMid62[26] , 
        \wAMid62[25] , \wAMid62[24] , \wAMid62[23] , \wAMid62[22] , 
        \wAMid62[21] , \wAMid62[20] , \wAMid62[19] , \wAMid62[18] , 
        \wAMid62[17] , \wAMid62[16] , \wAMid62[15] , \wAMid62[14] , 
        \wAMid62[13] , \wAMid62[12] , \wAMid62[11] , \wAMid62[10] , 
        \wAMid62[9] , \wAMid62[8] , \wAMid62[7] , \wAMid62[6] , \wAMid62[5] , 
        \wAMid62[4] , \wAMid62[3] , \wAMid62[2] , \wAMid62[1] , \wAMid62[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid52[31] , \wAMid52[30] , \wAMid52[29] , \wAMid52[28] , 
        \wAMid52[27] , \wAMid52[26] , \wAMid52[25] , \wAMid52[24] , 
        \wAMid52[23] , \wAMid52[22] , \wAMid52[21] , \wAMid52[20] , 
        \wAMid52[19] , \wAMid52[18] , \wAMid52[17] , \wAMid52[16] , 
        \wAMid52[15] , \wAMid52[14] , \wAMid52[13] , \wAMid52[12] , 
        \wAMid52[11] , \wAMid52[10] , \wAMid52[9] , \wAMid52[8] , \wAMid52[7] , 
        \wAMid52[6] , \wAMid52[5] , \wAMid52[4] , \wAMid52[3] , \wAMid52[2] , 
        \wAMid52[1] , \wAMid52[0] }), .BIn({\wBMid52[31] , \wBMid52[30] , 
        \wBMid52[29] , \wBMid52[28] , \wBMid52[27] , \wBMid52[26] , 
        \wBMid52[25] , \wBMid52[24] , \wBMid52[23] , \wBMid52[22] , 
        \wBMid52[21] , \wBMid52[20] , \wBMid52[19] , \wBMid52[18] , 
        \wBMid52[17] , \wBMid52[16] , \wBMid52[15] , \wBMid52[14] , 
        \wBMid52[13] , \wBMid52[12] , \wBMid52[11] , \wBMid52[10] , 
        \wBMid52[9] , \wBMid52[8] , \wBMid52[7] , \wBMid52[6] , \wBMid52[5] , 
        \wBMid52[4] , \wBMid52[3] , \wBMid52[2] , \wBMid52[1] , \wBMid52[0] }), 
        .HiOut({\wRegInB52[31] , \wRegInB52[30] , \wRegInB52[29] , 
        \wRegInB52[28] , \wRegInB52[27] , \wRegInB52[26] , \wRegInB52[25] , 
        \wRegInB52[24] , \wRegInB52[23] , \wRegInB52[22] , \wRegInB52[21] , 
        \wRegInB52[20] , \wRegInB52[19] , \wRegInB52[18] , \wRegInB52[17] , 
        \wRegInB52[16] , \wRegInB52[15] , \wRegInB52[14] , \wRegInB52[13] , 
        \wRegInB52[12] , \wRegInB52[11] , \wRegInB52[10] , \wRegInB52[9] , 
        \wRegInB52[8] , \wRegInB52[7] , \wRegInB52[6] , \wRegInB52[5] , 
        \wRegInB52[4] , \wRegInB52[3] , \wRegInB52[2] , \wRegInB52[1] , 
        \wRegInB52[0] }), .LoOut({\wRegInA53[31] , \wRegInA53[30] , 
        \wRegInA53[29] , \wRegInA53[28] , \wRegInA53[27] , \wRegInA53[26] , 
        \wRegInA53[25] , \wRegInA53[24] , \wRegInA53[23] , \wRegInA53[22] , 
        \wRegInA53[21] , \wRegInA53[20] , \wRegInA53[19] , \wRegInA53[18] , 
        \wRegInA53[17] , \wRegInA53[16] , \wRegInA53[15] , \wRegInA53[14] , 
        \wRegInA53[13] , \wRegInA53[12] , \wRegInA53[11] , \wRegInA53[10] , 
        \wRegInA53[9] , \wRegInA53[8] , \wRegInA53[7] , \wRegInA53[6] , 
        \wRegInA53[5] , \wRegInA53[4] , \wRegInA53[3] , \wRegInA53[2] , 
        \wRegInA53[1] , \wRegInA53[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_167 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink168[31] , \ScanLink168[30] , \ScanLink168[29] , 
        \ScanLink168[28] , \ScanLink168[27] , \ScanLink168[26] , 
        \ScanLink168[25] , \ScanLink168[24] , \ScanLink168[23] , 
        \ScanLink168[22] , \ScanLink168[21] , \ScanLink168[20] , 
        \ScanLink168[19] , \ScanLink168[18] , \ScanLink168[17] , 
        \ScanLink168[16] , \ScanLink168[15] , \ScanLink168[14] , 
        \ScanLink168[13] , \ScanLink168[12] , \ScanLink168[11] , 
        \ScanLink168[10] , \ScanLink168[9] , \ScanLink168[8] , 
        \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , \ScanLink168[4] , 
        \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , \ScanLink168[0] 
        }), .ScanOut({\ScanLink167[31] , \ScanLink167[30] , \ScanLink167[29] , 
        \ScanLink167[28] , \ScanLink167[27] , \ScanLink167[26] , 
        \ScanLink167[25] , \ScanLink167[24] , \ScanLink167[23] , 
        \ScanLink167[22] , \ScanLink167[21] , \ScanLink167[20] , 
        \ScanLink167[19] , \ScanLink167[18] , \ScanLink167[17] , 
        \ScanLink167[16] , \ScanLink167[15] , \ScanLink167[14] , 
        \ScanLink167[13] , \ScanLink167[12] , \ScanLink167[11] , 
        \ScanLink167[10] , \ScanLink167[9] , \ScanLink167[8] , 
        \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , \ScanLink167[4] , 
        \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , \ScanLink167[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA44[31] , \wRegInA44[30] , \wRegInA44[29] , 
        \wRegInA44[28] , \wRegInA44[27] , \wRegInA44[26] , \wRegInA44[25] , 
        \wRegInA44[24] , \wRegInA44[23] , \wRegInA44[22] , \wRegInA44[21] , 
        \wRegInA44[20] , \wRegInA44[19] , \wRegInA44[18] , \wRegInA44[17] , 
        \wRegInA44[16] , \wRegInA44[15] , \wRegInA44[14] , \wRegInA44[13] , 
        \wRegInA44[12] , \wRegInA44[11] , \wRegInA44[10] , \wRegInA44[9] , 
        \wRegInA44[8] , \wRegInA44[7] , \wRegInA44[6] , \wRegInA44[5] , 
        \wRegInA44[4] , \wRegInA44[3] , \wRegInA44[2] , \wRegInA44[1] , 
        \wRegInA44[0] }), .Out({\wAIn44[31] , \wAIn44[30] , \wAIn44[29] , 
        \wAIn44[28] , \wAIn44[27] , \wAIn44[26] , \wAIn44[25] , \wAIn44[24] , 
        \wAIn44[23] , \wAIn44[22] , \wAIn44[21] , \wAIn44[20] , \wAIn44[19] , 
        \wAIn44[18] , \wAIn44[17] , \wAIn44[16] , \wAIn44[15] , \wAIn44[14] , 
        \wAIn44[13] , \wAIn44[12] , \wAIn44[11] , \wAIn44[10] , \wAIn44[9] , 
        \wAIn44[8] , \wAIn44[7] , \wAIn44[6] , \wAIn44[5] , \wAIn44[4] , 
        \wAIn44[3] , \wAIn44[2] , \wAIn44[1] , \wAIn44[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_37 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink38[31] , \ScanLink38[30] , \ScanLink38[29] , 
        \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , \ScanLink38[25] , 
        \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , \ScanLink38[21] , 
        \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , \ScanLink38[17] , 
        \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , \ScanLink38[13] , 
        \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , \ScanLink38[9] , 
        \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , \ScanLink38[5] , 
        \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , \ScanLink38[1] , 
        \ScanLink38[0] }), .ScanOut({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA109[31] , \wRegInA109[30] , 
        \wRegInA109[29] , \wRegInA109[28] , \wRegInA109[27] , \wRegInA109[26] , 
        \wRegInA109[25] , \wRegInA109[24] , \wRegInA109[23] , \wRegInA109[22] , 
        \wRegInA109[21] , \wRegInA109[20] , \wRegInA109[19] , \wRegInA109[18] , 
        \wRegInA109[17] , \wRegInA109[16] , \wRegInA109[15] , \wRegInA109[14] , 
        \wRegInA109[13] , \wRegInA109[12] , \wRegInA109[11] , \wRegInA109[10] , 
        \wRegInA109[9] , \wRegInA109[8] , \wRegInA109[7] , \wRegInA109[6] , 
        \wRegInA109[5] , \wRegInA109[4] , \wRegInA109[3] , \wRegInA109[2] , 
        \wRegInA109[1] , \wRegInA109[0] }), .Out({\wAIn109[31] , \wAIn109[30] , 
        \wAIn109[29] , \wAIn109[28] , \wAIn109[27] , \wAIn109[26] , 
        \wAIn109[25] , \wAIn109[24] , \wAIn109[23] , \wAIn109[22] , 
        \wAIn109[21] , \wAIn109[20] , \wAIn109[19] , \wAIn109[18] , 
        \wAIn109[17] , \wAIn109[16] , \wAIn109[15] , \wAIn109[14] , 
        \wAIn109[13] , \wAIn109[12] , \wAIn109[11] , \wAIn109[10] , 
        \wAIn109[9] , \wAIn109[8] , \wAIn109[7] , \wAIn109[6] , \wAIn109[5] , 
        \wAIn109[4] , \wAIn109[3] , \wAIn109[2] , \wAIn109[1] , \wAIn109[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn79[31] , \wAIn79[30] , \wAIn79[29] , \wAIn79[28] , \wAIn79[27] , 
        \wAIn79[26] , \wAIn79[25] , \wAIn79[24] , \wAIn79[23] , \wAIn79[22] , 
        \wAIn79[21] , \wAIn79[20] , \wAIn79[19] , \wAIn79[18] , \wAIn79[17] , 
        \wAIn79[16] , \wAIn79[15] , \wAIn79[14] , \wAIn79[13] , \wAIn79[12] , 
        \wAIn79[11] , \wAIn79[10] , \wAIn79[9] , \wAIn79[8] , \wAIn79[7] , 
        \wAIn79[6] , \wAIn79[5] , \wAIn79[4] , \wAIn79[3] , \wAIn79[2] , 
        \wAIn79[1] , \wAIn79[0] }), .BIn({\wBIn79[31] , \wBIn79[30] , 
        \wBIn79[29] , \wBIn79[28] , \wBIn79[27] , \wBIn79[26] , \wBIn79[25] , 
        \wBIn79[24] , \wBIn79[23] , \wBIn79[22] , \wBIn79[21] , \wBIn79[20] , 
        \wBIn79[19] , \wBIn79[18] , \wBIn79[17] , \wBIn79[16] , \wBIn79[15] , 
        \wBIn79[14] , \wBIn79[13] , \wBIn79[12] , \wBIn79[11] , \wBIn79[10] , 
        \wBIn79[9] , \wBIn79[8] , \wBIn79[7] , \wBIn79[6] , \wBIn79[5] , 
        \wBIn79[4] , \wBIn79[3] , \wBIn79[2] , \wBIn79[1] , \wBIn79[0] }), 
        .HiOut({\wBMid78[31] , \wBMid78[30] , \wBMid78[29] , \wBMid78[28] , 
        \wBMid78[27] , \wBMid78[26] , \wBMid78[25] , \wBMid78[24] , 
        \wBMid78[23] , \wBMid78[22] , \wBMid78[21] , \wBMid78[20] , 
        \wBMid78[19] , \wBMid78[18] , \wBMid78[17] , \wBMid78[16] , 
        \wBMid78[15] , \wBMid78[14] , \wBMid78[13] , \wBMid78[12] , 
        \wBMid78[11] , \wBMid78[10] , \wBMid78[9] , \wBMid78[8] , \wBMid78[7] , 
        \wBMid78[6] , \wBMid78[5] , \wBMid78[4] , \wBMid78[3] , \wBMid78[2] , 
        \wBMid78[1] , \wBMid78[0] }), .LoOut({\wAMid79[31] , \wAMid79[30] , 
        \wAMid79[29] , \wAMid79[28] , \wAMid79[27] , \wAMid79[26] , 
        \wAMid79[25] , \wAMid79[24] , \wAMid79[23] , \wAMid79[22] , 
        \wAMid79[21] , \wAMid79[20] , \wAMid79[19] , \wAMid79[18] , 
        \wAMid79[17] , \wAMid79[16] , \wAMid79[15] , \wAMid79[14] , 
        \wAMid79[13] , \wAMid79[12] , \wAMid79[11] , \wAMid79[10] , 
        \wAMid79[9] , \wAMid79[8] , \wAMid79[7] , \wAMid79[6] , \wAMid79[5] , 
        \wAMid79[4] , \wAMid79[3] , \wAMid79[2] , \wAMid79[1] , \wAMid79[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn109[31] , \wAIn109[30] , \wAIn109[29] , \wAIn109[28] , 
        \wAIn109[27] , \wAIn109[26] , \wAIn109[25] , \wAIn109[24] , 
        \wAIn109[23] , \wAIn109[22] , \wAIn109[21] , \wAIn109[20] , 
        \wAIn109[19] , \wAIn109[18] , \wAIn109[17] , \wAIn109[16] , 
        \wAIn109[15] , \wAIn109[14] , \wAIn109[13] , \wAIn109[12] , 
        \wAIn109[11] , \wAIn109[10] , \wAIn109[9] , \wAIn109[8] , \wAIn109[7] , 
        \wAIn109[6] , \wAIn109[5] , \wAIn109[4] , \wAIn109[3] , \wAIn109[2] , 
        \wAIn109[1] , \wAIn109[0] }), .BIn({\wBIn109[31] , \wBIn109[30] , 
        \wBIn109[29] , \wBIn109[28] , \wBIn109[27] , \wBIn109[26] , 
        \wBIn109[25] , \wBIn109[24] , \wBIn109[23] , \wBIn109[22] , 
        \wBIn109[21] , \wBIn109[20] , \wBIn109[19] , \wBIn109[18] , 
        \wBIn109[17] , \wBIn109[16] , \wBIn109[15] , \wBIn109[14] , 
        \wBIn109[13] , \wBIn109[12] , \wBIn109[11] , \wBIn109[10] , 
        \wBIn109[9] , \wBIn109[8] , \wBIn109[7] , \wBIn109[6] , \wBIn109[5] , 
        \wBIn109[4] , \wBIn109[3] , \wBIn109[2] , \wBIn109[1] , \wBIn109[0] }), 
        .HiOut({\wBMid108[31] , \wBMid108[30] , \wBMid108[29] , \wBMid108[28] , 
        \wBMid108[27] , \wBMid108[26] , \wBMid108[25] , \wBMid108[24] , 
        \wBMid108[23] , \wBMid108[22] , \wBMid108[21] , \wBMid108[20] , 
        \wBMid108[19] , \wBMid108[18] , \wBMid108[17] , \wBMid108[16] , 
        \wBMid108[15] , \wBMid108[14] , \wBMid108[13] , \wBMid108[12] , 
        \wBMid108[11] , \wBMid108[10] , \wBMid108[9] , \wBMid108[8] , 
        \wBMid108[7] , \wBMid108[6] , \wBMid108[5] , \wBMid108[4] , 
        \wBMid108[3] , \wBMid108[2] , \wBMid108[1] , \wBMid108[0] }), .LoOut({
        \wAMid109[31] , \wAMid109[30] , \wAMid109[29] , \wAMid109[28] , 
        \wAMid109[27] , \wAMid109[26] , \wAMid109[25] , \wAMid109[24] , 
        \wAMid109[23] , \wAMid109[22] , \wAMid109[21] , \wAMid109[20] , 
        \wAMid109[19] , \wAMid109[18] , \wAMid109[17] , \wAMid109[16] , 
        \wAMid109[15] , \wAMid109[14] , \wAMid109[13] , \wAMid109[12] , 
        \wAMid109[11] , \wAMid109[10] , \wAMid109[9] , \wAMid109[8] , 
        \wAMid109[7] , \wAMid109[6] , \wAMid109[5] , \wAMid109[4] , 
        \wAMid109[3] , \wAMid109[2] , \wAMid109[1] , \wAMid109[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn112[31] , \wAIn112[30] , \wAIn112[29] , \wAIn112[28] , 
        \wAIn112[27] , \wAIn112[26] , \wAIn112[25] , \wAIn112[24] , 
        \wAIn112[23] , \wAIn112[22] , \wAIn112[21] , \wAIn112[20] , 
        \wAIn112[19] , \wAIn112[18] , \wAIn112[17] , \wAIn112[16] , 
        \wAIn112[15] , \wAIn112[14] , \wAIn112[13] , \wAIn112[12] , 
        \wAIn112[11] , \wAIn112[10] , \wAIn112[9] , \wAIn112[8] , \wAIn112[7] , 
        \wAIn112[6] , \wAIn112[5] , \wAIn112[4] , \wAIn112[3] , \wAIn112[2] , 
        \wAIn112[1] , \wAIn112[0] }), .BIn({\wBIn112[31] , \wBIn112[30] , 
        \wBIn112[29] , \wBIn112[28] , \wBIn112[27] , \wBIn112[26] , 
        \wBIn112[25] , \wBIn112[24] , \wBIn112[23] , \wBIn112[22] , 
        \wBIn112[21] , \wBIn112[20] , \wBIn112[19] , \wBIn112[18] , 
        \wBIn112[17] , \wBIn112[16] , \wBIn112[15] , \wBIn112[14] , 
        \wBIn112[13] , \wBIn112[12] , \wBIn112[11] , \wBIn112[10] , 
        \wBIn112[9] , \wBIn112[8] , \wBIn112[7] , \wBIn112[6] , \wBIn112[5] , 
        \wBIn112[4] , \wBIn112[3] , \wBIn112[2] , \wBIn112[1] , \wBIn112[0] }), 
        .HiOut({\wBMid111[31] , \wBMid111[30] , \wBMid111[29] , \wBMid111[28] , 
        \wBMid111[27] , \wBMid111[26] , \wBMid111[25] , \wBMid111[24] , 
        \wBMid111[23] , \wBMid111[22] , \wBMid111[21] , \wBMid111[20] , 
        \wBMid111[19] , \wBMid111[18] , \wBMid111[17] , \wBMid111[16] , 
        \wBMid111[15] , \wBMid111[14] , \wBMid111[13] , \wBMid111[12] , 
        \wBMid111[11] , \wBMid111[10] , \wBMid111[9] , \wBMid111[8] , 
        \wBMid111[7] , \wBMid111[6] , \wBMid111[5] , \wBMid111[4] , 
        \wBMid111[3] , \wBMid111[2] , \wBMid111[1] , \wBMid111[0] }), .LoOut({
        \wAMid112[31] , \wAMid112[30] , \wAMid112[29] , \wAMid112[28] , 
        \wAMid112[27] , \wAMid112[26] , \wAMid112[25] , \wAMid112[24] , 
        \wAMid112[23] , \wAMid112[22] , \wAMid112[21] , \wAMid112[20] , 
        \wAMid112[19] , \wAMid112[18] , \wAMid112[17] , \wAMid112[16] , 
        \wAMid112[15] , \wAMid112[14] , \wAMid112[13] , \wAMid112[12] , 
        \wAMid112[11] , \wAMid112[10] , \wAMid112[9] , \wAMid112[8] , 
        \wAMid112[7] , \wAMid112[6] , \wAMid112[5] , \wAMid112[4] , 
        \wAMid112[3] , \wAMid112[2] , \wAMid112[1] , \wAMid112[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid103[31] , \wAMid103[30] , \wAMid103[29] , \wAMid103[28] , 
        \wAMid103[27] , \wAMid103[26] , \wAMid103[25] , \wAMid103[24] , 
        \wAMid103[23] , \wAMid103[22] , \wAMid103[21] , \wAMid103[20] , 
        \wAMid103[19] , \wAMid103[18] , \wAMid103[17] , \wAMid103[16] , 
        \wAMid103[15] , \wAMid103[14] , \wAMid103[13] , \wAMid103[12] , 
        \wAMid103[11] , \wAMid103[10] , \wAMid103[9] , \wAMid103[8] , 
        \wAMid103[7] , \wAMid103[6] , \wAMid103[5] , \wAMid103[4] , 
        \wAMid103[3] , \wAMid103[2] , \wAMid103[1] , \wAMid103[0] }), .BIn({
        \wBMid103[31] , \wBMid103[30] , \wBMid103[29] , \wBMid103[28] , 
        \wBMid103[27] , \wBMid103[26] , \wBMid103[25] , \wBMid103[24] , 
        \wBMid103[23] , \wBMid103[22] , \wBMid103[21] , \wBMid103[20] , 
        \wBMid103[19] , \wBMid103[18] , \wBMid103[17] , \wBMid103[16] , 
        \wBMid103[15] , \wBMid103[14] , \wBMid103[13] , \wBMid103[12] , 
        \wBMid103[11] , \wBMid103[10] , \wBMid103[9] , \wBMid103[8] , 
        \wBMid103[7] , \wBMid103[6] , \wBMid103[5] , \wBMid103[4] , 
        \wBMid103[3] , \wBMid103[2] , \wBMid103[1] , \wBMid103[0] }), .HiOut({
        \wRegInB103[31] , \wRegInB103[30] , \wRegInB103[29] , \wRegInB103[28] , 
        \wRegInB103[27] , \wRegInB103[26] , \wRegInB103[25] , \wRegInB103[24] , 
        \wRegInB103[23] , \wRegInB103[22] , \wRegInB103[21] , \wRegInB103[20] , 
        \wRegInB103[19] , \wRegInB103[18] , \wRegInB103[17] , \wRegInB103[16] , 
        \wRegInB103[15] , \wRegInB103[14] , \wRegInB103[13] , \wRegInB103[12] , 
        \wRegInB103[11] , \wRegInB103[10] , \wRegInB103[9] , \wRegInB103[8] , 
        \wRegInB103[7] , \wRegInB103[6] , \wRegInB103[5] , \wRegInB103[4] , 
        \wRegInB103[3] , \wRegInB103[2] , \wRegInB103[1] , \wRegInB103[0] }), 
        .LoOut({\wRegInA104[31] , \wRegInA104[30] , \wRegInA104[29] , 
        \wRegInA104[28] , \wRegInA104[27] , \wRegInA104[26] , \wRegInA104[25] , 
        \wRegInA104[24] , \wRegInA104[23] , \wRegInA104[22] , \wRegInA104[21] , 
        \wRegInA104[20] , \wRegInA104[19] , \wRegInA104[18] , \wRegInA104[17] , 
        \wRegInA104[16] , \wRegInA104[15] , \wRegInA104[14] , \wRegInA104[13] , 
        \wRegInA104[12] , \wRegInA104[11] , \wRegInA104[10] , \wRegInA104[9] , 
        \wRegInA104[8] , \wRegInA104[7] , \wRegInA104[6] , \wRegInA104[5] , 
        \wRegInA104[4] , \wRegInA104[3] , \wRegInA104[2] , \wRegInA104[1] , 
        \wRegInA104[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid118[31] , \wAMid118[30] , \wAMid118[29] , \wAMid118[28] , 
        \wAMid118[27] , \wAMid118[26] , \wAMid118[25] , \wAMid118[24] , 
        \wAMid118[23] , \wAMid118[22] , \wAMid118[21] , \wAMid118[20] , 
        \wAMid118[19] , \wAMid118[18] , \wAMid118[17] , \wAMid118[16] , 
        \wAMid118[15] , \wAMid118[14] , \wAMid118[13] , \wAMid118[12] , 
        \wAMid118[11] , \wAMid118[10] , \wAMid118[9] , \wAMid118[8] , 
        \wAMid118[7] , \wAMid118[6] , \wAMid118[5] , \wAMid118[4] , 
        \wAMid118[3] , \wAMid118[2] , \wAMid118[1] , \wAMid118[0] }), .BIn({
        \wBMid118[31] , \wBMid118[30] , \wBMid118[29] , \wBMid118[28] , 
        \wBMid118[27] , \wBMid118[26] , \wBMid118[25] , \wBMid118[24] , 
        \wBMid118[23] , \wBMid118[22] , \wBMid118[21] , \wBMid118[20] , 
        \wBMid118[19] , \wBMid118[18] , \wBMid118[17] , \wBMid118[16] , 
        \wBMid118[15] , \wBMid118[14] , \wBMid118[13] , \wBMid118[12] , 
        \wBMid118[11] , \wBMid118[10] , \wBMid118[9] , \wBMid118[8] , 
        \wBMid118[7] , \wBMid118[6] , \wBMid118[5] , \wBMid118[4] , 
        \wBMid118[3] , \wBMid118[2] , \wBMid118[1] , \wBMid118[0] }), .HiOut({
        \wRegInB118[31] , \wRegInB118[30] , \wRegInB118[29] , \wRegInB118[28] , 
        \wRegInB118[27] , \wRegInB118[26] , \wRegInB118[25] , \wRegInB118[24] , 
        \wRegInB118[23] , \wRegInB118[22] , \wRegInB118[21] , \wRegInB118[20] , 
        \wRegInB118[19] , \wRegInB118[18] , \wRegInB118[17] , \wRegInB118[16] , 
        \wRegInB118[15] , \wRegInB118[14] , \wRegInB118[13] , \wRegInB118[12] , 
        \wRegInB118[11] , \wRegInB118[10] , \wRegInB118[9] , \wRegInB118[8] , 
        \wRegInB118[7] , \wRegInB118[6] , \wRegInB118[5] , \wRegInB118[4] , 
        \wRegInB118[3] , \wRegInB118[2] , \wRegInB118[1] , \wRegInB118[0] }), 
        .LoOut({\wRegInA119[31] , \wRegInA119[30] , \wRegInA119[29] , 
        \wRegInA119[28] , \wRegInA119[27] , \wRegInA119[26] , \wRegInA119[25] , 
        \wRegInA119[24] , \wRegInA119[23] , \wRegInA119[22] , \wRegInA119[21] , 
        \wRegInA119[20] , \wRegInA119[19] , \wRegInA119[18] , \wRegInA119[17] , 
        \wRegInA119[16] , \wRegInA119[15] , \wRegInA119[14] , \wRegInA119[13] , 
        \wRegInA119[12] , \wRegInA119[11] , \wRegInA119[10] , \wRegInA119[9] , 
        \wRegInA119[8] , \wRegInA119[7] , \wRegInA119[6] , \wRegInA119[5] , 
        \wRegInA119[4] , \wRegInA119[3] , \wRegInA119[2] , \wRegInA119[1] , 
        \wRegInA119[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid124[31] , \wAMid124[30] , \wAMid124[29] , \wAMid124[28] , 
        \wAMid124[27] , \wAMid124[26] , \wAMid124[25] , \wAMid124[24] , 
        \wAMid124[23] , \wAMid124[22] , \wAMid124[21] , \wAMid124[20] , 
        \wAMid124[19] , \wAMid124[18] , \wAMid124[17] , \wAMid124[16] , 
        \wAMid124[15] , \wAMid124[14] , \wAMid124[13] , \wAMid124[12] , 
        \wAMid124[11] , \wAMid124[10] , \wAMid124[9] , \wAMid124[8] , 
        \wAMid124[7] , \wAMid124[6] , \wAMid124[5] , \wAMid124[4] , 
        \wAMid124[3] , \wAMid124[2] , \wAMid124[1] , \wAMid124[0] }), .BIn({
        \wBMid124[31] , \wBMid124[30] , \wBMid124[29] , \wBMid124[28] , 
        \wBMid124[27] , \wBMid124[26] , \wBMid124[25] , \wBMid124[24] , 
        \wBMid124[23] , \wBMid124[22] , \wBMid124[21] , \wBMid124[20] , 
        \wBMid124[19] , \wBMid124[18] , \wBMid124[17] , \wBMid124[16] , 
        \wBMid124[15] , \wBMid124[14] , \wBMid124[13] , \wBMid124[12] , 
        \wBMid124[11] , \wBMid124[10] , \wBMid124[9] , \wBMid124[8] , 
        \wBMid124[7] , \wBMid124[6] , \wBMid124[5] , \wBMid124[4] , 
        \wBMid124[3] , \wBMid124[2] , \wBMid124[1] , \wBMid124[0] }), .HiOut({
        \wRegInB124[31] , \wRegInB124[30] , \wRegInB124[29] , \wRegInB124[28] , 
        \wRegInB124[27] , \wRegInB124[26] , \wRegInB124[25] , \wRegInB124[24] , 
        \wRegInB124[23] , \wRegInB124[22] , \wRegInB124[21] , \wRegInB124[20] , 
        \wRegInB124[19] , \wRegInB124[18] , \wRegInB124[17] , \wRegInB124[16] , 
        \wRegInB124[15] , \wRegInB124[14] , \wRegInB124[13] , \wRegInB124[12] , 
        \wRegInB124[11] , \wRegInB124[10] , \wRegInB124[9] , \wRegInB124[8] , 
        \wRegInB124[7] , \wRegInB124[6] , \wRegInB124[5] , \wRegInB124[4] , 
        \wRegInB124[3] , \wRegInB124[2] , \wRegInB124[1] , \wRegInB124[0] }), 
        .LoOut({\wRegInA125[31] , \wRegInA125[30] , \wRegInA125[29] , 
        \wRegInA125[28] , \wRegInA125[27] , \wRegInA125[26] , \wRegInA125[25] , 
        \wRegInA125[24] , \wRegInA125[23] , \wRegInA125[22] , \wRegInA125[21] , 
        \wRegInA125[20] , \wRegInA125[19] , \wRegInA125[18] , \wRegInA125[17] , 
        \wRegInA125[16] , \wRegInA125[15] , \wRegInA125[14] , \wRegInA125[13] , 
        \wRegInA125[12] , \wRegInA125[11] , \wRegInA125[10] , \wRegInA125[9] , 
        \wRegInA125[8] , \wRegInA125[7] , \wRegInA125[6] , \wRegInA125[5] , 
        \wRegInA125[4] , \wRegInA125[3] , \wRegInA125[2] , \wRegInA125[1] , 
        \wRegInA125[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_80 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink81[31] , \ScanLink81[30] , \ScanLink81[29] , 
        \ScanLink81[28] , \ScanLink81[27] , \ScanLink81[26] , \ScanLink81[25] , 
        \ScanLink81[24] , \ScanLink81[23] , \ScanLink81[22] , \ScanLink81[21] , 
        \ScanLink81[20] , \ScanLink81[19] , \ScanLink81[18] , \ScanLink81[17] , 
        \ScanLink81[16] , \ScanLink81[15] , \ScanLink81[14] , \ScanLink81[13] , 
        \ScanLink81[12] , \ScanLink81[11] , \ScanLink81[10] , \ScanLink81[9] , 
        \ScanLink81[8] , \ScanLink81[7] , \ScanLink81[6] , \ScanLink81[5] , 
        \ScanLink81[4] , \ScanLink81[3] , \ScanLink81[2] , \ScanLink81[1] , 
        \ScanLink81[0] }), .ScanOut({\ScanLink80[31] , \ScanLink80[30] , 
        \ScanLink80[29] , \ScanLink80[28] , \ScanLink80[27] , \ScanLink80[26] , 
        \ScanLink80[25] , \ScanLink80[24] , \ScanLink80[23] , \ScanLink80[22] , 
        \ScanLink80[21] , \ScanLink80[20] , \ScanLink80[19] , \ScanLink80[18] , 
        \ScanLink80[17] , \ScanLink80[16] , \ScanLink80[15] , \ScanLink80[14] , 
        \ScanLink80[13] , \ScanLink80[12] , \ScanLink80[11] , \ScanLink80[10] , 
        \ScanLink80[9] , \ScanLink80[8] , \ScanLink80[7] , \ScanLink80[6] , 
        \ScanLink80[5] , \ScanLink80[4] , \ScanLink80[3] , \ScanLink80[2] , 
        \ScanLink80[1] , \ScanLink80[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB87[31] , \wRegInB87[30] , 
        \wRegInB87[29] , \wRegInB87[28] , \wRegInB87[27] , \wRegInB87[26] , 
        \wRegInB87[25] , \wRegInB87[24] , \wRegInB87[23] , \wRegInB87[22] , 
        \wRegInB87[21] , \wRegInB87[20] , \wRegInB87[19] , \wRegInB87[18] , 
        \wRegInB87[17] , \wRegInB87[16] , \wRegInB87[15] , \wRegInB87[14] , 
        \wRegInB87[13] , \wRegInB87[12] , \wRegInB87[11] , \wRegInB87[10] , 
        \wRegInB87[9] , \wRegInB87[8] , \wRegInB87[7] , \wRegInB87[6] , 
        \wRegInB87[5] , \wRegInB87[4] , \wRegInB87[3] , \wRegInB87[2] , 
        \wRegInB87[1] , \wRegInB87[0] }), .Out({\wBIn87[31] , \wBIn87[30] , 
        \wBIn87[29] , \wBIn87[28] , \wBIn87[27] , \wBIn87[26] , \wBIn87[25] , 
        \wBIn87[24] , \wBIn87[23] , \wBIn87[22] , \wBIn87[21] , \wBIn87[20] , 
        \wBIn87[19] , \wBIn87[18] , \wBIn87[17] , \wBIn87[16] , \wBIn87[15] , 
        \wBIn87[14] , \wBIn87[13] , \wBIn87[12] , \wBIn87[11] , \wBIn87[10] , 
        \wBIn87[9] , \wBIn87[8] , \wBIn87[7] , \wBIn87[6] , \wBIn87[5] , 
        \wBIn87[4] , \wBIn87[3] , \wBIn87[2] , \wBIn87[1] , \wBIn87[0] }) );
    BubbleSort_Control_CWIDTH8_IDWIDTH1_WIDTH32_SCAN1 U_BSC ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink256[31] , 
        \ScanLink256[30] , \ScanLink256[29] , \ScanLink256[28] , 
        \ScanLink256[27] , \ScanLink256[26] , \ScanLink256[25] , 
        \ScanLink256[24] , \ScanLink256[23] , \ScanLink256[22] , 
        \ScanLink256[21] , \ScanLink256[20] , \ScanLink256[19] , 
        \ScanLink256[18] , \ScanLink256[17] , \ScanLink256[16] , 
        \ScanLink256[15] , \ScanLink256[14] , \ScanLink256[13] , 
        \ScanLink256[12] , \ScanLink256[11] , \ScanLink256[10] , 
        \ScanLink256[9] , \ScanLink256[8] , \ScanLink256[7] , \ScanLink256[6] , 
        \ScanLink256[5] , \ScanLink256[4] , \ScanLink256[3] , \ScanLink256[2] , 
        \ScanLink256[1] , \ScanLink256[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b0), .Id(1'b1), .Enable(\wEnable[0] ) );
    BubbleSort_Node_WIDTH32 BSN2_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid49[31] , \wAMid49[30] , \wAMid49[29] , \wAMid49[28] , 
        \wAMid49[27] , \wAMid49[26] , \wAMid49[25] , \wAMid49[24] , 
        \wAMid49[23] , \wAMid49[22] , \wAMid49[21] , \wAMid49[20] , 
        \wAMid49[19] , \wAMid49[18] , \wAMid49[17] , \wAMid49[16] , 
        \wAMid49[15] , \wAMid49[14] , \wAMid49[13] , \wAMid49[12] , 
        \wAMid49[11] , \wAMid49[10] , \wAMid49[9] , \wAMid49[8] , \wAMid49[7] , 
        \wAMid49[6] , \wAMid49[5] , \wAMid49[4] , \wAMid49[3] , \wAMid49[2] , 
        \wAMid49[1] , \wAMid49[0] }), .BIn({\wBMid49[31] , \wBMid49[30] , 
        \wBMid49[29] , \wBMid49[28] , \wBMid49[27] , \wBMid49[26] , 
        \wBMid49[25] , \wBMid49[24] , \wBMid49[23] , \wBMid49[22] , 
        \wBMid49[21] , \wBMid49[20] , \wBMid49[19] , \wBMid49[18] , 
        \wBMid49[17] , \wBMid49[16] , \wBMid49[15] , \wBMid49[14] , 
        \wBMid49[13] , \wBMid49[12] , \wBMid49[11] , \wBMid49[10] , 
        \wBMid49[9] , \wBMid49[8] , \wBMid49[7] , \wBMid49[6] , \wBMid49[5] , 
        \wBMid49[4] , \wBMid49[3] , \wBMid49[2] , \wBMid49[1] , \wBMid49[0] }), 
        .HiOut({\wRegInB49[31] , \wRegInB49[30] , \wRegInB49[29] , 
        \wRegInB49[28] , \wRegInB49[27] , \wRegInB49[26] , \wRegInB49[25] , 
        \wRegInB49[24] , \wRegInB49[23] , \wRegInB49[22] , \wRegInB49[21] , 
        \wRegInB49[20] , \wRegInB49[19] , \wRegInB49[18] , \wRegInB49[17] , 
        \wRegInB49[16] , \wRegInB49[15] , \wRegInB49[14] , \wRegInB49[13] , 
        \wRegInB49[12] , \wRegInB49[11] , \wRegInB49[10] , \wRegInB49[9] , 
        \wRegInB49[8] , \wRegInB49[7] , \wRegInB49[6] , \wRegInB49[5] , 
        \wRegInB49[4] , \wRegInB49[3] , \wRegInB49[2] , \wRegInB49[1] , 
        \wRegInB49[0] }), .LoOut({\wRegInA50[31] , \wRegInA50[30] , 
        \wRegInA50[29] , \wRegInA50[28] , \wRegInA50[27] , \wRegInA50[26] , 
        \wRegInA50[25] , \wRegInA50[24] , \wRegInA50[23] , \wRegInA50[22] , 
        \wRegInA50[21] , \wRegInA50[20] , \wRegInA50[19] , \wRegInA50[18] , 
        \wRegInA50[17] , \wRegInA50[16] , \wRegInA50[15] , \wRegInA50[14] , 
        \wRegInA50[13] , \wRegInA50[12] , \wRegInA50[11] , \wRegInA50[10] , 
        \wRegInA50[9] , \wRegInA50[8] , \wRegInA50[7] , \wRegInA50[6] , 
        \wRegInA50[5] , \wRegInA50[4] , \wRegInA50[3] , \wRegInA50[2] , 
        \wRegInA50[1] , \wRegInA50[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_222 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink223[31] , \ScanLink223[30] , \ScanLink223[29] , 
        \ScanLink223[28] , \ScanLink223[27] , \ScanLink223[26] , 
        \ScanLink223[25] , \ScanLink223[24] , \ScanLink223[23] , 
        \ScanLink223[22] , \ScanLink223[21] , \ScanLink223[20] , 
        \ScanLink223[19] , \ScanLink223[18] , \ScanLink223[17] , 
        \ScanLink223[16] , \ScanLink223[15] , \ScanLink223[14] , 
        \ScanLink223[13] , \ScanLink223[12] , \ScanLink223[11] , 
        \ScanLink223[10] , \ScanLink223[9] , \ScanLink223[8] , 
        \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , \ScanLink223[4] , 
        \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , \ScanLink223[0] 
        }), .ScanOut({\ScanLink222[31] , \ScanLink222[30] , \ScanLink222[29] , 
        \ScanLink222[28] , \ScanLink222[27] , \ScanLink222[26] , 
        \ScanLink222[25] , \ScanLink222[24] , \ScanLink222[23] , 
        \ScanLink222[22] , \ScanLink222[21] , \ScanLink222[20] , 
        \ScanLink222[19] , \ScanLink222[18] , \ScanLink222[17] , 
        \ScanLink222[16] , \ScanLink222[15] , \ScanLink222[14] , 
        \ScanLink222[13] , \ScanLink222[12] , \ScanLink222[11] , 
        \ScanLink222[10] , \ScanLink222[9] , \ScanLink222[8] , 
        \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , \ScanLink222[4] , 
        \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , \ScanLink222[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB16[31] , \wRegInB16[30] , \wRegInB16[29] , 
        \wRegInB16[28] , \wRegInB16[27] , \wRegInB16[26] , \wRegInB16[25] , 
        \wRegInB16[24] , \wRegInB16[23] , \wRegInB16[22] , \wRegInB16[21] , 
        \wRegInB16[20] , \wRegInB16[19] , \wRegInB16[18] , \wRegInB16[17] , 
        \wRegInB16[16] , \wRegInB16[15] , \wRegInB16[14] , \wRegInB16[13] , 
        \wRegInB16[12] , \wRegInB16[11] , \wRegInB16[10] , \wRegInB16[9] , 
        \wRegInB16[8] , \wRegInB16[7] , \wRegInB16[6] , \wRegInB16[5] , 
        \wRegInB16[4] , \wRegInB16[3] , \wRegInB16[2] , \wRegInB16[1] , 
        \wRegInB16[0] }), .Out({\wBIn16[31] , \wBIn16[30] , \wBIn16[29] , 
        \wBIn16[28] , \wBIn16[27] , \wBIn16[26] , \wBIn16[25] , \wBIn16[24] , 
        \wBIn16[23] , \wBIn16[22] , \wBIn16[21] , \wBIn16[20] , \wBIn16[19] , 
        \wBIn16[18] , \wBIn16[17] , \wBIn16[16] , \wBIn16[15] , \wBIn16[14] , 
        \wBIn16[13] , \wBIn16[12] , \wBIn16[11] , \wBIn16[10] , \wBIn16[9] , 
        \wBIn16[8] , \wBIn16[7] , \wBIn16[6] , \wBIn16[5] , \wBIn16[4] , 
        \wBIn16[3] , \wBIn16[2] , \wBIn16[1] , \wBIn16[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_205 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink206[31] , \ScanLink206[30] , \ScanLink206[29] , 
        \ScanLink206[28] , \ScanLink206[27] , \ScanLink206[26] , 
        \ScanLink206[25] , \ScanLink206[24] , \ScanLink206[23] , 
        \ScanLink206[22] , \ScanLink206[21] , \ScanLink206[20] , 
        \ScanLink206[19] , \ScanLink206[18] , \ScanLink206[17] , 
        \ScanLink206[16] , \ScanLink206[15] , \ScanLink206[14] , 
        \ScanLink206[13] , \ScanLink206[12] , \ScanLink206[11] , 
        \ScanLink206[10] , \ScanLink206[9] , \ScanLink206[8] , 
        \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , \ScanLink206[4] , 
        \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , \ScanLink206[0] 
        }), .ScanOut({\ScanLink205[31] , \ScanLink205[30] , \ScanLink205[29] , 
        \ScanLink205[28] , \ScanLink205[27] , \ScanLink205[26] , 
        \ScanLink205[25] , \ScanLink205[24] , \ScanLink205[23] , 
        \ScanLink205[22] , \ScanLink205[21] , \ScanLink205[20] , 
        \ScanLink205[19] , \ScanLink205[18] , \ScanLink205[17] , 
        \ScanLink205[16] , \ScanLink205[15] , \ScanLink205[14] , 
        \ScanLink205[13] , \ScanLink205[12] , \ScanLink205[11] , 
        \ScanLink205[10] , \ScanLink205[9] , \ScanLink205[8] , 
        \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , \ScanLink205[4] , 
        \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , \ScanLink205[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA25[31] , \wRegInA25[30] , \wRegInA25[29] , 
        \wRegInA25[28] , \wRegInA25[27] , \wRegInA25[26] , \wRegInA25[25] , 
        \wRegInA25[24] , \wRegInA25[23] , \wRegInA25[22] , \wRegInA25[21] , 
        \wRegInA25[20] , \wRegInA25[19] , \wRegInA25[18] , \wRegInA25[17] , 
        \wRegInA25[16] , \wRegInA25[15] , \wRegInA25[14] , \wRegInA25[13] , 
        \wRegInA25[12] , \wRegInA25[11] , \wRegInA25[10] , \wRegInA25[9] , 
        \wRegInA25[8] , \wRegInA25[7] , \wRegInA25[6] , \wRegInA25[5] , 
        \wRegInA25[4] , \wRegInA25[3] , \wRegInA25[2] , \wRegInA25[1] , 
        \wRegInA25[0] }), .Out({\wAIn25[31] , \wAIn25[30] , \wAIn25[29] , 
        \wAIn25[28] , \wAIn25[27] , \wAIn25[26] , \wAIn25[25] , \wAIn25[24] , 
        \wAIn25[23] , \wAIn25[22] , \wAIn25[21] , \wAIn25[20] , \wAIn25[19] , 
        \wAIn25[18] , \wAIn25[17] , \wAIn25[16] , \wAIn25[15] , \wAIn25[14] , 
        \wAIn25[13] , \wAIn25[12] , \wAIn25[11] , \wAIn25[10] , \wAIn25[9] , 
        \wAIn25[8] , \wAIn25[7] , \wAIn25[6] , \wAIn25[5] , \wAIn25[4] , 
        \wAIn25[3] , \wAIn25[2] , \wAIn25[1] , \wAIn25[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_135 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink136[31] , \ScanLink136[30] , \ScanLink136[29] , 
        \ScanLink136[28] , \ScanLink136[27] , \ScanLink136[26] , 
        \ScanLink136[25] , \ScanLink136[24] , \ScanLink136[23] , 
        \ScanLink136[22] , \ScanLink136[21] , \ScanLink136[20] , 
        \ScanLink136[19] , \ScanLink136[18] , \ScanLink136[17] , 
        \ScanLink136[16] , \ScanLink136[15] , \ScanLink136[14] , 
        \ScanLink136[13] , \ScanLink136[12] , \ScanLink136[11] , 
        \ScanLink136[10] , \ScanLink136[9] , \ScanLink136[8] , 
        \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , \ScanLink136[4] , 
        \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , \ScanLink136[0] 
        }), .ScanOut({\ScanLink135[31] , \ScanLink135[30] , \ScanLink135[29] , 
        \ScanLink135[28] , \ScanLink135[27] , \ScanLink135[26] , 
        \ScanLink135[25] , \ScanLink135[24] , \ScanLink135[23] , 
        \ScanLink135[22] , \ScanLink135[21] , \ScanLink135[20] , 
        \ScanLink135[19] , \ScanLink135[18] , \ScanLink135[17] , 
        \ScanLink135[16] , \ScanLink135[15] , \ScanLink135[14] , 
        \ScanLink135[13] , \ScanLink135[12] , \ScanLink135[11] , 
        \ScanLink135[10] , \ScanLink135[9] , \ScanLink135[8] , 
        \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , \ScanLink135[4] , 
        \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , \ScanLink135[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA60[31] , \wRegInA60[30] , \wRegInA60[29] , 
        \wRegInA60[28] , \wRegInA60[27] , \wRegInA60[26] , \wRegInA60[25] , 
        \wRegInA60[24] , \wRegInA60[23] , \wRegInA60[22] , \wRegInA60[21] , 
        \wRegInA60[20] , \wRegInA60[19] , \wRegInA60[18] , \wRegInA60[17] , 
        \wRegInA60[16] , \wRegInA60[15] , \wRegInA60[14] , \wRegInA60[13] , 
        \wRegInA60[12] , \wRegInA60[11] , \wRegInA60[10] , \wRegInA60[9] , 
        \wRegInA60[8] , \wRegInA60[7] , \wRegInA60[6] , \wRegInA60[5] , 
        \wRegInA60[4] , \wRegInA60[3] , \wRegInA60[2] , \wRegInA60[1] , 
        \wRegInA60[0] }), .Out({\wAIn60[31] , \wAIn60[30] , \wAIn60[29] , 
        \wAIn60[28] , \wAIn60[27] , \wAIn60[26] , \wAIn60[25] , \wAIn60[24] , 
        \wAIn60[23] , \wAIn60[22] , \wAIn60[21] , \wAIn60[20] , \wAIn60[19] , 
        \wAIn60[18] , \wAIn60[17] , \wAIn60[16] , \wAIn60[15] , \wAIn60[14] , 
        \wAIn60[13] , \wAIn60[12] , \wAIn60[11] , \wAIn60[10] , \wAIn60[9] , 
        \wAIn60[8] , \wAIn60[7] , \wAIn60[6] , \wAIn60[5] , \wAIn60[4] , 
        \wAIn60[3] , \wAIn60[2] , \wAIn60[1] , \wAIn60[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_65 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink66[31] , \ScanLink66[30] , \ScanLink66[29] , 
        \ScanLink66[28] , \ScanLink66[27] , \ScanLink66[26] , \ScanLink66[25] , 
        \ScanLink66[24] , \ScanLink66[23] , \ScanLink66[22] , \ScanLink66[21] , 
        \ScanLink66[20] , \ScanLink66[19] , \ScanLink66[18] , \ScanLink66[17] , 
        \ScanLink66[16] , \ScanLink66[15] , \ScanLink66[14] , \ScanLink66[13] , 
        \ScanLink66[12] , \ScanLink66[11] , \ScanLink66[10] , \ScanLink66[9] , 
        \ScanLink66[8] , \ScanLink66[7] , \ScanLink66[6] , \ScanLink66[5] , 
        \ScanLink66[4] , \ScanLink66[3] , \ScanLink66[2] , \ScanLink66[1] , 
        \ScanLink66[0] }), .ScanOut({\ScanLink65[31] , \ScanLink65[30] , 
        \ScanLink65[29] , \ScanLink65[28] , \ScanLink65[27] , \ScanLink65[26] , 
        \ScanLink65[25] , \ScanLink65[24] , \ScanLink65[23] , \ScanLink65[22] , 
        \ScanLink65[21] , \ScanLink65[20] , \ScanLink65[19] , \ScanLink65[18] , 
        \ScanLink65[17] , \ScanLink65[16] , \ScanLink65[15] , \ScanLink65[14] , 
        \ScanLink65[13] , \ScanLink65[12] , \ScanLink65[11] , \ScanLink65[10] , 
        \ScanLink65[9] , \ScanLink65[8] , \ScanLink65[7] , \ScanLink65[6] , 
        \ScanLink65[5] , \ScanLink65[4] , \ScanLink65[3] , \ScanLink65[2] , 
        \ScanLink65[1] , \ScanLink65[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA95[31] , \wRegInA95[30] , 
        \wRegInA95[29] , \wRegInA95[28] , \wRegInA95[27] , \wRegInA95[26] , 
        \wRegInA95[25] , \wRegInA95[24] , \wRegInA95[23] , \wRegInA95[22] , 
        \wRegInA95[21] , \wRegInA95[20] , \wRegInA95[19] , \wRegInA95[18] , 
        \wRegInA95[17] , \wRegInA95[16] , \wRegInA95[15] , \wRegInA95[14] , 
        \wRegInA95[13] , \wRegInA95[12] , \wRegInA95[11] , \wRegInA95[10] , 
        \wRegInA95[9] , \wRegInA95[8] , \wRegInA95[7] , \wRegInA95[6] , 
        \wRegInA95[5] , \wRegInA95[4] , \wRegInA95[3] , \wRegInA95[2] , 
        \wRegInA95[1] , \wRegInA95[0] }), .Out({\wAIn95[31] , \wAIn95[30] , 
        \wAIn95[29] , \wAIn95[28] , \wAIn95[27] , \wAIn95[26] , \wAIn95[25] , 
        \wAIn95[24] , \wAIn95[23] , \wAIn95[22] , \wAIn95[21] , \wAIn95[20] , 
        \wAIn95[19] , \wAIn95[18] , \wAIn95[17] , \wAIn95[16] , \wAIn95[15] , 
        \wAIn95[14] , \wAIn95[13] , \wAIn95[12] , \wAIn95[11] , \wAIn95[10] , 
        \wAIn95[9] , \wAIn95[8] , \wAIn95[7] , \wAIn95[6] , \wAIn95[5] , 
        \wAIn95[4] , \wAIn95[3] , \wAIn95[2] , \wAIn95[1] , \wAIn95[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_1 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA127[31] , \wRegInA127[30] , 
        \wRegInA127[29] , \wRegInA127[28] , \wRegInA127[27] , \wRegInA127[26] , 
        \wRegInA127[25] , \wRegInA127[24] , \wRegInA127[23] , \wRegInA127[22] , 
        \wRegInA127[21] , \wRegInA127[20] , \wRegInA127[19] , \wRegInA127[18] , 
        \wRegInA127[17] , \wRegInA127[16] , \wRegInA127[15] , \wRegInA127[14] , 
        \wRegInA127[13] , \wRegInA127[12] , \wRegInA127[11] , \wRegInA127[10] , 
        \wRegInA127[9] , \wRegInA127[8] , \wRegInA127[7] , \wRegInA127[6] , 
        \wRegInA127[5] , \wRegInA127[4] , \wRegInA127[3] , \wRegInA127[2] , 
        \wRegInA127[1] , \wRegInA127[0] }), .Out({\wAIn127[31] , \wAIn127[30] , 
        \wAIn127[29] , \wAIn127[28] , \wAIn127[27] , \wAIn127[26] , 
        \wAIn127[25] , \wAIn127[24] , \wAIn127[23] , \wAIn127[22] , 
        \wAIn127[21] , \wAIn127[20] , \wAIn127[19] , \wAIn127[18] , 
        \wAIn127[17] , \wAIn127[16] , \wAIn127[15] , \wAIn127[14] , 
        \wAIn127[13] , \wAIn127[12] , \wAIn127[11] , \wAIn127[10] , 
        \wAIn127[9] , \wAIn127[8] , \wAIn127[7] , \wAIn127[6] , \wAIn127[5] , 
        \wAIn127[4] , \wAIn127[3] , \wAIn127[2] , \wAIn127[1] , \wAIn127[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid20[31] , \wAMid20[30] , \wAMid20[29] , \wAMid20[28] , 
        \wAMid20[27] , \wAMid20[26] , \wAMid20[25] , \wAMid20[24] , 
        \wAMid20[23] , \wAMid20[22] , \wAMid20[21] , \wAMid20[20] , 
        \wAMid20[19] , \wAMid20[18] , \wAMid20[17] , \wAMid20[16] , 
        \wAMid20[15] , \wAMid20[14] , \wAMid20[13] , \wAMid20[12] , 
        \wAMid20[11] , \wAMid20[10] , \wAMid20[9] , \wAMid20[8] , \wAMid20[7] , 
        \wAMid20[6] , \wAMid20[5] , \wAMid20[4] , \wAMid20[3] , \wAMid20[2] , 
        \wAMid20[1] , \wAMid20[0] }), .BIn({\wBMid20[31] , \wBMid20[30] , 
        \wBMid20[29] , \wBMid20[28] , \wBMid20[27] , \wBMid20[26] , 
        \wBMid20[25] , \wBMid20[24] , \wBMid20[23] , \wBMid20[22] , 
        \wBMid20[21] , \wBMid20[20] , \wBMid20[19] , \wBMid20[18] , 
        \wBMid20[17] , \wBMid20[16] , \wBMid20[15] , \wBMid20[14] , 
        \wBMid20[13] , \wBMid20[12] , \wBMid20[11] , \wBMid20[10] , 
        \wBMid20[9] , \wBMid20[8] , \wBMid20[7] , \wBMid20[6] , \wBMid20[5] , 
        \wBMid20[4] , \wBMid20[3] , \wBMid20[2] , \wBMid20[1] , \wBMid20[0] }), 
        .HiOut({\wRegInB20[31] , \wRegInB20[30] , \wRegInB20[29] , 
        \wRegInB20[28] , \wRegInB20[27] , \wRegInB20[26] , \wRegInB20[25] , 
        \wRegInB20[24] , \wRegInB20[23] , \wRegInB20[22] , \wRegInB20[21] , 
        \wRegInB20[20] , \wRegInB20[19] , \wRegInB20[18] , \wRegInB20[17] , 
        \wRegInB20[16] , \wRegInB20[15] , \wRegInB20[14] , \wRegInB20[13] , 
        \wRegInB20[12] , \wRegInB20[11] , \wRegInB20[10] , \wRegInB20[9] , 
        \wRegInB20[8] , \wRegInB20[7] , \wRegInB20[6] , \wRegInB20[5] , 
        \wRegInB20[4] , \wRegInB20[3] , \wRegInB20[2] , \wRegInB20[1] , 
        \wRegInB20[0] }), .LoOut({\wRegInA21[31] , \wRegInA21[30] , 
        \wRegInA21[29] , \wRegInA21[28] , \wRegInA21[27] , \wRegInA21[26] , 
        \wRegInA21[25] , \wRegInA21[24] , \wRegInA21[23] , \wRegInA21[22] , 
        \wRegInA21[21] , \wRegInA21[20] , \wRegInA21[19] , \wRegInA21[18] , 
        \wRegInA21[17] , \wRegInA21[16] , \wRegInA21[15] , \wRegInA21[14] , 
        \wRegInA21[13] , \wRegInA21[12] , \wRegInA21[11] , \wRegInA21[10] , 
        \wRegInA21[9] , \wRegInA21[8] , \wRegInA21[7] , \wRegInA21[6] , 
        \wRegInA21[5] , \wRegInA21[4] , \wRegInA21[3] , \wRegInA21[2] , 
        \wRegInA21[1] , \wRegInA21[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid27[31] , \wAMid27[30] , \wAMid27[29] , \wAMid27[28] , 
        \wAMid27[27] , \wAMid27[26] , \wAMid27[25] , \wAMid27[24] , 
        \wAMid27[23] , \wAMid27[22] , \wAMid27[21] , \wAMid27[20] , 
        \wAMid27[19] , \wAMid27[18] , \wAMid27[17] , \wAMid27[16] , 
        \wAMid27[15] , \wAMid27[14] , \wAMid27[13] , \wAMid27[12] , 
        \wAMid27[11] , \wAMid27[10] , \wAMid27[9] , \wAMid27[8] , \wAMid27[7] , 
        \wAMid27[6] , \wAMid27[5] , \wAMid27[4] , \wAMid27[3] , \wAMid27[2] , 
        \wAMid27[1] , \wAMid27[0] }), .BIn({\wBMid27[31] , \wBMid27[30] , 
        \wBMid27[29] , \wBMid27[28] , \wBMid27[27] , \wBMid27[26] , 
        \wBMid27[25] , \wBMid27[24] , \wBMid27[23] , \wBMid27[22] , 
        \wBMid27[21] , \wBMid27[20] , \wBMid27[19] , \wBMid27[18] , 
        \wBMid27[17] , \wBMid27[16] , \wBMid27[15] , \wBMid27[14] , 
        \wBMid27[13] , \wBMid27[12] , \wBMid27[11] , \wBMid27[10] , 
        \wBMid27[9] , \wBMid27[8] , \wBMid27[7] , \wBMid27[6] , \wBMid27[5] , 
        \wBMid27[4] , \wBMid27[3] , \wBMid27[2] , \wBMid27[1] , \wBMid27[0] }), 
        .HiOut({\wRegInB27[31] , \wRegInB27[30] , \wRegInB27[29] , 
        \wRegInB27[28] , \wRegInB27[27] , \wRegInB27[26] , \wRegInB27[25] , 
        \wRegInB27[24] , \wRegInB27[23] , \wRegInB27[22] , \wRegInB27[21] , 
        \wRegInB27[20] , \wRegInB27[19] , \wRegInB27[18] , \wRegInB27[17] , 
        \wRegInB27[16] , \wRegInB27[15] , \wRegInB27[14] , \wRegInB27[13] , 
        \wRegInB27[12] , \wRegInB27[11] , \wRegInB27[10] , \wRegInB27[9] , 
        \wRegInB27[8] , \wRegInB27[7] , \wRegInB27[6] , \wRegInB27[5] , 
        \wRegInB27[4] , \wRegInB27[3] , \wRegInB27[2] , \wRegInB27[1] , 
        \wRegInB27[0] }), .LoOut({\wRegInA28[31] , \wRegInA28[30] , 
        \wRegInA28[29] , \wRegInA28[28] , \wRegInA28[27] , \wRegInA28[26] , 
        \wRegInA28[25] , \wRegInA28[24] , \wRegInA28[23] , \wRegInA28[22] , 
        \wRegInA28[21] , \wRegInA28[20] , \wRegInA28[19] , \wRegInA28[18] , 
        \wRegInA28[17] , \wRegInA28[16] , \wRegInA28[15] , \wRegInA28[14] , 
        \wRegInA28[13] , \wRegInA28[12] , \wRegInA28[11] , \wRegInA28[10] , 
        \wRegInA28[9] , \wRegInA28[8] , \wRegInA28[7] , \wRegInA28[6] , 
        \wRegInA28[5] , \wRegInA28[4] , \wRegInA28[3] , \wRegInA28[2] , 
        \wRegInA28[1] , \wRegInA28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_112 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink113[31] , \ScanLink113[30] , \ScanLink113[29] , 
        \ScanLink113[28] , \ScanLink113[27] , \ScanLink113[26] , 
        \ScanLink113[25] , \ScanLink113[24] , \ScanLink113[23] , 
        \ScanLink113[22] , \ScanLink113[21] , \ScanLink113[20] , 
        \ScanLink113[19] , \ScanLink113[18] , \ScanLink113[17] , 
        \ScanLink113[16] , \ScanLink113[15] , \ScanLink113[14] , 
        \ScanLink113[13] , \ScanLink113[12] , \ScanLink113[11] , 
        \ScanLink113[10] , \ScanLink113[9] , \ScanLink113[8] , 
        \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , \ScanLink113[4] , 
        \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , \ScanLink113[0] 
        }), .ScanOut({\ScanLink112[31] , \ScanLink112[30] , \ScanLink112[29] , 
        \ScanLink112[28] , \ScanLink112[27] , \ScanLink112[26] , 
        \ScanLink112[25] , \ScanLink112[24] , \ScanLink112[23] , 
        \ScanLink112[22] , \ScanLink112[21] , \ScanLink112[20] , 
        \ScanLink112[19] , \ScanLink112[18] , \ScanLink112[17] , 
        \ScanLink112[16] , \ScanLink112[15] , \ScanLink112[14] , 
        \ScanLink112[13] , \ScanLink112[12] , \ScanLink112[11] , 
        \ScanLink112[10] , \ScanLink112[9] , \ScanLink112[8] , 
        \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , \ScanLink112[4] , 
        \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , \ScanLink112[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB71[31] , \wRegInB71[30] , \wRegInB71[29] , 
        \wRegInB71[28] , \wRegInB71[27] , \wRegInB71[26] , \wRegInB71[25] , 
        \wRegInB71[24] , \wRegInB71[23] , \wRegInB71[22] , \wRegInB71[21] , 
        \wRegInB71[20] , \wRegInB71[19] , \wRegInB71[18] , \wRegInB71[17] , 
        \wRegInB71[16] , \wRegInB71[15] , \wRegInB71[14] , \wRegInB71[13] , 
        \wRegInB71[12] , \wRegInB71[11] , \wRegInB71[10] , \wRegInB71[9] , 
        \wRegInB71[8] , \wRegInB71[7] , \wRegInB71[6] , \wRegInB71[5] , 
        \wRegInB71[4] , \wRegInB71[3] , \wRegInB71[2] , \wRegInB71[1] , 
        \wRegInB71[0] }), .Out({\wBIn71[31] , \wBIn71[30] , \wBIn71[29] , 
        \wBIn71[28] , \wBIn71[27] , \wBIn71[26] , \wBIn71[25] , \wBIn71[24] , 
        \wBIn71[23] , \wBIn71[22] , \wBIn71[21] , \wBIn71[20] , \wBIn71[19] , 
        \wBIn71[18] , \wBIn71[17] , \wBIn71[16] , \wBIn71[15] , \wBIn71[14] , 
        \wBIn71[13] , \wBIn71[12] , \wBIn71[11] , \wBIn71[10] , \wBIn71[9] , 
        \wBIn71[8] , \wBIn71[7] , \wBIn71[6] , \wBIn71[5] , \wBIn71[4] , 
        \wBIn71[3] , \wBIn71[2] , \wBIn71[1] , \wBIn71[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_42 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink43[31] , \ScanLink43[30] , \ScanLink43[29] , 
        \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , \ScanLink43[25] , 
        \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , \ScanLink43[21] , 
        \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , \ScanLink43[17] , 
        \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , \ScanLink43[13] , 
        \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , \ScanLink43[9] , 
        \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , \ScanLink43[5] , 
        \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , \ScanLink43[1] , 
        \ScanLink43[0] }), .ScanOut({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB106[31] , \wRegInB106[30] , 
        \wRegInB106[29] , \wRegInB106[28] , \wRegInB106[27] , \wRegInB106[26] , 
        \wRegInB106[25] , \wRegInB106[24] , \wRegInB106[23] , \wRegInB106[22] , 
        \wRegInB106[21] , \wRegInB106[20] , \wRegInB106[19] , \wRegInB106[18] , 
        \wRegInB106[17] , \wRegInB106[16] , \wRegInB106[15] , \wRegInB106[14] , 
        \wRegInB106[13] , \wRegInB106[12] , \wRegInB106[11] , \wRegInB106[10] , 
        \wRegInB106[9] , \wRegInB106[8] , \wRegInB106[7] , \wRegInB106[6] , 
        \wRegInB106[5] , \wRegInB106[4] , \wRegInB106[3] , \wRegInB106[2] , 
        \wRegInB106[1] , \wRegInB106[0] }), .Out({\wBIn106[31] , \wBIn106[30] , 
        \wBIn106[29] , \wBIn106[28] , \wBIn106[27] , \wBIn106[26] , 
        \wBIn106[25] , \wBIn106[24] , \wBIn106[23] , \wBIn106[22] , 
        \wBIn106[21] , \wBIn106[20] , \wBIn106[19] , \wBIn106[18] , 
        \wBIn106[17] , \wBIn106[16] , \wBIn106[15] , \wBIn106[14] , 
        \wBIn106[13] , \wBIn106[12] , \wBIn106[11] , \wBIn106[10] , 
        \wBIn106[9] , \wBIn106[8] , \wBIn106[7] , \wBIn106[6] , \wBIn106[5] , 
        \wBIn106[4] , \wBIn106[3] , \wBIn106[2] , \wBIn106[1] , \wBIn106[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_199 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink200[31] , \ScanLink200[30] , \ScanLink200[29] , 
        \ScanLink200[28] , \ScanLink200[27] , \ScanLink200[26] , 
        \ScanLink200[25] , \ScanLink200[24] , \ScanLink200[23] , 
        \ScanLink200[22] , \ScanLink200[21] , \ScanLink200[20] , 
        \ScanLink200[19] , \ScanLink200[18] , \ScanLink200[17] , 
        \ScanLink200[16] , \ScanLink200[15] , \ScanLink200[14] , 
        \ScanLink200[13] , \ScanLink200[12] , \ScanLink200[11] , 
        \ScanLink200[10] , \ScanLink200[9] , \ScanLink200[8] , 
        \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , \ScanLink200[4] , 
        \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , \ScanLink200[0] 
        }), .ScanOut({\ScanLink199[31] , \ScanLink199[30] , \ScanLink199[29] , 
        \ScanLink199[28] , \ScanLink199[27] , \ScanLink199[26] , 
        \ScanLink199[25] , \ScanLink199[24] , \ScanLink199[23] , 
        \ScanLink199[22] , \ScanLink199[21] , \ScanLink199[20] , 
        \ScanLink199[19] , \ScanLink199[18] , \ScanLink199[17] , 
        \ScanLink199[16] , \ScanLink199[15] , \ScanLink199[14] , 
        \ScanLink199[13] , \ScanLink199[12] , \ScanLink199[11] , 
        \ScanLink199[10] , \ScanLink199[9] , \ScanLink199[8] , 
        \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , \ScanLink199[4] , 
        \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , \ScanLink199[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA28[31] , \wRegInA28[30] , \wRegInA28[29] , 
        \wRegInA28[28] , \wRegInA28[27] , \wRegInA28[26] , \wRegInA28[25] , 
        \wRegInA28[24] , \wRegInA28[23] , \wRegInA28[22] , \wRegInA28[21] , 
        \wRegInA28[20] , \wRegInA28[19] , \wRegInA28[18] , \wRegInA28[17] , 
        \wRegInA28[16] , \wRegInA28[15] , \wRegInA28[14] , \wRegInA28[13] , 
        \wRegInA28[12] , \wRegInA28[11] , \wRegInA28[10] , \wRegInA28[9] , 
        \wRegInA28[8] , \wRegInA28[7] , \wRegInA28[6] , \wRegInA28[5] , 
        \wRegInA28[4] , \wRegInA28[3] , \wRegInA28[2] , \wRegInA28[1] , 
        \wRegInA28[0] }), .Out({\wAIn28[31] , \wAIn28[30] , \wAIn28[29] , 
        \wAIn28[28] , \wAIn28[27] , \wAIn28[26] , \wAIn28[25] , \wAIn28[24] , 
        \wAIn28[23] , \wAIn28[22] , \wAIn28[21] , \wAIn28[20] , \wAIn28[19] , 
        \wAIn28[18] , \wAIn28[17] , \wAIn28[16] , \wAIn28[15] , \wAIn28[14] , 
        \wAIn28[13] , \wAIn28[12] , \wAIn28[11] , \wAIn28[10] , \wAIn28[9] , 
        \wAIn28[8] , \wAIn28[7] , \wAIn28[6] , \wAIn28[5] , \wAIn28[4] , 
        \wAIn28[3] , \wAIn28[2] , \wAIn28[1] , \wAIn28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_45 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink46[31] , \ScanLink46[30] , \ScanLink46[29] , 
        \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , \ScanLink46[25] , 
        \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , \ScanLink46[21] , 
        \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , \ScanLink46[17] , 
        \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , \ScanLink46[13] , 
        \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , \ScanLink46[9] , 
        \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , \ScanLink46[5] , 
        \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , \ScanLink46[1] , 
        \ScanLink46[0] }), .ScanOut({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA105[31] , \wRegInA105[30] , 
        \wRegInA105[29] , \wRegInA105[28] , \wRegInA105[27] , \wRegInA105[26] , 
        \wRegInA105[25] , \wRegInA105[24] , \wRegInA105[23] , \wRegInA105[22] , 
        \wRegInA105[21] , \wRegInA105[20] , \wRegInA105[19] , \wRegInA105[18] , 
        \wRegInA105[17] , \wRegInA105[16] , \wRegInA105[15] , \wRegInA105[14] , 
        \wRegInA105[13] , \wRegInA105[12] , \wRegInA105[11] , \wRegInA105[10] , 
        \wRegInA105[9] , \wRegInA105[8] , \wRegInA105[7] , \wRegInA105[6] , 
        \wRegInA105[5] , \wRegInA105[4] , \wRegInA105[3] , \wRegInA105[2] , 
        \wRegInA105[1] , \wRegInA105[0] }), .Out({\wAIn105[31] , \wAIn105[30] , 
        \wAIn105[29] , \wAIn105[28] , \wAIn105[27] , \wAIn105[26] , 
        \wAIn105[25] , \wAIn105[24] , \wAIn105[23] , \wAIn105[22] , 
        \wAIn105[21] , \wAIn105[20] , \wAIn105[19] , \wAIn105[18] , 
        \wAIn105[17] , \wAIn105[16] , \wAIn105[15] , \wAIn105[14] , 
        \wAIn105[13] , \wAIn105[12] , \wAIn105[11] , \wAIn105[10] , 
        \wAIn105[9] , \wAIn105[8] , \wAIn105[7] , \wAIn105[6] , \wAIn105[5] , 
        \wAIn105[4] , \wAIn105[3] , \wAIn105[2] , \wAIn105[1] , \wAIn105[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_115 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink116[31] , \ScanLink116[30] , \ScanLink116[29] , 
        \ScanLink116[28] , \ScanLink116[27] , \ScanLink116[26] , 
        \ScanLink116[25] , \ScanLink116[24] , \ScanLink116[23] , 
        \ScanLink116[22] , \ScanLink116[21] , \ScanLink116[20] , 
        \ScanLink116[19] , \ScanLink116[18] , \ScanLink116[17] , 
        \ScanLink116[16] , \ScanLink116[15] , \ScanLink116[14] , 
        \ScanLink116[13] , \ScanLink116[12] , \ScanLink116[11] , 
        \ScanLink116[10] , \ScanLink116[9] , \ScanLink116[8] , 
        \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , \ScanLink116[4] , 
        \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , \ScanLink116[0] 
        }), .ScanOut({\ScanLink115[31] , \ScanLink115[30] , \ScanLink115[29] , 
        \ScanLink115[28] , \ScanLink115[27] , \ScanLink115[26] , 
        \ScanLink115[25] , \ScanLink115[24] , \ScanLink115[23] , 
        \ScanLink115[22] , \ScanLink115[21] , \ScanLink115[20] , 
        \ScanLink115[19] , \ScanLink115[18] , \ScanLink115[17] , 
        \ScanLink115[16] , \ScanLink115[15] , \ScanLink115[14] , 
        \ScanLink115[13] , \ScanLink115[12] , \ScanLink115[11] , 
        \ScanLink115[10] , \ScanLink115[9] , \ScanLink115[8] , 
        \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , \ScanLink115[4] , 
        \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , \ScanLink115[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA70[31] , \wRegInA70[30] , \wRegInA70[29] , 
        \wRegInA70[28] , \wRegInA70[27] , \wRegInA70[26] , \wRegInA70[25] , 
        \wRegInA70[24] , \wRegInA70[23] , \wRegInA70[22] , \wRegInA70[21] , 
        \wRegInA70[20] , \wRegInA70[19] , \wRegInA70[18] , \wRegInA70[17] , 
        \wRegInA70[16] , \wRegInA70[15] , \wRegInA70[14] , \wRegInA70[13] , 
        \wRegInA70[12] , \wRegInA70[11] , \wRegInA70[10] , \wRegInA70[9] , 
        \wRegInA70[8] , \wRegInA70[7] , \wRegInA70[6] , \wRegInA70[5] , 
        \wRegInA70[4] , \wRegInA70[3] , \wRegInA70[2] , \wRegInA70[1] , 
        \wRegInA70[0] }), .Out({\wAIn70[31] , \wAIn70[30] , \wAIn70[29] , 
        \wAIn70[28] , \wAIn70[27] , \wAIn70[26] , \wAIn70[25] , \wAIn70[24] , 
        \wAIn70[23] , \wAIn70[22] , \wAIn70[21] , \wAIn70[20] , \wAIn70[19] , 
        \wAIn70[18] , \wAIn70[17] , \wAIn70[16] , \wAIn70[15] , \wAIn70[14] , 
        \wAIn70[13] , \wAIn70[12] , \wAIn70[11] , \wAIn70[10] , \wAIn70[9] , 
        \wAIn70[8] , \wAIn70[7] , \wAIn70[6] , \wAIn70[5] , \wAIn70[4] , 
        \wAIn70[3] , \wAIn70[2] , \wAIn70[1] , \wAIn70[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn37[31] , \wAIn37[30] , \wAIn37[29] , \wAIn37[28] , \wAIn37[27] , 
        \wAIn37[26] , \wAIn37[25] , \wAIn37[24] , \wAIn37[23] , \wAIn37[22] , 
        \wAIn37[21] , \wAIn37[20] , \wAIn37[19] , \wAIn37[18] , \wAIn37[17] , 
        \wAIn37[16] , \wAIn37[15] , \wAIn37[14] , \wAIn37[13] , \wAIn37[12] , 
        \wAIn37[11] , \wAIn37[10] , \wAIn37[9] , \wAIn37[8] , \wAIn37[7] , 
        \wAIn37[6] , \wAIn37[5] , \wAIn37[4] , \wAIn37[3] , \wAIn37[2] , 
        \wAIn37[1] , \wAIn37[0] }), .BIn({\wBIn37[31] , \wBIn37[30] , 
        \wBIn37[29] , \wBIn37[28] , \wBIn37[27] , \wBIn37[26] , \wBIn37[25] , 
        \wBIn37[24] , \wBIn37[23] , \wBIn37[22] , \wBIn37[21] , \wBIn37[20] , 
        \wBIn37[19] , \wBIn37[18] , \wBIn37[17] , \wBIn37[16] , \wBIn37[15] , 
        \wBIn37[14] , \wBIn37[13] , \wBIn37[12] , \wBIn37[11] , \wBIn37[10] , 
        \wBIn37[9] , \wBIn37[8] , \wBIn37[7] , \wBIn37[6] , \wBIn37[5] , 
        \wBIn37[4] , \wBIn37[3] , \wBIn37[2] , \wBIn37[1] , \wBIn37[0] }), 
        .HiOut({\wBMid36[31] , \wBMid36[30] , \wBMid36[29] , \wBMid36[28] , 
        \wBMid36[27] , \wBMid36[26] , \wBMid36[25] , \wBMid36[24] , 
        \wBMid36[23] , \wBMid36[22] , \wBMid36[21] , \wBMid36[20] , 
        \wBMid36[19] , \wBMid36[18] , \wBMid36[17] , \wBMid36[16] , 
        \wBMid36[15] , \wBMid36[14] , \wBMid36[13] , \wBMid36[12] , 
        \wBMid36[11] , \wBMid36[10] , \wBMid36[9] , \wBMid36[8] , \wBMid36[7] , 
        \wBMid36[6] , \wBMid36[5] , \wBMid36[4] , \wBMid36[3] , \wBMid36[2] , 
        \wBMid36[1] , \wBMid36[0] }), .LoOut({\wAMid37[31] , \wAMid37[30] , 
        \wAMid37[29] , \wAMid37[28] , \wAMid37[27] , \wAMid37[26] , 
        \wAMid37[25] , \wAMid37[24] , \wAMid37[23] , \wAMid37[22] , 
        \wAMid37[21] , \wAMid37[20] , \wAMid37[19] , \wAMid37[18] , 
        \wAMid37[17] , \wAMid37[16] , \wAMid37[15] , \wAMid37[14] , 
        \wAMid37[13] , \wAMid37[12] , \wAMid37[11] , \wAMid37[10] , 
        \wAMid37[9] , \wAMid37[8] , \wAMid37[7] , \wAMid37[6] , \wAMid37[5] , 
        \wAMid37[4] , \wAMid37[3] , \wAMid37[2] , \wAMid37[1] , \wAMid37[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_225 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink226[31] , \ScanLink226[30] , \ScanLink226[29] , 
        \ScanLink226[28] , \ScanLink226[27] , \ScanLink226[26] , 
        \ScanLink226[25] , \ScanLink226[24] , \ScanLink226[23] , 
        \ScanLink226[22] , \ScanLink226[21] , \ScanLink226[20] , 
        \ScanLink226[19] , \ScanLink226[18] , \ScanLink226[17] , 
        \ScanLink226[16] , \ScanLink226[15] , \ScanLink226[14] , 
        \ScanLink226[13] , \ScanLink226[12] , \ScanLink226[11] , 
        \ScanLink226[10] , \ScanLink226[9] , \ScanLink226[8] , 
        \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , \ScanLink226[4] , 
        \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , \ScanLink226[0] 
        }), .ScanOut({\ScanLink225[31] , \ScanLink225[30] , \ScanLink225[29] , 
        \ScanLink225[28] , \ScanLink225[27] , \ScanLink225[26] , 
        \ScanLink225[25] , \ScanLink225[24] , \ScanLink225[23] , 
        \ScanLink225[22] , \ScanLink225[21] , \ScanLink225[20] , 
        \ScanLink225[19] , \ScanLink225[18] , \ScanLink225[17] , 
        \ScanLink225[16] , \ScanLink225[15] , \ScanLink225[14] , 
        \ScanLink225[13] , \ScanLink225[12] , \ScanLink225[11] , 
        \ScanLink225[10] , \ScanLink225[9] , \ScanLink225[8] , 
        \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , \ScanLink225[4] , 
        \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , \ScanLink225[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA15[31] , \wRegInA15[30] , \wRegInA15[29] , 
        \wRegInA15[28] , \wRegInA15[27] , \wRegInA15[26] , \wRegInA15[25] , 
        \wRegInA15[24] , \wRegInA15[23] , \wRegInA15[22] , \wRegInA15[21] , 
        \wRegInA15[20] , \wRegInA15[19] , \wRegInA15[18] , \wRegInA15[17] , 
        \wRegInA15[16] , \wRegInA15[15] , \wRegInA15[14] , \wRegInA15[13] , 
        \wRegInA15[12] , \wRegInA15[11] , \wRegInA15[10] , \wRegInA15[9] , 
        \wRegInA15[8] , \wRegInA15[7] , \wRegInA15[6] , \wRegInA15[5] , 
        \wRegInA15[4] , \wRegInA15[3] , \wRegInA15[2] , \wRegInA15[1] , 
        \wRegInA15[0] }), .Out({\wAIn15[31] , \wAIn15[30] , \wAIn15[29] , 
        \wAIn15[28] , \wAIn15[27] , \wAIn15[26] , \wAIn15[25] , \wAIn15[24] , 
        \wAIn15[23] , \wAIn15[22] , \wAIn15[21] , \wAIn15[20] , \wAIn15[19] , 
        \wAIn15[18] , \wAIn15[17] , \wAIn15[16] , \wAIn15[15] , \wAIn15[14] , 
        \wAIn15[13] , \wAIn15[12] , \wAIn15[11] , \wAIn15[10] , \wAIn15[9] , 
        \wAIn15[8] , \wAIn15[7] , \wAIn15[6] , \wAIn15[5] , \wAIn15[4] , 
        \wAIn15[3] , \wAIn15[2] , \wAIn15[1] , \wAIn15[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_202 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink203[31] , \ScanLink203[30] , \ScanLink203[29] , 
        \ScanLink203[28] , \ScanLink203[27] , \ScanLink203[26] , 
        \ScanLink203[25] , \ScanLink203[24] , \ScanLink203[23] , 
        \ScanLink203[22] , \ScanLink203[21] , \ScanLink203[20] , 
        \ScanLink203[19] , \ScanLink203[18] , \ScanLink203[17] , 
        \ScanLink203[16] , \ScanLink203[15] , \ScanLink203[14] , 
        \ScanLink203[13] , \ScanLink203[12] , \ScanLink203[11] , 
        \ScanLink203[10] , \ScanLink203[9] , \ScanLink203[8] , 
        \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , \ScanLink203[4] , 
        \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , \ScanLink203[0] 
        }), .ScanOut({\ScanLink202[31] , \ScanLink202[30] , \ScanLink202[29] , 
        \ScanLink202[28] , \ScanLink202[27] , \ScanLink202[26] , 
        \ScanLink202[25] , \ScanLink202[24] , \ScanLink202[23] , 
        \ScanLink202[22] , \ScanLink202[21] , \ScanLink202[20] , 
        \ScanLink202[19] , \ScanLink202[18] , \ScanLink202[17] , 
        \ScanLink202[16] , \ScanLink202[15] , \ScanLink202[14] , 
        \ScanLink202[13] , \ScanLink202[12] , \ScanLink202[11] , 
        \ScanLink202[10] , \ScanLink202[9] , \ScanLink202[8] , 
        \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , \ScanLink202[4] , 
        \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , \ScanLink202[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB26[31] , \wRegInB26[30] , \wRegInB26[29] , 
        \wRegInB26[28] , \wRegInB26[27] , \wRegInB26[26] , \wRegInB26[25] , 
        \wRegInB26[24] , \wRegInB26[23] , \wRegInB26[22] , \wRegInB26[21] , 
        \wRegInB26[20] , \wRegInB26[19] , \wRegInB26[18] , \wRegInB26[17] , 
        \wRegInB26[16] , \wRegInB26[15] , \wRegInB26[14] , \wRegInB26[13] , 
        \wRegInB26[12] , \wRegInB26[11] , \wRegInB26[10] , \wRegInB26[9] , 
        \wRegInB26[8] , \wRegInB26[7] , \wRegInB26[6] , \wRegInB26[5] , 
        \wRegInB26[4] , \wRegInB26[3] , \wRegInB26[2] , \wRegInB26[1] , 
        \wRegInB26[0] }), .Out({\wBIn26[31] , \wBIn26[30] , \wBIn26[29] , 
        \wBIn26[28] , \wBIn26[27] , \wBIn26[26] , \wBIn26[25] , \wBIn26[24] , 
        \wBIn26[23] , \wBIn26[22] , \wBIn26[21] , \wBIn26[20] , \wBIn26[19] , 
        \wBIn26[18] , \wBIn26[17] , \wBIn26[16] , \wBIn26[15] , \wBIn26[14] , 
        \wBIn26[13] , \wBIn26[12] , \wBIn26[11] , \wBIn26[10] , \wBIn26[9] , 
        \wBIn26[8] , \wBIn26[7] , \wBIn26[6] , \wBIn26[5] , \wBIn26[4] , 
        \wBIn26[3] , \wBIn26[2] , \wBIn26[1] , \wBIn26[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_132 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink133[31] , \ScanLink133[30] , \ScanLink133[29] , 
        \ScanLink133[28] , \ScanLink133[27] , \ScanLink133[26] , 
        \ScanLink133[25] , \ScanLink133[24] , \ScanLink133[23] , 
        \ScanLink133[22] , \ScanLink133[21] , \ScanLink133[20] , 
        \ScanLink133[19] , \ScanLink133[18] , \ScanLink133[17] , 
        \ScanLink133[16] , \ScanLink133[15] , \ScanLink133[14] , 
        \ScanLink133[13] , \ScanLink133[12] , \ScanLink133[11] , 
        \ScanLink133[10] , \ScanLink133[9] , \ScanLink133[8] , 
        \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , \ScanLink133[4] , 
        \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , \ScanLink133[0] 
        }), .ScanOut({\ScanLink132[31] , \ScanLink132[30] , \ScanLink132[29] , 
        \ScanLink132[28] , \ScanLink132[27] , \ScanLink132[26] , 
        \ScanLink132[25] , \ScanLink132[24] , \ScanLink132[23] , 
        \ScanLink132[22] , \ScanLink132[21] , \ScanLink132[20] , 
        \ScanLink132[19] , \ScanLink132[18] , \ScanLink132[17] , 
        \ScanLink132[16] , \ScanLink132[15] , \ScanLink132[14] , 
        \ScanLink132[13] , \ScanLink132[12] , \ScanLink132[11] , 
        \ScanLink132[10] , \ScanLink132[9] , \ScanLink132[8] , 
        \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , \ScanLink132[4] , 
        \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , \ScanLink132[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB61[31] , \wRegInB61[30] , \wRegInB61[29] , 
        \wRegInB61[28] , \wRegInB61[27] , \wRegInB61[26] , \wRegInB61[25] , 
        \wRegInB61[24] , \wRegInB61[23] , \wRegInB61[22] , \wRegInB61[21] , 
        \wRegInB61[20] , \wRegInB61[19] , \wRegInB61[18] , \wRegInB61[17] , 
        \wRegInB61[16] , \wRegInB61[15] , \wRegInB61[14] , \wRegInB61[13] , 
        \wRegInB61[12] , \wRegInB61[11] , \wRegInB61[10] , \wRegInB61[9] , 
        \wRegInB61[8] , \wRegInB61[7] , \wRegInB61[6] , \wRegInB61[5] , 
        \wRegInB61[4] , \wRegInB61[3] , \wRegInB61[2] , \wRegInB61[1] , 
        \wRegInB61[0] }), .Out({\wBIn61[31] , \wBIn61[30] , \wBIn61[29] , 
        \wBIn61[28] , \wBIn61[27] , \wBIn61[26] , \wBIn61[25] , \wBIn61[24] , 
        \wBIn61[23] , \wBIn61[22] , \wBIn61[21] , \wBIn61[20] , \wBIn61[19] , 
        \wBIn61[18] , \wBIn61[17] , \wBIn61[16] , \wBIn61[15] , \wBIn61[14] , 
        \wBIn61[13] , \wBIn61[12] , \wBIn61[11] , \wBIn61[10] , \wBIn61[9] , 
        \wBIn61[8] , \wBIn61[7] , \wBIn61[6] , \wBIn61[5] , \wBIn61[4] , 
        \wBIn61[3] , \wBIn61[2] , \wBIn61[1] , \wBIn61[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_62 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink63[31] , \ScanLink63[30] , \ScanLink63[29] , 
        \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , \ScanLink63[25] , 
        \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , \ScanLink63[21] , 
        \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , \ScanLink63[17] , 
        \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , \ScanLink63[13] , 
        \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , \ScanLink63[9] , 
        \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , \ScanLink63[5] , 
        \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , \ScanLink63[1] , 
        \ScanLink63[0] }), .ScanOut({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB96[31] , \wRegInB96[30] , 
        \wRegInB96[29] , \wRegInB96[28] , \wRegInB96[27] , \wRegInB96[26] , 
        \wRegInB96[25] , \wRegInB96[24] , \wRegInB96[23] , \wRegInB96[22] , 
        \wRegInB96[21] , \wRegInB96[20] , \wRegInB96[19] , \wRegInB96[18] , 
        \wRegInB96[17] , \wRegInB96[16] , \wRegInB96[15] , \wRegInB96[14] , 
        \wRegInB96[13] , \wRegInB96[12] , \wRegInB96[11] , \wRegInB96[10] , 
        \wRegInB96[9] , \wRegInB96[8] , \wRegInB96[7] , \wRegInB96[6] , 
        \wRegInB96[5] , \wRegInB96[4] , \wRegInB96[3] , \wRegInB96[2] , 
        \wRegInB96[1] , \wRegInB96[0] }), .Out({\wBIn96[31] , \wBIn96[30] , 
        \wBIn96[29] , \wBIn96[28] , \wBIn96[27] , \wBIn96[26] , \wBIn96[25] , 
        \wBIn96[24] , \wBIn96[23] , \wBIn96[22] , \wBIn96[21] , \wBIn96[20] , 
        \wBIn96[19] , \wBIn96[18] , \wBIn96[17] , \wBIn96[16] , \wBIn96[15] , 
        \wBIn96[14] , \wBIn96[13] , \wBIn96[12] , \wBIn96[11] , \wBIn96[10] , 
        \wBIn96[9] , \wBIn96[8] , \wBIn96[7] , \wBIn96[6] , \wBIn96[5] , 
        \wBIn96[4] , \wBIn96[3] , \wBIn96[2] , \wBIn96[1] , \wBIn96[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_6 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[31] , \ScanLink7[30] , \ScanLink7[29] , 
        \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , \ScanLink7[25] , 
        \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , \ScanLink7[21] , 
        \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , \ScanLink7[17] , 
        \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , \ScanLink7[13] , 
        \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , \ScanLink7[9] , 
        \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB124[31] , \wRegInB124[30] , 
        \wRegInB124[29] , \wRegInB124[28] , \wRegInB124[27] , \wRegInB124[26] , 
        \wRegInB124[25] , \wRegInB124[24] , \wRegInB124[23] , \wRegInB124[22] , 
        \wRegInB124[21] , \wRegInB124[20] , \wRegInB124[19] , \wRegInB124[18] , 
        \wRegInB124[17] , \wRegInB124[16] , \wRegInB124[15] , \wRegInB124[14] , 
        \wRegInB124[13] , \wRegInB124[12] , \wRegInB124[11] , \wRegInB124[10] , 
        \wRegInB124[9] , \wRegInB124[8] , \wRegInB124[7] , \wRegInB124[6] , 
        \wRegInB124[5] , \wRegInB124[4] , \wRegInB124[3] , \wRegInB124[2] , 
        \wRegInB124[1] , \wRegInB124[0] }), .Out({\wBIn124[31] , \wBIn124[30] , 
        \wBIn124[29] , \wBIn124[28] , \wBIn124[27] , \wBIn124[26] , 
        \wBIn124[25] , \wBIn124[24] , \wBIn124[23] , \wBIn124[22] , 
        \wBIn124[21] , \wBIn124[20] , \wBIn124[19] , \wBIn124[18] , 
        \wBIn124[17] , \wBIn124[16] , \wBIn124[15] , \wBIn124[14] , 
        \wBIn124[13] , \wBIn124[12] , \wBIn124[11] , \wBIn124[10] , 
        \wBIn124[9] , \wBIn124[8] , \wBIn124[7] , \wBIn124[6] , \wBIn124[5] , 
        \wBIn124[4] , \wBIn124[3] , \wBIn124[2] , \wBIn124[1] , \wBIn124[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn42[31] , \wAIn42[30] , \wAIn42[29] , \wAIn42[28] , \wAIn42[27] , 
        \wAIn42[26] , \wAIn42[25] , \wAIn42[24] , \wAIn42[23] , \wAIn42[22] , 
        \wAIn42[21] , \wAIn42[20] , \wAIn42[19] , \wAIn42[18] , \wAIn42[17] , 
        \wAIn42[16] , \wAIn42[15] , \wAIn42[14] , \wAIn42[13] , \wAIn42[12] , 
        \wAIn42[11] , \wAIn42[10] , \wAIn42[9] , \wAIn42[8] , \wAIn42[7] , 
        \wAIn42[6] , \wAIn42[5] , \wAIn42[4] , \wAIn42[3] , \wAIn42[2] , 
        \wAIn42[1] , \wAIn42[0] }), .BIn({\wBIn42[31] , \wBIn42[30] , 
        \wBIn42[29] , \wBIn42[28] , \wBIn42[27] , \wBIn42[26] , \wBIn42[25] , 
        \wBIn42[24] , \wBIn42[23] , \wBIn42[22] , \wBIn42[21] , \wBIn42[20] , 
        \wBIn42[19] , \wBIn42[18] , \wBIn42[17] , \wBIn42[16] , \wBIn42[15] , 
        \wBIn42[14] , \wBIn42[13] , \wBIn42[12] , \wBIn42[11] , \wBIn42[10] , 
        \wBIn42[9] , \wBIn42[8] , \wBIn42[7] , \wBIn42[6] , \wBIn42[5] , 
        \wBIn42[4] , \wBIn42[3] , \wBIn42[2] , \wBIn42[1] , \wBIn42[0] }), 
        .HiOut({\wBMid41[31] , \wBMid41[30] , \wBMid41[29] , \wBMid41[28] , 
        \wBMid41[27] , \wBMid41[26] , \wBMid41[25] , \wBMid41[24] , 
        \wBMid41[23] , \wBMid41[22] , \wBMid41[21] , \wBMid41[20] , 
        \wBMid41[19] , \wBMid41[18] , \wBMid41[17] , \wBMid41[16] , 
        \wBMid41[15] , \wBMid41[14] , \wBMid41[13] , \wBMid41[12] , 
        \wBMid41[11] , \wBMid41[10] , \wBMid41[9] , \wBMid41[8] , \wBMid41[7] , 
        \wBMid41[6] , \wBMid41[5] , \wBMid41[4] , \wBMid41[3] , \wBMid41[2] , 
        \wBMid41[1] , \wBMid41[0] }), .LoOut({\wAMid42[31] , \wAMid42[30] , 
        \wAMid42[29] , \wAMid42[28] , \wAMid42[27] , \wAMid42[26] , 
        \wAMid42[25] , \wAMid42[24] , \wAMid42[23] , \wAMid42[22] , 
        \wAMid42[21] , \wAMid42[20] , \wAMid42[19] , \wAMid42[18] , 
        \wAMid42[17] , \wAMid42[16] , \wAMid42[15] , \wAMid42[14] , 
        \wAMid42[13] , \wAMid42[12] , \wAMid42[11] , \wAMid42[10] , 
        \wAMid42[9] , \wAMid42[8] , \wAMid42[7] , \wAMid42[6] , \wAMid42[5] , 
        \wAMid42[4] , \wAMid42[3] , \wAMid42[2] , \wAMid42[1] , \wAMid42[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn59[31] , \wAIn59[30] , \wAIn59[29] , \wAIn59[28] , \wAIn59[27] , 
        \wAIn59[26] , \wAIn59[25] , \wAIn59[24] , \wAIn59[23] , \wAIn59[22] , 
        \wAIn59[21] , \wAIn59[20] , \wAIn59[19] , \wAIn59[18] , \wAIn59[17] , 
        \wAIn59[16] , \wAIn59[15] , \wAIn59[14] , \wAIn59[13] , \wAIn59[12] , 
        \wAIn59[11] , \wAIn59[10] , \wAIn59[9] , \wAIn59[8] , \wAIn59[7] , 
        \wAIn59[6] , \wAIn59[5] , \wAIn59[4] , \wAIn59[3] , \wAIn59[2] , 
        \wAIn59[1] , \wAIn59[0] }), .BIn({\wBIn59[31] , \wBIn59[30] , 
        \wBIn59[29] , \wBIn59[28] , \wBIn59[27] , \wBIn59[26] , \wBIn59[25] , 
        \wBIn59[24] , \wBIn59[23] , \wBIn59[22] , \wBIn59[21] , \wBIn59[20] , 
        \wBIn59[19] , \wBIn59[18] , \wBIn59[17] , \wBIn59[16] , \wBIn59[15] , 
        \wBIn59[14] , \wBIn59[13] , \wBIn59[12] , \wBIn59[11] , \wBIn59[10] , 
        \wBIn59[9] , \wBIn59[8] , \wBIn59[7] , \wBIn59[6] , \wBIn59[5] , 
        \wBIn59[4] , \wBIn59[3] , \wBIn59[2] , \wBIn59[1] , \wBIn59[0] }), 
        .HiOut({\wBMid58[31] , \wBMid58[30] , \wBMid58[29] , \wBMid58[28] , 
        \wBMid58[27] , \wBMid58[26] , \wBMid58[25] , \wBMid58[24] , 
        \wBMid58[23] , \wBMid58[22] , \wBMid58[21] , \wBMid58[20] , 
        \wBMid58[19] , \wBMid58[18] , \wBMid58[17] , \wBMid58[16] , 
        \wBMid58[15] , \wBMid58[14] , \wBMid58[13] , \wBMid58[12] , 
        \wBMid58[11] , \wBMid58[10] , \wBMid58[9] , \wBMid58[8] , \wBMid58[7] , 
        \wBMid58[6] , \wBMid58[5] , \wBMid58[4] , \wBMid58[3] , \wBMid58[2] , 
        \wBMid58[1] , \wBMid58[0] }), .LoOut({\wAMid59[31] , \wAMid59[30] , 
        \wAMid59[29] , \wAMid59[28] , \wAMid59[27] , \wAMid59[26] , 
        \wAMid59[25] , \wAMid59[24] , \wAMid59[23] , \wAMid59[22] , 
        \wAMid59[21] , \wAMid59[20] , \wAMid59[19] , \wAMid59[18] , 
        \wAMid59[17] , \wAMid59[16] , \wAMid59[15] , \wAMid59[14] , 
        \wAMid59[13] , \wAMid59[12] , \wAMid59[11] , \wAMid59[10] , 
        \wAMid59[9] , \wAMid59[8] , \wAMid59[7] , \wAMid59[6] , \wAMid59[5] , 
        \wAMid59[4] , \wAMid59[3] , \wAMid59[2] , \wAMid59[1] , \wAMid59[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid69[31] , \wAMid69[30] , \wAMid69[29] , \wAMid69[28] , 
        \wAMid69[27] , \wAMid69[26] , \wAMid69[25] , \wAMid69[24] , 
        \wAMid69[23] , \wAMid69[22] , \wAMid69[21] , \wAMid69[20] , 
        \wAMid69[19] , \wAMid69[18] , \wAMid69[17] , \wAMid69[16] , 
        \wAMid69[15] , \wAMid69[14] , \wAMid69[13] , \wAMid69[12] , 
        \wAMid69[11] , \wAMid69[10] , \wAMid69[9] , \wAMid69[8] , \wAMid69[7] , 
        \wAMid69[6] , \wAMid69[5] , \wAMid69[4] , \wAMid69[3] , \wAMid69[2] , 
        \wAMid69[1] , \wAMid69[0] }), .BIn({\wBMid69[31] , \wBMid69[30] , 
        \wBMid69[29] , \wBMid69[28] , \wBMid69[27] , \wBMid69[26] , 
        \wBMid69[25] , \wBMid69[24] , \wBMid69[23] , \wBMid69[22] , 
        \wBMid69[21] , \wBMid69[20] , \wBMid69[19] , \wBMid69[18] , 
        \wBMid69[17] , \wBMid69[16] , \wBMid69[15] , \wBMid69[14] , 
        \wBMid69[13] , \wBMid69[12] , \wBMid69[11] , \wBMid69[10] , 
        \wBMid69[9] , \wBMid69[8] , \wBMid69[7] , \wBMid69[6] , \wBMid69[5] , 
        \wBMid69[4] , \wBMid69[3] , \wBMid69[2] , \wBMid69[1] , \wBMid69[0] }), 
        .HiOut({\wRegInB69[31] , \wRegInB69[30] , \wRegInB69[29] , 
        \wRegInB69[28] , \wRegInB69[27] , \wRegInB69[26] , \wRegInB69[25] , 
        \wRegInB69[24] , \wRegInB69[23] , \wRegInB69[22] , \wRegInB69[21] , 
        \wRegInB69[20] , \wRegInB69[19] , \wRegInB69[18] , \wRegInB69[17] , 
        \wRegInB69[16] , \wRegInB69[15] , \wRegInB69[14] , \wRegInB69[13] , 
        \wRegInB69[12] , \wRegInB69[11] , \wRegInB69[10] , \wRegInB69[9] , 
        \wRegInB69[8] , \wRegInB69[7] , \wRegInB69[6] , \wRegInB69[5] , 
        \wRegInB69[4] , \wRegInB69[3] , \wRegInB69[2] , \wRegInB69[1] , 
        \wRegInB69[0] }), .LoOut({\wRegInA70[31] , \wRegInA70[30] , 
        \wRegInA70[29] , \wRegInA70[28] , \wRegInA70[27] , \wRegInA70[26] , 
        \wRegInA70[25] , \wRegInA70[24] , \wRegInA70[23] , \wRegInA70[22] , 
        \wRegInA70[21] , \wRegInA70[20] , \wRegInA70[19] , \wRegInA70[18] , 
        \wRegInA70[17] , \wRegInA70[16] , \wRegInA70[15] , \wRegInA70[14] , 
        \wRegInA70[13] , \wRegInA70[12] , \wRegInA70[11] , \wRegInA70[10] , 
        \wRegInA70[9] , \wRegInA70[8] , \wRegInA70[7] , \wRegInA70[6] , 
        \wRegInA70[5] , \wRegInA70[4] , \wRegInA70[3] , \wRegInA70[2] , 
        \wRegInA70[1] , \wRegInA70[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid104[31] , \wAMid104[30] , \wAMid104[29] , \wAMid104[28] , 
        \wAMid104[27] , \wAMid104[26] , \wAMid104[25] , \wAMid104[24] , 
        \wAMid104[23] , \wAMid104[22] , \wAMid104[21] , \wAMid104[20] , 
        \wAMid104[19] , \wAMid104[18] , \wAMid104[17] , \wAMid104[16] , 
        \wAMid104[15] , \wAMid104[14] , \wAMid104[13] , \wAMid104[12] , 
        \wAMid104[11] , \wAMid104[10] , \wAMid104[9] , \wAMid104[8] , 
        \wAMid104[7] , \wAMid104[6] , \wAMid104[5] , \wAMid104[4] , 
        \wAMid104[3] , \wAMid104[2] , \wAMid104[1] , \wAMid104[0] }), .BIn({
        \wBMid104[31] , \wBMid104[30] , \wBMid104[29] , \wBMid104[28] , 
        \wBMid104[27] , \wBMid104[26] , \wBMid104[25] , \wBMid104[24] , 
        \wBMid104[23] , \wBMid104[22] , \wBMid104[21] , \wBMid104[20] , 
        \wBMid104[19] , \wBMid104[18] , \wBMid104[17] , \wBMid104[16] , 
        \wBMid104[15] , \wBMid104[14] , \wBMid104[13] , \wBMid104[12] , 
        \wBMid104[11] , \wBMid104[10] , \wBMid104[9] , \wBMid104[8] , 
        \wBMid104[7] , \wBMid104[6] , \wBMid104[5] , \wBMid104[4] , 
        \wBMid104[3] , \wBMid104[2] , \wBMid104[1] , \wBMid104[0] }), .HiOut({
        \wRegInB104[31] , \wRegInB104[30] , \wRegInB104[29] , \wRegInB104[28] , 
        \wRegInB104[27] , \wRegInB104[26] , \wRegInB104[25] , \wRegInB104[24] , 
        \wRegInB104[23] , \wRegInB104[22] , \wRegInB104[21] , \wRegInB104[20] , 
        \wRegInB104[19] , \wRegInB104[18] , \wRegInB104[17] , \wRegInB104[16] , 
        \wRegInB104[15] , \wRegInB104[14] , \wRegInB104[13] , \wRegInB104[12] , 
        \wRegInB104[11] , \wRegInB104[10] , \wRegInB104[9] , \wRegInB104[8] , 
        \wRegInB104[7] , \wRegInB104[6] , \wRegInB104[5] , \wRegInB104[4] , 
        \wRegInB104[3] , \wRegInB104[2] , \wRegInB104[1] , \wRegInB104[0] }), 
        .LoOut({\wRegInA105[31] , \wRegInA105[30] , \wRegInA105[29] , 
        \wRegInA105[28] , \wRegInA105[27] , \wRegInA105[26] , \wRegInA105[25] , 
        \wRegInA105[24] , \wRegInA105[23] , \wRegInA105[22] , \wRegInA105[21] , 
        \wRegInA105[20] , \wRegInA105[19] , \wRegInA105[18] , \wRegInA105[17] , 
        \wRegInA105[16] , \wRegInA105[15] , \wRegInA105[14] , \wRegInA105[13] , 
        \wRegInA105[12] , \wRegInA105[11] , \wRegInA105[10] , \wRegInA105[9] , 
        \wRegInA105[8] , \wRegInA105[7] , \wRegInA105[6] , \wRegInA105[5] , 
        \wRegInA105[4] , \wRegInA105[3] , \wRegInA105[2] , \wRegInA105[1] , 
        \wRegInA105[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid123[31] , \wAMid123[30] , \wAMid123[29] , \wAMid123[28] , 
        \wAMid123[27] , \wAMid123[26] , \wAMid123[25] , \wAMid123[24] , 
        \wAMid123[23] , \wAMid123[22] , \wAMid123[21] , \wAMid123[20] , 
        \wAMid123[19] , \wAMid123[18] , \wAMid123[17] , \wAMid123[16] , 
        \wAMid123[15] , \wAMid123[14] , \wAMid123[13] , \wAMid123[12] , 
        \wAMid123[11] , \wAMid123[10] , \wAMid123[9] , \wAMid123[8] , 
        \wAMid123[7] , \wAMid123[6] , \wAMid123[5] , \wAMid123[4] , 
        \wAMid123[3] , \wAMid123[2] , \wAMid123[1] , \wAMid123[0] }), .BIn({
        \wBMid123[31] , \wBMid123[30] , \wBMid123[29] , \wBMid123[28] , 
        \wBMid123[27] , \wBMid123[26] , \wBMid123[25] , \wBMid123[24] , 
        \wBMid123[23] , \wBMid123[22] , \wBMid123[21] , \wBMid123[20] , 
        \wBMid123[19] , \wBMid123[18] , \wBMid123[17] , \wBMid123[16] , 
        \wBMid123[15] , \wBMid123[14] , \wBMid123[13] , \wBMid123[12] , 
        \wBMid123[11] , \wBMid123[10] , \wBMid123[9] , \wBMid123[8] , 
        \wBMid123[7] , \wBMid123[6] , \wBMid123[5] , \wBMid123[4] , 
        \wBMid123[3] , \wBMid123[2] , \wBMid123[1] , \wBMid123[0] }), .HiOut({
        \wRegInB123[31] , \wRegInB123[30] , \wRegInB123[29] , \wRegInB123[28] , 
        \wRegInB123[27] , \wRegInB123[26] , \wRegInB123[25] , \wRegInB123[24] , 
        \wRegInB123[23] , \wRegInB123[22] , \wRegInB123[21] , \wRegInB123[20] , 
        \wRegInB123[19] , \wRegInB123[18] , \wRegInB123[17] , \wRegInB123[16] , 
        \wRegInB123[15] , \wRegInB123[14] , \wRegInB123[13] , \wRegInB123[12] , 
        \wRegInB123[11] , \wRegInB123[10] , \wRegInB123[9] , \wRegInB123[8] , 
        \wRegInB123[7] , \wRegInB123[6] , \wRegInB123[5] , \wRegInB123[4] , 
        \wRegInB123[3] , \wRegInB123[2] , \wRegInB123[1] , \wRegInB123[0] }), 
        .LoOut({\wRegInA124[31] , \wRegInA124[30] , \wRegInA124[29] , 
        \wRegInA124[28] , \wRegInA124[27] , \wRegInA124[26] , \wRegInA124[25] , 
        \wRegInA124[24] , \wRegInA124[23] , \wRegInA124[22] , \wRegInA124[21] , 
        \wRegInA124[20] , \wRegInA124[19] , \wRegInA124[18] , \wRegInA124[17] , 
        \wRegInA124[16] , \wRegInA124[15] , \wRegInA124[14] , \wRegInA124[13] , 
        \wRegInA124[12] , \wRegInA124[11] , \wRegInA124[10] , \wRegInA124[9] , 
        \wRegInA124[8] , \wRegInA124[7] , \wRegInA124[6] , \wRegInA124[5] , 
        \wRegInA124[4] , \wRegInA124[3] , \wRegInA124[2] , \wRegInA124[1] , 
        \wRegInA124[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_87 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink88[31] , \ScanLink88[30] , \ScanLink88[29] , 
        \ScanLink88[28] , \ScanLink88[27] , \ScanLink88[26] , \ScanLink88[25] , 
        \ScanLink88[24] , \ScanLink88[23] , \ScanLink88[22] , \ScanLink88[21] , 
        \ScanLink88[20] , \ScanLink88[19] , \ScanLink88[18] , \ScanLink88[17] , 
        \ScanLink88[16] , \ScanLink88[15] , \ScanLink88[14] , \ScanLink88[13] , 
        \ScanLink88[12] , \ScanLink88[11] , \ScanLink88[10] , \ScanLink88[9] , 
        \ScanLink88[8] , \ScanLink88[7] , \ScanLink88[6] , \ScanLink88[5] , 
        \ScanLink88[4] , \ScanLink88[3] , \ScanLink88[2] , \ScanLink88[1] , 
        \ScanLink88[0] }), .ScanOut({\ScanLink87[31] , \ScanLink87[30] , 
        \ScanLink87[29] , \ScanLink87[28] , \ScanLink87[27] , \ScanLink87[26] , 
        \ScanLink87[25] , \ScanLink87[24] , \ScanLink87[23] , \ScanLink87[22] , 
        \ScanLink87[21] , \ScanLink87[20] , \ScanLink87[19] , \ScanLink87[18] , 
        \ScanLink87[17] , \ScanLink87[16] , \ScanLink87[15] , \ScanLink87[14] , 
        \ScanLink87[13] , \ScanLink87[12] , \ScanLink87[11] , \ScanLink87[10] , 
        \ScanLink87[9] , \ScanLink87[8] , \ScanLink87[7] , \ScanLink87[6] , 
        \ScanLink87[5] , \ScanLink87[4] , \ScanLink87[3] , \ScanLink87[2] , 
        \ScanLink87[1] , \ScanLink87[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA84[31] , \wRegInA84[30] , 
        \wRegInA84[29] , \wRegInA84[28] , \wRegInA84[27] , \wRegInA84[26] , 
        \wRegInA84[25] , \wRegInA84[24] , \wRegInA84[23] , \wRegInA84[22] , 
        \wRegInA84[21] , \wRegInA84[20] , \wRegInA84[19] , \wRegInA84[18] , 
        \wRegInA84[17] , \wRegInA84[16] , \wRegInA84[15] , \wRegInA84[14] , 
        \wRegInA84[13] , \wRegInA84[12] , \wRegInA84[11] , \wRegInA84[10] , 
        \wRegInA84[9] , \wRegInA84[8] , \wRegInA84[7] , \wRegInA84[6] , 
        \wRegInA84[5] , \wRegInA84[4] , \wRegInA84[3] , \wRegInA84[2] , 
        \wRegInA84[1] , \wRegInA84[0] }), .Out({\wAIn84[31] , \wAIn84[30] , 
        \wAIn84[29] , \wAIn84[28] , \wAIn84[27] , \wAIn84[26] , \wAIn84[25] , 
        \wAIn84[24] , \wAIn84[23] , \wAIn84[22] , \wAIn84[21] , \wAIn84[20] , 
        \wAIn84[19] , \wAIn84[18] , \wAIn84[17] , \wAIn84[16] , \wAIn84[15] , 
        \wAIn84[14] , \wAIn84[13] , \wAIn84[12] , \wAIn84[11] , \wAIn84[10] , 
        \wAIn84[9] , \wAIn84[8] , \wAIn84[7] , \wAIn84[6] , \wAIn84[5] , 
        \wAIn84[4] , \wAIn84[3] , \wAIn84[2] , \wAIn84[1] , \wAIn84[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn65[31] , \wAIn65[30] , \wAIn65[29] , \wAIn65[28] , \wAIn65[27] , 
        \wAIn65[26] , \wAIn65[25] , \wAIn65[24] , \wAIn65[23] , \wAIn65[22] , 
        \wAIn65[21] , \wAIn65[20] , \wAIn65[19] , \wAIn65[18] , \wAIn65[17] , 
        \wAIn65[16] , \wAIn65[15] , \wAIn65[14] , \wAIn65[13] , \wAIn65[12] , 
        \wAIn65[11] , \wAIn65[10] , \wAIn65[9] , \wAIn65[8] , \wAIn65[7] , 
        \wAIn65[6] , \wAIn65[5] , \wAIn65[4] , \wAIn65[3] , \wAIn65[2] , 
        \wAIn65[1] , \wAIn65[0] }), .BIn({\wBIn65[31] , \wBIn65[30] , 
        \wBIn65[29] , \wBIn65[28] , \wBIn65[27] , \wBIn65[26] , \wBIn65[25] , 
        \wBIn65[24] , \wBIn65[23] , \wBIn65[22] , \wBIn65[21] , \wBIn65[20] , 
        \wBIn65[19] , \wBIn65[18] , \wBIn65[17] , \wBIn65[16] , \wBIn65[15] , 
        \wBIn65[14] , \wBIn65[13] , \wBIn65[12] , \wBIn65[11] , \wBIn65[10] , 
        \wBIn65[9] , \wBIn65[8] , \wBIn65[7] , \wBIn65[6] , \wBIn65[5] , 
        \wBIn65[4] , \wBIn65[3] , \wBIn65[2] , \wBIn65[1] , \wBIn65[0] }), 
        .HiOut({\wBMid64[31] , \wBMid64[30] , \wBMid64[29] , \wBMid64[28] , 
        \wBMid64[27] , \wBMid64[26] , \wBMid64[25] , \wBMid64[24] , 
        \wBMid64[23] , \wBMid64[22] , \wBMid64[21] , \wBMid64[20] , 
        \wBMid64[19] , \wBMid64[18] , \wBMid64[17] , \wBMid64[16] , 
        \wBMid64[15] , \wBMid64[14] , \wBMid64[13] , \wBMid64[12] , 
        \wBMid64[11] , \wBMid64[10] , \wBMid64[9] , \wBMid64[8] , \wBMid64[7] , 
        \wBMid64[6] , \wBMid64[5] , \wBMid64[4] , \wBMid64[3] , \wBMid64[2] , 
        \wBMid64[1] , \wBMid64[0] }), .LoOut({\wAMid65[31] , \wAMid65[30] , 
        \wAMid65[29] , \wAMid65[28] , \wAMid65[27] , \wAMid65[26] , 
        \wAMid65[25] , \wAMid65[24] , \wAMid65[23] , \wAMid65[22] , 
        \wAMid65[21] , \wAMid65[20] , \wAMid65[19] , \wAMid65[18] , 
        \wAMid65[17] , \wAMid65[16] , \wAMid65[15] , \wAMid65[14] , 
        \wAMid65[13] , \wAMid65[12] , \wAMid65[11] , \wAMid65[10] , 
        \wAMid65[9] , \wAMid65[8] , \wAMid65[7] , \wAMid65[6] , \wAMid65[5] , 
        \wAMid65[4] , \wAMid65[3] , \wAMid65[2] , \wAMid65[1] , \wAMid65[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn115[31] , \wAIn115[30] , \wAIn115[29] , \wAIn115[28] , 
        \wAIn115[27] , \wAIn115[26] , \wAIn115[25] , \wAIn115[24] , 
        \wAIn115[23] , \wAIn115[22] , \wAIn115[21] , \wAIn115[20] , 
        \wAIn115[19] , \wAIn115[18] , \wAIn115[17] , \wAIn115[16] , 
        \wAIn115[15] , \wAIn115[14] , \wAIn115[13] , \wAIn115[12] , 
        \wAIn115[11] , \wAIn115[10] , \wAIn115[9] , \wAIn115[8] , \wAIn115[7] , 
        \wAIn115[6] , \wAIn115[5] , \wAIn115[4] , \wAIn115[3] , \wAIn115[2] , 
        \wAIn115[1] , \wAIn115[0] }), .BIn({\wBIn115[31] , \wBIn115[30] , 
        \wBIn115[29] , \wBIn115[28] , \wBIn115[27] , \wBIn115[26] , 
        \wBIn115[25] , \wBIn115[24] , \wBIn115[23] , \wBIn115[22] , 
        \wBIn115[21] , \wBIn115[20] , \wBIn115[19] , \wBIn115[18] , 
        \wBIn115[17] , \wBIn115[16] , \wBIn115[15] , \wBIn115[14] , 
        \wBIn115[13] , \wBIn115[12] , \wBIn115[11] , \wBIn115[10] , 
        \wBIn115[9] , \wBIn115[8] , \wBIn115[7] , \wBIn115[6] , \wBIn115[5] , 
        \wBIn115[4] , \wBIn115[3] , \wBIn115[2] , \wBIn115[1] , \wBIn115[0] }), 
        .HiOut({\wBMid114[31] , \wBMid114[30] , \wBMid114[29] , \wBMid114[28] , 
        \wBMid114[27] , \wBMid114[26] , \wBMid114[25] , \wBMid114[24] , 
        \wBMid114[23] , \wBMid114[22] , \wBMid114[21] , \wBMid114[20] , 
        \wBMid114[19] , \wBMid114[18] , \wBMid114[17] , \wBMid114[16] , 
        \wBMid114[15] , \wBMid114[14] , \wBMid114[13] , \wBMid114[12] , 
        \wBMid114[11] , \wBMid114[10] , \wBMid114[9] , \wBMid114[8] , 
        \wBMid114[7] , \wBMid114[6] , \wBMid114[5] , \wBMid114[4] , 
        \wBMid114[3] , \wBMid114[2] , \wBMid114[1] , \wBMid114[0] }), .LoOut({
        \wAMid115[31] , \wAMid115[30] , \wAMid115[29] , \wAMid115[28] , 
        \wAMid115[27] , \wAMid115[26] , \wAMid115[25] , \wAMid115[24] , 
        \wAMid115[23] , \wAMid115[22] , \wAMid115[21] , \wAMid115[20] , 
        \wAMid115[19] , \wAMid115[18] , \wAMid115[17] , \wAMid115[16] , 
        \wAMid115[15] , \wAMid115[14] , \wAMid115[13] , \wAMid115[12] , 
        \wAMid115[11] , \wAMid115[10] , \wAMid115[9] , \wAMid115[8] , 
        \wAMid115[7] , \wAMid115[6] , \wAMid115[5] , \wAMid115[4] , 
        \wAMid115[3] , \wAMid115[2] , \wAMid115[1] , \wAMid115[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_250 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink251[31] , \ScanLink251[30] , \ScanLink251[29] , 
        \ScanLink251[28] , \ScanLink251[27] , \ScanLink251[26] , 
        \ScanLink251[25] , \ScanLink251[24] , \ScanLink251[23] , 
        \ScanLink251[22] , \ScanLink251[21] , \ScanLink251[20] , 
        \ScanLink251[19] , \ScanLink251[18] , \ScanLink251[17] , 
        \ScanLink251[16] , \ScanLink251[15] , \ScanLink251[14] , 
        \ScanLink251[13] , \ScanLink251[12] , \ScanLink251[11] , 
        \ScanLink251[10] , \ScanLink251[9] , \ScanLink251[8] , 
        \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , \ScanLink251[4] , 
        \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , \ScanLink251[0] 
        }), .ScanOut({\ScanLink250[31] , \ScanLink250[30] , \ScanLink250[29] , 
        \ScanLink250[28] , \ScanLink250[27] , \ScanLink250[26] , 
        \ScanLink250[25] , \ScanLink250[24] , \ScanLink250[23] , 
        \ScanLink250[22] , \ScanLink250[21] , \ScanLink250[20] , 
        \ScanLink250[19] , \ScanLink250[18] , \ScanLink250[17] , 
        \ScanLink250[16] , \ScanLink250[15] , \ScanLink250[14] , 
        \ScanLink250[13] , \ScanLink250[12] , \ScanLink250[11] , 
        \ScanLink250[10] , \ScanLink250[9] , \ScanLink250[8] , 
        \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , \ScanLink250[4] , 
        \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , \ScanLink250[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB2[31] , \wRegInB2[30] , \wRegInB2[29] , \wRegInB2[28] , 
        \wRegInB2[27] , \wRegInB2[26] , \wRegInB2[25] , \wRegInB2[24] , 
        \wRegInB2[23] , \wRegInB2[22] , \wRegInB2[21] , \wRegInB2[20] , 
        \wRegInB2[19] , \wRegInB2[18] , \wRegInB2[17] , \wRegInB2[16] , 
        \wRegInB2[15] , \wRegInB2[14] , \wRegInB2[13] , \wRegInB2[12] , 
        \wRegInB2[11] , \wRegInB2[10] , \wRegInB2[9] , \wRegInB2[8] , 
        \wRegInB2[7] , \wRegInB2[6] , \wRegInB2[5] , \wRegInB2[4] , 
        \wRegInB2[3] , \wRegInB2[2] , \wRegInB2[1] , \wRegInB2[0] }), .Out({
        \wBIn2[31] , \wBIn2[30] , \wBIn2[29] , \wBIn2[28] , \wBIn2[27] , 
        \wBIn2[26] , \wBIn2[25] , \wBIn2[24] , \wBIn2[23] , \wBIn2[22] , 
        \wBIn2[21] , \wBIn2[20] , \wBIn2[19] , \wBIn2[18] , \wBIn2[17] , 
        \wBIn2[16] , \wBIn2[15] , \wBIn2[14] , \wBIn2[13] , \wBIn2[12] , 
        \wBIn2[11] , \wBIn2[10] , \wBIn2[9] , \wBIn2[8] , \wBIn2[7] , 
        \wBIn2[6] , \wBIn2[5] , \wBIn2[4] , \wBIn2[3] , \wBIn2[2] , \wBIn2[1] , 
        \wBIn2[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid55[31] , \wAMid55[30] , \wAMid55[29] , \wAMid55[28] , 
        \wAMid55[27] , \wAMid55[26] , \wAMid55[25] , \wAMid55[24] , 
        \wAMid55[23] , \wAMid55[22] , \wAMid55[21] , \wAMid55[20] , 
        \wAMid55[19] , \wAMid55[18] , \wAMid55[17] , \wAMid55[16] , 
        \wAMid55[15] , \wAMid55[14] , \wAMid55[13] , \wAMid55[12] , 
        \wAMid55[11] , \wAMid55[10] , \wAMid55[9] , \wAMid55[8] , \wAMid55[7] , 
        \wAMid55[6] , \wAMid55[5] , \wAMid55[4] , \wAMid55[3] , \wAMid55[2] , 
        \wAMid55[1] , \wAMid55[0] }), .BIn({\wBMid55[31] , \wBMid55[30] , 
        \wBMid55[29] , \wBMid55[28] , \wBMid55[27] , \wBMid55[26] , 
        \wBMid55[25] , \wBMid55[24] , \wBMid55[23] , \wBMid55[22] , 
        \wBMid55[21] , \wBMid55[20] , \wBMid55[19] , \wBMid55[18] , 
        \wBMid55[17] , \wBMid55[16] , \wBMid55[15] , \wBMid55[14] , 
        \wBMid55[13] , \wBMid55[12] , \wBMid55[11] , \wBMid55[10] , 
        \wBMid55[9] , \wBMid55[8] , \wBMid55[7] , \wBMid55[6] , \wBMid55[5] , 
        \wBMid55[4] , \wBMid55[3] , \wBMid55[2] , \wBMid55[1] , \wBMid55[0] }), 
        .HiOut({\wRegInB55[31] , \wRegInB55[30] , \wRegInB55[29] , 
        \wRegInB55[28] , \wRegInB55[27] , \wRegInB55[26] , \wRegInB55[25] , 
        \wRegInB55[24] , \wRegInB55[23] , \wRegInB55[22] , \wRegInB55[21] , 
        \wRegInB55[20] , \wRegInB55[19] , \wRegInB55[18] , \wRegInB55[17] , 
        \wRegInB55[16] , \wRegInB55[15] , \wRegInB55[14] , \wRegInB55[13] , 
        \wRegInB55[12] , \wRegInB55[11] , \wRegInB55[10] , \wRegInB55[9] , 
        \wRegInB55[8] , \wRegInB55[7] , \wRegInB55[6] , \wRegInB55[5] , 
        \wRegInB55[4] , \wRegInB55[3] , \wRegInB55[2] , \wRegInB55[1] , 
        \wRegInB55[0] }), .LoOut({\wRegInA56[31] , \wRegInA56[30] , 
        \wRegInA56[29] , \wRegInA56[28] , \wRegInA56[27] , \wRegInA56[26] , 
        \wRegInA56[25] , \wRegInA56[24] , \wRegInA56[23] , \wRegInA56[22] , 
        \wRegInA56[21] , \wRegInA56[20] , \wRegInA56[19] , \wRegInA56[18] , 
        \wRegInA56[17] , \wRegInA56[16] , \wRegInA56[15] , \wRegInA56[14] , 
        \wRegInA56[13] , \wRegInA56[12] , \wRegInA56[11] , \wRegInA56[10] , 
        \wRegInA56[9] , \wRegInA56[8] , \wRegInA56[7] , \wRegInA56[6] , 
        \wRegInA56[5] , \wRegInA56[4] , \wRegInA56[3] , \wRegInA56[2] , 
        \wRegInA56[1] , \wRegInA56[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_30 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink31[31] , \ScanLink31[30] , \ScanLink31[29] , 
        \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , \ScanLink31[25] , 
        \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , \ScanLink31[21] , 
        \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , \ScanLink31[17] , 
        \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , \ScanLink31[13] , 
        \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , \ScanLink31[9] , 
        \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , \ScanLink31[5] , 
        \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , \ScanLink31[1] , 
        \ScanLink31[0] }), .ScanOut({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB112[31] , \wRegInB112[30] , 
        \wRegInB112[29] , \wRegInB112[28] , \wRegInB112[27] , \wRegInB112[26] , 
        \wRegInB112[25] , \wRegInB112[24] , \wRegInB112[23] , \wRegInB112[22] , 
        \wRegInB112[21] , \wRegInB112[20] , \wRegInB112[19] , \wRegInB112[18] , 
        \wRegInB112[17] , \wRegInB112[16] , \wRegInB112[15] , \wRegInB112[14] , 
        \wRegInB112[13] , \wRegInB112[12] , \wRegInB112[11] , \wRegInB112[10] , 
        \wRegInB112[9] , \wRegInB112[8] , \wRegInB112[7] , \wRegInB112[6] , 
        \wRegInB112[5] , \wRegInB112[4] , \wRegInB112[3] , \wRegInB112[2] , 
        \wRegInB112[1] , \wRegInB112[0] }), .Out({\wBIn112[31] , \wBIn112[30] , 
        \wBIn112[29] , \wBIn112[28] , \wBIn112[27] , \wBIn112[26] , 
        \wBIn112[25] , \wBIn112[24] , \wBIn112[23] , \wBIn112[22] , 
        \wBIn112[21] , \wBIn112[20] , \wBIn112[19] , \wBIn112[18] , 
        \wBIn112[17] , \wBIn112[16] , \wBIn112[15] , \wBIn112[14] , 
        \wBIn112[13] , \wBIn112[12] , \wBIn112[11] , \wBIn112[10] , 
        \wBIn112[9] , \wBIn112[8] , \wBIn112[7] , \wBIn112[6] , \wBIn112[5] , 
        \wBIn112[4] , \wBIn112[3] , \wBIn112[2] , \wBIn112[1] , \wBIn112[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_160 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink161[31] , \ScanLink161[30] , \ScanLink161[29] , 
        \ScanLink161[28] , \ScanLink161[27] , \ScanLink161[26] , 
        \ScanLink161[25] , \ScanLink161[24] , \ScanLink161[23] , 
        \ScanLink161[22] , \ScanLink161[21] , \ScanLink161[20] , 
        \ScanLink161[19] , \ScanLink161[18] , \ScanLink161[17] , 
        \ScanLink161[16] , \ScanLink161[15] , \ScanLink161[14] , 
        \ScanLink161[13] , \ScanLink161[12] , \ScanLink161[11] , 
        \ScanLink161[10] , \ScanLink161[9] , \ScanLink161[8] , 
        \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , \ScanLink161[4] , 
        \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , \ScanLink161[0] 
        }), .ScanOut({\ScanLink160[31] , \ScanLink160[30] , \ScanLink160[29] , 
        \ScanLink160[28] , \ScanLink160[27] , \ScanLink160[26] , 
        \ScanLink160[25] , \ScanLink160[24] , \ScanLink160[23] , 
        \ScanLink160[22] , \ScanLink160[21] , \ScanLink160[20] , 
        \ScanLink160[19] , \ScanLink160[18] , \ScanLink160[17] , 
        \ScanLink160[16] , \ScanLink160[15] , \ScanLink160[14] , 
        \ScanLink160[13] , \ScanLink160[12] , \ScanLink160[11] , 
        \ScanLink160[10] , \ScanLink160[9] , \ScanLink160[8] , 
        \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , \ScanLink160[4] , 
        \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , \ScanLink160[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB47[31] , \wRegInB47[30] , \wRegInB47[29] , 
        \wRegInB47[28] , \wRegInB47[27] , \wRegInB47[26] , \wRegInB47[25] , 
        \wRegInB47[24] , \wRegInB47[23] , \wRegInB47[22] , \wRegInB47[21] , 
        \wRegInB47[20] , \wRegInB47[19] , \wRegInB47[18] , \wRegInB47[17] , 
        \wRegInB47[16] , \wRegInB47[15] , \wRegInB47[14] , \wRegInB47[13] , 
        \wRegInB47[12] , \wRegInB47[11] , \wRegInB47[10] , \wRegInB47[9] , 
        \wRegInB47[8] , \wRegInB47[7] , \wRegInB47[6] , \wRegInB47[5] , 
        \wRegInB47[4] , \wRegInB47[3] , \wRegInB47[2] , \wRegInB47[1] , 
        \wRegInB47[0] }), .Out({\wBIn47[31] , \wBIn47[30] , \wBIn47[29] , 
        \wBIn47[28] , \wBIn47[27] , \wBIn47[26] , \wBIn47[25] , \wBIn47[24] , 
        \wBIn47[23] , \wBIn47[22] , \wBIn47[21] , \wBIn47[20] , \wBIn47[19] , 
        \wBIn47[18] , \wBIn47[17] , \wBIn47[16] , \wBIn47[15] , \wBIn47[14] , 
        \wBIn47[13] , \wBIn47[12] , \wBIn47[11] , \wBIn47[10] , \wBIn47[9] , 
        \wBIn47[8] , \wBIn47[7] , \wBIn47[6] , \wBIn47[5] , \wBIn47[4] , 
        \wBIn47[3] , \wBIn47[2] , \wBIn47[1] , \wBIn47[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid72[31] , \wAMid72[30] , \wAMid72[29] , \wAMid72[28] , 
        \wAMid72[27] , \wAMid72[26] , \wAMid72[25] , \wAMid72[24] , 
        \wAMid72[23] , \wAMid72[22] , \wAMid72[21] , \wAMid72[20] , 
        \wAMid72[19] , \wAMid72[18] , \wAMid72[17] , \wAMid72[16] , 
        \wAMid72[15] , \wAMid72[14] , \wAMid72[13] , \wAMid72[12] , 
        \wAMid72[11] , \wAMid72[10] , \wAMid72[9] , \wAMid72[8] , \wAMid72[7] , 
        \wAMid72[6] , \wAMid72[5] , \wAMid72[4] , \wAMid72[3] , \wAMid72[2] , 
        \wAMid72[1] , \wAMid72[0] }), .BIn({\wBMid72[31] , \wBMid72[30] , 
        \wBMid72[29] , \wBMid72[28] , \wBMid72[27] , \wBMid72[26] , 
        \wBMid72[25] , \wBMid72[24] , \wBMid72[23] , \wBMid72[22] , 
        \wBMid72[21] , \wBMid72[20] , \wBMid72[19] , \wBMid72[18] , 
        \wBMid72[17] , \wBMid72[16] , \wBMid72[15] , \wBMid72[14] , 
        \wBMid72[13] , \wBMid72[12] , \wBMid72[11] , \wBMid72[10] , 
        \wBMid72[9] , \wBMid72[8] , \wBMid72[7] , \wBMid72[6] , \wBMid72[5] , 
        \wBMid72[4] , \wBMid72[3] , \wBMid72[2] , \wBMid72[1] , \wBMid72[0] }), 
        .HiOut({\wRegInB72[31] , \wRegInB72[30] , \wRegInB72[29] , 
        \wRegInB72[28] , \wRegInB72[27] , \wRegInB72[26] , \wRegInB72[25] , 
        \wRegInB72[24] , \wRegInB72[23] , \wRegInB72[22] , \wRegInB72[21] , 
        \wRegInB72[20] , \wRegInB72[19] , \wRegInB72[18] , \wRegInB72[17] , 
        \wRegInB72[16] , \wRegInB72[15] , \wRegInB72[14] , \wRegInB72[13] , 
        \wRegInB72[12] , \wRegInB72[11] , \wRegInB72[10] , \wRegInB72[9] , 
        \wRegInB72[8] , \wRegInB72[7] , \wRegInB72[6] , \wRegInB72[5] , 
        \wRegInB72[4] , \wRegInB72[3] , \wRegInB72[2] , \wRegInB72[1] , 
        \wRegInB72[0] }), .LoOut({\wRegInA73[31] , \wRegInA73[30] , 
        \wRegInA73[29] , \wRegInA73[28] , \wRegInA73[27] , \wRegInA73[26] , 
        \wRegInA73[25] , \wRegInA73[24] , \wRegInA73[23] , \wRegInA73[22] , 
        \wRegInA73[21] , \wRegInA73[20] , \wRegInA73[19] , \wRegInA73[18] , 
        \wRegInA73[17] , \wRegInA73[16] , \wRegInA73[15] , \wRegInA73[14] , 
        \wRegInA73[13] , \wRegInA73[12] , \wRegInA73[11] , \wRegInA73[10] , 
        \wRegInA73[9] , \wRegInA73[8] , \wRegInA73[7] , \wRegInA73[6] , 
        \wRegInA73[5] , \wRegInA73[4] , \wRegInA73[3] , \wRegInA73[2] , 
        \wRegInA73[1] , \wRegInA73[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid97[31] , \wAMid97[30] , \wAMid97[29] , \wAMid97[28] , 
        \wAMid97[27] , \wAMid97[26] , \wAMid97[25] , \wAMid97[24] , 
        \wAMid97[23] , \wAMid97[22] , \wAMid97[21] , \wAMid97[20] , 
        \wAMid97[19] , \wAMid97[18] , \wAMid97[17] , \wAMid97[16] , 
        \wAMid97[15] , \wAMid97[14] , \wAMid97[13] , \wAMid97[12] , 
        \wAMid97[11] , \wAMid97[10] , \wAMid97[9] , \wAMid97[8] , \wAMid97[7] , 
        \wAMid97[6] , \wAMid97[5] , \wAMid97[4] , \wAMid97[3] , \wAMid97[2] , 
        \wAMid97[1] , \wAMid97[0] }), .BIn({\wBMid97[31] , \wBMid97[30] , 
        \wBMid97[29] , \wBMid97[28] , \wBMid97[27] , \wBMid97[26] , 
        \wBMid97[25] , \wBMid97[24] , \wBMid97[23] , \wBMid97[22] , 
        \wBMid97[21] , \wBMid97[20] , \wBMid97[19] , \wBMid97[18] , 
        \wBMid97[17] , \wBMid97[16] , \wBMid97[15] , \wBMid97[14] , 
        \wBMid97[13] , \wBMid97[12] , \wBMid97[11] , \wBMid97[10] , 
        \wBMid97[9] , \wBMid97[8] , \wBMid97[7] , \wBMid97[6] , \wBMid97[5] , 
        \wBMid97[4] , \wBMid97[3] , \wBMid97[2] , \wBMid97[1] , \wBMid97[0] }), 
        .HiOut({\wRegInB97[31] , \wRegInB97[30] , \wRegInB97[29] , 
        \wRegInB97[28] , \wRegInB97[27] , \wRegInB97[26] , \wRegInB97[25] , 
        \wRegInB97[24] , \wRegInB97[23] , \wRegInB97[22] , \wRegInB97[21] , 
        \wRegInB97[20] , \wRegInB97[19] , \wRegInB97[18] , \wRegInB97[17] , 
        \wRegInB97[16] , \wRegInB97[15] , \wRegInB97[14] , \wRegInB97[13] , 
        \wRegInB97[12] , \wRegInB97[11] , \wRegInB97[10] , \wRegInB97[9] , 
        \wRegInB97[8] , \wRegInB97[7] , \wRegInB97[6] , \wRegInB97[5] , 
        \wRegInB97[4] , \wRegInB97[3] , \wRegInB97[2] , \wRegInB97[1] , 
        \wRegInB97[0] }), .LoOut({\wRegInA98[31] , \wRegInA98[30] , 
        \wRegInA98[29] , \wRegInA98[28] , \wRegInA98[27] , \wRegInA98[26] , 
        \wRegInA98[25] , \wRegInA98[24] , \wRegInA98[23] , \wRegInA98[22] , 
        \wRegInA98[21] , \wRegInA98[20] , \wRegInA98[19] , \wRegInA98[18] , 
        \wRegInA98[17] , \wRegInA98[16] , \wRegInA98[15] , \wRegInA98[14] , 
        \wRegInA98[13] , \wRegInA98[12] , \wRegInA98[11] , \wRegInA98[10] , 
        \wRegInA98[9] , \wRegInA98[8] , \wRegInA98[7] , \wRegInA98[6] , 
        \wRegInA98[5] , \wRegInA98[4] , \wRegInA98[3] , \wRegInA98[2] , 
        \wRegInA98[1] , \wRegInA98[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_147 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink148[31] , \ScanLink148[30] , \ScanLink148[29] , 
        \ScanLink148[28] , \ScanLink148[27] , \ScanLink148[26] , 
        \ScanLink148[25] , \ScanLink148[24] , \ScanLink148[23] , 
        \ScanLink148[22] , \ScanLink148[21] , \ScanLink148[20] , 
        \ScanLink148[19] , \ScanLink148[18] , \ScanLink148[17] , 
        \ScanLink148[16] , \ScanLink148[15] , \ScanLink148[14] , 
        \ScanLink148[13] , \ScanLink148[12] , \ScanLink148[11] , 
        \ScanLink148[10] , \ScanLink148[9] , \ScanLink148[8] , 
        \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , \ScanLink148[4] , 
        \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , \ScanLink148[0] 
        }), .ScanOut({\ScanLink147[31] , \ScanLink147[30] , \ScanLink147[29] , 
        \ScanLink147[28] , \ScanLink147[27] , \ScanLink147[26] , 
        \ScanLink147[25] , \ScanLink147[24] , \ScanLink147[23] , 
        \ScanLink147[22] , \ScanLink147[21] , \ScanLink147[20] , 
        \ScanLink147[19] , \ScanLink147[18] , \ScanLink147[17] , 
        \ScanLink147[16] , \ScanLink147[15] , \ScanLink147[14] , 
        \ScanLink147[13] , \ScanLink147[12] , \ScanLink147[11] , 
        \ScanLink147[10] , \ScanLink147[9] , \ScanLink147[8] , 
        \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , \ScanLink147[4] , 
        \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , \ScanLink147[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA54[31] , \wRegInA54[30] , \wRegInA54[29] , 
        \wRegInA54[28] , \wRegInA54[27] , \wRegInA54[26] , \wRegInA54[25] , 
        \wRegInA54[24] , \wRegInA54[23] , \wRegInA54[22] , \wRegInA54[21] , 
        \wRegInA54[20] , \wRegInA54[19] , \wRegInA54[18] , \wRegInA54[17] , 
        \wRegInA54[16] , \wRegInA54[15] , \wRegInA54[14] , \wRegInA54[13] , 
        \wRegInA54[12] , \wRegInA54[11] , \wRegInA54[10] , \wRegInA54[9] , 
        \wRegInA54[8] , \wRegInA54[7] , \wRegInA54[6] , \wRegInA54[5] , 
        \wRegInA54[4] , \wRegInA54[3] , \wRegInA54[2] , \wRegInA54[1] , 
        \wRegInA54[0] }), .Out({\wAIn54[31] , \wAIn54[30] , \wAIn54[29] , 
        \wAIn54[28] , \wAIn54[27] , \wAIn54[26] , \wAIn54[25] , \wAIn54[24] , 
        \wAIn54[23] , \wAIn54[22] , \wAIn54[21] , \wAIn54[20] , \wAIn54[19] , 
        \wAIn54[18] , \wAIn54[17] , \wAIn54[16] , \wAIn54[15] , \wAIn54[14] , 
        \wAIn54[13] , \wAIn54[12] , \wAIn54[11] , \wAIn54[10] , \wAIn54[9] , 
        \wAIn54[8] , \wAIn54[7] , \wAIn54[6] , \wAIn54[5] , \wAIn54[4] , 
        \wAIn54[3] , \wAIn54[2] , \wAIn54[1] , \wAIn54[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_17 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink18[31] , \ScanLink18[30] , \ScanLink18[29] , 
        \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , \ScanLink18[25] , 
        \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , \ScanLink18[21] , 
        \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , \ScanLink18[17] , 
        \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , \ScanLink18[13] , 
        \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , \ScanLink18[9] , 
        \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , \ScanLink18[5] , 
        \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , \ScanLink18[1] , 
        \ScanLink18[0] }), .ScanOut({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA119[31] , \wRegInA119[30] , 
        \wRegInA119[29] , \wRegInA119[28] , \wRegInA119[27] , \wRegInA119[26] , 
        \wRegInA119[25] , \wRegInA119[24] , \wRegInA119[23] , \wRegInA119[22] , 
        \wRegInA119[21] , \wRegInA119[20] , \wRegInA119[19] , \wRegInA119[18] , 
        \wRegInA119[17] , \wRegInA119[16] , \wRegInA119[15] , \wRegInA119[14] , 
        \wRegInA119[13] , \wRegInA119[12] , \wRegInA119[11] , \wRegInA119[10] , 
        \wRegInA119[9] , \wRegInA119[8] , \wRegInA119[7] , \wRegInA119[6] , 
        \wRegInA119[5] , \wRegInA119[4] , \wRegInA119[3] , \wRegInA119[2] , 
        \wRegInA119[1] , \wRegInA119[0] }), .Out({\wAIn119[31] , \wAIn119[30] , 
        \wAIn119[29] , \wAIn119[28] , \wAIn119[27] , \wAIn119[26] , 
        \wAIn119[25] , \wAIn119[24] , \wAIn119[23] , \wAIn119[22] , 
        \wAIn119[21] , \wAIn119[20] , \wAIn119[19] , \wAIn119[18] , 
        \wAIn119[17] , \wAIn119[16] , \wAIn119[15] , \wAIn119[14] , 
        \wAIn119[13] , \wAIn119[12] , \wAIn119[11] , \wAIn119[10] , 
        \wAIn119[9] , \wAIn119[8] , \wAIn119[7] , \wAIn119[6] , \wAIn119[5] , 
        \wAIn119[4] , \wAIn119[3] , \wAIn119[2] , \wAIn119[1] , \wAIn119[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn19[31] , \wAIn19[30] , \wAIn19[29] , \wAIn19[28] , \wAIn19[27] , 
        \wAIn19[26] , \wAIn19[25] , \wAIn19[24] , \wAIn19[23] , \wAIn19[22] , 
        \wAIn19[21] , \wAIn19[20] , \wAIn19[19] , \wAIn19[18] , \wAIn19[17] , 
        \wAIn19[16] , \wAIn19[15] , \wAIn19[14] , \wAIn19[13] , \wAIn19[12] , 
        \wAIn19[11] , \wAIn19[10] , \wAIn19[9] , \wAIn19[8] , \wAIn19[7] , 
        \wAIn19[6] , \wAIn19[5] , \wAIn19[4] , \wAIn19[3] , \wAIn19[2] , 
        \wAIn19[1] , \wAIn19[0] }), .BIn({\wBIn19[31] , \wBIn19[30] , 
        \wBIn19[29] , \wBIn19[28] , \wBIn19[27] , \wBIn19[26] , \wBIn19[25] , 
        \wBIn19[24] , \wBIn19[23] , \wBIn19[22] , \wBIn19[21] , \wBIn19[20] , 
        \wBIn19[19] , \wBIn19[18] , \wBIn19[17] , \wBIn19[16] , \wBIn19[15] , 
        \wBIn19[14] , \wBIn19[13] , \wBIn19[12] , \wBIn19[11] , \wBIn19[10] , 
        \wBIn19[9] , \wBIn19[8] , \wBIn19[7] , \wBIn19[6] , \wBIn19[5] , 
        \wBIn19[4] , \wBIn19[3] , \wBIn19[2] , \wBIn19[1] , \wBIn19[0] }), 
        .HiOut({\wBMid18[31] , \wBMid18[30] , \wBMid18[29] , \wBMid18[28] , 
        \wBMid18[27] , \wBMid18[26] , \wBMid18[25] , \wBMid18[24] , 
        \wBMid18[23] , \wBMid18[22] , \wBMid18[21] , \wBMid18[20] , 
        \wBMid18[19] , \wBMid18[18] , \wBMid18[17] , \wBMid18[16] , 
        \wBMid18[15] , \wBMid18[14] , \wBMid18[13] , \wBMid18[12] , 
        \wBMid18[11] , \wBMid18[10] , \wBMid18[9] , \wBMid18[8] , \wBMid18[7] , 
        \wBMid18[6] , \wBMid18[5] , \wBMid18[4] , \wBMid18[3] , \wBMid18[2] , 
        \wBMid18[1] , \wBMid18[0] }), .LoOut({\wAMid19[31] , \wAMid19[30] , 
        \wAMid19[29] , \wAMid19[28] , \wAMid19[27] , \wAMid19[26] , 
        \wAMid19[25] , \wAMid19[24] , \wAMid19[23] , \wAMid19[22] , 
        \wAMid19[21] , \wAMid19[20] , \wAMid19[19] , \wAMid19[18] , 
        \wAMid19[17] , \wAMid19[16] , \wAMid19[15] , \wAMid19[14] , 
        \wAMid19[13] , \wAMid19[12] , \wAMid19[11] , \wAMid19[10] , 
        \wAMid19[9] , \wAMid19[8] , \wAMid19[7] , \wAMid19[6] , \wAMid19[5] , 
        \wAMid19[4] , \wAMid19[3] , \wAMid19[2] , \wAMid19[1] , \wAMid19[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn80[31] , \wAIn80[30] , \wAIn80[29] , \wAIn80[28] , \wAIn80[27] , 
        \wAIn80[26] , \wAIn80[25] , \wAIn80[24] , \wAIn80[23] , \wAIn80[22] , 
        \wAIn80[21] , \wAIn80[20] , \wAIn80[19] , \wAIn80[18] , \wAIn80[17] , 
        \wAIn80[16] , \wAIn80[15] , \wAIn80[14] , \wAIn80[13] , \wAIn80[12] , 
        \wAIn80[11] , \wAIn80[10] , \wAIn80[9] , \wAIn80[8] , \wAIn80[7] , 
        \wAIn80[6] , \wAIn80[5] , \wAIn80[4] , \wAIn80[3] , \wAIn80[2] , 
        \wAIn80[1] , \wAIn80[0] }), .BIn({\wBIn80[31] , \wBIn80[30] , 
        \wBIn80[29] , \wBIn80[28] , \wBIn80[27] , \wBIn80[26] , \wBIn80[25] , 
        \wBIn80[24] , \wBIn80[23] , \wBIn80[22] , \wBIn80[21] , \wBIn80[20] , 
        \wBIn80[19] , \wBIn80[18] , \wBIn80[17] , \wBIn80[16] , \wBIn80[15] , 
        \wBIn80[14] , \wBIn80[13] , \wBIn80[12] , \wBIn80[11] , \wBIn80[10] , 
        \wBIn80[9] , \wBIn80[8] , \wBIn80[7] , \wBIn80[6] , \wBIn80[5] , 
        \wBIn80[4] , \wBIn80[3] , \wBIn80[2] , \wBIn80[1] , \wBIn80[0] }), 
        .HiOut({\wBMid79[31] , \wBMid79[30] , \wBMid79[29] , \wBMid79[28] , 
        \wBMid79[27] , \wBMid79[26] , \wBMid79[25] , \wBMid79[24] , 
        \wBMid79[23] , \wBMid79[22] , \wBMid79[21] , \wBMid79[20] , 
        \wBMid79[19] , \wBMid79[18] , \wBMid79[17] , \wBMid79[16] , 
        \wBMid79[15] , \wBMid79[14] , \wBMid79[13] , \wBMid79[12] , 
        \wBMid79[11] , \wBMid79[10] , \wBMid79[9] , \wBMid79[8] , \wBMid79[7] , 
        \wBMid79[6] , \wBMid79[5] , \wBMid79[4] , \wBMid79[3] , \wBMid79[2] , 
        \wBMid79[1] , \wBMid79[0] }), .LoOut({\wAMid80[31] , \wAMid80[30] , 
        \wAMid80[29] , \wAMid80[28] , \wAMid80[27] , \wAMid80[26] , 
        \wAMid80[25] , \wAMid80[24] , \wAMid80[23] , \wAMid80[22] , 
        \wAMid80[21] , \wAMid80[20] , \wAMid80[19] , \wAMid80[18] , 
        \wAMid80[17] , \wAMid80[16] , \wAMid80[15] , \wAMid80[14] , 
        \wAMid80[13] , \wAMid80[12] , \wAMid80[11] , \wAMid80[10] , 
        \wAMid80[9] , \wAMid80[8] , \wAMid80[7] , \wAMid80[6] , \wAMid80[5] , 
        \wAMid80[4] , \wAMid80[3] , \wAMid80[2] , \wAMid80[1] , \wAMid80[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_185 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink186[31] , \ScanLink186[30] , \ScanLink186[29] , 
        \ScanLink186[28] , \ScanLink186[27] , \ScanLink186[26] , 
        \ScanLink186[25] , \ScanLink186[24] , \ScanLink186[23] , 
        \ScanLink186[22] , \ScanLink186[21] , \ScanLink186[20] , 
        \ScanLink186[19] , \ScanLink186[18] , \ScanLink186[17] , 
        \ScanLink186[16] , \ScanLink186[15] , \ScanLink186[14] , 
        \ScanLink186[13] , \ScanLink186[12] , \ScanLink186[11] , 
        \ScanLink186[10] , \ScanLink186[9] , \ScanLink186[8] , 
        \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , \ScanLink186[4] , 
        \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , \ScanLink186[0] 
        }), .ScanOut({\ScanLink185[31] , \ScanLink185[30] , \ScanLink185[29] , 
        \ScanLink185[28] , \ScanLink185[27] , \ScanLink185[26] , 
        \ScanLink185[25] , \ScanLink185[24] , \ScanLink185[23] , 
        \ScanLink185[22] , \ScanLink185[21] , \ScanLink185[20] , 
        \ScanLink185[19] , \ScanLink185[18] , \ScanLink185[17] , 
        \ScanLink185[16] , \ScanLink185[15] , \ScanLink185[14] , 
        \ScanLink185[13] , \ScanLink185[12] , \ScanLink185[11] , 
        \ScanLink185[10] , \ScanLink185[9] , \ScanLink185[8] , 
        \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , \ScanLink185[4] , 
        \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , \ScanLink185[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA35[31] , \wRegInA35[30] , \wRegInA35[29] , 
        \wRegInA35[28] , \wRegInA35[27] , \wRegInA35[26] , \wRegInA35[25] , 
        \wRegInA35[24] , \wRegInA35[23] , \wRegInA35[22] , \wRegInA35[21] , 
        \wRegInA35[20] , \wRegInA35[19] , \wRegInA35[18] , \wRegInA35[17] , 
        \wRegInA35[16] , \wRegInA35[15] , \wRegInA35[14] , \wRegInA35[13] , 
        \wRegInA35[12] , \wRegInA35[11] , \wRegInA35[10] , \wRegInA35[9] , 
        \wRegInA35[8] , \wRegInA35[7] , \wRegInA35[6] , \wRegInA35[5] , 
        \wRegInA35[4] , \wRegInA35[3] , \wRegInA35[2] , \wRegInA35[1] , 
        \wRegInA35[0] }), .Out({\wAIn35[31] , \wAIn35[30] , \wAIn35[29] , 
        \wAIn35[28] , \wAIn35[27] , \wAIn35[26] , \wAIn35[25] , \wAIn35[24] , 
        \wAIn35[23] , \wAIn35[22] , \wAIn35[21] , \wAIn35[20] , \wAIn35[19] , 
        \wAIn35[18] , \wAIn35[17] , \wAIn35[16] , \wAIn35[15] , \wAIn35[14] , 
        \wAIn35[13] , \wAIn35[12] , \wAIn35[11] , \wAIn35[10] , \wAIn35[9] , 
        \wAIn35[8] , \wAIn35[7] , \wAIn35[6] , \wAIn35[5] , \wAIn35[4] , 
        \wAIn35[3] , \wAIn35[2] , \wAIn35[1] , \wAIn35[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_219 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink220[31] , \ScanLink220[30] , \ScanLink220[29] , 
        \ScanLink220[28] , \ScanLink220[27] , \ScanLink220[26] , 
        \ScanLink220[25] , \ScanLink220[24] , \ScanLink220[23] , 
        \ScanLink220[22] , \ScanLink220[21] , \ScanLink220[20] , 
        \ScanLink220[19] , \ScanLink220[18] , \ScanLink220[17] , 
        \ScanLink220[16] , \ScanLink220[15] , \ScanLink220[14] , 
        \ScanLink220[13] , \ScanLink220[12] , \ScanLink220[11] , 
        \ScanLink220[10] , \ScanLink220[9] , \ScanLink220[8] , 
        \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , \ScanLink220[4] , 
        \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , \ScanLink220[0] 
        }), .ScanOut({\ScanLink219[31] , \ScanLink219[30] , \ScanLink219[29] , 
        \ScanLink219[28] , \ScanLink219[27] , \ScanLink219[26] , 
        \ScanLink219[25] , \ScanLink219[24] , \ScanLink219[23] , 
        \ScanLink219[22] , \ScanLink219[21] , \ScanLink219[20] , 
        \ScanLink219[19] , \ScanLink219[18] , \ScanLink219[17] , 
        \ScanLink219[16] , \ScanLink219[15] , \ScanLink219[14] , 
        \ScanLink219[13] , \ScanLink219[12] , \ScanLink219[11] , 
        \ScanLink219[10] , \ScanLink219[9] , \ScanLink219[8] , 
        \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , \ScanLink219[4] , 
        \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , \ScanLink219[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA18[31] , \wRegInA18[30] , \wRegInA18[29] , 
        \wRegInA18[28] , \wRegInA18[27] , \wRegInA18[26] , \wRegInA18[25] , 
        \wRegInA18[24] , \wRegInA18[23] , \wRegInA18[22] , \wRegInA18[21] , 
        \wRegInA18[20] , \wRegInA18[19] , \wRegInA18[18] , \wRegInA18[17] , 
        \wRegInA18[16] , \wRegInA18[15] , \wRegInA18[14] , \wRegInA18[13] , 
        \wRegInA18[12] , \wRegInA18[11] , \wRegInA18[10] , \wRegInA18[9] , 
        \wRegInA18[8] , \wRegInA18[7] , \wRegInA18[6] , \wRegInA18[5] , 
        \wRegInA18[4] , \wRegInA18[3] , \wRegInA18[2] , \wRegInA18[1] , 
        \wRegInA18[0] }), .Out({\wAIn18[31] , \wAIn18[30] , \wAIn18[29] , 
        \wAIn18[28] , \wAIn18[27] , \wAIn18[26] , \wAIn18[25] , \wAIn18[24] , 
        \wAIn18[23] , \wAIn18[22] , \wAIn18[21] , \wAIn18[20] , \wAIn18[19] , 
        \wAIn18[18] , \wAIn18[17] , \wAIn18[16] , \wAIn18[15] , \wAIn18[14] , 
        \wAIn18[13] , \wAIn18[12] , \wAIn18[11] , \wAIn18[10] , \wAIn18[9] , 
        \wAIn18[8] , \wAIn18[7] , \wAIn18[6] , \wAIn18[5] , \wAIn18[4] , 
        \wAIn18[3] , \wAIn18[2] , \wAIn18[1] , \wAIn18[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_129 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink130[31] , \ScanLink130[30] , \ScanLink130[29] , 
        \ScanLink130[28] , \ScanLink130[27] , \ScanLink130[26] , 
        \ScanLink130[25] , \ScanLink130[24] , \ScanLink130[23] , 
        \ScanLink130[22] , \ScanLink130[21] , \ScanLink130[20] , 
        \ScanLink130[19] , \ScanLink130[18] , \ScanLink130[17] , 
        \ScanLink130[16] , \ScanLink130[15] , \ScanLink130[14] , 
        \ScanLink130[13] , \ScanLink130[12] , \ScanLink130[11] , 
        \ScanLink130[10] , \ScanLink130[9] , \ScanLink130[8] , 
        \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , \ScanLink130[4] , 
        \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , \ScanLink130[0] 
        }), .ScanOut({\ScanLink129[31] , \ScanLink129[30] , \ScanLink129[29] , 
        \ScanLink129[28] , \ScanLink129[27] , \ScanLink129[26] , 
        \ScanLink129[25] , \ScanLink129[24] , \ScanLink129[23] , 
        \ScanLink129[22] , \ScanLink129[21] , \ScanLink129[20] , 
        \ScanLink129[19] , \ScanLink129[18] , \ScanLink129[17] , 
        \ScanLink129[16] , \ScanLink129[15] , \ScanLink129[14] , 
        \ScanLink129[13] , \ScanLink129[12] , \ScanLink129[11] , 
        \ScanLink129[10] , \ScanLink129[9] , \ScanLink129[8] , 
        \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , \ScanLink129[4] , 
        \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , \ScanLink129[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA63[31] , \wRegInA63[30] , \wRegInA63[29] , 
        \wRegInA63[28] , \wRegInA63[27] , \wRegInA63[26] , \wRegInA63[25] , 
        \wRegInA63[24] , \wRegInA63[23] , \wRegInA63[22] , \wRegInA63[21] , 
        \wRegInA63[20] , \wRegInA63[19] , \wRegInA63[18] , \wRegInA63[17] , 
        \wRegInA63[16] , \wRegInA63[15] , \wRegInA63[14] , \wRegInA63[13] , 
        \wRegInA63[12] , \wRegInA63[11] , \wRegInA63[10] , \wRegInA63[9] , 
        \wRegInA63[8] , \wRegInA63[7] , \wRegInA63[6] , \wRegInA63[5] , 
        \wRegInA63[4] , \wRegInA63[3] , \wRegInA63[2] , \wRegInA63[1] , 
        \wRegInA63[0] }), .Out({\wAIn63[31] , \wAIn63[30] , \wAIn63[29] , 
        \wAIn63[28] , \wAIn63[27] , \wAIn63[26] , \wAIn63[25] , \wAIn63[24] , 
        \wAIn63[23] , \wAIn63[22] , \wAIn63[21] , \wAIn63[20] , \wAIn63[19] , 
        \wAIn63[18] , \wAIn63[17] , \wAIn63[16] , \wAIn63[15] , \wAIn63[14] , 
        \wAIn63[13] , \wAIn63[12] , \wAIn63[11] , \wAIn63[10] , \wAIn63[9] , 
        \wAIn63[8] , \wAIn63[7] , \wAIn63[6] , \wAIn63[5] , \wAIn63[4] , 
        \wAIn63[3] , \wAIn63[2] , \wAIn63[1] , \wAIn63[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_79 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink80[31] , \ScanLink80[30] , \ScanLink80[29] , 
        \ScanLink80[28] , \ScanLink80[27] , \ScanLink80[26] , \ScanLink80[25] , 
        \ScanLink80[24] , \ScanLink80[23] , \ScanLink80[22] , \ScanLink80[21] , 
        \ScanLink80[20] , \ScanLink80[19] , \ScanLink80[18] , \ScanLink80[17] , 
        \ScanLink80[16] , \ScanLink80[15] , \ScanLink80[14] , \ScanLink80[13] , 
        \ScanLink80[12] , \ScanLink80[11] , \ScanLink80[10] , \ScanLink80[9] , 
        \ScanLink80[8] , \ScanLink80[7] , \ScanLink80[6] , \ScanLink80[5] , 
        \ScanLink80[4] , \ScanLink80[3] , \ScanLink80[2] , \ScanLink80[1] , 
        \ScanLink80[0] }), .ScanOut({\ScanLink79[31] , \ScanLink79[30] , 
        \ScanLink79[29] , \ScanLink79[28] , \ScanLink79[27] , \ScanLink79[26] , 
        \ScanLink79[25] , \ScanLink79[24] , \ScanLink79[23] , \ScanLink79[22] , 
        \ScanLink79[21] , \ScanLink79[20] , \ScanLink79[19] , \ScanLink79[18] , 
        \ScanLink79[17] , \ScanLink79[16] , \ScanLink79[15] , \ScanLink79[14] , 
        \ScanLink79[13] , \ScanLink79[12] , \ScanLink79[11] , \ScanLink79[10] , 
        \ScanLink79[9] , \ScanLink79[8] , \ScanLink79[7] , \ScanLink79[6] , 
        \ScanLink79[5] , \ScanLink79[4] , \ScanLink79[3] , \ScanLink79[2] , 
        \ScanLink79[1] , \ScanLink79[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA88[31] , \wRegInA88[30] , 
        \wRegInA88[29] , \wRegInA88[28] , \wRegInA88[27] , \wRegInA88[26] , 
        \wRegInA88[25] , \wRegInA88[24] , \wRegInA88[23] , \wRegInA88[22] , 
        \wRegInA88[21] , \wRegInA88[20] , \wRegInA88[19] , \wRegInA88[18] , 
        \wRegInA88[17] , \wRegInA88[16] , \wRegInA88[15] , \wRegInA88[14] , 
        \wRegInA88[13] , \wRegInA88[12] , \wRegInA88[11] , \wRegInA88[10] , 
        \wRegInA88[9] , \wRegInA88[8] , \wRegInA88[7] , \wRegInA88[6] , 
        \wRegInA88[5] , \wRegInA88[4] , \wRegInA88[3] , \wRegInA88[2] , 
        \wRegInA88[1] , \wRegInA88[0] }), .Out({\wAIn88[31] , \wAIn88[30] , 
        \wAIn88[29] , \wAIn88[28] , \wAIn88[27] , \wAIn88[26] , \wAIn88[25] , 
        \wAIn88[24] , \wAIn88[23] , \wAIn88[22] , \wAIn88[21] , \wAIn88[20] , 
        \wAIn88[19] , \wAIn88[18] , \wAIn88[17] , \wAIn88[16] , \wAIn88[15] , 
        \wAIn88[14] , \wAIn88[13] , \wAIn88[12] , \wAIn88[11] , \wAIn88[10] , 
        \wAIn88[9] , \wAIn88[8] , \wAIn88[7] , \wAIn88[6] , \wAIn88[5] , 
        \wAIn88[4] , \wAIn88[3] , \wAIn88[2] , \wAIn88[1] , \wAIn88[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn25[31] , \wAIn25[30] , \wAIn25[29] , \wAIn25[28] , \wAIn25[27] , 
        \wAIn25[26] , \wAIn25[25] , \wAIn25[24] , \wAIn25[23] , \wAIn25[22] , 
        \wAIn25[21] , \wAIn25[20] , \wAIn25[19] , \wAIn25[18] , \wAIn25[17] , 
        \wAIn25[16] , \wAIn25[15] , \wAIn25[14] , \wAIn25[13] , \wAIn25[12] , 
        \wAIn25[11] , \wAIn25[10] , \wAIn25[9] , \wAIn25[8] , \wAIn25[7] , 
        \wAIn25[6] , \wAIn25[5] , \wAIn25[4] , \wAIn25[3] , \wAIn25[2] , 
        \wAIn25[1] , \wAIn25[0] }), .BIn({\wBIn25[31] , \wBIn25[30] , 
        \wBIn25[29] , \wBIn25[28] , \wBIn25[27] , \wBIn25[26] , \wBIn25[25] , 
        \wBIn25[24] , \wBIn25[23] , \wBIn25[22] , \wBIn25[21] , \wBIn25[20] , 
        \wBIn25[19] , \wBIn25[18] , \wBIn25[17] , \wBIn25[16] , \wBIn25[15] , 
        \wBIn25[14] , \wBIn25[13] , \wBIn25[12] , \wBIn25[11] , \wBIn25[10] , 
        \wBIn25[9] , \wBIn25[8] , \wBIn25[7] , \wBIn25[6] , \wBIn25[5] , 
        \wBIn25[4] , \wBIn25[3] , \wBIn25[2] , \wBIn25[1] , \wBIn25[0] }), 
        .HiOut({\wBMid24[31] , \wBMid24[30] , \wBMid24[29] , \wBMid24[28] , 
        \wBMid24[27] , \wBMid24[26] , \wBMid24[25] , \wBMid24[24] , 
        \wBMid24[23] , \wBMid24[22] , \wBMid24[21] , \wBMid24[20] , 
        \wBMid24[19] , \wBMid24[18] , \wBMid24[17] , \wBMid24[16] , 
        \wBMid24[15] , \wBMid24[14] , \wBMid24[13] , \wBMid24[12] , 
        \wBMid24[11] , \wBMid24[10] , \wBMid24[9] , \wBMid24[8] , \wBMid24[7] , 
        \wBMid24[6] , \wBMid24[5] , \wBMid24[4] , \wBMid24[3] , \wBMid24[2] , 
        \wBMid24[1] , \wBMid24[0] }), .LoOut({\wAMid25[31] , \wAMid25[30] , 
        \wAMid25[29] , \wAMid25[28] , \wAMid25[27] , \wAMid25[26] , 
        \wAMid25[25] , \wAMid25[24] , \wAMid25[23] , \wAMid25[22] , 
        \wAMid25[21] , \wAMid25[20] , \wAMid25[19] , \wAMid25[18] , 
        \wAMid25[17] , \wAMid25[16] , \wAMid25[15] , \wAMid25[14] , 
        \wAMid25[13] , \wAMid25[12] , \wAMid25[11] , \wAMid25[10] , 
        \wAMid25[9] , \wAMid25[8] , \wAMid25[7] , \wAMid25[6] , \wAMid25[5] , 
        \wAMid25[4] , \wAMid25[3] , \wAMid25[2] , \wAMid25[1] , \wAMid25[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn50[31] , \wAIn50[30] , \wAIn50[29] , \wAIn50[28] , \wAIn50[27] , 
        \wAIn50[26] , \wAIn50[25] , \wAIn50[24] , \wAIn50[23] , \wAIn50[22] , 
        \wAIn50[21] , \wAIn50[20] , \wAIn50[19] , \wAIn50[18] , \wAIn50[17] , 
        \wAIn50[16] , \wAIn50[15] , \wAIn50[14] , \wAIn50[13] , \wAIn50[12] , 
        \wAIn50[11] , \wAIn50[10] , \wAIn50[9] , \wAIn50[8] , \wAIn50[7] , 
        \wAIn50[6] , \wAIn50[5] , \wAIn50[4] , \wAIn50[3] , \wAIn50[2] , 
        \wAIn50[1] , \wAIn50[0] }), .BIn({\wBIn50[31] , \wBIn50[30] , 
        \wBIn50[29] , \wBIn50[28] , \wBIn50[27] , \wBIn50[26] , \wBIn50[25] , 
        \wBIn50[24] , \wBIn50[23] , \wBIn50[22] , \wBIn50[21] , \wBIn50[20] , 
        \wBIn50[19] , \wBIn50[18] , \wBIn50[17] , \wBIn50[16] , \wBIn50[15] , 
        \wBIn50[14] , \wBIn50[13] , \wBIn50[12] , \wBIn50[11] , \wBIn50[10] , 
        \wBIn50[9] , \wBIn50[8] , \wBIn50[7] , \wBIn50[6] , \wBIn50[5] , 
        \wBIn50[4] , \wBIn50[3] , \wBIn50[2] , \wBIn50[1] , \wBIn50[0] }), 
        .HiOut({\wBMid49[31] , \wBMid49[30] , \wBMid49[29] , \wBMid49[28] , 
        \wBMid49[27] , \wBMid49[26] , \wBMid49[25] , \wBMid49[24] , 
        \wBMid49[23] , \wBMid49[22] , \wBMid49[21] , \wBMid49[20] , 
        \wBMid49[19] , \wBMid49[18] , \wBMid49[17] , \wBMid49[16] , 
        \wBMid49[15] , \wBMid49[14] , \wBMid49[13] , \wBMid49[12] , 
        \wBMid49[11] , \wBMid49[10] , \wBMid49[9] , \wBMid49[8] , \wBMid49[7] , 
        \wBMid49[6] , \wBMid49[5] , \wBMid49[4] , \wBMid49[3] , \wBMid49[2] , 
        \wBMid49[1] , \wBMid49[0] }), .LoOut({\wAMid50[31] , \wAMid50[30] , 
        \wAMid50[29] , \wAMid50[28] , \wAMid50[27] , \wAMid50[26] , 
        \wAMid50[25] , \wAMid50[24] , \wAMid50[23] , \wAMid50[22] , 
        \wAMid50[21] , \wAMid50[20] , \wAMid50[19] , \wAMid50[18] , 
        \wAMid50[17] , \wAMid50[16] , \wAMid50[15] , \wAMid50[14] , 
        \wAMid50[13] , \wAMid50[12] , \wAMid50[11] , \wAMid50[10] , 
        \wAMid50[9] , \wAMid50[8] , \wAMid50[7] , \wAMid50[6] , \wAMid50[5] , 
        \wAMid50[4] , \wAMid50[3] , \wAMid50[2] , \wAMid50[1] , \wAMid50[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn77[31] , \wAIn77[30] , \wAIn77[29] , \wAIn77[28] , \wAIn77[27] , 
        \wAIn77[26] , \wAIn77[25] , \wAIn77[24] , \wAIn77[23] , \wAIn77[22] , 
        \wAIn77[21] , \wAIn77[20] , \wAIn77[19] , \wAIn77[18] , \wAIn77[17] , 
        \wAIn77[16] , \wAIn77[15] , \wAIn77[14] , \wAIn77[13] , \wAIn77[12] , 
        \wAIn77[11] , \wAIn77[10] , \wAIn77[9] , \wAIn77[8] , \wAIn77[7] , 
        \wAIn77[6] , \wAIn77[5] , \wAIn77[4] , \wAIn77[3] , \wAIn77[2] , 
        \wAIn77[1] , \wAIn77[0] }), .BIn({\wBIn77[31] , \wBIn77[30] , 
        \wBIn77[29] , \wBIn77[28] , \wBIn77[27] , \wBIn77[26] , \wBIn77[25] , 
        \wBIn77[24] , \wBIn77[23] , \wBIn77[22] , \wBIn77[21] , \wBIn77[20] , 
        \wBIn77[19] , \wBIn77[18] , \wBIn77[17] , \wBIn77[16] , \wBIn77[15] , 
        \wBIn77[14] , \wBIn77[13] , \wBIn77[12] , \wBIn77[11] , \wBIn77[10] , 
        \wBIn77[9] , \wBIn77[8] , \wBIn77[7] , \wBIn77[6] , \wBIn77[5] , 
        \wBIn77[4] , \wBIn77[3] , \wBIn77[2] , \wBIn77[1] , \wBIn77[0] }), 
        .HiOut({\wBMid76[31] , \wBMid76[30] , \wBMid76[29] , \wBMid76[28] , 
        \wBMid76[27] , \wBMid76[26] , \wBMid76[25] , \wBMid76[24] , 
        \wBMid76[23] , \wBMid76[22] , \wBMid76[21] , \wBMid76[20] , 
        \wBMid76[19] , \wBMid76[18] , \wBMid76[17] , \wBMid76[16] , 
        \wBMid76[15] , \wBMid76[14] , \wBMid76[13] , \wBMid76[12] , 
        \wBMid76[11] , \wBMid76[10] , \wBMid76[9] , \wBMid76[8] , \wBMid76[7] , 
        \wBMid76[6] , \wBMid76[5] , \wBMid76[4] , \wBMid76[3] , \wBMid76[2] , 
        \wBMid76[1] , \wBMid76[0] }), .LoOut({\wAMid77[31] , \wAMid77[30] , 
        \wAMid77[29] , \wAMid77[28] , \wAMid77[27] , \wAMid77[26] , 
        \wAMid77[25] , \wAMid77[24] , \wAMid77[23] , \wAMid77[22] , 
        \wAMid77[21] , \wAMid77[20] , \wAMid77[19] , \wAMid77[18] , 
        \wAMid77[17] , \wAMid77[16] , \wAMid77[15] , \wAMid77[14] , 
        \wAMid77[13] , \wAMid77[12] , \wAMid77[11] , \wAMid77[10] , 
        \wAMid77[9] , \wAMid77[8] , \wAMid77[7] , \wAMid77[6] , \wAMid77[5] , 
        \wAMid77[4] , \wAMid77[3] , \wAMid77[2] , \wAMid77[1] , \wAMid77[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn92[31] , \wAIn92[30] , \wAIn92[29] , \wAIn92[28] , \wAIn92[27] , 
        \wAIn92[26] , \wAIn92[25] , \wAIn92[24] , \wAIn92[23] , \wAIn92[22] , 
        \wAIn92[21] , \wAIn92[20] , \wAIn92[19] , \wAIn92[18] , \wAIn92[17] , 
        \wAIn92[16] , \wAIn92[15] , \wAIn92[14] , \wAIn92[13] , \wAIn92[12] , 
        \wAIn92[11] , \wAIn92[10] , \wAIn92[9] , \wAIn92[8] , \wAIn92[7] , 
        \wAIn92[6] , \wAIn92[5] , \wAIn92[4] , \wAIn92[3] , \wAIn92[2] , 
        \wAIn92[1] , \wAIn92[0] }), .BIn({\wBIn92[31] , \wBIn92[30] , 
        \wBIn92[29] , \wBIn92[28] , \wBIn92[27] , \wBIn92[26] , \wBIn92[25] , 
        \wBIn92[24] , \wBIn92[23] , \wBIn92[22] , \wBIn92[21] , \wBIn92[20] , 
        \wBIn92[19] , \wBIn92[18] , \wBIn92[17] , \wBIn92[16] , \wBIn92[15] , 
        \wBIn92[14] , \wBIn92[13] , \wBIn92[12] , \wBIn92[11] , \wBIn92[10] , 
        \wBIn92[9] , \wBIn92[8] , \wBIn92[7] , \wBIn92[6] , \wBIn92[5] , 
        \wBIn92[4] , \wBIn92[3] , \wBIn92[2] , \wBIn92[1] , \wBIn92[0] }), 
        .HiOut({\wBMid91[31] , \wBMid91[30] , \wBMid91[29] , \wBMid91[28] , 
        \wBMid91[27] , \wBMid91[26] , \wBMid91[25] , \wBMid91[24] , 
        \wBMid91[23] , \wBMid91[22] , \wBMid91[21] , \wBMid91[20] , 
        \wBMid91[19] , \wBMid91[18] , \wBMid91[17] , \wBMid91[16] , 
        \wBMid91[15] , \wBMid91[14] , \wBMid91[13] , \wBMid91[12] , 
        \wBMid91[11] , \wBMid91[10] , \wBMid91[9] , \wBMid91[8] , \wBMid91[7] , 
        \wBMid91[6] , \wBMid91[5] , \wBMid91[4] , \wBMid91[3] , \wBMid91[2] , 
        \wBMid91[1] , \wBMid91[0] }), .LoOut({\wAMid92[31] , \wAMid92[30] , 
        \wAMid92[29] , \wAMid92[28] , \wAMid92[27] , \wAMid92[26] , 
        \wAMid92[25] , \wAMid92[24] , \wAMid92[23] , \wAMid92[22] , 
        \wAMid92[21] , \wAMid92[20] , \wAMid92[19] , \wAMid92[18] , 
        \wAMid92[17] , \wAMid92[16] , \wAMid92[15] , \wAMid92[14] , 
        \wAMid92[13] , \wAMid92[12] , \wAMid92[11] , \wAMid92[10] , 
        \wAMid92[9] , \wAMid92[8] , \wAMid92[7] , \wAMid92[6] , \wAMid92[5] , 
        \wAMid92[4] , \wAMid92[3] , \wAMid92[2] , \wAMid92[1] , \wAMid92[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid3[31] , 
        \wAMid3[30] , \wAMid3[29] , \wAMid3[28] , \wAMid3[27] , \wAMid3[26] , 
        \wAMid3[25] , \wAMid3[24] , \wAMid3[23] , \wAMid3[22] , \wAMid3[21] , 
        \wAMid3[20] , \wAMid3[19] , \wAMid3[18] , \wAMid3[17] , \wAMid3[16] , 
        \wAMid3[15] , \wAMid3[14] , \wAMid3[13] , \wAMid3[12] , \wAMid3[11] , 
        \wAMid3[10] , \wAMid3[9] , \wAMid3[8] , \wAMid3[7] , \wAMid3[6] , 
        \wAMid3[5] , \wAMid3[4] , \wAMid3[3] , \wAMid3[2] , \wAMid3[1] , 
        \wAMid3[0] }), .BIn({\wBMid3[31] , \wBMid3[30] , \wBMid3[29] , 
        \wBMid3[28] , \wBMid3[27] , \wBMid3[26] , \wBMid3[25] , \wBMid3[24] , 
        \wBMid3[23] , \wBMid3[22] , \wBMid3[21] , \wBMid3[20] , \wBMid3[19] , 
        \wBMid3[18] , \wBMid3[17] , \wBMid3[16] , \wBMid3[15] , \wBMid3[14] , 
        \wBMid3[13] , \wBMid3[12] , \wBMid3[11] , \wBMid3[10] , \wBMid3[9] , 
        \wBMid3[8] , \wBMid3[7] , \wBMid3[6] , \wBMid3[5] , \wBMid3[4] , 
        \wBMid3[3] , \wBMid3[2] , \wBMid3[1] , \wBMid3[0] }), .HiOut({
        \wRegInB3[31] , \wRegInB3[30] , \wRegInB3[29] , \wRegInB3[28] , 
        \wRegInB3[27] , \wRegInB3[26] , \wRegInB3[25] , \wRegInB3[24] , 
        \wRegInB3[23] , \wRegInB3[22] , \wRegInB3[21] , \wRegInB3[20] , 
        \wRegInB3[19] , \wRegInB3[18] , \wRegInB3[17] , \wRegInB3[16] , 
        \wRegInB3[15] , \wRegInB3[14] , \wRegInB3[13] , \wRegInB3[12] , 
        \wRegInB3[11] , \wRegInB3[10] , \wRegInB3[9] , \wRegInB3[8] , 
        \wRegInB3[7] , \wRegInB3[6] , \wRegInB3[5] , \wRegInB3[4] , 
        \wRegInB3[3] , \wRegInB3[2] , \wRegInB3[1] , \wRegInB3[0] }), .LoOut({
        \wRegInA4[31] , \wRegInA4[30] , \wRegInA4[29] , \wRegInA4[28] , 
        \wRegInA4[27] , \wRegInA4[26] , \wRegInA4[25] , \wRegInA4[24] , 
        \wRegInA4[23] , \wRegInA4[22] , \wRegInA4[21] , \wRegInA4[20] , 
        \wRegInA4[19] , \wRegInA4[18] , \wRegInA4[17] , \wRegInA4[16] , 
        \wRegInA4[15] , \wRegInA4[14] , \wRegInA4[13] , \wRegInA4[12] , 
        \wRegInA4[11] , \wRegInA4[10] , \wRegInA4[9] , \wRegInA4[8] , 
        \wRegInA4[7] , \wRegInA4[6] , \wRegInA4[5] , \wRegInA4[4] , 
        \wRegInA4[3] , \wRegInA4[2] , \wRegInA4[1] , \wRegInA4[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid29[31] , \wAMid29[30] , \wAMid29[29] , \wAMid29[28] , 
        \wAMid29[27] , \wAMid29[26] , \wAMid29[25] , \wAMid29[24] , 
        \wAMid29[23] , \wAMid29[22] , \wAMid29[21] , \wAMid29[20] , 
        \wAMid29[19] , \wAMid29[18] , \wAMid29[17] , \wAMid29[16] , 
        \wAMid29[15] , \wAMid29[14] , \wAMid29[13] , \wAMid29[12] , 
        \wAMid29[11] , \wAMid29[10] , \wAMid29[9] , \wAMid29[8] , \wAMid29[7] , 
        \wAMid29[6] , \wAMid29[5] , \wAMid29[4] , \wAMid29[3] , \wAMid29[2] , 
        \wAMid29[1] , \wAMid29[0] }), .BIn({\wBMid29[31] , \wBMid29[30] , 
        \wBMid29[29] , \wBMid29[28] , \wBMid29[27] , \wBMid29[26] , 
        \wBMid29[25] , \wBMid29[24] , \wBMid29[23] , \wBMid29[22] , 
        \wBMid29[21] , \wBMid29[20] , \wBMid29[19] , \wBMid29[18] , 
        \wBMid29[17] , \wBMid29[16] , \wBMid29[15] , \wBMid29[14] , 
        \wBMid29[13] , \wBMid29[12] , \wBMid29[11] , \wBMid29[10] , 
        \wBMid29[9] , \wBMid29[8] , \wBMid29[7] , \wBMid29[6] , \wBMid29[5] , 
        \wBMid29[4] , \wBMid29[3] , \wBMid29[2] , \wBMid29[1] , \wBMid29[0] }), 
        .HiOut({\wRegInB29[31] , \wRegInB29[30] , \wRegInB29[29] , 
        \wRegInB29[28] , \wRegInB29[27] , \wRegInB29[26] , \wRegInB29[25] , 
        \wRegInB29[24] , \wRegInB29[23] , \wRegInB29[22] , \wRegInB29[21] , 
        \wRegInB29[20] , \wRegInB29[19] , \wRegInB29[18] , \wRegInB29[17] , 
        \wRegInB29[16] , \wRegInB29[15] , \wRegInB29[14] , \wRegInB29[13] , 
        \wRegInB29[12] , \wRegInB29[11] , \wRegInB29[10] , \wRegInB29[9] , 
        \wRegInB29[8] , \wRegInB29[7] , \wRegInB29[6] , \wRegInB29[5] , 
        \wRegInB29[4] , \wRegInB29[3] , \wRegInB29[2] , \wRegInB29[1] , 
        \wRegInB29[0] }), .LoOut({\wRegInA30[31] , \wRegInA30[30] , 
        \wRegInA30[29] , \wRegInA30[28] , \wRegInA30[27] , \wRegInA30[26] , 
        \wRegInA30[25] , \wRegInA30[24] , \wRegInA30[23] , \wRegInA30[22] , 
        \wRegInA30[21] , \wRegInA30[20] , \wRegInA30[19] , \wRegInA30[18] , 
        \wRegInA30[17] , \wRegInA30[16] , \wRegInA30[15] , \wRegInA30[14] , 
        \wRegInA30[13] , \wRegInA30[12] , \wRegInA30[11] , \wRegInA30[10] , 
        \wRegInA30[9] , \wRegInA30[8] , \wRegInA30[7] , \wRegInA30[6] , 
        \wRegInA30[5] , \wRegInA30[4] , \wRegInA30[3] , \wRegInA30[2] , 
        \wRegInA30[1] , \wRegInA30[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid85[31] , \wAMid85[30] , \wAMid85[29] , \wAMid85[28] , 
        \wAMid85[27] , \wAMid85[26] , \wAMid85[25] , \wAMid85[24] , 
        \wAMid85[23] , \wAMid85[22] , \wAMid85[21] , \wAMid85[20] , 
        \wAMid85[19] , \wAMid85[18] , \wAMid85[17] , \wAMid85[16] , 
        \wAMid85[15] , \wAMid85[14] , \wAMid85[13] , \wAMid85[12] , 
        \wAMid85[11] , \wAMid85[10] , \wAMid85[9] , \wAMid85[8] , \wAMid85[7] , 
        \wAMid85[6] , \wAMid85[5] , \wAMid85[4] , \wAMid85[3] , \wAMid85[2] , 
        \wAMid85[1] , \wAMid85[0] }), .BIn({\wBMid85[31] , \wBMid85[30] , 
        \wBMid85[29] , \wBMid85[28] , \wBMid85[27] , \wBMid85[26] , 
        \wBMid85[25] , \wBMid85[24] , \wBMid85[23] , \wBMid85[22] , 
        \wBMid85[21] , \wBMid85[20] , \wBMid85[19] , \wBMid85[18] , 
        \wBMid85[17] , \wBMid85[16] , \wBMid85[15] , \wBMid85[14] , 
        \wBMid85[13] , \wBMid85[12] , \wBMid85[11] , \wBMid85[10] , 
        \wBMid85[9] , \wBMid85[8] , \wBMid85[7] , \wBMid85[6] , \wBMid85[5] , 
        \wBMid85[4] , \wBMid85[3] , \wBMid85[2] , \wBMid85[1] , \wBMid85[0] }), 
        .HiOut({\wRegInB85[31] , \wRegInB85[30] , \wRegInB85[29] , 
        \wRegInB85[28] , \wRegInB85[27] , \wRegInB85[26] , \wRegInB85[25] , 
        \wRegInB85[24] , \wRegInB85[23] , \wRegInB85[22] , \wRegInB85[21] , 
        \wRegInB85[20] , \wRegInB85[19] , \wRegInB85[18] , \wRegInB85[17] , 
        \wRegInB85[16] , \wRegInB85[15] , \wRegInB85[14] , \wRegInB85[13] , 
        \wRegInB85[12] , \wRegInB85[11] , \wRegInB85[10] , \wRegInB85[9] , 
        \wRegInB85[8] , \wRegInB85[7] , \wRegInB85[6] , \wRegInB85[5] , 
        \wRegInB85[4] , \wRegInB85[3] , \wRegInB85[2] , \wRegInB85[1] , 
        \wRegInB85[0] }), .LoOut({\wRegInA86[31] , \wRegInA86[30] , 
        \wRegInA86[29] , \wRegInA86[28] , \wRegInA86[27] , \wRegInA86[26] , 
        \wRegInA86[25] , \wRegInA86[24] , \wRegInA86[23] , \wRegInA86[22] , 
        \wRegInA86[21] , \wRegInA86[20] , \wRegInA86[19] , \wRegInA86[18] , 
        \wRegInA86[17] , \wRegInA86[16] , \wRegInA86[15] , \wRegInA86[14] , 
        \wRegInA86[13] , \wRegInA86[12] , \wRegInA86[11] , \wRegInA86[10] , 
        \wRegInA86[9] , \wRegInA86[8] , \wRegInA86[7] , \wRegInA86[6] , 
        \wRegInA86[5] , \wRegInA86[4] , \wRegInA86[3] , \wRegInA86[2] , 
        \wRegInA86[1] , \wRegInA86[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_197 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink198[31] , \ScanLink198[30] , \ScanLink198[29] , 
        \ScanLink198[28] , \ScanLink198[27] , \ScanLink198[26] , 
        \ScanLink198[25] , \ScanLink198[24] , \ScanLink198[23] , 
        \ScanLink198[22] , \ScanLink198[21] , \ScanLink198[20] , 
        \ScanLink198[19] , \ScanLink198[18] , \ScanLink198[17] , 
        \ScanLink198[16] , \ScanLink198[15] , \ScanLink198[14] , 
        \ScanLink198[13] , \ScanLink198[12] , \ScanLink198[11] , 
        \ScanLink198[10] , \ScanLink198[9] , \ScanLink198[8] , 
        \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , \ScanLink198[4] , 
        \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , \ScanLink198[0] 
        }), .ScanOut({\ScanLink197[31] , \ScanLink197[30] , \ScanLink197[29] , 
        \ScanLink197[28] , \ScanLink197[27] , \ScanLink197[26] , 
        \ScanLink197[25] , \ScanLink197[24] , \ScanLink197[23] , 
        \ScanLink197[22] , \ScanLink197[21] , \ScanLink197[20] , 
        \ScanLink197[19] , \ScanLink197[18] , \ScanLink197[17] , 
        \ScanLink197[16] , \ScanLink197[15] , \ScanLink197[14] , 
        \ScanLink197[13] , \ScanLink197[12] , \ScanLink197[11] , 
        \ScanLink197[10] , \ScanLink197[9] , \ScanLink197[8] , 
        \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , \ScanLink197[4] , 
        \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , \ScanLink197[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA29[31] , \wRegInA29[30] , \wRegInA29[29] , 
        \wRegInA29[28] , \wRegInA29[27] , \wRegInA29[26] , \wRegInA29[25] , 
        \wRegInA29[24] , \wRegInA29[23] , \wRegInA29[22] , \wRegInA29[21] , 
        \wRegInA29[20] , \wRegInA29[19] , \wRegInA29[18] , \wRegInA29[17] , 
        \wRegInA29[16] , \wRegInA29[15] , \wRegInA29[14] , \wRegInA29[13] , 
        \wRegInA29[12] , \wRegInA29[11] , \wRegInA29[10] , \wRegInA29[9] , 
        \wRegInA29[8] , \wRegInA29[7] , \wRegInA29[6] , \wRegInA29[5] , 
        \wRegInA29[4] , \wRegInA29[3] , \wRegInA29[2] , \wRegInA29[1] , 
        \wRegInA29[0] }), .Out({\wAIn29[31] , \wAIn29[30] , \wAIn29[29] , 
        \wAIn29[28] , \wAIn29[27] , \wAIn29[26] , \wAIn29[25] , \wAIn29[24] , 
        \wAIn29[23] , \wAIn29[22] , \wAIn29[21] , \wAIn29[20] , \wAIn29[19] , 
        \wAIn29[18] , \wAIn29[17] , \wAIn29[16] , \wAIn29[15] , \wAIn29[14] , 
        \wAIn29[13] , \wAIn29[12] , \wAIn29[11] , \wAIn29[10] , \wAIn29[9] , 
        \wAIn29[8] , \wAIn29[7] , \wAIn29[6] , \wAIn29[5] , \wAIn29[4] , 
        \wAIn29[3] , \wAIn29[2] , \wAIn29[1] , \wAIn29[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn107[31] , \wAIn107[30] , \wAIn107[29] , \wAIn107[28] , 
        \wAIn107[27] , \wAIn107[26] , \wAIn107[25] , \wAIn107[24] , 
        \wAIn107[23] , \wAIn107[22] , \wAIn107[21] , \wAIn107[20] , 
        \wAIn107[19] , \wAIn107[18] , \wAIn107[17] , \wAIn107[16] , 
        \wAIn107[15] , \wAIn107[14] , \wAIn107[13] , \wAIn107[12] , 
        \wAIn107[11] , \wAIn107[10] , \wAIn107[9] , \wAIn107[8] , \wAIn107[7] , 
        \wAIn107[6] , \wAIn107[5] , \wAIn107[4] , \wAIn107[3] , \wAIn107[2] , 
        \wAIn107[1] , \wAIn107[0] }), .BIn({\wBIn107[31] , \wBIn107[30] , 
        \wBIn107[29] , \wBIn107[28] , \wBIn107[27] , \wBIn107[26] , 
        \wBIn107[25] , \wBIn107[24] , \wBIn107[23] , \wBIn107[22] , 
        \wBIn107[21] , \wBIn107[20] , \wBIn107[19] , \wBIn107[18] , 
        \wBIn107[17] , \wBIn107[16] , \wBIn107[15] , \wBIn107[14] , 
        \wBIn107[13] , \wBIn107[12] , \wBIn107[11] , \wBIn107[10] , 
        \wBIn107[9] , \wBIn107[8] , \wBIn107[7] , \wBIn107[6] , \wBIn107[5] , 
        \wBIn107[4] , \wBIn107[3] , \wBIn107[2] , \wBIn107[1] , \wBIn107[0] }), 
        .HiOut({\wBMid106[31] , \wBMid106[30] , \wBMid106[29] , \wBMid106[28] , 
        \wBMid106[27] , \wBMid106[26] , \wBMid106[25] , \wBMid106[24] , 
        \wBMid106[23] , \wBMid106[22] , \wBMid106[21] , \wBMid106[20] , 
        \wBMid106[19] , \wBMid106[18] , \wBMid106[17] , \wBMid106[16] , 
        \wBMid106[15] , \wBMid106[14] , \wBMid106[13] , \wBMid106[12] , 
        \wBMid106[11] , \wBMid106[10] , \wBMid106[9] , \wBMid106[8] , 
        \wBMid106[7] , \wBMid106[6] , \wBMid106[5] , \wBMid106[4] , 
        \wBMid106[3] , \wBMid106[2] , \wBMid106[1] , \wBMid106[0] }), .LoOut({
        \wAMid107[31] , \wAMid107[30] , \wAMid107[29] , \wAMid107[28] , 
        \wAMid107[27] , \wAMid107[26] , \wAMid107[25] , \wAMid107[24] , 
        \wAMid107[23] , \wAMid107[22] , \wAMid107[21] , \wAMid107[20] , 
        \wAMid107[19] , \wAMid107[18] , \wAMid107[17] , \wAMid107[16] , 
        \wAMid107[15] , \wAMid107[14] , \wAMid107[13] , \wAMid107[12] , 
        \wAMid107[11] , \wAMid107[10] , \wAMid107[9] , \wAMid107[8] , 
        \wAMid107[7] , \wAMid107[6] , \wAMid107[5] , \wAMid107[4] , 
        \wAMid107[3] , \wAMid107[2] , \wAMid107[1] , \wAMid107[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_242 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink243[31] , \ScanLink243[30] , \ScanLink243[29] , 
        \ScanLink243[28] , \ScanLink243[27] , \ScanLink243[26] , 
        \ScanLink243[25] , \ScanLink243[24] , \ScanLink243[23] , 
        \ScanLink243[22] , \ScanLink243[21] , \ScanLink243[20] , 
        \ScanLink243[19] , \ScanLink243[18] , \ScanLink243[17] , 
        \ScanLink243[16] , \ScanLink243[15] , \ScanLink243[14] , 
        \ScanLink243[13] , \ScanLink243[12] , \ScanLink243[11] , 
        \ScanLink243[10] , \ScanLink243[9] , \ScanLink243[8] , 
        \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , \ScanLink243[4] , 
        \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , \ScanLink243[0] 
        }), .ScanOut({\ScanLink242[31] , \ScanLink242[30] , \ScanLink242[29] , 
        \ScanLink242[28] , \ScanLink242[27] , \ScanLink242[26] , 
        \ScanLink242[25] , \ScanLink242[24] , \ScanLink242[23] , 
        \ScanLink242[22] , \ScanLink242[21] , \ScanLink242[20] , 
        \ScanLink242[19] , \ScanLink242[18] , \ScanLink242[17] , 
        \ScanLink242[16] , \ScanLink242[15] , \ScanLink242[14] , 
        \ScanLink242[13] , \ScanLink242[12] , \ScanLink242[11] , 
        \ScanLink242[10] , \ScanLink242[9] , \ScanLink242[8] , 
        \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , \ScanLink242[4] , 
        \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , \ScanLink242[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB6[31] , \wRegInB6[30] , \wRegInB6[29] , \wRegInB6[28] , 
        \wRegInB6[27] , \wRegInB6[26] , \wRegInB6[25] , \wRegInB6[24] , 
        \wRegInB6[23] , \wRegInB6[22] , \wRegInB6[21] , \wRegInB6[20] , 
        \wRegInB6[19] , \wRegInB6[18] , \wRegInB6[17] , \wRegInB6[16] , 
        \wRegInB6[15] , \wRegInB6[14] , \wRegInB6[13] , \wRegInB6[12] , 
        \wRegInB6[11] , \wRegInB6[10] , \wRegInB6[9] , \wRegInB6[8] , 
        \wRegInB6[7] , \wRegInB6[6] , \wRegInB6[5] , \wRegInB6[4] , 
        \wRegInB6[3] , \wRegInB6[2] , \wRegInB6[1] , \wRegInB6[0] }), .Out({
        \wBIn6[31] , \wBIn6[30] , \wBIn6[29] , \wBIn6[28] , \wBIn6[27] , 
        \wBIn6[26] , \wBIn6[25] , \wBIn6[24] , \wBIn6[23] , \wBIn6[22] , 
        \wBIn6[21] , \wBIn6[20] , \wBIn6[19] , \wBIn6[18] , \wBIn6[17] , 
        \wBIn6[16] , \wBIn6[15] , \wBIn6[14] , \wBIn6[13] , \wBIn6[12] , 
        \wBIn6[11] , \wBIn6[10] , \wBIn6[9] , \wBIn6[8] , \wBIn6[7] , 
        \wBIn6[6] , \wBIn6[5] , \wBIn6[4] , \wBIn6[3] , \wBIn6[2] , \wBIn6[1] , 
        \wBIn6[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid47[31] , \wAMid47[30] , \wAMid47[29] , \wAMid47[28] , 
        \wAMid47[27] , \wAMid47[26] , \wAMid47[25] , \wAMid47[24] , 
        \wAMid47[23] , \wAMid47[22] , \wAMid47[21] , \wAMid47[20] , 
        \wAMid47[19] , \wAMid47[18] , \wAMid47[17] , \wAMid47[16] , 
        \wAMid47[15] , \wAMid47[14] , \wAMid47[13] , \wAMid47[12] , 
        \wAMid47[11] , \wAMid47[10] , \wAMid47[9] , \wAMid47[8] , \wAMid47[7] , 
        \wAMid47[6] , \wAMid47[5] , \wAMid47[4] , \wAMid47[3] , \wAMid47[2] , 
        \wAMid47[1] , \wAMid47[0] }), .BIn({\wBMid47[31] , \wBMid47[30] , 
        \wBMid47[29] , \wBMid47[28] , \wBMid47[27] , \wBMid47[26] , 
        \wBMid47[25] , \wBMid47[24] , \wBMid47[23] , \wBMid47[22] , 
        \wBMid47[21] , \wBMid47[20] , \wBMid47[19] , \wBMid47[18] , 
        \wBMid47[17] , \wBMid47[16] , \wBMid47[15] , \wBMid47[14] , 
        \wBMid47[13] , \wBMid47[12] , \wBMid47[11] , \wBMid47[10] , 
        \wBMid47[9] , \wBMid47[8] , \wBMid47[7] , \wBMid47[6] , \wBMid47[5] , 
        \wBMid47[4] , \wBMid47[3] , \wBMid47[2] , \wBMid47[1] , \wBMid47[0] }), 
        .HiOut({\wRegInB47[31] , \wRegInB47[30] , \wRegInB47[29] , 
        \wRegInB47[28] , \wRegInB47[27] , \wRegInB47[26] , \wRegInB47[25] , 
        \wRegInB47[24] , \wRegInB47[23] , \wRegInB47[22] , \wRegInB47[21] , 
        \wRegInB47[20] , \wRegInB47[19] , \wRegInB47[18] , \wRegInB47[17] , 
        \wRegInB47[16] , \wRegInB47[15] , \wRegInB47[14] , \wRegInB47[13] , 
        \wRegInB47[12] , \wRegInB47[11] , \wRegInB47[10] , \wRegInB47[9] , 
        \wRegInB47[8] , \wRegInB47[7] , \wRegInB47[6] , \wRegInB47[5] , 
        \wRegInB47[4] , \wRegInB47[3] , \wRegInB47[2] , \wRegInB47[1] , 
        \wRegInB47[0] }), .LoOut({\wRegInA48[31] , \wRegInA48[30] , 
        \wRegInA48[29] , \wRegInA48[28] , \wRegInA48[27] , \wRegInA48[26] , 
        \wRegInA48[25] , \wRegInA48[24] , \wRegInA48[23] , \wRegInA48[22] , 
        \wRegInA48[21] , \wRegInA48[20] , \wRegInA48[19] , \wRegInA48[18] , 
        \wRegInA48[17] , \wRegInA48[16] , \wRegInA48[15] , \wRegInA48[14] , 
        \wRegInA48[13] , \wRegInA48[12] , \wRegInA48[11] , \wRegInA48[10] , 
        \wRegInA48[9] , \wRegInA48[8] , \wRegInA48[7] , \wRegInA48[6] , 
        \wRegInA48[5] , \wRegInA48[4] , \wRegInA48[3] , \wRegInA48[2] , 
        \wRegInA48[1] , \wRegInA48[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_172 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink173[31] , \ScanLink173[30] , \ScanLink173[29] , 
        \ScanLink173[28] , \ScanLink173[27] , \ScanLink173[26] , 
        \ScanLink173[25] , \ScanLink173[24] , \ScanLink173[23] , 
        \ScanLink173[22] , \ScanLink173[21] , \ScanLink173[20] , 
        \ScanLink173[19] , \ScanLink173[18] , \ScanLink173[17] , 
        \ScanLink173[16] , \ScanLink173[15] , \ScanLink173[14] , 
        \ScanLink173[13] , \ScanLink173[12] , \ScanLink173[11] , 
        \ScanLink173[10] , \ScanLink173[9] , \ScanLink173[8] , 
        \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , \ScanLink173[4] , 
        \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , \ScanLink173[0] 
        }), .ScanOut({\ScanLink172[31] , \ScanLink172[30] , \ScanLink172[29] , 
        \ScanLink172[28] , \ScanLink172[27] , \ScanLink172[26] , 
        \ScanLink172[25] , \ScanLink172[24] , \ScanLink172[23] , 
        \ScanLink172[22] , \ScanLink172[21] , \ScanLink172[20] , 
        \ScanLink172[19] , \ScanLink172[18] , \ScanLink172[17] , 
        \ScanLink172[16] , \ScanLink172[15] , \ScanLink172[14] , 
        \ScanLink172[13] , \ScanLink172[12] , \ScanLink172[11] , 
        \ScanLink172[10] , \ScanLink172[9] , \ScanLink172[8] , 
        \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , \ScanLink172[4] , 
        \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , \ScanLink172[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB41[31] , \wRegInB41[30] , \wRegInB41[29] , 
        \wRegInB41[28] , \wRegInB41[27] , \wRegInB41[26] , \wRegInB41[25] , 
        \wRegInB41[24] , \wRegInB41[23] , \wRegInB41[22] , \wRegInB41[21] , 
        \wRegInB41[20] , \wRegInB41[19] , \wRegInB41[18] , \wRegInB41[17] , 
        \wRegInB41[16] , \wRegInB41[15] , \wRegInB41[14] , \wRegInB41[13] , 
        \wRegInB41[12] , \wRegInB41[11] , \wRegInB41[10] , \wRegInB41[9] , 
        \wRegInB41[8] , \wRegInB41[7] , \wRegInB41[6] , \wRegInB41[5] , 
        \wRegInB41[4] , \wRegInB41[3] , \wRegInB41[2] , \wRegInB41[1] , 
        \wRegInB41[0] }), .Out({\wBIn41[31] , \wBIn41[30] , \wBIn41[29] , 
        \wBIn41[28] , \wBIn41[27] , \wBIn41[26] , \wBIn41[25] , \wBIn41[24] , 
        \wBIn41[23] , \wBIn41[22] , \wBIn41[21] , \wBIn41[20] , \wBIn41[19] , 
        \wBIn41[18] , \wBIn41[17] , \wBIn41[16] , \wBIn41[15] , \wBIn41[14] , 
        \wBIn41[13] , \wBIn41[12] , \wBIn41[11] , \wBIn41[10] , \wBIn41[9] , 
        \wBIn41[8] , \wBIn41[7] , \wBIn41[6] , \wBIn41[5] , \wBIn41[4] , 
        \wBIn41[3] , \wBIn41[2] , \wBIn41[1] , \wBIn41[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_22 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink23[31] , \ScanLink23[30] , \ScanLink23[29] , 
        \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , \ScanLink23[25] , 
        \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , \ScanLink23[21] , 
        \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , \ScanLink23[17] , 
        \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , \ScanLink23[13] , 
        \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , \ScanLink23[9] , 
        \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , \ScanLink23[5] , 
        \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , \ScanLink23[1] , 
        \ScanLink23[0] }), .ScanOut({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB116[31] , \wRegInB116[30] , 
        \wRegInB116[29] , \wRegInB116[28] , \wRegInB116[27] , \wRegInB116[26] , 
        \wRegInB116[25] , \wRegInB116[24] , \wRegInB116[23] , \wRegInB116[22] , 
        \wRegInB116[21] , \wRegInB116[20] , \wRegInB116[19] , \wRegInB116[18] , 
        \wRegInB116[17] , \wRegInB116[16] , \wRegInB116[15] , \wRegInB116[14] , 
        \wRegInB116[13] , \wRegInB116[12] , \wRegInB116[11] , \wRegInB116[10] , 
        \wRegInB116[9] , \wRegInB116[8] , \wRegInB116[7] , \wRegInB116[6] , 
        \wRegInB116[5] , \wRegInB116[4] , \wRegInB116[3] , \wRegInB116[2] , 
        \wRegInB116[1] , \wRegInB116[0] }), .Out({\wBIn116[31] , \wBIn116[30] , 
        \wBIn116[29] , \wBIn116[28] , \wBIn116[27] , \wBIn116[26] , 
        \wBIn116[25] , \wBIn116[24] , \wBIn116[23] , \wBIn116[22] , 
        \wBIn116[21] , \wBIn116[20] , \wBIn116[19] , \wBIn116[18] , 
        \wBIn116[17] , \wBIn116[16] , \wBIn116[15] , \wBIn116[14] , 
        \wBIn116[13] , \wBIn116[12] , \wBIn116[11] , \wBIn116[10] , 
        \wBIn116[9] , \wBIn116[8] , \wBIn116[7] , \wBIn116[6] , \wBIn116[5] , 
        \wBIn116[4] , \wBIn116[3] , \wBIn116[2] , \wBIn116[1] , \wBIn116[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn89[31] , \wAIn89[30] , \wAIn89[29] , \wAIn89[28] , \wAIn89[27] , 
        \wAIn89[26] , \wAIn89[25] , \wAIn89[24] , \wAIn89[23] , \wAIn89[22] , 
        \wAIn89[21] , \wAIn89[20] , \wAIn89[19] , \wAIn89[18] , \wAIn89[17] , 
        \wAIn89[16] , \wAIn89[15] , \wAIn89[14] , \wAIn89[13] , \wAIn89[12] , 
        \wAIn89[11] , \wAIn89[10] , \wAIn89[9] , \wAIn89[8] , \wAIn89[7] , 
        \wAIn89[6] , \wAIn89[5] , \wAIn89[4] , \wAIn89[3] , \wAIn89[2] , 
        \wAIn89[1] , \wAIn89[0] }), .BIn({\wBIn89[31] , \wBIn89[30] , 
        \wBIn89[29] , \wBIn89[28] , \wBIn89[27] , \wBIn89[26] , \wBIn89[25] , 
        \wBIn89[24] , \wBIn89[23] , \wBIn89[22] , \wBIn89[21] , \wBIn89[20] , 
        \wBIn89[19] , \wBIn89[18] , \wBIn89[17] , \wBIn89[16] , \wBIn89[15] , 
        \wBIn89[14] , \wBIn89[13] , \wBIn89[12] , \wBIn89[11] , \wBIn89[10] , 
        \wBIn89[9] , \wBIn89[8] , \wBIn89[7] , \wBIn89[6] , \wBIn89[5] , 
        \wBIn89[4] , \wBIn89[3] , \wBIn89[2] , \wBIn89[1] , \wBIn89[0] }), 
        .HiOut({\wBMid88[31] , \wBMid88[30] , \wBMid88[29] , \wBMid88[28] , 
        \wBMid88[27] , \wBMid88[26] , \wBMid88[25] , \wBMid88[24] , 
        \wBMid88[23] , \wBMid88[22] , \wBMid88[21] , \wBMid88[20] , 
        \wBMid88[19] , \wBMid88[18] , \wBMid88[17] , \wBMid88[16] , 
        \wBMid88[15] , \wBMid88[14] , \wBMid88[13] , \wBMid88[12] , 
        \wBMid88[11] , \wBMid88[10] , \wBMid88[9] , \wBMid88[8] , \wBMid88[7] , 
        \wBMid88[6] , \wBMid88[5] , \wBMid88[4] , \wBMid88[3] , \wBMid88[2] , 
        \wBMid88[1] , \wBMid88[0] }), .LoOut({\wAMid89[31] , \wAMid89[30] , 
        \wAMid89[29] , \wAMid89[28] , \wAMid89[27] , \wAMid89[26] , 
        \wAMid89[25] , \wAMid89[24] , \wAMid89[23] , \wAMid89[22] , 
        \wAMid89[21] , \wAMid89[20] , \wAMid89[19] , \wAMid89[18] , 
        \wAMid89[17] , \wAMid89[16] , \wAMid89[15] , \wAMid89[14] , 
        \wAMid89[13] , \wAMid89[12] , \wAMid89[11] , \wAMid89[10] , 
        \wAMid89[9] , \wAMid89[8] , \wAMid89[7] , \wAMid89[6] , \wAMid89[5] , 
        \wAMid89[4] , \wAMid89[3] , \wAMid89[2] , \wAMid89[1] , \wAMid89[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn120[31] , \wAIn120[30] , \wAIn120[29] , \wAIn120[28] , 
        \wAIn120[27] , \wAIn120[26] , \wAIn120[25] , \wAIn120[24] , 
        \wAIn120[23] , \wAIn120[22] , \wAIn120[21] , \wAIn120[20] , 
        \wAIn120[19] , \wAIn120[18] , \wAIn120[17] , \wAIn120[16] , 
        \wAIn120[15] , \wAIn120[14] , \wAIn120[13] , \wAIn120[12] , 
        \wAIn120[11] , \wAIn120[10] , \wAIn120[9] , \wAIn120[8] , \wAIn120[7] , 
        \wAIn120[6] , \wAIn120[5] , \wAIn120[4] , \wAIn120[3] , \wAIn120[2] , 
        \wAIn120[1] , \wAIn120[0] }), .BIn({\wBIn120[31] , \wBIn120[30] , 
        \wBIn120[29] , \wBIn120[28] , \wBIn120[27] , \wBIn120[26] , 
        \wBIn120[25] , \wBIn120[24] , \wBIn120[23] , \wBIn120[22] , 
        \wBIn120[21] , \wBIn120[20] , \wBIn120[19] , \wBIn120[18] , 
        \wBIn120[17] , \wBIn120[16] , \wBIn120[15] , \wBIn120[14] , 
        \wBIn120[13] , \wBIn120[12] , \wBIn120[11] , \wBIn120[10] , 
        \wBIn120[9] , \wBIn120[8] , \wBIn120[7] , \wBIn120[6] , \wBIn120[5] , 
        \wBIn120[4] , \wBIn120[3] , \wBIn120[2] , \wBIn120[1] , \wBIn120[0] }), 
        .HiOut({\wBMid119[31] , \wBMid119[30] , \wBMid119[29] , \wBMid119[28] , 
        \wBMid119[27] , \wBMid119[26] , \wBMid119[25] , \wBMid119[24] , 
        \wBMid119[23] , \wBMid119[22] , \wBMid119[21] , \wBMid119[20] , 
        \wBMid119[19] , \wBMid119[18] , \wBMid119[17] , \wBMid119[16] , 
        \wBMid119[15] , \wBMid119[14] , \wBMid119[13] , \wBMid119[12] , 
        \wBMid119[11] , \wBMid119[10] , \wBMid119[9] , \wBMid119[8] , 
        \wBMid119[7] , \wBMid119[6] , \wBMid119[5] , \wBMid119[4] , 
        \wBMid119[3] , \wBMid119[2] , \wBMid119[1] , \wBMid119[0] }), .LoOut({
        \wAMid120[31] , \wAMid120[30] , \wAMid120[29] , \wAMid120[28] , 
        \wAMid120[27] , \wAMid120[26] , \wAMid120[25] , \wAMid120[24] , 
        \wAMid120[23] , \wAMid120[22] , \wAMid120[21] , \wAMid120[20] , 
        \wAMid120[19] , \wAMid120[18] , \wAMid120[17] , \wAMid120[16] , 
        \wAMid120[15] , \wAMid120[14] , \wAMid120[13] , \wAMid120[12] , 
        \wAMid120[11] , \wAMid120[10] , \wAMid120[9] , \wAMid120[8] , 
        \wAMid120[7] , \wAMid120[6] , \wAMid120[5] , \wAMid120[4] , 
        \wAMid120[3] , \wAMid120[2] , \wAMid120[1] , \wAMid120[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid60[31] , \wAMid60[30] , \wAMid60[29] , \wAMid60[28] , 
        \wAMid60[27] , \wAMid60[26] , \wAMid60[25] , \wAMid60[24] , 
        \wAMid60[23] , \wAMid60[22] , \wAMid60[21] , \wAMid60[20] , 
        \wAMid60[19] , \wAMid60[18] , \wAMid60[17] , \wAMid60[16] , 
        \wAMid60[15] , \wAMid60[14] , \wAMid60[13] , \wAMid60[12] , 
        \wAMid60[11] , \wAMid60[10] , \wAMid60[9] , \wAMid60[8] , \wAMid60[7] , 
        \wAMid60[6] , \wAMid60[5] , \wAMid60[4] , \wAMid60[3] , \wAMid60[2] , 
        \wAMid60[1] , \wAMid60[0] }), .BIn({\wBMid60[31] , \wBMid60[30] , 
        \wBMid60[29] , \wBMid60[28] , \wBMid60[27] , \wBMid60[26] , 
        \wBMid60[25] , \wBMid60[24] , \wBMid60[23] , \wBMid60[22] , 
        \wBMid60[21] , \wBMid60[20] , \wBMid60[19] , \wBMid60[18] , 
        \wBMid60[17] , \wBMid60[16] , \wBMid60[15] , \wBMid60[14] , 
        \wBMid60[13] , \wBMid60[12] , \wBMid60[11] , \wBMid60[10] , 
        \wBMid60[9] , \wBMid60[8] , \wBMid60[7] , \wBMid60[6] , \wBMid60[5] , 
        \wBMid60[4] , \wBMid60[3] , \wBMid60[2] , \wBMid60[1] , \wBMid60[0] }), 
        .HiOut({\wRegInB60[31] , \wRegInB60[30] , \wRegInB60[29] , 
        \wRegInB60[28] , \wRegInB60[27] , \wRegInB60[26] , \wRegInB60[25] , 
        \wRegInB60[24] , \wRegInB60[23] , \wRegInB60[22] , \wRegInB60[21] , 
        \wRegInB60[20] , \wRegInB60[19] , \wRegInB60[18] , \wRegInB60[17] , 
        \wRegInB60[16] , \wRegInB60[15] , \wRegInB60[14] , \wRegInB60[13] , 
        \wRegInB60[12] , \wRegInB60[11] , \wRegInB60[10] , \wRegInB60[9] , 
        \wRegInB60[8] , \wRegInB60[7] , \wRegInB60[6] , \wRegInB60[5] , 
        \wRegInB60[4] , \wRegInB60[3] , \wRegInB60[2] , \wRegInB60[1] , 
        \wRegInB60[0] }), .LoOut({\wRegInA61[31] , \wRegInA61[30] , 
        \wRegInA61[29] , \wRegInA61[28] , \wRegInA61[27] , \wRegInA61[26] , 
        \wRegInA61[25] , \wRegInA61[24] , \wRegInA61[23] , \wRegInA61[22] , 
        \wRegInA61[21] , \wRegInA61[20] , \wRegInA61[19] , \wRegInA61[18] , 
        \wRegInA61[17] , \wRegInA61[16] , \wRegInA61[15] , \wRegInA61[14] , 
        \wRegInA61[13] , \wRegInA61[12] , \wRegInA61[11] , \wRegInA61[10] , 
        \wRegInA61[9] , \wRegInA61[8] , \wRegInA61[7] , \wRegInA61[6] , 
        \wRegInA61[5] , \wRegInA61[4] , \wRegInA61[3] , \wRegInA61[2] , 
        \wRegInA61[1] , \wRegInA61[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_155 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink156[31] , \ScanLink156[30] , \ScanLink156[29] , 
        \ScanLink156[28] , \ScanLink156[27] , \ScanLink156[26] , 
        \ScanLink156[25] , \ScanLink156[24] , \ScanLink156[23] , 
        \ScanLink156[22] , \ScanLink156[21] , \ScanLink156[20] , 
        \ScanLink156[19] , \ScanLink156[18] , \ScanLink156[17] , 
        \ScanLink156[16] , \ScanLink156[15] , \ScanLink156[14] , 
        \ScanLink156[13] , \ScanLink156[12] , \ScanLink156[11] , 
        \ScanLink156[10] , \ScanLink156[9] , \ScanLink156[8] , 
        \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , \ScanLink156[4] , 
        \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , \ScanLink156[0] 
        }), .ScanOut({\ScanLink155[31] , \ScanLink155[30] , \ScanLink155[29] , 
        \ScanLink155[28] , \ScanLink155[27] , \ScanLink155[26] , 
        \ScanLink155[25] , \ScanLink155[24] , \ScanLink155[23] , 
        \ScanLink155[22] , \ScanLink155[21] , \ScanLink155[20] , 
        \ScanLink155[19] , \ScanLink155[18] , \ScanLink155[17] , 
        \ScanLink155[16] , \ScanLink155[15] , \ScanLink155[14] , 
        \ScanLink155[13] , \ScanLink155[12] , \ScanLink155[11] , 
        \ScanLink155[10] , \ScanLink155[9] , \ScanLink155[8] , 
        \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , \ScanLink155[4] , 
        \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , \ScanLink155[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA50[31] , \wRegInA50[30] , \wRegInA50[29] , 
        \wRegInA50[28] , \wRegInA50[27] , \wRegInA50[26] , \wRegInA50[25] , 
        \wRegInA50[24] , \wRegInA50[23] , \wRegInA50[22] , \wRegInA50[21] , 
        \wRegInA50[20] , \wRegInA50[19] , \wRegInA50[18] , \wRegInA50[17] , 
        \wRegInA50[16] , \wRegInA50[15] , \wRegInA50[14] , \wRegInA50[13] , 
        \wRegInA50[12] , \wRegInA50[11] , \wRegInA50[10] , \wRegInA50[9] , 
        \wRegInA50[8] , \wRegInA50[7] , \wRegInA50[6] , \wRegInA50[5] , 
        \wRegInA50[4] , \wRegInA50[3] , \wRegInA50[2] , \wRegInA50[1] , 
        \wRegInA50[0] }), .Out({\wAIn50[31] , \wAIn50[30] , \wAIn50[29] , 
        \wAIn50[28] , \wAIn50[27] , \wAIn50[26] , \wAIn50[25] , \wAIn50[24] , 
        \wAIn50[23] , \wAIn50[22] , \wAIn50[21] , \wAIn50[20] , \wAIn50[19] , 
        \wAIn50[18] , \wAIn50[17] , \wAIn50[16] , \wAIn50[15] , \wAIn50[14] , 
        \wAIn50[13] , \wAIn50[12] , \wAIn50[11] , \wAIn50[10] , \wAIn50[9] , 
        \wAIn50[8] , \wAIn50[7] , \wAIn50[6] , \wAIn50[5] , \wAIn50[4] , 
        \wAIn50[3] , \wAIn50[2] , \wAIn50[1] , \wAIn50[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid116[31] , \wAMid116[30] , \wAMid116[29] , \wAMid116[28] , 
        \wAMid116[27] , \wAMid116[26] , \wAMid116[25] , \wAMid116[24] , 
        \wAMid116[23] , \wAMid116[22] , \wAMid116[21] , \wAMid116[20] , 
        \wAMid116[19] , \wAMid116[18] , \wAMid116[17] , \wAMid116[16] , 
        \wAMid116[15] , \wAMid116[14] , \wAMid116[13] , \wAMid116[12] , 
        \wAMid116[11] , \wAMid116[10] , \wAMid116[9] , \wAMid116[8] , 
        \wAMid116[7] , \wAMid116[6] , \wAMid116[5] , \wAMid116[4] , 
        \wAMid116[3] , \wAMid116[2] , \wAMid116[1] , \wAMid116[0] }), .BIn({
        \wBMid116[31] , \wBMid116[30] , \wBMid116[29] , \wBMid116[28] , 
        \wBMid116[27] , \wBMid116[26] , \wBMid116[25] , \wBMid116[24] , 
        \wBMid116[23] , \wBMid116[22] , \wBMid116[21] , \wBMid116[20] , 
        \wBMid116[19] , \wBMid116[18] , \wBMid116[17] , \wBMid116[16] , 
        \wBMid116[15] , \wBMid116[14] , \wBMid116[13] , \wBMid116[12] , 
        \wBMid116[11] , \wBMid116[10] , \wBMid116[9] , \wBMid116[8] , 
        \wBMid116[7] , \wBMid116[6] , \wBMid116[5] , \wBMid116[4] , 
        \wBMid116[3] , \wBMid116[2] , \wBMid116[1] , \wBMid116[0] }), .HiOut({
        \wRegInB116[31] , \wRegInB116[30] , \wRegInB116[29] , \wRegInB116[28] , 
        \wRegInB116[27] , \wRegInB116[26] , \wRegInB116[25] , \wRegInB116[24] , 
        \wRegInB116[23] , \wRegInB116[22] , \wRegInB116[21] , \wRegInB116[20] , 
        \wRegInB116[19] , \wRegInB116[18] , \wRegInB116[17] , \wRegInB116[16] , 
        \wRegInB116[15] , \wRegInB116[14] , \wRegInB116[13] , \wRegInB116[12] , 
        \wRegInB116[11] , \wRegInB116[10] , \wRegInB116[9] , \wRegInB116[8] , 
        \wRegInB116[7] , \wRegInB116[6] , \wRegInB116[5] , \wRegInB116[4] , 
        \wRegInB116[3] , \wRegInB116[2] , \wRegInB116[1] , \wRegInB116[0] }), 
        .LoOut({\wRegInA117[31] , \wRegInA117[30] , \wRegInA117[29] , 
        \wRegInA117[28] , \wRegInA117[27] , \wRegInA117[26] , \wRegInA117[25] , 
        \wRegInA117[24] , \wRegInA117[23] , \wRegInA117[22] , \wRegInA117[21] , 
        \wRegInA117[20] , \wRegInA117[19] , \wRegInA117[18] , \wRegInA117[17] , 
        \wRegInA117[16] , \wRegInA117[15] , \wRegInA117[14] , \wRegInA117[13] , 
        \wRegInA117[12] , \wRegInA117[11] , \wRegInA117[10] , \wRegInA117[9] , 
        \wRegInA117[8] , \wRegInA117[7] , \wRegInA117[6] , \wRegInA117[5] , 
        \wRegInA117[4] , \wRegInA117[3] , \wRegInA117[2] , \wRegInA117[1] , 
        \wRegInA117[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_169 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink170[31] , \ScanLink170[30] , \ScanLink170[29] , 
        \ScanLink170[28] , \ScanLink170[27] , \ScanLink170[26] , 
        \ScanLink170[25] , \ScanLink170[24] , \ScanLink170[23] , 
        \ScanLink170[22] , \ScanLink170[21] , \ScanLink170[20] , 
        \ScanLink170[19] , \ScanLink170[18] , \ScanLink170[17] , 
        \ScanLink170[16] , \ScanLink170[15] , \ScanLink170[14] , 
        \ScanLink170[13] , \ScanLink170[12] , \ScanLink170[11] , 
        \ScanLink170[10] , \ScanLink170[9] , \ScanLink170[8] , 
        \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , \ScanLink170[4] , 
        \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , \ScanLink170[0] 
        }), .ScanOut({\ScanLink169[31] , \ScanLink169[30] , \ScanLink169[29] , 
        \ScanLink169[28] , \ScanLink169[27] , \ScanLink169[26] , 
        \ScanLink169[25] , \ScanLink169[24] , \ScanLink169[23] , 
        \ScanLink169[22] , \ScanLink169[21] , \ScanLink169[20] , 
        \ScanLink169[19] , \ScanLink169[18] , \ScanLink169[17] , 
        \ScanLink169[16] , \ScanLink169[15] , \ScanLink169[14] , 
        \ScanLink169[13] , \ScanLink169[12] , \ScanLink169[11] , 
        \ScanLink169[10] , \ScanLink169[9] , \ScanLink169[8] , 
        \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , \ScanLink169[4] , 
        \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , \ScanLink169[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA43[31] , \wRegInA43[30] , \wRegInA43[29] , 
        \wRegInA43[28] , \wRegInA43[27] , \wRegInA43[26] , \wRegInA43[25] , 
        \wRegInA43[24] , \wRegInA43[23] , \wRegInA43[22] , \wRegInA43[21] , 
        \wRegInA43[20] , \wRegInA43[19] , \wRegInA43[18] , \wRegInA43[17] , 
        \wRegInA43[16] , \wRegInA43[15] , \wRegInA43[14] , \wRegInA43[13] , 
        \wRegInA43[12] , \wRegInA43[11] , \wRegInA43[10] , \wRegInA43[9] , 
        \wRegInA43[8] , \wRegInA43[7] , \wRegInA43[6] , \wRegInA43[5] , 
        \wRegInA43[4] , \wRegInA43[3] , \wRegInA43[2] , \wRegInA43[1] , 
        \wRegInA43[0] }), .Out({\wAIn43[31] , \wAIn43[30] , \wAIn43[29] , 
        \wAIn43[28] , \wAIn43[27] , \wAIn43[26] , \wAIn43[25] , \wAIn43[24] , 
        \wAIn43[23] , \wAIn43[22] , \wAIn43[21] , \wAIn43[20] , \wAIn43[19] , 
        \wAIn43[18] , \wAIn43[17] , \wAIn43[16] , \wAIn43[15] , \wAIn43[14] , 
        \wAIn43[13] , \wAIn43[12] , \wAIn43[11] , \wAIn43[10] , \wAIn43[9] , 
        \wAIn43[8] , \wAIn43[7] , \wAIn43[6] , \wAIn43[5] , \wAIn43[4] , 
        \wAIn43[3] , \wAIn43[2] , \wAIn43[1] , \wAIn43[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_39 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink40[31] , \ScanLink40[30] , \ScanLink40[29] , 
        \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , \ScanLink40[25] , 
        \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , \ScanLink40[21] , 
        \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , \ScanLink40[17] , 
        \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , \ScanLink40[13] , 
        \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , \ScanLink40[9] , 
        \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , \ScanLink40[5] , 
        \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , \ScanLink40[1] , 
        \ScanLink40[0] }), .ScanOut({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA108[31] , \wRegInA108[30] , 
        \wRegInA108[29] , \wRegInA108[28] , \wRegInA108[27] , \wRegInA108[26] , 
        \wRegInA108[25] , \wRegInA108[24] , \wRegInA108[23] , \wRegInA108[22] , 
        \wRegInA108[21] , \wRegInA108[20] , \wRegInA108[19] , \wRegInA108[18] , 
        \wRegInA108[17] , \wRegInA108[16] , \wRegInA108[15] , \wRegInA108[14] , 
        \wRegInA108[13] , \wRegInA108[12] , \wRegInA108[11] , \wRegInA108[10] , 
        \wRegInA108[9] , \wRegInA108[8] , \wRegInA108[7] , \wRegInA108[6] , 
        \wRegInA108[5] , \wRegInA108[4] , \wRegInA108[3] , \wRegInA108[2] , 
        \wRegInA108[1] , \wRegInA108[0] }), .Out({\wAIn108[31] , \wAIn108[30] , 
        \wAIn108[29] , \wAIn108[28] , \wAIn108[27] , \wAIn108[26] , 
        \wAIn108[25] , \wAIn108[24] , \wAIn108[23] , \wAIn108[22] , 
        \wAIn108[21] , \wAIn108[20] , \wAIn108[19] , \wAIn108[18] , 
        \wAIn108[17] , \wAIn108[16] , \wAIn108[15] , \wAIn108[14] , 
        \wAIn108[13] , \wAIn108[12] , \wAIn108[11] , \wAIn108[10] , 
        \wAIn108[9] , \wAIn108[8] , \wAIn108[7] , \wAIn108[6] , \wAIn108[5] , 
        \wAIn108[4] , \wAIn108[3] , \wAIn108[2] , \wAIn108[1] , \wAIn108[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_95 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink96[31] , \ScanLink96[30] , \ScanLink96[29] , 
        \ScanLink96[28] , \ScanLink96[27] , \ScanLink96[26] , \ScanLink96[25] , 
        \ScanLink96[24] , \ScanLink96[23] , \ScanLink96[22] , \ScanLink96[21] , 
        \ScanLink96[20] , \ScanLink96[19] , \ScanLink96[18] , \ScanLink96[17] , 
        \ScanLink96[16] , \ScanLink96[15] , \ScanLink96[14] , \ScanLink96[13] , 
        \ScanLink96[12] , \ScanLink96[11] , \ScanLink96[10] , \ScanLink96[9] , 
        \ScanLink96[8] , \ScanLink96[7] , \ScanLink96[6] , \ScanLink96[5] , 
        \ScanLink96[4] , \ScanLink96[3] , \ScanLink96[2] , \ScanLink96[1] , 
        \ScanLink96[0] }), .ScanOut({\ScanLink95[31] , \ScanLink95[30] , 
        \ScanLink95[29] , \ScanLink95[28] , \ScanLink95[27] , \ScanLink95[26] , 
        \ScanLink95[25] , \ScanLink95[24] , \ScanLink95[23] , \ScanLink95[22] , 
        \ScanLink95[21] , \ScanLink95[20] , \ScanLink95[19] , \ScanLink95[18] , 
        \ScanLink95[17] , \ScanLink95[16] , \ScanLink95[15] , \ScanLink95[14] , 
        \ScanLink95[13] , \ScanLink95[12] , \ScanLink95[11] , \ScanLink95[10] , 
        \ScanLink95[9] , \ScanLink95[8] , \ScanLink95[7] , \ScanLink95[6] , 
        \ScanLink95[5] , \ScanLink95[4] , \ScanLink95[3] , \ScanLink95[2] , 
        \ScanLink95[1] , \ScanLink95[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA80[31] , \wRegInA80[30] , 
        \wRegInA80[29] , \wRegInA80[28] , \wRegInA80[27] , \wRegInA80[26] , 
        \wRegInA80[25] , \wRegInA80[24] , \wRegInA80[23] , \wRegInA80[22] , 
        \wRegInA80[21] , \wRegInA80[20] , \wRegInA80[19] , \wRegInA80[18] , 
        \wRegInA80[17] , \wRegInA80[16] , \wRegInA80[15] , \wRegInA80[14] , 
        \wRegInA80[13] , \wRegInA80[12] , \wRegInA80[11] , \wRegInA80[10] , 
        \wRegInA80[9] , \wRegInA80[8] , \wRegInA80[7] , \wRegInA80[6] , 
        \wRegInA80[5] , \wRegInA80[4] , \wRegInA80[3] , \wRegInA80[2] , 
        \wRegInA80[1] , \wRegInA80[0] }), .Out({\wAIn80[31] , \wAIn80[30] , 
        \wAIn80[29] , \wAIn80[28] , \wAIn80[27] , \wAIn80[26] , \wAIn80[25] , 
        \wAIn80[24] , \wAIn80[23] , \wAIn80[22] , \wAIn80[21] , \wAIn80[20] , 
        \wAIn80[19] , \wAIn80[18] , \wAIn80[17] , \wAIn80[16] , \wAIn80[15] , 
        \wAIn80[14] , \wAIn80[13] , \wAIn80[12] , \wAIn80[11] , \wAIn80[10] , 
        \wAIn80[9] , \wAIn80[8] , \wAIn80[7] , \wAIn80[6] , \wAIn80[5] , 
        \wAIn80[4] , \wAIn80[3] , \wAIn80[2] , \wAIn80[1] , \wAIn80[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid15[31] , \wAMid15[30] , \wAMid15[29] , \wAMid15[28] , 
        \wAMid15[27] , \wAMid15[26] , \wAMid15[25] , \wAMid15[24] , 
        \wAMid15[23] , \wAMid15[22] , \wAMid15[21] , \wAMid15[20] , 
        \wAMid15[19] , \wAMid15[18] , \wAMid15[17] , \wAMid15[16] , 
        \wAMid15[15] , \wAMid15[14] , \wAMid15[13] , \wAMid15[12] , 
        \wAMid15[11] , \wAMid15[10] , \wAMid15[9] , \wAMid15[8] , \wAMid15[7] , 
        \wAMid15[6] , \wAMid15[5] , \wAMid15[4] , \wAMid15[3] , \wAMid15[2] , 
        \wAMid15[1] , \wAMid15[0] }), .BIn({\wBMid15[31] , \wBMid15[30] , 
        \wBMid15[29] , \wBMid15[28] , \wBMid15[27] , \wBMid15[26] , 
        \wBMid15[25] , \wBMid15[24] , \wBMid15[23] , \wBMid15[22] , 
        \wBMid15[21] , \wBMid15[20] , \wBMid15[19] , \wBMid15[18] , 
        \wBMid15[17] , \wBMid15[16] , \wBMid15[15] , \wBMid15[14] , 
        \wBMid15[13] , \wBMid15[12] , \wBMid15[11] , \wBMid15[10] , 
        \wBMid15[9] , \wBMid15[8] , \wBMid15[7] , \wBMid15[6] , \wBMid15[5] , 
        \wBMid15[4] , \wBMid15[3] , \wBMid15[2] , \wBMid15[1] , \wBMid15[0] }), 
        .HiOut({\wRegInB15[31] , \wRegInB15[30] , \wRegInB15[29] , 
        \wRegInB15[28] , \wRegInB15[27] , \wRegInB15[26] , \wRegInB15[25] , 
        \wRegInB15[24] , \wRegInB15[23] , \wRegInB15[22] , \wRegInB15[21] , 
        \wRegInB15[20] , \wRegInB15[19] , \wRegInB15[18] , \wRegInB15[17] , 
        \wRegInB15[16] , \wRegInB15[15] , \wRegInB15[14] , \wRegInB15[13] , 
        \wRegInB15[12] , \wRegInB15[11] , \wRegInB15[10] , \wRegInB15[9] , 
        \wRegInB15[8] , \wRegInB15[7] , \wRegInB15[6] , \wRegInB15[5] , 
        \wRegInB15[4] , \wRegInB15[3] , \wRegInB15[2] , \wRegInB15[1] , 
        \wRegInB15[0] }), .LoOut({\wRegInA16[31] , \wRegInA16[30] , 
        \wRegInA16[29] , \wRegInA16[28] , \wRegInA16[27] , \wRegInA16[26] , 
        \wRegInA16[25] , \wRegInA16[24] , \wRegInA16[23] , \wRegInA16[22] , 
        \wRegInA16[21] , \wRegInA16[20] , \wRegInA16[19] , \wRegInA16[18] , 
        \wRegInA16[17] , \wRegInA16[16] , \wRegInA16[15] , \wRegInA16[14] , 
        \wRegInA16[13] , \wRegInA16[12] , \wRegInA16[11] , \wRegInA16[10] , 
        \wRegInA16[9] , \wRegInA16[8] , \wRegInA16[7] , \wRegInA16[6] , 
        \wRegInA16[5] , \wRegInA16[4] , \wRegInA16[3] , \wRegInA16[2] , 
        \wRegInA16[1] , \wRegInA16[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid32[31] , \wAMid32[30] , \wAMid32[29] , \wAMid32[28] , 
        \wAMid32[27] , \wAMid32[26] , \wAMid32[25] , \wAMid32[24] , 
        \wAMid32[23] , \wAMid32[22] , \wAMid32[21] , \wAMid32[20] , 
        \wAMid32[19] , \wAMid32[18] , \wAMid32[17] , \wAMid32[16] , 
        \wAMid32[15] , \wAMid32[14] , \wAMid32[13] , \wAMid32[12] , 
        \wAMid32[11] , \wAMid32[10] , \wAMid32[9] , \wAMid32[8] , \wAMid32[7] , 
        \wAMid32[6] , \wAMid32[5] , \wAMid32[4] , \wAMid32[3] , \wAMid32[2] , 
        \wAMid32[1] , \wAMid32[0] }), .BIn({\wBMid32[31] , \wBMid32[30] , 
        \wBMid32[29] , \wBMid32[28] , \wBMid32[27] , \wBMid32[26] , 
        \wBMid32[25] , \wBMid32[24] , \wBMid32[23] , \wBMid32[22] , 
        \wBMid32[21] , \wBMid32[20] , \wBMid32[19] , \wBMid32[18] , 
        \wBMid32[17] , \wBMid32[16] , \wBMid32[15] , \wBMid32[14] , 
        \wBMid32[13] , \wBMid32[12] , \wBMid32[11] , \wBMid32[10] , 
        \wBMid32[9] , \wBMid32[8] , \wBMid32[7] , \wBMid32[6] , \wBMid32[5] , 
        \wBMid32[4] , \wBMid32[3] , \wBMid32[2] , \wBMid32[1] , \wBMid32[0] }), 
        .HiOut({\wRegInB32[31] , \wRegInB32[30] , \wRegInB32[29] , 
        \wRegInB32[28] , \wRegInB32[27] , \wRegInB32[26] , \wRegInB32[25] , 
        \wRegInB32[24] , \wRegInB32[23] , \wRegInB32[22] , \wRegInB32[21] , 
        \wRegInB32[20] , \wRegInB32[19] , \wRegInB32[18] , \wRegInB32[17] , 
        \wRegInB32[16] , \wRegInB32[15] , \wRegInB32[14] , \wRegInB32[13] , 
        \wRegInB32[12] , \wRegInB32[11] , \wRegInB32[10] , \wRegInB32[9] , 
        \wRegInB32[8] , \wRegInB32[7] , \wRegInB32[6] , \wRegInB32[5] , 
        \wRegInB32[4] , \wRegInB32[3] , \wRegInB32[2] , \wRegInB32[1] , 
        \wRegInB32[0] }), .LoOut({\wRegInA33[31] , \wRegInA33[30] , 
        \wRegInA33[29] , \wRegInA33[28] , \wRegInA33[27] , \wRegInA33[26] , 
        \wRegInA33[25] , \wRegInA33[24] , \wRegInA33[23] , \wRegInA33[22] , 
        \wRegInA33[21] , \wRegInA33[20] , \wRegInA33[19] , \wRegInA33[18] , 
        \wRegInA33[17] , \wRegInA33[16] , \wRegInA33[15] , \wRegInA33[14] , 
        \wRegInA33[13] , \wRegInA33[12] , \wRegInA33[11] , \wRegInA33[10] , 
        \wRegInA33[9] , \wRegInA33[8] , \wRegInA33[7] , \wRegInA33[6] , 
        \wRegInA33[5] , \wRegInA33[4] , \wRegInA33[3] , \wRegInA33[2] , 
        \wRegInA33[1] , \wRegInA33[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_107 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink108[31] , \ScanLink108[30] , \ScanLink108[29] , 
        \ScanLink108[28] , \ScanLink108[27] , \ScanLink108[26] , 
        \ScanLink108[25] , \ScanLink108[24] , \ScanLink108[23] , 
        \ScanLink108[22] , \ScanLink108[21] , \ScanLink108[20] , 
        \ScanLink108[19] , \ScanLink108[18] , \ScanLink108[17] , 
        \ScanLink108[16] , \ScanLink108[15] , \ScanLink108[14] , 
        \ScanLink108[13] , \ScanLink108[12] , \ScanLink108[11] , 
        \ScanLink108[10] , \ScanLink108[9] , \ScanLink108[8] , 
        \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , \ScanLink108[4] , 
        \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , \ScanLink108[0] 
        }), .ScanOut({\ScanLink107[31] , \ScanLink107[30] , \ScanLink107[29] , 
        \ScanLink107[28] , \ScanLink107[27] , \ScanLink107[26] , 
        \ScanLink107[25] , \ScanLink107[24] , \ScanLink107[23] , 
        \ScanLink107[22] , \ScanLink107[21] , \ScanLink107[20] , 
        \ScanLink107[19] , \ScanLink107[18] , \ScanLink107[17] , 
        \ScanLink107[16] , \ScanLink107[15] , \ScanLink107[14] , 
        \ScanLink107[13] , \ScanLink107[12] , \ScanLink107[11] , 
        \ScanLink107[10] , \ScanLink107[9] , \ScanLink107[8] , 
        \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , \ScanLink107[4] , 
        \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , \ScanLink107[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA74[31] , \wRegInA74[30] , \wRegInA74[29] , 
        \wRegInA74[28] , \wRegInA74[27] , \wRegInA74[26] , \wRegInA74[25] , 
        \wRegInA74[24] , \wRegInA74[23] , \wRegInA74[22] , \wRegInA74[21] , 
        \wRegInA74[20] , \wRegInA74[19] , \wRegInA74[18] , \wRegInA74[17] , 
        \wRegInA74[16] , \wRegInA74[15] , \wRegInA74[14] , \wRegInA74[13] , 
        \wRegInA74[12] , \wRegInA74[11] , \wRegInA74[10] , \wRegInA74[9] , 
        \wRegInA74[8] , \wRegInA74[7] , \wRegInA74[6] , \wRegInA74[5] , 
        \wRegInA74[4] , \wRegInA74[3] , \wRegInA74[2] , \wRegInA74[1] , 
        \wRegInA74[0] }), .Out({\wAIn74[31] , \wAIn74[30] , \wAIn74[29] , 
        \wAIn74[28] , \wAIn74[27] , \wAIn74[26] , \wAIn74[25] , \wAIn74[24] , 
        \wAIn74[23] , \wAIn74[22] , \wAIn74[21] , \wAIn74[20] , \wAIn74[19] , 
        \wAIn74[18] , \wAIn74[17] , \wAIn74[16] , \wAIn74[15] , \wAIn74[14] , 
        \wAIn74[13] , \wAIn74[12] , \wAIn74[11] , \wAIn74[10] , \wAIn74[9] , 
        \wAIn74[8] , \wAIn74[7] , \wAIn74[6] , \wAIn74[5] , \wAIn74[4] , 
        \wAIn74[3] , \wAIn74[2] , \wAIn74[1] , \wAIn74[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_57 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink58[31] , \ScanLink58[30] , \ScanLink58[29] , 
        \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , \ScanLink58[25] , 
        \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , \ScanLink58[21] , 
        \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , \ScanLink58[17] , 
        \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , \ScanLink58[13] , 
        \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , \ScanLink58[9] , 
        \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , \ScanLink58[5] , 
        \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , \ScanLink58[1] , 
        \ScanLink58[0] }), .ScanOut({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA99[31] , \wRegInA99[30] , 
        \wRegInA99[29] , \wRegInA99[28] , \wRegInA99[27] , \wRegInA99[26] , 
        \wRegInA99[25] , \wRegInA99[24] , \wRegInA99[23] , \wRegInA99[22] , 
        \wRegInA99[21] , \wRegInA99[20] , \wRegInA99[19] , \wRegInA99[18] , 
        \wRegInA99[17] , \wRegInA99[16] , \wRegInA99[15] , \wRegInA99[14] , 
        \wRegInA99[13] , \wRegInA99[12] , \wRegInA99[11] , \wRegInA99[10] , 
        \wRegInA99[9] , \wRegInA99[8] , \wRegInA99[7] , \wRegInA99[6] , 
        \wRegInA99[5] , \wRegInA99[4] , \wRegInA99[3] , \wRegInA99[2] , 
        \wRegInA99[1] , \wRegInA99[0] }), .Out({\wAIn99[31] , \wAIn99[30] , 
        \wAIn99[29] , \wAIn99[28] , \wAIn99[27] , \wAIn99[26] , \wAIn99[25] , 
        \wAIn99[24] , \wAIn99[23] , \wAIn99[22] , \wAIn99[21] , \wAIn99[20] , 
        \wAIn99[19] , \wAIn99[18] , \wAIn99[17] , \wAIn99[16] , \wAIn99[15] , 
        \wAIn99[14] , \wAIn99[13] , \wAIn99[12] , \wAIn99[11] , \wAIn99[10] , 
        \wAIn99[9] , \wAIn99[8] , \wAIn99[7] , \wAIn99[6] , \wAIn99[5] , 
        \wAIn99[4] , \wAIn99[3] , \wAIn99[2] , \wAIn99[1] , \wAIn99[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_237 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink238[31] , \ScanLink238[30] , \ScanLink238[29] , 
        \ScanLink238[28] , \ScanLink238[27] , \ScanLink238[26] , 
        \ScanLink238[25] , \ScanLink238[24] , \ScanLink238[23] , 
        \ScanLink238[22] , \ScanLink238[21] , \ScanLink238[20] , 
        \ScanLink238[19] , \ScanLink238[18] , \ScanLink238[17] , 
        \ScanLink238[16] , \ScanLink238[15] , \ScanLink238[14] , 
        \ScanLink238[13] , \ScanLink238[12] , \ScanLink238[11] , 
        \ScanLink238[10] , \ScanLink238[9] , \ScanLink238[8] , 
        \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , \ScanLink238[4] , 
        \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , \ScanLink238[0] 
        }), .ScanOut({\ScanLink237[31] , \ScanLink237[30] , \ScanLink237[29] , 
        \ScanLink237[28] , \ScanLink237[27] , \ScanLink237[26] , 
        \ScanLink237[25] , \ScanLink237[24] , \ScanLink237[23] , 
        \ScanLink237[22] , \ScanLink237[21] , \ScanLink237[20] , 
        \ScanLink237[19] , \ScanLink237[18] , \ScanLink237[17] , 
        \ScanLink237[16] , \ScanLink237[15] , \ScanLink237[14] , 
        \ScanLink237[13] , \ScanLink237[12] , \ScanLink237[11] , 
        \ScanLink237[10] , \ScanLink237[9] , \ScanLink237[8] , 
        \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , \ScanLink237[4] , 
        \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , \ScanLink237[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInA9[31] , \wRegInA9[30] , \wRegInA9[29] , \wRegInA9[28] , 
        \wRegInA9[27] , \wRegInA9[26] , \wRegInA9[25] , \wRegInA9[24] , 
        \wRegInA9[23] , \wRegInA9[22] , \wRegInA9[21] , \wRegInA9[20] , 
        \wRegInA9[19] , \wRegInA9[18] , \wRegInA9[17] , \wRegInA9[16] , 
        \wRegInA9[15] , \wRegInA9[14] , \wRegInA9[13] , \wRegInA9[12] , 
        \wRegInA9[11] , \wRegInA9[10] , \wRegInA9[9] , \wRegInA9[8] , 
        \wRegInA9[7] , \wRegInA9[6] , \wRegInA9[5] , \wRegInA9[4] , 
        \wRegInA9[3] , \wRegInA9[2] , \wRegInA9[1] , \wRegInA9[0] }), .Out({
        \wAIn9[31] , \wAIn9[30] , \wAIn9[29] , \wAIn9[28] , \wAIn9[27] , 
        \wAIn9[26] , \wAIn9[25] , \wAIn9[24] , \wAIn9[23] , \wAIn9[22] , 
        \wAIn9[21] , \wAIn9[20] , \wAIn9[19] , \wAIn9[18] , \wAIn9[17] , 
        \wAIn9[16] , \wAIn9[15] , \wAIn9[14] , \wAIn9[13] , \wAIn9[12] , 
        \wAIn9[11] , \wAIn9[10] , \wAIn9[9] , \wAIn9[8] , \wAIn9[7] , 
        \wAIn9[6] , \wAIn9[5] , \wAIn9[4] , \wAIn9[3] , \wAIn9[2] , \wAIn9[1] , 
        \wAIn9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_210 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink211[31] , \ScanLink211[30] , \ScanLink211[29] , 
        \ScanLink211[28] , \ScanLink211[27] , \ScanLink211[26] , 
        \ScanLink211[25] , \ScanLink211[24] , \ScanLink211[23] , 
        \ScanLink211[22] , \ScanLink211[21] , \ScanLink211[20] , 
        \ScanLink211[19] , \ScanLink211[18] , \ScanLink211[17] , 
        \ScanLink211[16] , \ScanLink211[15] , \ScanLink211[14] , 
        \ScanLink211[13] , \ScanLink211[12] , \ScanLink211[11] , 
        \ScanLink211[10] , \ScanLink211[9] , \ScanLink211[8] , 
        \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , \ScanLink211[4] , 
        \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , \ScanLink211[0] 
        }), .ScanOut({\ScanLink210[31] , \ScanLink210[30] , \ScanLink210[29] , 
        \ScanLink210[28] , \ScanLink210[27] , \ScanLink210[26] , 
        \ScanLink210[25] , \ScanLink210[24] , \ScanLink210[23] , 
        \ScanLink210[22] , \ScanLink210[21] , \ScanLink210[20] , 
        \ScanLink210[19] , \ScanLink210[18] , \ScanLink210[17] , 
        \ScanLink210[16] , \ScanLink210[15] , \ScanLink210[14] , 
        \ScanLink210[13] , \ScanLink210[12] , \ScanLink210[11] , 
        \ScanLink210[10] , \ScanLink210[9] , \ScanLink210[8] , 
        \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , \ScanLink210[4] , 
        \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , \ScanLink210[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB22[31] , \wRegInB22[30] , \wRegInB22[29] , 
        \wRegInB22[28] , \wRegInB22[27] , \wRegInB22[26] , \wRegInB22[25] , 
        \wRegInB22[24] , \wRegInB22[23] , \wRegInB22[22] , \wRegInB22[21] , 
        \wRegInB22[20] , \wRegInB22[19] , \wRegInB22[18] , \wRegInB22[17] , 
        \wRegInB22[16] , \wRegInB22[15] , \wRegInB22[14] , \wRegInB22[13] , 
        \wRegInB22[12] , \wRegInB22[11] , \wRegInB22[10] , \wRegInB22[9] , 
        \wRegInB22[8] , \wRegInB22[7] , \wRegInB22[6] , \wRegInB22[5] , 
        \wRegInB22[4] , \wRegInB22[3] , \wRegInB22[2] , \wRegInB22[1] , 
        \wRegInB22[0] }), .Out({\wBIn22[31] , \wBIn22[30] , \wBIn22[29] , 
        \wBIn22[28] , \wBIn22[27] , \wBIn22[26] , \wBIn22[25] , \wBIn22[24] , 
        \wBIn22[23] , \wBIn22[22] , \wBIn22[21] , \wBIn22[20] , \wBIn22[19] , 
        \wBIn22[18] , \wBIn22[17] , \wBIn22[16] , \wBIn22[15] , \wBIn22[14] , 
        \wBIn22[13] , \wBIn22[12] , \wBIn22[11] , \wBIn22[10] , \wBIn22[9] , 
        \wBIn22[8] , \wBIn22[7] , \wBIn22[6] , \wBIn22[5] , \wBIn22[4] , 
        \wBIn22[3] , \wBIn22[2] , \wBIn22[1] , \wBIn22[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_120 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink121[31] , \ScanLink121[30] , \ScanLink121[29] , 
        \ScanLink121[28] , \ScanLink121[27] , \ScanLink121[26] , 
        \ScanLink121[25] , \ScanLink121[24] , \ScanLink121[23] , 
        \ScanLink121[22] , \ScanLink121[21] , \ScanLink121[20] , 
        \ScanLink121[19] , \ScanLink121[18] , \ScanLink121[17] , 
        \ScanLink121[16] , \ScanLink121[15] , \ScanLink121[14] , 
        \ScanLink121[13] , \ScanLink121[12] , \ScanLink121[11] , 
        \ScanLink121[10] , \ScanLink121[9] , \ScanLink121[8] , 
        \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , \ScanLink121[4] , 
        \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , \ScanLink121[0] 
        }), .ScanOut({\ScanLink120[31] , \ScanLink120[30] , \ScanLink120[29] , 
        \ScanLink120[28] , \ScanLink120[27] , \ScanLink120[26] , 
        \ScanLink120[25] , \ScanLink120[24] , \ScanLink120[23] , 
        \ScanLink120[22] , \ScanLink120[21] , \ScanLink120[20] , 
        \ScanLink120[19] , \ScanLink120[18] , \ScanLink120[17] , 
        \ScanLink120[16] , \ScanLink120[15] , \ScanLink120[14] , 
        \ScanLink120[13] , \ScanLink120[12] , \ScanLink120[11] , 
        \ScanLink120[10] , \ScanLink120[9] , \ScanLink120[8] , 
        \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , \ScanLink120[4] , 
        \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , \ScanLink120[0] 
        }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Enable(\wEnable[0] ), 
        .In({\wRegInB67[31] , \wRegInB67[30] , \wRegInB67[29] , 
        \wRegInB67[28] , \wRegInB67[27] , \wRegInB67[26] , \wRegInB67[25] , 
        \wRegInB67[24] , \wRegInB67[23] , \wRegInB67[22] , \wRegInB67[21] , 
        \wRegInB67[20] , \wRegInB67[19] , \wRegInB67[18] , \wRegInB67[17] , 
        \wRegInB67[16] , \wRegInB67[15] , \wRegInB67[14] , \wRegInB67[13] , 
        \wRegInB67[12] , \wRegInB67[11] , \wRegInB67[10] , \wRegInB67[9] , 
        \wRegInB67[8] , \wRegInB67[7] , \wRegInB67[6] , \wRegInB67[5] , 
        \wRegInB67[4] , \wRegInB67[3] , \wRegInB67[2] , \wRegInB67[1] , 
        \wRegInB67[0] }), .Out({\wBIn67[31] , \wBIn67[30] , \wBIn67[29] , 
        \wBIn67[28] , \wBIn67[27] , \wBIn67[26] , \wBIn67[25] , \wBIn67[24] , 
        \wBIn67[23] , \wBIn67[22] , \wBIn67[21] , \wBIn67[20] , \wBIn67[19] , 
        \wBIn67[18] , \wBIn67[17] , \wBIn67[16] , \wBIn67[15] , \wBIn67[14] , 
        \wBIn67[13] , \wBIn67[12] , \wBIn67[11] , \wBIn67[10] , \wBIn67[9] , 
        \wBIn67[8] , \wBIn67[7] , \wBIn67[6] , \wBIn67[5] , \wBIn67[4] , 
        \wBIn67[3] , \wBIn67[2] , \wBIn67[1] , \wBIn67[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_70 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink71[31] , \ScanLink71[30] , \ScanLink71[29] , 
        \ScanLink71[28] , \ScanLink71[27] , \ScanLink71[26] , \ScanLink71[25] , 
        \ScanLink71[24] , \ScanLink71[23] , \ScanLink71[22] , \ScanLink71[21] , 
        \ScanLink71[20] , \ScanLink71[19] , \ScanLink71[18] , \ScanLink71[17] , 
        \ScanLink71[16] , \ScanLink71[15] , \ScanLink71[14] , \ScanLink71[13] , 
        \ScanLink71[12] , \ScanLink71[11] , \ScanLink71[10] , \ScanLink71[9] , 
        \ScanLink71[8] , \ScanLink71[7] , \ScanLink71[6] , \ScanLink71[5] , 
        \ScanLink71[4] , \ScanLink71[3] , \ScanLink71[2] , \ScanLink71[1] , 
        \ScanLink71[0] }), .ScanOut({\ScanLink70[31] , \ScanLink70[30] , 
        \ScanLink70[29] , \ScanLink70[28] , \ScanLink70[27] , \ScanLink70[26] , 
        \ScanLink70[25] , \ScanLink70[24] , \ScanLink70[23] , \ScanLink70[22] , 
        \ScanLink70[21] , \ScanLink70[20] , \ScanLink70[19] , \ScanLink70[18] , 
        \ScanLink70[17] , \ScanLink70[16] , \ScanLink70[15] , \ScanLink70[14] , 
        \ScanLink70[13] , \ScanLink70[12] , \ScanLink70[11] , \ScanLink70[10] , 
        \ScanLink70[9] , \ScanLink70[8] , \ScanLink70[7] , \ScanLink70[6] , 
        \ScanLink70[5] , \ScanLink70[4] , \ScanLink70[3] , \ScanLink70[2] , 
        \ScanLink70[1] , \ScanLink70[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB92[31] , \wRegInB92[30] , 
        \wRegInB92[29] , \wRegInB92[28] , \wRegInB92[27] , \wRegInB92[26] , 
        \wRegInB92[25] , \wRegInB92[24] , \wRegInB92[23] , \wRegInB92[22] , 
        \wRegInB92[21] , \wRegInB92[20] , \wRegInB92[19] , \wRegInB92[18] , 
        \wRegInB92[17] , \wRegInB92[16] , \wRegInB92[15] , \wRegInB92[14] , 
        \wRegInB92[13] , \wRegInB92[12] , \wRegInB92[11] , \wRegInB92[10] , 
        \wRegInB92[9] , \wRegInB92[8] , \wRegInB92[7] , \wRegInB92[6] , 
        \wRegInB92[5] , \wRegInB92[4] , \wRegInB92[3] , \wRegInB92[2] , 
        \wRegInB92[1] , \wRegInB92[0] }), .Out({\wBIn92[31] , \wBIn92[30] , 
        \wBIn92[29] , \wBIn92[28] , \wBIn92[27] , \wBIn92[26] , \wBIn92[25] , 
        \wBIn92[24] , \wBIn92[23] , \wBIn92[22] , \wBIn92[21] , \wBIn92[20] , 
        \wBIn92[19] , \wBIn92[18] , \wBIn92[17] , \wBIn92[16] , \wBIn92[15] , 
        \wBIn92[14] , \wBIn92[13] , \wBIn92[12] , \wBIn92[11] , \wBIn92[10] , 
        \wBIn92[9] , \wBIn92[8] , \wBIn92[7] , \wBIn92[6] , \wBIn92[5] , 
        \wBIn92[4] , \wBIn92[3] , \wBIn92[2] , \wBIn92[1] , \wBIn92[0] }) );
endmodule

