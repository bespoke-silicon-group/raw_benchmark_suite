
module BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, Out, Enable1, Enable2, In1, In2
     );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  Clk, Reset, RD, WR, ScanEnable, Enable1, Enable2;
    wire \ScanOut[31] , n288, \ScanOut[5]1 , \ScanOut[4]1 , n245, n287, n262, 
        n279, n217, n230, \ScanOut[10]1 , n302, n222, n305, n257, n270, n295, 
        n239, n292, \ScanOut[23]1 , \ScanOut[8]1 , n219, n225, n250, n277, 
        n289, n237, n259, \ScanOut[22]1 , \ScanOut[11]1 , n265, n242, 
        \ScanOut[9]1 , n310, n280, n224, n276, n303, n251, n293, 
        \ScanOut[19]1 , n218, n311, n281, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , n264, \ScanOut[0]1 , n243, n258, \ScanOut[15]1 , n236, 
        n216, n231, n278, \ScanOut[27]1 , n244, \ScanOut[14]1 , n263, n316, 
        n286, n304, n294, n271, n238, n256, n223, n233, n228, n314, n284, n214, 
        n246, n261, \ScanOut[28]1 , n221, \ScanOut[3]1 , n268, \ScanOut[30]1 , 
        \ScanOut[29]1 , \ScanOut[2]1 , n254, n273, n306, n296, n301, n291, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, n274, 
        \ScanOut[16]1 , n226, n234, n308, n298, n241, n313, n266, n283, 
        \ScanOut[6]1 , n227, n249, \ScanOut[7]1 , n312, n300, n252, n290, n275, 
        n282, n215, n309, n235, n240, n267, n299, \ScanOut[13]1 , n232, n247, 
        n260, \ScanOut[21]1 , n315, n285, n229, n307, n297, \ScanOut[12]1 , 
        n272, n255, n269, \ScanOut[20]1 , n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_OR2 U54 ( .A(n258), .B(n259), .Z(n294) );
    VMW_AO22 U73 ( .A(In1[7]), .B(n281), .C(In2[7]), .D(n280), .Z(n228) );
    VMW_AO22 U113 ( .A(In1[18]), .B(n281), .C(In2[18]), .D(n280), .Z(n250) );
    VMW_INV U134 ( .A(Enable1), .Z(n282) );
    VMW_NOR4 U68 ( .A(Enable1), .B(Enable2), .C(ScanEnable), .D(Reset), .Z(
        n279) );
    VMW_AO22 U96 ( .A(\ScanOut[26]1 ), .B(n279), .C(ScanIn[26]), .D(n283), .Z(
        n267) );
    VMW_AO22 U108 ( .A(\ScanOut[20]1 ), .B(n279), .C(ScanIn[20]), .D(n283), 
        .Z(n255) );
    VMW_OR2 U33 ( .A(n216), .B(n217), .Z(n315) );
    VMW_OR2 U34 ( .A(n218), .B(n219), .Z(n314) );
    VMW_OR2 U41 ( .A(n232), .B(n233), .Z(n307) );
    VMW_OR2 U46 ( .A(n242), .B(n243), .Z(n302) );
    VMW_OR2 U61 ( .A(n272), .B(n273), .Z(n287) );
    VMW_AO22 U84 ( .A(\ScanOut[31] ), .B(n279), .C(ScanIn[31]), .D(n283), .Z(
        n277) );
    VMW_AO22 U101 ( .A(In1[23]), .B(n281), .C(In2[23]), .D(n280), .Z(n260) );
    VMW_AO22 U126 ( .A(\ScanOut[12]1 ), .B(n279), .C(ScanIn[12]), .D(n283), 
        .Z(n239) );
    VMW_NOR2 U66 ( .A(n278), .B(n282), .Z(n281) );
    VMW_AO22 U106 ( .A(\ScanOut[21]1 ), .B(n279), .C(ScanIn[21]), .D(n283), 
        .Z(n257) );
    VMW_AO22 U121 ( .A(In1[14]), .B(n281), .C(In2[14]), .D(n280), .Z(n242) );
    VMW_AO22 U83 ( .A(In1[31]), .B(n281), .C(In2[31]), .D(n280), .Z(n276) );
    VMW_AO22 U98 ( .A(\ScanOut[25]1 ), .B(n279), .C(ScanIn[25]), .D(n283), .Z(
        n265) );
    VMW_OR2 U35 ( .A(n220), .B(n221), .Z(n313) );
    VMW_OR2 U48 ( .A(n246), .B(n247), .Z(n300) );
    VMW_AO22 U128 ( .A(\ScanOut[11]1 ), .B(n279), .C(ScanIn[11]), .D(n283), 
        .Z(n237) );
    VMW_OR2 U53 ( .A(n256), .B(n257), .Z(n295) );
    VMW_AO22 U91 ( .A(In1[28]), .B(n281), .C(In2[28]), .D(n280), .Z(n270) );
    VMW_AO22 U74 ( .A(\ScanOut[7]1 ), .B(n279), .C(ScanIn[7]), .D(n283), .Z(
        n229) );
    VMW_AO22 U114 ( .A(\ScanOut[18]1 ), .B(n279), .C(ScanIn[18]), .D(n283), 
        .Z(n251) );
    VMW_INV U133 ( .A(ScanEnable), .Z(n284) );
    VMW_AO22 U99 ( .A(In1[24]), .B(n281), .C(In2[24]), .D(n280), .Z(n262) );
    VMW_FD \Out_reg[25]  ( .D(n291), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n300), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_OR2 U32 ( .A(n214), .B(n215), .Z(n316) );
    VMW_OR2 U40 ( .A(n230), .B(n231), .Z(n308) );
    VMW_AO22 U82 ( .A(\ScanOut[3]1 ), .B(n279), .C(ScanIn[3]), .D(n283), .Z(
        n221) );
    VMW_FD \Out_reg[5]  ( .D(n311), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_OR2 U47 ( .A(n244), .B(n245), .Z(n301) );
    VMW_OR2 U49 ( .A(n248), .B(n249), .Z(n299) );
    VMW_OR2 U52 ( .A(n254), .B(n255), .Z(n296) );
    VMW_NOR2 U67 ( .A(n284), .B(Reset), .Z(n283) );
    VMW_AO22 U107 ( .A(In1[20]), .B(n281), .C(In2[20]), .D(n280), .Z(n254) );
    VMW_AO22 U120 ( .A(\ScanOut[15]1 ), .B(n279), .C(ScanIn[15]), .D(n283), 
        .Z(n245) );
    VMW_AO22 U75 ( .A(In1[6]), .B(n281), .C(In2[6]), .D(n280), .Z(n226) );
    VMW_AO22 U115 ( .A(In1[17]), .B(n281), .C(In2[17]), .D(n280), .Z(n248) );
    VMW_AO22 U132 ( .A(\ScanOut[0]1 ), .B(n279), .C(ScanIn[0]), .D(n283), .Z(
        n215) );
    VMW_FD \Out_reg[12]  ( .D(n304), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(\ScanOut[29]1 ), .B(n279), .C(ScanIn[29]), .D(n283), .Z(
        n273) );
    VMW_FD \Out_reg[21]  ( .D(n295), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_AO22 U129 ( .A(In1[10]), .B(n281), .C(In2[10]), .D(n280), .Z(n234) );
    VMW_FD \Out_reg[31]  ( .D(n285), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n288), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n308), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n315), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_OR2 U55 ( .A(n260), .B(n261), .Z(n293) );
    VMW_AO22 U69 ( .A(In1[9]), .B(n281), .C(In2[9]), .D(n280), .Z(n232) );
    VMW_AO22 U109 ( .A(In1[1]), .B(n281), .C(In2[1]), .D(n280), .Z(n216) );
    VMW_FD \Out_reg[19]  ( .D(n297), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(\ScanOut[8]1 ), .B(n279), .C(ScanIn[8]), .D(n283), .Z(
        n231) );
    VMW_AO22 U97 ( .A(In1[25]), .B(n281), .C(In2[25]), .D(n280), .Z(n264) );
    VMW_FD \Out_reg[3]  ( .D(n313), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_AO22 U112 ( .A(\ScanOut[19]1 ), .B(n279), .C(ScanIn[19]), .D(n283), 
        .Z(n253) );
    VMW_FD \Out_reg[23]  ( .D(n293), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n306), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_OR2 U60 ( .A(n270), .B(n271), .Z(n288) );
    VMW_FD \Out_reg[7]  ( .D(n309), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO22 U100 ( .A(\ScanOut[24]1 ), .B(n279), .C(ScanIn[24]), .D(n283), 
        .Z(n263) );
    VMW_AO22 U127 ( .A(In1[11]), .B(n281), .C(In2[11]), .D(n280), .Z(n236) );
    VMW_AO22 U85 ( .A(In1[30]), .B(n281), .C(In2[30]), .D(n280), .Z(n274) );
    VMW_FD \Out_reg[27]  ( .D(n289), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n302), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_OR2 U36 ( .A(n222), .B(n223), .Z(n312) );
    VMW_OR2 U37 ( .A(n224), .B(n225), .Z(n311) );
    VMW_OR2 U39 ( .A(n228), .B(n229), .Z(n309) );
    VMW_OR2 U57 ( .A(n264), .B(n265), .Z(n291) );
    VMW_FD \Out_reg[6]  ( .D(n310), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(\ScanOut[9]1 ), .B(n279), .C(ScanIn[9]), .D(n283), .Z(
        n233) );
    VMW_AO22 U110 ( .A(\ScanOut[1]1 ), .B(n279), .C(ScanIn[1]), .D(n283), .Z(
        n217) );
    VMW_OR2 U42 ( .A(n234), .B(n235), .Z(n306) );
    VMW_OR2 U45 ( .A(n240), .B(n241), .Z(n303) );
    VMW_AO22 U79 ( .A(In1[4]), .B(n281), .C(In2[4]), .D(n280), .Z(n222) );
    VMW_AO22 U95 ( .A(In1[26]), .B(n281), .C(In2[26]), .D(n280), .Z(n266) );
    VMW_AO22 U119 ( .A(In1[15]), .B(n281), .C(In2[15]), .D(n280), .Z(n244) );
    VMW_FD \Out_reg[26]  ( .D(n290), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n301), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n298), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO22 U87 ( .A(In1[2]), .B(n281), .C(In2[2]), .D(n280), .Z(n218) );
    VMW_FD \Out_reg[2]  ( .D(n314), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_AO22 U125 ( .A(In1[12]), .B(n281), .C(In2[12]), .D(n280), .Z(n238) );
    VMW_FD \Out_reg[11]  ( .D(n305), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_OR2 U62 ( .A(n274), .B(n275), .Z(n286) );
    VMW_FD \Out_reg[22]  ( .D(n294), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_NOR2 U65 ( .A(Enable1), .B(n278), .Z(n280) );
    VMW_AO22 U102 ( .A(\ScanOut[23]1 ), .B(n279), .C(ScanIn[23]), .D(n283), 
        .Z(n261) );
    VMW_AO22 U105 ( .A(In1[21]), .B(n281), .C(In2[21]), .D(n280), .Z(n256) );
    VMW_FD \Out_reg[20]  ( .D(n296), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n303), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(\ScanOut[4]1 ), .B(n279), .C(ScanIn[4]), .D(n283), .Z(
        n223) );
    VMW_AO22 U122 ( .A(\ScanOut[14]1 ), .B(n279), .C(ScanIn[14]), .D(n283), 
        .Z(n243) );
    VMW_FD \Out_reg[9]  ( .D(n307), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_OR2 U50 ( .A(n250), .B(n251), .Z(n298) );
    VMW_OR2 U59 ( .A(n268), .B(n269), .Z(n289) );
    VMW_FD \Out_reg[30]  ( .D(n286), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n316), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n287), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(In1[5]), .B(n281), .C(In2[5]), .D(n280), .Z(n224) );
    VMW_AO22 U89 ( .A(In1[29]), .B(n281), .C(In2[29]), .D(n280), .Z(n272) );
    VMW_AO22 U92 ( .A(\ScanOut[28]1 ), .B(n279), .C(ScanIn[28]), .D(n283), .Z(
        n271) );
    VMW_FD \Out_reg[24]  ( .D(n292), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n299), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_AO22 U117 ( .A(In1[16]), .B(n281), .C(In2[16]), .D(n280), .Z(n246) );
    VMW_FD \Out_reg[4]  ( .D(n312), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_OR2 U58 ( .A(n266), .B(n267), .Z(n290) );
    VMW_AO22 U130 ( .A(\ScanOut[10]1 ), .B(n279), .C(ScanIn[10]), .D(n283), 
        .Z(n235) );
    VMW_OR2 U38 ( .A(n226), .B(n227), .Z(n310) );
    VMW_OR2 U43 ( .A(n236), .B(n237), .Z(n305) );
    VMW_OR3 U64 ( .A(Reset), .B(ScanEnable), .C(n279), .Z(n278) );
    VMW_AO22 U81 ( .A(In1[3]), .B(n281), .C(In2[3]), .D(n280), .Z(n220) );
    VMW_AO22 U104 ( .A(\ScanOut[22]1 ), .B(n279), .C(ScanIn[22]), .D(n283), 
        .Z(n259) );
    VMW_OR2 U51 ( .A(n252), .B(n253), .Z(n297) );
    VMW_AO22 U76 ( .A(\ScanOut[6]1 ), .B(n279), .C(ScanIn[6]), .D(n283), .Z(
        n227) );
    VMW_AO22 U116 ( .A(\ScanOut[17]1 ), .B(n279), .C(ScanIn[17]), .D(n283), 
        .Z(n249) );
    VMW_AO22 U123 ( .A(In1[13]), .B(n281), .C(In2[13]), .D(n280), .Z(n240) );
    VMW_AO22 U88 ( .A(\ScanOut[2]1 ), .B(n279), .C(ScanIn[2]), .D(n283), .Z(
        n219) );
    VMW_AO22 U93 ( .A(In1[27]), .B(n281), .C(In2[27]), .D(n280), .Z(n268) );
    VMW_AO22 U131 ( .A(In1[0]), .B(n281), .C(In2[0]), .D(n280), .Z(n214) );
    VMW_OR2 U44 ( .A(n238), .B(n239), .Z(n304) );
    VMW_OR2 U56 ( .A(n262), .B(n263), .Z(n292) );
    VMW_AO22 U94 ( .A(\ScanOut[27]1 ), .B(n279), .C(ScanIn[27]), .D(n283), .Z(
        n269) );
    VMW_AO22 U71 ( .A(In1[8]), .B(n281), .C(In2[8]), .D(n280), .Z(n230) );
    VMW_AO22 U111 ( .A(In1[19]), .B(n281), .C(In2[19]), .D(n280), .Z(n252) );
    VMW_AO22 U124 ( .A(\ScanOut[13]1 ), .B(n279), .C(ScanIn[13]), .D(n283), 
        .Z(n241) );
    VMW_OR2 U63 ( .A(n276), .B(n277), .Z(n285) );
    VMW_AO22 U78 ( .A(\ScanOut[5]1 ), .B(n279), .C(ScanIn[5]), .D(n283), .Z(
        n225) );
    VMW_AO22 U86 ( .A(\ScanOut[30]1 ), .B(n279), .C(ScanIn[30]), .D(n283), .Z(
        n275) );
    VMW_AO22 U103 ( .A(In1[22]), .B(n281), .C(In2[22]), .D(n280), .Z(n258) );
    VMW_AO22 U118 ( .A(\ScanOut[16]1 ), .B(n279), .C(ScanIn[16]), .D(n283), 
        .Z(n247) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_3 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n115, n107, n52, n75, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, n118, n94, 
        n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, 
        n116, n104, n18, n24, n88, n37, n51, n93, n59, n76, n117, n80, n42, 
        n65, n19, n50, n77, n89, n25, n102, n105, n22, n39, n95, n45, n57, n70, 
        n62, n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n99), .Z(n103) );
    VMW_INV U73 ( .A(B[27]), .Z(n109) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n117) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n114), .B(A[29]), .Z(n115) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n91), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n102), .C(n96), .D(n89), .Z(n101) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n99) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n114) );
    VMW_NAND2 U52 ( .A(n99), .B(B[26]), .Z(n97) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n94), .C(n88), .D(n83), .Z(n93) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n105), .C(n103), .D(n101), .Z(n104) );
    VMW_INV U72 ( .A(A[27]), .Z(n112) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n114), .C(n111), .D(n106), .Z(n113) );
    VMW_INV U100 ( .A(B[23]), .Z(n94) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n109), .C(n104), .D(n97), .Z(n108) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n117), .C(n115), .D(n113), .Z(n116) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n112), .C(n110), .D(n108), .Z(n111) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n94), .B(A[23]), .Z(n95) );
    VMW_INV U77 ( .A(A[25]), .Z(n105) );
    VMW_INV U92 ( .A(A[28]), .Z(n107) );
    VMW_OR2 U58 ( .A(B[28]), .B(n107), .Z(n110) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n116), .B(n118), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n91), .C(n95), .D(n93), .Z(n96) );
    VMW_INV U76 ( .A(B[25]), .Z(n102) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n107), .B(B[28]), .Z(n106) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n117), .B(B[30]), .Z(n118) );
    VMW_INV U86 ( .A(A[24]), .Z(n91) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n217, n135, n205, n199, n140, n167, 
        n182, n120, n129, n185, n147, n160, n132, n202, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n218, n154, n196, n168, 
        n173, n211, n216, n126, n148, n153, n174, n183, n191, n166, n141, n134, 
        n204, n151, n193, n198, n176, n124, n214, n188, n206, n136, n143, n158, 
        n144, n164, n163, n181, n186, n178, n123, n131, n201, n213, n171, n156, 
        n130, n138, n194, n208, n179, n200, n145, n162, n187, n195, n122, n139, 
        n209, n170, n157, n125, n212, n215, n189, n150, n177, n192, n119, n142, 
        n180, n165, n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n119), .C(n120), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n124), .B(B[0]), .C(n125), .D(B[1]), .Z(n123) );
    VMW_OR2 U6 ( .A(B[2]), .B(n122), .Z(n126) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_OR2 U54 ( .A(B[26]), .B(n200), .Z(n203) );
    VMW_INV U73 ( .A(B[27]), .Z(n209) );
    VMW_INV U96 ( .A(B[31]), .Z(n119) );
    VMW_INV U68 ( .A(A[30]), .Z(n217) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n170), .C(n166), .D(n161), .Z(n169) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n125), .C(n126), .D(n123), .Z(n127) );
    VMW_NAND2 U8 ( .A(n129), .B(B[4]), .Z(n128) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n128), .Z(n137) );
    VMW_OR2 U34 ( .A(B[16]), .B(n168), .Z(n171) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n184), .C(n179), .D(n174), .Z(n183) );
    VMW_NAND2 U46 ( .A(n190), .B(A[21]), .Z(n191) );
    VMW_NAND2 U61 ( .A(n214), .B(A[29]), .Z(n215) );
    VMW_INV U84 ( .A(B[15]), .Z(n170) );
    VMW_INV U101 ( .A(A[6]), .Z(n136) );
    VMW_INV U66 ( .A(B[7]), .Z(n145) );
    VMW_INV U83 ( .A(A[15]), .Z(n173) );
    VMW_INV U98 ( .A(B[13]), .Z(n164) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_NAND2 U48 ( .A(n194), .B(B[24]), .Z(n193) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n131), .C(n127), .D(n121), .Z(n130) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n173), .C(n171), .D(n169), .Z(n172) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n202), .C(n198), .D(n193), .Z(n201) );
    VMW_INV U91 ( .A(B[11]), .Z(n158) );
    VMW_INV U74 ( .A(A[3]), .Z(n134) );
    VMW_INV U99 ( .A(A[26]), .Z(n200) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U40 ( .A(n182), .B(B[20]), .Z(n181) );
    VMW_INV U82 ( .A(B[29]), .Z(n214) );
    VMW_NAND2 U52 ( .A(n200), .B(B[26]), .Z(n199) );
    VMW_INV U67 ( .A(A[7]), .Z(n148) );
    VMW_INV U75 ( .A(B[3]), .Z(n131) );
    VMW_INV U90 ( .A(A[14]), .Z(n162) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U69 ( .A(B[17]), .Z(n177) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n205), .C(n203), .D(n201), .Z(n204) );
    VMW_INV U72 ( .A(A[27]), .Z(n212) );
    VMW_INV U97 ( .A(A[16]), .Z(n168) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n214), .C(n211), .D(n206), .Z(n213) );
    VMW_INV U100 ( .A(B[23]), .Z(n196) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_INV U85 ( .A(A[4]), .Z(n129) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_NAND2 U32 ( .A(n168), .B(B[16]), .Z(n167) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n180), .C(n178), .D(n176), .Z(n179) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n209), .C(n204), .D(n199), .Z(n208) );
    VMW_INV U70 ( .A(A[17]), .Z(n180) );
    VMW_INV U95 ( .A(A[1]), .Z(n125) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_INV U79 ( .A(B[19]), .Z(n184) );
    VMW_INV U87 ( .A(A[8]), .Z(n143) );
    VMW_OR2 U10 ( .A(B[4]), .B(n129), .Z(n132) );
    VMW_NAND2 U42 ( .A(n184), .B(A[19]), .Z(n185) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n217), .C(n215), .D(n213), .Z(n216) );
    VMW_INV U65 ( .A(A[12]), .Z(n156) );
    VMW_INV U102 ( .A(A[2]), .Z(n122) );
    VMW_INV U80 ( .A(A[10]), .Z(n150) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n132), .D(n130), .Z(n133) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n177), .C(n172), .D(n167), .Z(n176) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U89 ( .A(A[18]), .Z(n175) );
    VMW_NAND2 U50 ( .A(n196), .B(A[23]), .Z(n197) );
    VMW_INV U77 ( .A(A[25]), .Z(n205) );
    VMW_INV U92 ( .A(A[28]), .Z(n207) );
    VMW_OR2 U58 ( .A(B[28]), .B(n207), .Z(n210) );
    VMW_NAND2 U36 ( .A(n175), .B(B[18]), .Z(n174) );
    VMW_INV U81 ( .A(B[9]), .Z(n152) );
    VMW_NAND2 U4 ( .A(n122), .B(B[2]), .Z(n121) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_AO22 U64 ( .A(n216), .B(n218), .C(A[31]), .D(n119), .Z(n120) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n194), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U76 ( .A(B[25]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_INV U88 ( .A(B[21]), .Z(n190) );
    VMW_INV U93 ( .A(A[5]), .Z(n141) );
    VMW_OR2 U38 ( .A(B[18]), .B(n175), .Z(n178) );
    VMW_NAND2 U44 ( .A(n188), .B(B[22]), .Z(n187) );
    VMW_NAND2 U56 ( .A(n207), .B(B[28]), .Z(n206) );
    VMW_INV U94 ( .A(B[5]), .Z(n138) );
    VMW_INV U71 ( .A(A[22]), .Z(n188) );
    VMW_NAND2 U63 ( .A(n217), .B(B[30]), .Z(n218) );
    VMW_INV U86 ( .A(A[24]), .Z(n194) );
    VMW_INV U103 ( .A(A[0]), .Z(n124) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_INV U78 ( .A(A[20]), .Z(n182) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n287, n317, n245, n262, n279, n222, n230, n257, n270, n239, n295, 
        n305, n219, n292, n302, n250, n277, n225, n237, n289, n259, n265, n242, 
        n280, n310, n224, n288, n318, n276, n236, n243, n251, n264, n281, n293, 
        n303, n311, n258, n231, n238, n244, n278, n263, n286, n316, n294, n304, 
        n256, n271, n223, n228, n284, n314, n261, n246, n233, n221, n248, n253, 
        n254, n268, n273, n291, n296, n301, n306, n274, n226, n234, n298, n308, 
        n241, n266, n227, n283, n313, n249, n252, n275, n290, n300, n282, n312, 
        n240, n267, n232, n235, n299, n309, n247, n260, n229, n285, n315, n255, 
        n272, n297, n307, n269, n220;
    VMW_OAI21 U3 ( .A(A[31]), .B(n219), .C(n220), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_OR2 U54 ( .A(B[26]), .B(n300), .Z(n303) );
    VMW_INV U73 ( .A(B[27]), .Z(n309) );
    VMW_INV U96 ( .A(B[31]), .Z(n219) );
    VMW_INV U68 ( .A(A[30]), .Z(n317) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n270), .C(n266), .D(n261), .Z(n269) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U34 ( .A(B[16]), .B(n268), .Z(n271) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n284), .C(n279), .D(n274), .Z(n283) );
    VMW_NAND2 U46 ( .A(n290), .B(A[21]), .Z(n291) );
    VMW_NAND2 U61 ( .A(n314), .B(A[29]), .Z(n315) );
    VMW_INV U84 ( .A(B[15]), .Z(n270) );
    VMW_INV U101 ( .A(A[6]), .Z(n236) );
    VMW_INV U66 ( .A(B[7]), .Z(n245) );
    VMW_INV U83 ( .A(A[15]), .Z(n273) );
    VMW_INV U98 ( .A(B[13]), .Z(n264) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_NAND2 U48 ( .A(n294), .B(B[24]), .Z(n293) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n273), .C(n271), .D(n269), .Z(n272) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n302), .C(n298), .D(n293), .Z(n301) );
    VMW_INV U91 ( .A(B[11]), .Z(n258) );
    VMW_INV U74 ( .A(A[3]), .Z(n234) );
    VMW_INV U99 ( .A(A[26]), .Z(n300) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U40 ( .A(n282), .B(B[20]), .Z(n281) );
    VMW_INV U82 ( .A(B[29]), .Z(n314) );
    VMW_NAND2 U52 ( .A(n300), .B(B[26]), .Z(n299) );
    VMW_INV U67 ( .A(A[7]), .Z(n248) );
    VMW_INV U75 ( .A(B[3]), .Z(n231) );
    VMW_INV U90 ( .A(A[14]), .Z(n262) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n296), .C(n292), .D(n287), .Z(n295) );
    VMW_INV U69 ( .A(B[17]), .Z(n277) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n288), .C(n291), .D(n289), .Z(n292) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n305), .C(n303), .D(n301), .Z(n304) );
    VMW_INV U72 ( .A(A[27]), .Z(n312) );
    VMW_INV U97 ( .A(A[16]), .Z(n268) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n314), .C(n311), .D(n306), .Z(n313) );
    VMW_INV U100 ( .A(B[23]), .Z(n296) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_INV U85 ( .A(A[4]), .Z(n229) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_NAND2 U32 ( .A(n268), .B(B[16]), .Z(n267) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n280), .C(n278), .D(n276), .Z(n279) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n309), .C(n304), .D(n299), .Z(n308) );
    VMW_INV U70 ( .A(A[17]), .Z(n280) );
    VMW_INV U95 ( .A(A[1]), .Z(n225) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_INV U79 ( .A(B[19]), .Z(n284) );
    VMW_INV U87 ( .A(A[8]), .Z(n243) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_NAND2 U42 ( .A(n284), .B(A[19]), .Z(n285) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n290), .C(n286), .D(n281), .Z(n289) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n317), .C(n315), .D(n313), .Z(n316) );
    VMW_INV U65 ( .A(A[12]), .Z(n256) );
    VMW_INV U102 ( .A(A[2]), .Z(n222) );
    VMW_INV U80 ( .A(A[10]), .Z(n250) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n277), .C(n272), .D(n267), .Z(n276) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n312), .C(n310), .D(n308), .Z(n311) );
    VMW_INV U89 ( .A(A[18]), .Z(n275) );
    VMW_NAND2 U50 ( .A(n296), .B(A[23]), .Z(n297) );
    VMW_INV U77 ( .A(A[25]), .Z(n305) );
    VMW_INV U92 ( .A(A[28]), .Z(n307) );
    VMW_OR2 U58 ( .A(B[28]), .B(n307), .Z(n310) );
    VMW_NAND2 U36 ( .A(n275), .B(B[18]), .Z(n274) );
    VMW_INV U81 ( .A(B[9]), .Z(n252) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n282), .C(n285), .D(n283), .Z(n286) );
    VMW_AO22 U64 ( .A(n316), .B(n318), .C(A[31]), .D(n219), .Z(n220) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n294), .C(n297), .D(n295), .Z(n298) );
    VMW_INV U76 ( .A(B[25]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_INV U88 ( .A(B[21]), .Z(n290) );
    VMW_INV U93 ( .A(A[5]), .Z(n241) );
    VMW_OR2 U38 ( .A(B[18]), .B(n275), .Z(n278) );
    VMW_NAND2 U44 ( .A(n288), .B(B[22]), .Z(n287) );
    VMW_NAND2 U56 ( .A(n307), .B(B[28]), .Z(n306) );
    VMW_INV U94 ( .A(B[5]), .Z(n238) );
    VMW_INV U71 ( .A(A[22]), .Z(n288) );
    VMW_NAND2 U63 ( .A(n317), .B(B[30]), .Z(n318) );
    VMW_INV U86 ( .A(A[24]), .Z(n294) );
    VMW_INV U103 ( .A(A[0]), .Z(n224) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_INV U78 ( .A(A[20]), .Z(n282) );
endmodule


module BHeap_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n330, n379, n362, n339, n345, n387, n395, n406, n414, n370, n357, 
        n322, n319, n325, n389, n408, n350, n377, n392, n413, n342, n380, n401, 
        n359, n365, n337, n351, n393, n412, n376, n324, n336, n388, n409, n343, 
        n358, n364, n381, n400, n386, n407, n323, n331, n344, n363, n378, n356, 
        n371, n333, n338, n394, n415, n328, n346, n361, n384, n405, n396, n321, 
        n354, n368, n373, n326, n348, n353, n374, n383, n391, n410, n402, n341, 
        n366, n334, n390, n398, n411, n349, n352, n375, n327, n335, n399, n340, 
        n367, n329, n382, n403, n385, n404, n347, n360, n332, n320, n369, n355, 
        n372, n397, n416;
    VMW_OAI21 U3 ( .A(A[31]), .B(n319), .C(n320), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n322), .C(B[0]), .Z(n323) );
    VMW_AO22 U6 ( .A(A[2]), .B(n325), .C(n323), .D(A[0]), .Z(n324) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_OR2 U54 ( .A(B[26]), .B(n398), .Z(n401) );
    VMW_INV U73 ( .A(B[27]), .Z(n407) );
    VMW_INV U96 ( .A(A[16]), .Z(n366) );
    VMW_INV U68 ( .A(A[30]), .Z(n415) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n368), .C(n364), .D(n359), .Z(n367) );
    VMW_OAI22 U7 ( .A(n321), .B(n324), .C(A[2]), .D(n325), .Z(n326) );
    VMW_NAND2 U8 ( .A(n328), .B(B[4]), .Z(n327) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n332), .D(n327), .Z(n335) );
    VMW_OR2 U34 ( .A(B[16]), .B(n366), .Z(n369) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n382), .C(n377), .D(n372), .Z(n381) );
    VMW_NAND2 U46 ( .A(n388), .B(A[21]), .Z(n389) );
    VMW_NAND2 U61 ( .A(n412), .B(A[29]), .Z(n413) );
    VMW_INV U84 ( .A(A[4]), .Z(n328) );
    VMW_INV U101 ( .A(B[2]), .Z(n325) );
    VMW_INV U66 ( .A(B[7]), .Z(n343) );
    VMW_INV U83 ( .A(B[15]), .Z(n368) );
    VMW_INV U98 ( .A(A[26]), .Z(n398) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_NAND2 U48 ( .A(n392), .B(B[24]), .Z(n391) );
    VMW_AO21 U9 ( .A(B[3]), .B(n330), .C(n326), .Z(n329) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n371), .C(n369), .D(n367), .Z(n370) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n400), .C(n396), .D(n391), .Z(n399) );
    VMW_INV U91 ( .A(A[28]), .Z(n405) );
    VMW_INV U74 ( .A(A[3]), .Z(n330) );
    VMW_INV U99 ( .A(B[23]), .Z(n394) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U40 ( .A(n380), .B(B[20]), .Z(n379) );
    VMW_INV U82 ( .A(A[15]), .Z(n371) );
    VMW_NAND2 U52 ( .A(n398), .B(B[26]), .Z(n397) );
    VMW_INV U67 ( .A(A[7]), .Z(n346) );
    VMW_INV U75 ( .A(B[25]), .Z(n400) );
    VMW_INV U90 ( .A(B[11]), .Z(n356) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n394), .C(n390), .D(n385), .Z(n393) );
    VMW_INV U69 ( .A(B[17]), .Z(n375) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n386), .C(n389), .D(n387), .Z(n390) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n403), .C(n401), .D(n399), .Z(n402) );
    VMW_INV U72 ( .A(A[27]), .Z(n410) );
    VMW_INV U97 ( .A(B[13]), .Z(n362) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n412), .C(n409), .D(n404), .Z(n411) );
    VMW_INV U100 ( .A(A[6]), .Z(n334) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_INV U85 ( .A(A[24]), .Z(n392) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_NAND2 U32 ( .A(n366), .B(B[16]), .Z(n365) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n378), .C(n376), .D(n374), .Z(n377) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n407), .C(n402), .D(n397), .Z(n406) );
    VMW_INV U70 ( .A(A[17]), .Z(n378) );
    VMW_INV U95 ( .A(B[31]), .Z(n319) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_INV U79 ( .A(A[10]), .Z(n348) );
    VMW_INV U87 ( .A(B[21]), .Z(n388) );
    VMW_OR2 U10 ( .A(B[4]), .B(n328), .Z(n331) );
    VMW_NAND2 U42 ( .A(n382), .B(A[19]), .Z(n383) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n388), .C(n384), .D(n379), .Z(n387) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n415), .C(n413), .D(n411), .Z(n414) );
    VMW_INV U65 ( .A(A[12]), .Z(n354) );
    VMW_INV U80 ( .A(B[9]), .Z(n350) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n330), .C(n331), .D(n329), .Z(n332) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n375), .C(n370), .D(n365), .Z(n374) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n410), .C(n408), .D(n406), .Z(n409) );
    VMW_INV U89 ( .A(A[14]), .Z(n360) );
    VMW_NAND2 U50 ( .A(n394), .B(A[23]), .Z(n395) );
    VMW_INV U77 ( .A(A[20]), .Z(n380) );
    VMW_INV U92 ( .A(A[5]), .Z(n339) );
    VMW_OR2 U58 ( .A(B[28]), .B(n405), .Z(n408) );
    VMW_NAND2 U36 ( .A(n373), .B(B[18]), .Z(n372) );
    VMW_INV U81 ( .A(B[29]), .Z(n412) );
    VMW_NOR2 U4 ( .A(n322), .B(B[1]), .Z(n321) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n380), .C(n383), .D(n381), .Z(n384) );
    VMW_AO22 U64 ( .A(n414), .B(n416), .C(A[31]), .D(n319), .Z(n320) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n392), .C(n395), .D(n393), .Z(n396) );
    VMW_INV U76 ( .A(A[25]), .Z(n403) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_INV U88 ( .A(A[18]), .Z(n373) );
    VMW_INV U93 ( .A(B[5]), .Z(n336) );
    VMW_OR2 U38 ( .A(B[18]), .B(n373), .Z(n376) );
    VMW_NAND2 U44 ( .A(n386), .B(B[22]), .Z(n385) );
    VMW_NAND2 U56 ( .A(n405), .B(B[28]), .Z(n404) );
    VMW_INV U94 ( .A(A[1]), .Z(n322) );
    VMW_INV U71 ( .A(A[22]), .Z(n386) );
    VMW_NAND2 U63 ( .A(n415), .B(B[30]), .Z(n416) );
    VMW_INV U86 ( .A(A[8]), .Z(n341) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_INV U78 ( .A(B[19]), .Z(n382) );
endmodule


module BHeap_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Enable, 
    P_WR, P_In, P_Out, L_WR, L_In, L_Out, R_WR, R_In, R_Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] P_Out;
output [31:0] L_Out;
input  [31:0] R_In;
input  [31:0] P_In;
input  [31:0] L_In;
output [31:0] R_Out;
input  Clk, Reset, RD, WR, Enable;
output P_WR, L_WR, R_WR;
    wire n454, n100, n421, n433, n446, n428, n441, n434, n426, n448, n90, n453, 
        n435, n449, n98, n440, n452, n427, n420, n429, n447, n439, n432, n422, 
        n417, n430, n445, n442, n437, n425, n450, n419, n436, n443, n418, n451, 
        n92, n424, n423, n438, n444, n431;
    tri \P_Out[31] , \R_Out[25]1 , \R_Out[16]1 , \R_Out[24]1 , \R_Out[17]1 , 
        \P_Out[21]1 , \P_Out[12]1 , \P_Out[20]1 , \P_Out[13]1 , \P_Out[7]1 , 
        \R_Out[2]1 , \L_Out[20]1 , \L_Out[13]1 , \L_Out[6]1 , \R_Out[3]1 , 
        \R_Out[30]1 , \R_Out[29]1 , \P_Out[6]1 , \L_Out[7]1 , \R_Out[28]1 , 
        \L_Out[21]1 , \L_Out[12]1 , \P_Out[24]1 , \P_Out[17]1 , \P_Out[25]1 , 
        \P_Out[16]1 , \L_Out[30]1 , \R_Out[20]1 , \R_Out[13]1 , \L_Out[29]1 , 
        \L_Out[28]1 , \R_Out[21]1 , \R_Out[12]1 , \L_Out[3]1 , \P_Out[2]1 , 
        \L_Out[25]1 , \L_Out[16]1 , \P_Out[3]1 , \L_Out[2]1 , \L_Out[24]1 , 
        \L_Out[17]1 , \R_Out[7]1 , \P_Out[28]1 , \P_Out[30]1 , \P_Out[29]1 , 
        \R_Out[6]1 , \P_Out[26]1 , \P_Out[15]1 , \R_Out[9]1 , \R_Out[8]1 , 
        \P_Out[27]1 , \P_Out[14]1 , \L_Out[18]1 , \R_Out[22]1 , \R_Out[11]1 , 
        \P_Out[0]1 , \L_Out[27]1 , \L_Out[19]1 , \R_Out[23]1 , \R_Out[10]1 , 
        \L_Out[1]1 , \L_Out[14]1 , \L_Out[0]1 , \P_Out[1]1 , \L_Out[26]1 , 
        \L_Out[15]1 , \R_Out[5]1 , \P_Out[19]1 , \P_Out[18]1 , \L_Out[31] , 
        \P_Out[9]1 , \L_Out[8]1 , \R_Out[4]1 , \R_Out[27]1 , \R_Out[14]1 , 
        \P_Out[23]1 , \P_Out[10]1 , \P_Out[8]1 , \L_Out[9]1 , \R_Out[26]1 , 
        \R_Out[15]1 , \P_Out[22]1 , \P_Out[11]1 , \P_Out[5]1 , \R_Out[0]1 , 
        \R_Out[1]1 , \L_Out[22]1 , \L_Out[11]1 , \L_Out[4]1 , \R_Out[18]1 , 
        \R_Out[31] , \P_Out[4]1 , \L_Out[5]1 , \R_Out[19]1 , \L_Out[23]1 , 
        \L_Out[10]1 ;
    assign P_Out[31] = \P_Out[31] ;
    assign P_Out[30] = \P_Out[30]1 ;
    assign P_Out[29] = \P_Out[29]1 ;
    assign P_Out[28] = \P_Out[28]1 ;
    assign P_Out[27] = \P_Out[27]1 ;
    assign P_Out[26] = \P_Out[26]1 ;
    assign P_Out[25] = \P_Out[25]1 ;
    assign P_Out[24] = \P_Out[24]1 ;
    assign P_Out[23] = \P_Out[23]1 ;
    assign P_Out[22] = \P_Out[22]1 ;
    assign P_Out[21] = \P_Out[21]1 ;
    assign P_Out[20] = \P_Out[20]1 ;
    assign P_Out[19] = \P_Out[19]1 ;
    assign P_Out[18] = \P_Out[18]1 ;
    assign P_Out[17] = \P_Out[17]1 ;
    assign P_Out[16] = \P_Out[16]1 ;
    assign P_Out[15] = \P_Out[15]1 ;
    assign P_Out[14] = \P_Out[14]1 ;
    assign P_Out[13] = \P_Out[13]1 ;
    assign P_Out[12] = \P_Out[12]1 ;
    assign P_Out[11] = \P_Out[11]1 ;
    assign P_Out[10] = \P_Out[10]1 ;
    assign P_Out[9] = \P_Out[9]1 ;
    assign P_Out[8] = \P_Out[8]1 ;
    assign P_Out[7] = \P_Out[7]1 ;
    assign P_Out[6] = \P_Out[6]1 ;
    assign P_Out[5] = \P_Out[5]1 ;
    assign P_Out[4] = \P_Out[4]1 ;
    assign P_Out[3] = \P_Out[3]1 ;
    assign P_Out[2] = \P_Out[2]1 ;
    assign P_Out[1] = \P_Out[1]1 ;
    assign P_Out[0] = \P_Out[0]1 ;
    assign L_Out[31] = \L_Out[31] ;
    assign L_Out[30] = \L_Out[30]1 ;
    assign L_Out[29] = \L_Out[29]1 ;
    assign L_Out[28] = \L_Out[28]1 ;
    assign L_Out[27] = \L_Out[27]1 ;
    assign L_Out[26] = \L_Out[26]1 ;
    assign L_Out[25] = \L_Out[25]1 ;
    assign L_Out[24] = \L_Out[24]1 ;
    assign L_Out[23] = \L_Out[23]1 ;
    assign L_Out[22] = \L_Out[22]1 ;
    assign L_Out[21] = \L_Out[21]1 ;
    assign L_Out[20] = \L_Out[20]1 ;
    assign L_Out[19] = \L_Out[19]1 ;
    assign L_Out[18] = \L_Out[18]1 ;
    assign L_Out[17] = \L_Out[17]1 ;
    assign L_Out[16] = \L_Out[16]1 ;
    assign L_Out[15] = \L_Out[15]1 ;
    assign L_Out[14] = \L_Out[14]1 ;
    assign L_Out[13] = \L_Out[13]1 ;
    assign L_Out[12] = \L_Out[12]1 ;
    assign L_Out[11] = \L_Out[11]1 ;
    assign L_Out[10] = \L_Out[10]1 ;
    assign L_Out[9] = \L_Out[9]1 ;
    assign L_Out[8] = \L_Out[8]1 ;
    assign L_Out[7] = \L_Out[7]1 ;
    assign L_Out[6] = \L_Out[6]1 ;
    assign L_Out[5] = \L_Out[5]1 ;
    assign L_Out[4] = \L_Out[4]1 ;
    assign L_Out[3] = \L_Out[3]1 ;
    assign L_Out[2] = \L_Out[2]1 ;
    assign L_Out[1] = \L_Out[1]1 ;
    assign L_Out[0] = \L_Out[0]1 ;
    assign R_Out[31] = \R_Out[31] ;
    assign R_Out[30] = \R_Out[30]1 ;
    assign R_Out[29] = \R_Out[29]1 ;
    assign R_Out[28] = \R_Out[28]1 ;
    assign R_Out[27] = \R_Out[27]1 ;
    assign R_Out[26] = \R_Out[26]1 ;
    assign R_Out[25] = \R_Out[25]1 ;
    assign R_Out[24] = \R_Out[24]1 ;
    assign R_Out[23] = \R_Out[23]1 ;
    assign R_Out[22] = \R_Out[22]1 ;
    assign R_Out[21] = \R_Out[21]1 ;
    assign R_Out[20] = \R_Out[20]1 ;
    assign R_Out[19] = \R_Out[19]1 ;
    assign R_Out[18] = \R_Out[18]1 ;
    assign R_Out[17] = \R_Out[17]1 ;
    assign R_Out[16] = \R_Out[16]1 ;
    assign R_Out[15] = \R_Out[15]1 ;
    assign R_Out[14] = \R_Out[14]1 ;
    assign R_Out[13] = \R_Out[13]1 ;
    assign R_Out[12] = \R_Out[12]1 ;
    assign R_Out[11] = \R_Out[11]1 ;
    assign R_Out[10] = \R_Out[10]1 ;
    assign R_Out[9] = \R_Out[9]1 ;
    assign R_Out[8] = \R_Out[8]1 ;
    assign R_Out[7] = \R_Out[7]1 ;
    assign R_Out[6] = \R_Out[6]1 ;
    assign R_Out[5] = \R_Out[5]1 ;
    assign R_Out[4] = \R_Out[4]1 ;
    assign R_Out[3] = \R_Out[3]1 ;
    assign R_Out[2] = \R_Out[2]1 ;
    assign R_Out[1] = \R_Out[1]1 ;
    assign R_Out[0] = \R_Out[0]1 ;
    VMW_AO22 U54 ( .A(R_In[26]), .B(n417), .C(L_In[26]), .D(L_WR), .Z(n431) );
    VMW_AND3 U73 ( .A(n92), .B(Enable), .C(n90), .Z(L_WR) );
    VMW_BUFIZ U113 ( .A(P_In[3]), .E(L_WR), .Z(\L_Out[3]1 ) );
    VMW_BUFIZ U134 ( .A(P_In[22]), .E(R_WR), .Z(\R_Out[22]1 ) );
    VMW_AO22 U68 ( .A(R_In[13]), .B(n417), .C(L_In[13]), .D(L_WR), .Z(n426) );
    VMW_BUFIZ U96 ( .A(n421), .E(P_WR), .Z(\P_Out[17]1 ) );
    VMW_BUFIZ U108 ( .A(P_In[12]), .E(R_WR), .Z(\R_Out[12]1 ) );
    VMW_BUFIZ U141 ( .A(n444), .E(P_WR), .Z(\P_Out[3]1 ) );
    VMW_BUFIZ U166 ( .A(P_In[4]), .E(R_WR), .Z(\R_Out[4]1 ) );
    VMW_PULLDOWN U35 ( .Z(n451) );
    VMW_AO22 U41 ( .A(R_In[9]), .B(n417), .C(L_In[9]), .D(L_WR), .Z(n429) );
    VMW_AO22 U46 ( .A(R_In[4]), .B(n417), .C(L_In[4]), .D(L_WR), .Z(n433) );
    VMW_AO22 U61 ( .A(R_In[1]), .B(n417), .C(L_In[1]), .D(L_WR), .Z(n443) );
    VMW_BUFIZ U84 ( .A(P_In[24]), .E(L_WR), .Z(\L_Out[24]1 ) );
    VMW_BUFIZ U148 ( .A(P_In[13]), .E(R_WR), .Z(\R_Out[13]1 ) );
    VMW_BUFIZ U153 ( .A(n449), .E(P_WR), .Z(\P_Out[16]1 ) );
    VMW_BUFIZ U101 ( .A(n424), .E(P_WR), .Z(\P_Out[20]1 ) );
    VMW_BUFIZ U126 ( .A(n434), .E(P_WR), .Z(\P_Out[27]1 ) );
    VMW_AO22 U48 ( .A(R_In[31]), .B(n417), .C(L_In[31]), .D(L_WR), .Z(n440) );
    VMW_AO22 U66 ( .A(R_In[15]), .B(n417), .C(L_In[15]), .D(L_WR), .Z(n432) );
    VMW_BUFIZ U106 ( .A(P_In[28]), .E(R_WR), .Z(\R_Out[28]1 ) );
    VMW_BUFIZ U121 ( .A(n432), .E(P_WR), .Z(\P_Out[15]1 ) );
    VMW_BUFIZ U83 ( .A(P_In[15]), .E(L_WR), .Z(\L_Out[15]1 ) );
    VMW_BUFIZ U168 ( .A(P_In[9]), .E(R_WR), .Z(\R_Out[9]1 ) );
    VMW_BUFIZ U98 ( .A(P_In[16]), .E(R_WR), .Z(\R_Out[16]1 ) );
    VMW_BUFIZ U128 ( .A(n436), .E(P_WR), .Z(\P_Out[14]1 ) );
    VMW_BUFIZ U154 ( .A(P_In[24]), .E(R_WR), .Z(\R_Out[24]1 ) );
    VMW_AO22 U53 ( .A(R_In[27]), .B(n417), .C(L_In[27]), .D(L_WR), .Z(n434) );
    VMW_BUFIZ U91 ( .A(n420), .E(P_WR), .Z(\P_Out[6]1 ) );
    VMW_BUFIZ U146 ( .A(P_In[9]), .E(L_WR), .Z(\L_Out[9]1 ) );
    VMW_BUFIZ U161 ( .A(P_In[25]), .E(L_WR), .Z(\L_Out[25]1 ) );
    VMW_AND3 U74 ( .A(n98), .B(n100), .C(Enable), .Z(R_WR) );
    VMW_BUFIZ U114 ( .A(P_In[23]), .E(R_WR), .Z(\R_Out[23]1 ) );
    VMW_BUFIZ U133 ( .A(P_In[2]), .E(L_WR), .Z(\L_Out[2]1 ) );
    VMW_BUFIZ U99 ( .A(n422), .E(P_WR), .Z(\P_Out[29]1 ) );
    VMW_BUFIZ U155 ( .A(P_In[17]), .E(R_WR), .Z(\R_Out[17]1 ) );
    VMW_OR2 U40 ( .A(L_WR), .B(R_WR), .Z(P_WR) );
    VMW_BUFIZ U82 ( .A(P_In[26]), .E(L_WR), .Z(\L_Out[26]1 ) );
    VMW_BUFIZ U169 ( .A(P_In[23]), .E(L_WR), .Z(\L_Out[23]1 ) );
    VMW_AO22 U47 ( .A(R_In[3]), .B(n417), .C(L_In[3]), .D(L_WR), .Z(n444) );
    VMW_AO22 U49 ( .A(R_In[30]), .B(n417), .C(L_In[30]), .D(L_WR), .Z(n418) );
    VMW_AO22 U52 ( .A(R_In[28]), .B(n417), .C(L_In[28]), .D(L_WR), .Z(n441) );
    VMW_AO22 U67 ( .A(R_In[14]), .B(n417), .C(L_In[14]), .D(L_WR), .Z(n436) );
    VMW_BUFIZ U107 ( .A(P_In[21]), .E(R_WR), .Z(\R_Out[21]1 ) );
    VMW_BUFIZ U120 ( .A(n431), .E(P_WR), .Z(\P_Out[26]1 ) );
    VMW_INV U75 ( .A(L_WR), .Z(n417) );
    VMW_BUFIZ U115 ( .A(P_In[10]), .E(R_WR), .Z(\R_Out[10]1 ) );
    VMW_BUFIZ U132 ( .A(n439), .E(P_WR), .Z(\P_Out[8]1 ) );
    VMW_BUFIZ U90 ( .A(n419), .E(P_WR), .Z(\P_Out[24]1 ) );
    VMW_BUFIZ U129 ( .A(n437), .E(P_WR), .Z(\P_Out[5]1 ) );
    VMW_BUFIZ U147 ( .A(P_In[20]), .E(R_WR), .Z(\R_Out[20]1 ) );
    VMW_BUFIZ U160 ( .A(P_In[28]), .E(L_WR), .Z(\L_Out[28]1 ) );
    VMW_AO22 U55 ( .A(R_In[25]), .B(n417), .C(L_In[25]), .D(L_WR), .Z(n448) );
    VMW_AO22 U69 ( .A(R_In[12]), .B(n417), .C(L_In[12]), .D(L_WR), .Z(n446) );
    VMW_BUFIZ U109 ( .A(n426), .E(P_WR), .Z(\P_Out[13]1 ) );
    VMW_AO22 U72 ( .A(R_In[0]), .B(n417), .C(L_In[0]), .D(L_WR), .Z(n430) );
    VMW_BUFIZ U97 ( .A(P_In[25]), .E(R_WR), .Z(\R_Out[25]1 ) );
    VMW_BUFIZ U140 ( .A(n443), .E(P_WR), .Z(\P_Out[1]1 ) );
    VMW_BUFIZ U167 ( .A(P_In[19]), .E(L_WR), .Z(\L_Out[19]1 ) );
    VMW_BUFIZ U112 ( .A(n429), .E(P_WR), .Z(\P_Out[9]1 ) );
    VMW_BUFIZ U135 ( .A(P_In[11]), .E(R_WR), .Z(\R_Out[11]1 ) );
    VMW_AO22 U60 ( .A(R_In[20]), .B(n417), .C(L_In[20]), .D(L_WR), .Z(n424) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_1 gt_48_1 ( .A(L_In), .B(R_In), .LEQ(n452), 
        .TC(n452), .LT_LE(n100) );
    VMW_BUFIZ U100 ( .A(n423), .E(P_WR), .Z(\P_Out[22]1 ) );
    VMW_BUFIZ U127 ( .A(n435), .E(P_WR), .Z(\P_Out[23]1 ) );
    VMW_BUFIZ U85 ( .A(P_In[17]), .E(L_WR), .Z(\L_Out[17]1 ) );
    VMW_BUFIZ U149 ( .A(n446), .E(P_WR), .Z(\P_Out[12]1 ) );
    VMW_BUFIZ U152 ( .A(n448), .E(P_WR), .Z(\P_Out[25]1 ) );
    VMW_PULLUP U36 ( .Z(n450) );
    VMW_PULLDOWN U37 ( .Z(n452) );
    VMW_PULLDOWN U39 ( .Z(n454) );
    VMW_AO22 U57 ( .A(R_In[23]), .B(n417), .C(L_In[23]), .D(L_WR), .Z(n435) );
    VMW_BUFIZ U137 ( .A(n441), .E(P_WR), .Z(\P_Out[28]1 ) );
    VMW_AO22 U70 ( .A(R_In[11]), .B(n417), .C(L_In[11]), .D(L_WR), .Z(n428) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_2 gt_48 ( .A(P_In), .B(R_In), .LEQ(n453), 
        .TC(n453), .LT_LE(n98) );
    VMW_BUFIZ U110 ( .A(n427), .E(P_WR), .Z(\P_Out[18]1 ) );
    VMW_BUFIZ U159 ( .A(P_In[12]), .E(L_WR), .Z(\L_Out[12]1 ) );
    VMW_AO22 U42 ( .A(R_In[8]), .B(n417), .C(L_In[8]), .D(L_WR), .Z(n439) );
    VMW_AO22 U45 ( .A(R_In[5]), .B(n417), .C(L_In[5]), .D(L_WR), .Z(n437) );
    VMW_BUFIZ U79 ( .A(P_In[11]), .E(L_WR), .Z(\L_Out[11]1 ) );
    VMW_BUFIZ U95 ( .A(P_In[5]), .E(L_WR), .Z(\L_Out[5]1 ) );
    VMW_BUFIZ U119 ( .A(P_In[14]), .E(R_WR), .Z(\R_Out[14]1 ) );
    VMW_BUFIZ U142 ( .A(P_In[0]), .E(L_WR), .Z(\L_Out[0]1 ) );
    VMW_BUFIZ U165 ( .A(P_In[14]), .E(L_WR), .Z(\L_Out[14]1 ) );
    VMW_BUFIZ U87 ( .A(P_In[13]), .E(L_WR), .Z(\L_Out[13]1 ) );
    VMW_BUFIZ U150 ( .A(n447), .E(P_WR), .Z(\P_Out[7]1 ) );
    VMW_BUFIZ U125 ( .A(P_In[15]), .E(R_WR), .Z(\R_Out[15]1 ) );
    VMW_AO22 U62 ( .A(R_In[19]), .B(n417), .C(L_In[19]), .D(L_WR), .Z(n442) );
    VMW_AO22 U65 ( .A(R_In[16]), .B(n417), .C(L_In[16]), .D(L_WR), .Z(n449) );
    VMW_BUFIZ U102 ( .A(n425), .E(P_WR), .Z(\P_Out[2]1 ) );
    VMW_BUFIZ U105 ( .A(P_In[31]), .E(R_WR), .Z(\R_Out[31] ) );
    VMW_BUFIZ U80 ( .A(P_In[5]), .E(R_WR), .Z(\R_Out[5]1 ) );
    VMW_BUFIZ U122 ( .A(n433), .E(P_WR), .Z(\P_Out[4]1 ) );
    VMW_BUFIZ U157 ( .A(P_In[31]), .E(L_WR), .Z(\L_Out[31] ) );
    VMW_BUFIZ U170 ( .A(P_In[10]), .E(L_WR), .Z(\L_Out[10]1 ) );
    VMW_AO22 U50 ( .A(R_In[2]), .B(n417), .C(L_In[2]), .D(L_WR), .Z(n425) );
    VMW_AO22 U59 ( .A(R_In[21]), .B(n417), .C(L_In[21]), .D(L_WR), .Z(n445) );
    VMW_BUFIZ U139 ( .A(P_In[18]), .E(R_WR), .Z(\R_Out[18]1 ) );
    VMW_BUFIZ U77 ( .A(P_In[18]), .E(L_WR), .Z(\L_Out[18]1 ) );
    VMW_BUFIZ U89 ( .A(n418), .E(P_WR), .Z(\P_Out[30]1 ) );
    VMW_BUFIZ U92 ( .A(P_In[30]), .E(L_WR), .Z(\L_Out[30]1 ) );
    VMW_BUFIZ U145 ( .A(n445), .E(P_WR), .Z(\P_Out[21]1 ) );
    VMW_BUFIZ U162 ( .A(P_In[16]), .E(L_WR), .Z(\L_Out[16]1 ) );
    VMW_BUFIZ U117 ( .A(n430), .E(P_WR), .Z(\P_Out[0]1 ) );
    VMW_AO22 U58 ( .A(R_In[22]), .B(n417), .C(L_In[22]), .D(L_WR), .Z(n423) );
    VMW_BUFIZ U130 ( .A(P_In[6]), .E(L_WR), .Z(\L_Out[6]1 ) );
    VMW_BUFIZ U138 ( .A(n442), .E(P_WR), .Z(\P_Out[19]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_3 gt_47 ( .A(P_In), .B(L_In), .LEQ(n454), 
        .TC(n454), .LT_LE(n90) );
    VMW_BUFIZ U156 ( .A(P_In[2]), .E(R_WR), .Z(\R_Out[2]1 ) );
    VMW_BUFIZ U171 ( .A(P_In[0]), .E(R_WR), .Z(\R_Out[0]1 ) );
    VMW_PULLDOWN U38 ( .Z(n453) );
    VMW_AO22 U43 ( .A(R_In[7]), .B(n417), .C(L_In[7]), .D(L_WR), .Z(n447) );
    VMW_AO22 U64 ( .A(R_In[17]), .B(n417), .C(L_In[17]), .D(L_WR), .Z(n421) );
    VMW_BUFIZ U81 ( .A(P_In[1]), .E(R_WR), .Z(\R_Out[1]1 ) );
    BHeap_Node_WIDTH32_DW01_cmp2_32_0 gte_47 ( .A(R_In), .B(L_In), .LEQ(n450), 
        .TC(n451), .LT_LE(n92) );
    VMW_BUFIZ U104 ( .A(P_In[1]), .E(L_WR), .Z(\L_Out[1]1 ) );
    VMW_AO22 U51 ( .A(R_In[29]), .B(n417), .C(L_In[29]), .D(L_WR), .Z(n422) );
    VMW_BUFIZ U76 ( .A(P_In[22]), .E(L_WR), .Z(\L_Out[22]1 ) );
    VMW_BUFIZ U116 ( .A(P_In[19]), .E(R_WR), .Z(\R_Out[19]1 ) );
    VMW_BUFIZ U123 ( .A(P_In[7]), .E(L_WR), .Z(\L_Out[7]1 ) );
    VMW_BUFIZ U88 ( .A(P_In[3]), .E(R_WR), .Z(\R_Out[3]1 ) );
    VMW_BUFIZ U93 ( .A(P_In[29]), .E(L_WR), .Z(\L_Out[29]1 ) );
    VMW_BUFIZ U131 ( .A(n438), .E(P_WR), .Z(\P_Out[10]1 ) );
    VMW_BUFIZ U143 ( .A(P_In[30]), .E(R_WR), .Z(\R_Out[30]1 ) );
    VMW_BUFIZ U144 ( .A(P_In[29]), .E(R_WR), .Z(\R_Out[29]1 ) );
    VMW_BUFIZ U163 ( .A(P_In[6]), .E(R_WR), .Z(\R_Out[6]1 ) );
    VMW_BUFIZ U158 ( .A(P_In[21]), .E(L_WR), .Z(\L_Out[21]1 ) );
    VMW_BUFIZ U164 ( .A(P_In[27]), .E(L_WR), .Z(\L_Out[27]1 ) );
    VMW_AO22 U44 ( .A(R_In[6]), .B(n417), .C(L_In[6]), .D(L_WR), .Z(n420) );
    VMW_AO22 U56 ( .A(R_In[24]), .B(n417), .C(L_In[24]), .D(L_WR), .Z(n419) );
    VMW_BUFIZ U94 ( .A(P_In[20]), .E(L_WR), .Z(\L_Out[20]1 ) );
    VMW_BUFIZ U136 ( .A(n440), .E(P_WR), .Z(\P_Out[31] ) );
    VMW_AO22 U71 ( .A(R_In[10]), .B(n417), .C(L_In[10]), .D(L_WR), .Z(n438) );
    VMW_BUFIZ U111 ( .A(n428), .E(P_WR), .Z(\P_Out[11]1 ) );
    VMW_BUFIZ U124 ( .A(P_In[26]), .E(R_WR), .Z(\R_Out[26]1 ) );
    VMW_AO22 U63 ( .A(R_In[18]), .B(n417), .C(L_In[18]), .D(L_WR), .Z(n427) );
    VMW_BUFIZ U78 ( .A(P_In[8]), .E(R_WR), .Z(\R_Out[8]1 ) );
    VMW_BUFIZ U86 ( .A(P_In[7]), .E(R_WR), .Z(\R_Out[7]1 ) );
    VMW_BUFIZ U103 ( .A(P_In[8]), .E(L_WR), .Z(\L_Out[8]1 ) );
    VMW_BUFIZ U118 ( .A(P_In[27]), .E(R_WR), .Z(\R_Out[27]1 ) );
    VMW_BUFIZ U151 ( .A(P_In[4]), .E(L_WR), .Z(\L_Out[4]1 ) );
endmodule


module BHeap_CtrlReg_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, In, 
    Out, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR, In;
output Out, Enable;
    wire n77, Out70;
    assign Enable = Out;
    VMW_NOR2 U12 ( .A(n77), .B(Reset), .Z(Out70) );
    VMW_INV U13 ( .A(In), .Z(n77) );
    VMW_FD Out_reg ( .D(Out70), .CP(Clk), .Q(Out) );
endmodule


module BHeap_Control_CWIDTH2_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Go, Done );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR, Done;
output ScanEnable, Go;
    wire n379, \Count[0] , n362, n345, n339, n370, n357, n377, n350, n380, 
        n342, n365, n359, n356, n376, n351, \ScanReg[15] , \ScanReg[26] , 
        \ScanReg[2] , \ScanReg[18] , n358, n364, n343, n381, \ScanReg[11] , 
        \ScanReg[6] , \ScanReg[22] , n386, \ScanReg[20] , \ScanReg[13] , 
        \ScanReg[4] , n363, n344, n378, \ScanReg[29] , \ScanReg[30] , 
        \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , n371, \ScanReg[9] , n338, 
        \ScanReg[16] , \ScanReg[25] , Go259, \ScanReg[1] , \ScanReg[8] , n361, 
        n346, \ScanReg[7] , n384, \ScanReg[5] , n373, \ScanReg[21] , 
        \ScanReg[12] , n354, n368, \ScanReg[28] , \ScanReg[31] , \ScanReg[19] , 
        n348, n374, n353, \ScanReg[10] , \ScanReg[23] , n383, n341, n366, 
        \ScanReg[14] , \ScanReg[27] , \ScanReg[3] , n375, n352, n349, n360, 
        n340, n367, n382, n385, n347, n369, \Count[1] , n372, n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U68 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_AND2 U73 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_NOR2 U96 ( .A(n341), .B(Reset), .Z(n385) );
    VMW_AND2 U113 ( .A(\ScanReg[28] ), .B(n342), .Z(n367) );
    VMW_XNOR2 U134 ( .A(n350), .B(\Count[1] ), .Z(n349) );
    VMW_FD \Count_reg[0]  ( .D(n386), .CP(Clk), .Q(\Count[0] ) );
    VMW_AND2 U108 ( .A(\ScanReg[20] ), .B(n342), .Z(n372) );
    VMW_MUX2I U141 ( .A(n349), .B(DataIn[1]), .S(n351), .Z(n341) );
    VMW_BUFIZ U166 ( .A(n374), .E(n357), .Z(\arr[24] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U66 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U84 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_BUFIZ U148 ( .A(n355), .E(n357), .Z(\arr[10] ) );
    VMW_BUFIZ U153 ( .A(n361), .E(n357), .Z(\arr[25] ) );
    VMW_BUFIZ U174 ( .A(n382), .E(n357), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U101 ( .A(\ScanReg[15] ), .B(n342), .Z(n379) );
    VMW_AND2 U106 ( .A(\ScanReg[24] ), .B(n342), .Z(n374) );
    VMW_AND2 U121 ( .A(\ScanReg[27] ), .B(n342), .Z(n359) );
    VMW_AO21 U126 ( .A(RD), .B(ScanEnable), .C(n343), .Z(n357) );
    VMW_AND2 U74 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U83 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_BUFIZ U168 ( .A(n376), .E(n357), .Z(\arr[7] ) );
    VMW_AND2 U91 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AND2 U98 ( .A(\ScanReg[11] ), .B(n342), .Z(n382) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_XNOR2 U128 ( .A(Addr[0]), .B(Id), .Z(n343) );
    VMW_BUFIZ U154 ( .A(n362), .E(n357), .Z(\arr[16] ) );
    VMW_BUFIZ U173 ( .A(n381), .E(n357), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n353), .E(n357), .Z(\arr[0] ) );
    VMW_BUFIZ U161 ( .A(n369), .E(n357), .Z(\arr[13] ) );
    VMW_AND2 U114 ( .A(\ScanReg[21] ), .B(n342), .Z(n366) );
    VMW_AO22 U133 ( .A(\ScanReg[0] ), .B(n342), .C(\Count[0] ), .D(n343), .Z(
        n353) );
    VMW_AND2 U99 ( .A(\ScanReg[22] ), .B(n342), .Z(n381) );
    VMW_BUFIZ U155 ( .A(n363), .E(n357), .Z(\arr[6] ) );
    VMW_BUFIZ U172 ( .A(n380), .E(n357), .Z(\arr[18] ) );
    VMW_AND2 U67 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U82 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_BUFIZ U169 ( .A(n377), .E(n357), .Z(\arr[5] ) );
    VMW_AND2 U107 ( .A(\ScanReg[3] ), .B(n342), .Z(n373) );
    VMW_AND2 U120 ( .A(\ScanReg[14] ), .B(n342), .Z(n360) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_AND2 U69 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U75 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U115 ( .A(\ScanReg[31] ), .B(n342), .Z(n365) );
    VMW_AO22 U132 ( .A(\ScanReg[1] ), .B(n342), .C(\Count[1] ), .D(n343), .Z(
        n383) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U90 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U109 ( .A(\ScanReg[29] ), .B(n342), .Z(n371) );
    VMW_OAI21 U129 ( .A(RD), .B(WR), .C(n345), .Z(n344) );
    VMW_BUFIZ U147 ( .A(n354), .E(n357), .Z(\arr[23] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n368), .E(n357), .Z(\arr[2] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U97 ( .A(\ScanReg[8] ), .B(n342), .Z(n384) );
    VMW_MUX2I U140 ( .A(n348), .B(DataIn[1]), .S(n351), .Z(n338) );
    VMW_BUFIZ U167 ( .A(n375), .E(n357), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD Go_reg ( .D(Go259), .CP(Clk), .Q(Go) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AND2 U85 ( .A(WR), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AND2 U100 ( .A(\ScanReg[18] ), .B(n342), .Z(n380) );
    VMW_AND2 U112 ( .A(\ScanReg[2] ), .B(n342), .Z(n368) );
    VMW_AND2 U135 ( .A(WR), .B(n343), .Z(n351) );
    VMW_AND2 U127 ( .A(\ScanReg[19] ), .B(n342), .Z(n352) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n356), .E(n357), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n360), .E(n357), .Z(\arr[14] ) );
    VMW_BUFIZ U175 ( .A(n383), .E(n357), .Z(\arr[1] ) );
    VMW_AOI21 U62 ( .A(n338), .B(n339), .C(Reset), .Z(Go259) );
    VMW_AND2 U70 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_OR3 U137 ( .A(n351), .B(Done), .C(n347), .Z(n340) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AOI21 U95 ( .A(n339), .B(n340), .C(Reset), .Z(n386) );
    VMW_AND2 U110 ( .A(\ScanReg[30] ), .B(n342), .Z(n370) );
    VMW_BUFIZ U159 ( .A(n367), .E(n357), .Z(\arr[28] ) );
    VMW_AND2 U119 ( .A(\ScanReg[25] ), .B(n342), .Z(n361) );
    VMW_INV U142 ( .A(n343), .Z(n342) );
    VMW_BUFIZ U165 ( .A(n373), .E(n357), .Z(\arr[3] ) );
    VMW_AND2 U87 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_BUFIZ U150 ( .A(n358), .E(n357), .Z(\arr[4] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AND2 U125 ( .A(\ScanReg[23] ), .B(n342), .Z(n354) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U63 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U64 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U65 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U102 ( .A(\ScanReg[26] ), .B(n342), .Z(n378) );
    VMW_AND2 U105 ( .A(\ScanReg[17] ), .B(n342), .Z(n375) );
    VMW_AND2 U77 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U80 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U122 ( .A(\ScanReg[4] ), .B(n342), .Z(n358) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_AND2 U89 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_MUX2I U139 ( .A(n346), .B(DataIn[0]), .S(n351), .Z(n339) );
    VMW_BUFIZ U157 ( .A(n365), .E(n357), .Z(\arr[31] ) );
    VMW_BUFIZ U170 ( .A(n378), .E(n357), .Z(\arr[26] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AND2 U92 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U145 ( .A(n352), .E(n357), .Z(\arr[19] ) );
    VMW_BUFIZ U162 ( .A(n370), .E(n357), .Z(\arr[30] ) );
    VMW_AND2 U117 ( .A(\ScanReg[6] ), .B(n342), .Z(n363) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AND2 U81 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_AND2 U130 ( .A(Done), .B(n347), .Z(n346) );
    VMW_XNOR2 U138 ( .A(Addr[0]), .B(ScanId), .Z(n345) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_BUFIZ U156 ( .A(n364), .E(n357), .Z(\arr[12] ) );
    VMW_BUFIZ U171 ( .A(n379), .E(n357), .Z(\arr[15] ) );
    VMW_AND2 U104 ( .A(\ScanReg[7] ), .B(n342), .Z(n376) );
    VMW_AND2 U71 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U76 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U116 ( .A(\ScanReg[12] ), .B(n342), .Z(n364) );
    VMW_AND2 U123 ( .A(\ScanReg[9] ), .B(n342), .Z(n356) );
    VMW_AND2 U88 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AND2 U93 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_AND2 U131 ( .A(\Count[1] ), .B(Done), .Z(n348) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_INV U143 ( .A(\Count[0] ), .Z(n347) );
    VMW_INV U144 ( .A(n344), .Z(ScanEnable) );
    VMW_BUFIZ U163 ( .A(n371), .E(n357), .Z(\arr[29] ) );
    VMW_BUFIZ U158 ( .A(n366), .E(n357), .Z(\arr[21] ) );
    VMW_BUFIZ U164 ( .A(n372), .E(n357), .Z(\arr[20] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_NAND2 U136 ( .A(n347), .B(Done), .Z(n350) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U111 ( .A(\ScanReg[13] ), .B(n342), .Z(n369) );
    VMW_AND2 U124 ( .A(\ScanReg[10] ), .B(n342), .Z(n355) );
    VMW_AND2 U78 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AND2 U86 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U103 ( .A(\ScanReg[5] ), .B(n342), .Z(n377) );
    VMW_FD \Count_reg[1]  ( .D(n385), .CP(Clk), .Q(\Count[1] ) );
    VMW_AND2 U118 ( .A(\ScanReg[16] ), .B(n342), .Z(n362) );
    VMW_BUFIZ U151 ( .A(n359), .E(n357), .Z(\arr[27] ) );
    VMW_BUFIZ U176 ( .A(n384), .E(n357), .Z(\arr[8] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \ScanLink0[13] , \wRegInTop_1_0[15] , \wRegInTop_1_0[26] , 
        \ScanLink1[19] , \ScanLink0[20] , \wRegOut_1_0[0] , \wRegOut_0_0[6] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[20] , 
        \wRegOut_1_0[9] , \wRegInBot_0_0[13] , \ScanLink1[23] , 
        \ScanLink1[10] , \ScanLink1[7] , \ScanLink2[4] , \wRegInTop_1_1[16] , 
        \wRegInTop_1_1[25] , \ScanLink0[30] , \ScanLink0[29] , 
        \wRegInTop_1_0[4] , \ScanLink0[17] , \ScanEnable[0] , \wRegOut_1_0[4] , 
        \ScanLink2[9] , \wRegInTop_1_1[31] , \wRegInTop_1_1[28] , 
        \wRegInTop_1_0[11] , \wRegInTop_1_0[9] , \ScanLink0[24] , 
        \wRegInTop_1_0[22] , \wRegOut_0_0[2] , \wRegInTop_1_0[18] , 
        \wRegInTop_1_0[0] , \ScanLink1[27] , \ScanLink1[14] , \ScanLink1[3] , 
        \ScanLink2[0] , \wRegInTop_1_1[12] , \wRegInTop_1_1[21] , 
        \wRegInBot_0_0[26] , \wRegInBot_0_0[24] , \wRegInBot_0_0[17] , 
        \ScanLink1[25] , \ScanLink1[16] , \ScanLink1[1] , \ScanLink2[2] , 
        \wRegInTop_1_1[10] , \wRegInTop_1_1[23] , \wRegInBot_0_0[15] , 
        \wRegInTop_1_0[30] , \wRegInTop_1_0[29] , \wRegOut_0_0[9] , 
        \wRegOut_0_0[0] , \wRegInTop_1_0[2] , \wCtrlOut_1[0] , \ScanLink0[15] , 
        \wRegInTop_1_0[13] , \wRegInTop_1_0[20] , \ScanLink0[26] , 
        \wRegOut_0_0[4] , \ScanLink1[8] , \wRegOut_1_0[6] , 
        \wRegInTop_1_1[19] , \ScanLink0[18] , \wRegInTop_1_0[6] , 
        \wRegInBot_0_0[22] , \wRegInBot_0_0[18] , \wRegInBot_0_0[11] , 
        \ScanLink1[31] , \ScanLink1[28] , \ScanLink1[21] , \ScanLink1[12] , 
        \ScanLink1[5] , \ScanLink2[6] , \wRegInTop_1_1[14] , 
        \wRegInTop_1_1[27] , \wRegOut_1_0[2] , \ScanLink0[11] , 
        \wRegInTop_1_0[17] , \ScanLink0[22] , \wRegInTop_1_0[24] , 
        \ScanLink2[24] , \ScanLink2[17] , \wRegOut_1_1[22] , \wRegOut_1_1[11] , 
        \wRegInTop_1_1[2] , \ScanLink0[1] , \wRegOut_1_0[31] , 
        \wRegOut_1_0[28] , \ScanLink3[2] , \wRegOut_0_0[16] , 
        \wRegOut_0_0[25] , \wRegInBot_0_0[2] , \ScanLink0[8] , 
        \wRegOut_1_0[21] , \wRegOut_1_0[12] , \wRegOut_1_1[6] , 
        \ScanLink3[27] , \wRegOut_0_0[12] , \wRegOut_1_1[18] , \ScanLink3[14] , 
        \wCtrlOut_0[0] , \ScanLink3[19] , \wRegOut_0_0[21] , \ScanLink0[5] , 
        \ScanLink3[6] , \wRegOut_0_0[31] , \wRegOut_0_0[28] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[20] , \wRegOut_1_1[26] , \wRegOut_1_1[15] , 
        \wRegInTop_1_1[6] , \ScanLink2[13] , \ScanLink3[23] , \ScanLink3[10] , 
        \wRegInBot_0_0[6] , \wRegOut_1_1[2] , \wRegOut_1_0[16] , 
        \wRegOut_1_0[25] , \wRegOut_1_1[0] , \ScanLink3[21] , 
        \wRegOut_0_0[19] , \wRegInBot_0_0[4] , \ScanLink3[12] , 
        \wRegOut_1_0[27] , \wRegOut_1_0[14] , \ScanLink2[18] , 
        \wRegOut_1_1[17] , \wRegInTop_1_1[4] , \ScanLink2[22] , 
        \wRegOut_1_1[24] , \wEnable_0[0] , \ScanLink2[11] , \wRegOut_0_0[10] , 
        \wRegOut_1_1[9] , \wRegOut_0_0[23] , \ScanLink3[31] , \ScanLink3[28] , 
        \wRegInBot_0_0[0] , \ScanLink0[7] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[10] , \wRegOut_1_1[30] , \ScanLink3[4] , 
        \wRegOut_1_1[29] , \wRegInTop_1_1[9] , \ScanLink3[9] , \ScanLink3[25] , 
        \ScanLink3[16] , \wRegOut_1_1[4] , \ScanLink0[3] , \wRegOut_1_0[19] , 
        \ScanLink3[0] , \wRegOut_0_0[14] , \wRegOut_0_0[27] , 
        \wRegInBot_0_0[9] , \ScanLink2[26] , \ScanLink2[15] , 
        \wRegOut_1_1[20] , \wRegOut_1_1[13] , \wRegInTop_1_1[0] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[11] , \wRegOut_1_1[31] , 
        \wRegOut_1_1[28] , \wRegInTop_1_1[8] , \ScanLink3[8] , 
        \wRegOut_1_1[5] , \ScanLink3[24] , \ScanLink3[17] , \wRegInBot_0_0[8] , 
        \wRegInBot_0_0[1] , \ScanLink0[2] , \wRegOut_1_0[18] , \ScanLink3[1] , 
        \wRegOut_0_0[15] , \wRegOut_0_0[26] , \ScanLink2[27] , \ScanLink2[14] , 
        \wRegOut_0_0[18] , \wRegInBot_0_0[5] , \wRegOut_1_1[21] , 
        \wRegOut_1_1[12] , \wRegInTop_1_1[1] , \ScanLink3[20] , 
        \wRegOut_1_0[26] , \wRegOut_1_0[15] , \wRegOut_1_1[1] , 
        \ScanLink3[13] , \ScanLink2[19] , \wRegOut_1_1[25] , \wRegOut_1_1[16] , 
        \wRegInTop_1_1[5] , \wRegOut_0_0[11] , \ScanLink2[23] , 
        \ScanLink2[10] , \wRegOut_0_0[22] , \wRegOut_1_1[8] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink0[6] , \ScanLink3[5] , \wRegOut_0_0[13] , 
        \ScanLink3[18] , \wRegOut_0_0[20] , \ScanLink0[4] , \wRegOut_1_1[27] , 
        \wRegOut_1_1[14] , \wRegInTop_1_1[7] , \ScanLink3[7] , 
        \wRegEnTop_1_1[0] , \ScanLink2[31] , \ScanLink2[21] , \ScanLink2[12] , 
        \ScanLink2[28] , \wRegOut_0_0[30] , \wRegInBot_0_0[7] , 
        \wRegOut_0_0[29] , \wRegOut_1_1[3] , \ScanLink3[22] , \ScanLink3[11] , 
        \wRegEnBot_0_0[0] , \wRegOut_1_0[24] , \wRegOut_1_0[17] , 
        \ScanLink2[25] , \ScanLink2[16] , \wRegOut_0_0[17] , \ScanLink0[0] , 
        \wRegOut_1_0[30] , \wRegOut_1_1[23] , \wRegOut_1_1[10] , 
        \wRegInTop_1_1[3] , \wRegOut_1_0[29] , \ScanLink3[3] , 
        \wRegOut_0_0[24] , \ScanLink0[9] , \wRegOut_1_0[13] , 
        \wRegOut_1_0[20] , \ScanLink3[26] , \wRegOut_0_0[5] , 
        \wRegInBot_0_0[3] , \wRegOut_1_1[7] , \ScanLink3[15] , \ScanLink0[19] , 
        \wRegOut_1_1[19] , \wRegEnTop_1_0[0] , \wRegInTop_1_0[7] , 
        \wRegInBot_0_0[23] , \ScanLink1[20] , \ScanLink1[13] , \ScanLink2[7] , 
        \ScanLink1[4] , \wRegInTop_1_1[15] , \wRegInTop_1_1[26] , 
        \wRegInBot_0_0[19] , \wRegInBot_0_0[10] , \wRegOut_1_0[3] , 
        \ScanLink1[30] , \ScanLink1[29] , \wRegInTop_1_0[16] , \ScanLink0[10] , 
        \wRegInBot_0_0[27] , \ScanLink0[23] , \wRegInTop_1_0[25] , 
        \wRegInBot_0_0[14] , \ScanLink1[24] , \ScanLink1[17] , \ScanLink1[0] , 
        \wRegInTop_1_1[11] , \ScanLink2[3] , \wRegInTop_1_1[22] , 
        \wRegOut_0_0[1] , \wRegInTop_1_0[31] , \wRegInTop_1_0[28] , 
        \wRegInTop_1_0[3] , \ScanLink0[14] , \ScanLink0[27] , 
        \wRegInTop_1_0[12] , \wRegInTop_1_0[21] , \wRegOut_0_0[8] , 
        \ScanLink1[9] , \wRegInTop_1_1[18] , \wRegOut_1_0[7] , \ScanLink2[8] , 
        \wRegInTop_1_1[30] , \wRegInTop_1_1[29] , \wRegOut_1_0[5] , 
        \wRegInTop_1_0[10] , \ScanLink0[16] , \wRegInTop_1_0[8] , 
        \wRegOut_0_0[3] , \ScanLink0[25] , \wRegInTop_1_0[23] , 
        \wRegInBot_0_0[25] , \wRegInTop_1_0[19] , \wRegInTop_1_0[1] , 
        \wRegInBot_0_0[16] , \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , 
        \ScanLink1[2] , \wRegInTop_1_1[13] , \ScanLink0[12] , 
        \wRegInTop_1_1[20] , \ScanLink0[21] , \wRegInTop_1_0[14] , 
        \wRegInTop_1_0[27] , \wRegInBot_0_0[31] , \wRegInBot_0_0[28] , 
        \wRegOut_1_0[1] , \wRegOut_0_0[7] , \wRegInBot_0_0[21] , 
        \ScanLink1[22] , \ScanLink1[18] , \ScanLink1[11] , \ScanLink1[6] , 
        \wRegOut_1_0[8] , \wRegInTop_1_1[17] , \ScanLink2[5] , 
        \wRegInTop_1_1[24] , \wRegInBot_0_0[12] , \ScanLink0[31] , 
        \ScanLink0[28] , \wRegInTop_1_0[5] ;
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_0_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_0_0[31] , \wRegOut_0_0[30] , \wRegOut_0_0[29] , 
        \wRegOut_0_0[28] , \wRegOut_0_0[27] , \wRegOut_0_0[26] , 
        \wRegOut_0_0[25] , \wRegOut_0_0[24] , \wRegOut_0_0[23] , 
        \wRegOut_0_0[22] , \wRegOut_0_0[21] , \wRegOut_0_0[20] , 
        \wRegOut_0_0[19] , \wRegOut_0_0[18] , \wRegOut_0_0[17] , 
        \wRegOut_0_0[16] , \wRegOut_0_0[15] , \wRegOut_0_0[14] , 
        \wRegOut_0_0[13] , \wRegOut_0_0[12] , \wRegOut_0_0[11] , 
        \wRegOut_0_0[10] , \wRegOut_0_0[9] , \wRegOut_0_0[8] , 
        \wRegOut_0_0[7] , \wRegOut_0_0[6] , \wRegOut_0_0[5] , \wRegOut_0_0[4] , 
        \wRegOut_0_0[3] , \wRegOut_0_0[2] , \wRegOut_0_0[1] , \wRegOut_0_0[0] 
        }), .Enable1(1'b0), .Enable2(\wRegEnBot_0_0[0] ), .In1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .In2({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .Enable1(\wRegEnTop_1_0[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_1_0[31] , \wRegInTop_1_0[30] , \wRegInTop_1_0[29] , 
        \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , \wRegInTop_1_0[26] , 
        \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , \wRegInTop_1_0[23] , 
        \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , \wRegInTop_1_0[20] , 
        \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , \wRegInTop_1_0[17] , 
        \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , \wRegInTop_1_0[14] , 
        \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , \wRegInTop_1_0[11] , 
        \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , \wRegInTop_1_0[8] , 
        \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , \wRegInTop_1_0[5] , 
        \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , \wRegInTop_1_0[2] , 
        \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Reg_WIDTH32_IDWIDTH1_SCAN1 BHR_1_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Out({\wRegOut_1_1[31] , \wRegOut_1_1[30] , \wRegOut_1_1[29] , 
        \wRegOut_1_1[28] , \wRegOut_1_1[27] , \wRegOut_1_1[26] , 
        \wRegOut_1_1[25] , \wRegOut_1_1[24] , \wRegOut_1_1[23] , 
        \wRegOut_1_1[22] , \wRegOut_1_1[21] , \wRegOut_1_1[20] , 
        \wRegOut_1_1[19] , \wRegOut_1_1[18] , \wRegOut_1_1[17] , 
        \wRegOut_1_1[16] , \wRegOut_1_1[15] , \wRegOut_1_1[14] , 
        \wRegOut_1_1[13] , \wRegOut_1_1[12] , \wRegOut_1_1[11] , 
        \wRegOut_1_1[10] , \wRegOut_1_1[9] , \wRegOut_1_1[8] , 
        \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , \wRegOut_1_1[4] , 
        \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , \wRegOut_1_1[0] 
        }), .Enable1(\wRegEnTop_1_1[0] ), .Enable2(1'b0), .In1({
        \wRegInTop_1_1[31] , \wRegInTop_1_1[30] , \wRegInTop_1_1[29] , 
        \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , \wRegInTop_1_1[26] , 
        \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , \wRegInTop_1_1[23] , 
        \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , \wRegInTop_1_1[20] , 
        \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , \wRegInTop_1_1[17] , 
        \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , \wRegInTop_1_1[14] , 
        \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , \wRegInTop_1_1[11] , 
        \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , \wRegInTop_1_1[8] , 
        \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , \wRegInTop_1_1[5] , 
        \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , \wRegInTop_1_1[2] , 
        \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }), .In2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
    BHeap_Node_WIDTH32 BHN_0_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(
        \wEnable_0[0] ), .P_WR(\wRegEnBot_0_0[0] ), .P_In({\wRegOut_0_0[31] , 
        \wRegOut_0_0[30] , \wRegOut_0_0[29] , \wRegOut_0_0[28] , 
        \wRegOut_0_0[27] , \wRegOut_0_0[26] , \wRegOut_0_0[25] , 
        \wRegOut_0_0[24] , \wRegOut_0_0[23] , \wRegOut_0_0[22] , 
        \wRegOut_0_0[21] , \wRegOut_0_0[20] , \wRegOut_0_0[19] , 
        \wRegOut_0_0[18] , \wRegOut_0_0[17] , \wRegOut_0_0[16] , 
        \wRegOut_0_0[15] , \wRegOut_0_0[14] , \wRegOut_0_0[13] , 
        \wRegOut_0_0[12] , \wRegOut_0_0[11] , \wRegOut_0_0[10] , 
        \wRegOut_0_0[9] , \wRegOut_0_0[8] , \wRegOut_0_0[7] , \wRegOut_0_0[6] , 
        \wRegOut_0_0[5] , \wRegOut_0_0[4] , \wRegOut_0_0[3] , \wRegOut_0_0[2] , 
        \wRegOut_0_0[1] , \wRegOut_0_0[0] }), .P_Out({\wRegInBot_0_0[31] , 
        \wRegInBot_0_0[30] , \wRegInBot_0_0[29] , \wRegInBot_0_0[28] , 
        \wRegInBot_0_0[27] , \wRegInBot_0_0[26] , \wRegInBot_0_0[25] , 
        \wRegInBot_0_0[24] , \wRegInBot_0_0[23] , \wRegInBot_0_0[22] , 
        \wRegInBot_0_0[21] , \wRegInBot_0_0[20] , \wRegInBot_0_0[19] , 
        \wRegInBot_0_0[18] , \wRegInBot_0_0[17] , \wRegInBot_0_0[16] , 
        \wRegInBot_0_0[15] , \wRegInBot_0_0[14] , \wRegInBot_0_0[13] , 
        \wRegInBot_0_0[12] , \wRegInBot_0_0[11] , \wRegInBot_0_0[10] , 
        \wRegInBot_0_0[9] , \wRegInBot_0_0[8] , \wRegInBot_0_0[7] , 
        \wRegInBot_0_0[6] , \wRegInBot_0_0[5] , \wRegInBot_0_0[4] , 
        \wRegInBot_0_0[3] , \wRegInBot_0_0[2] , \wRegInBot_0_0[1] , 
        \wRegInBot_0_0[0] }), .L_WR(\wRegEnTop_1_0[0] ), .L_In({
        \wRegOut_1_0[31] , \wRegOut_1_0[30] , \wRegOut_1_0[29] , 
        \wRegOut_1_0[28] , \wRegOut_1_0[27] , \wRegOut_1_0[26] , 
        \wRegOut_1_0[25] , \wRegOut_1_0[24] , \wRegOut_1_0[23] , 
        \wRegOut_1_0[22] , \wRegOut_1_0[21] , \wRegOut_1_0[20] , 
        \wRegOut_1_0[19] , \wRegOut_1_0[18] , \wRegOut_1_0[17] , 
        \wRegOut_1_0[16] , \wRegOut_1_0[15] , \wRegOut_1_0[14] , 
        \wRegOut_1_0[13] , \wRegOut_1_0[12] , \wRegOut_1_0[11] , 
        \wRegOut_1_0[10] , \wRegOut_1_0[9] , \wRegOut_1_0[8] , 
        \wRegOut_1_0[7] , \wRegOut_1_0[6] , \wRegOut_1_0[5] , \wRegOut_1_0[4] , 
        \wRegOut_1_0[3] , \wRegOut_1_0[2] , \wRegOut_1_0[1] , \wRegOut_1_0[0] 
        }), .L_Out({\wRegInTop_1_0[31] , \wRegInTop_1_0[30] , 
        \wRegInTop_1_0[29] , \wRegInTop_1_0[28] , \wRegInTop_1_0[27] , 
        \wRegInTop_1_0[26] , \wRegInTop_1_0[25] , \wRegInTop_1_0[24] , 
        \wRegInTop_1_0[23] , \wRegInTop_1_0[22] , \wRegInTop_1_0[21] , 
        \wRegInTop_1_0[20] , \wRegInTop_1_0[19] , \wRegInTop_1_0[18] , 
        \wRegInTop_1_0[17] , \wRegInTop_1_0[16] , \wRegInTop_1_0[15] , 
        \wRegInTop_1_0[14] , \wRegInTop_1_0[13] , \wRegInTop_1_0[12] , 
        \wRegInTop_1_0[11] , \wRegInTop_1_0[10] , \wRegInTop_1_0[9] , 
        \wRegInTop_1_0[8] , \wRegInTop_1_0[7] , \wRegInTop_1_0[6] , 
        \wRegInTop_1_0[5] , \wRegInTop_1_0[4] , \wRegInTop_1_0[3] , 
        \wRegInTop_1_0[2] , \wRegInTop_1_0[1] , \wRegInTop_1_0[0] }), .R_WR(
        \wRegEnTop_1_1[0] ), .R_In({\wRegOut_1_1[31] , \wRegOut_1_1[30] , 
        \wRegOut_1_1[29] , \wRegOut_1_1[28] , \wRegOut_1_1[27] , 
        \wRegOut_1_1[26] , \wRegOut_1_1[25] , \wRegOut_1_1[24] , 
        \wRegOut_1_1[23] , \wRegOut_1_1[22] , \wRegOut_1_1[21] , 
        \wRegOut_1_1[20] , \wRegOut_1_1[19] , \wRegOut_1_1[18] , 
        \wRegOut_1_1[17] , \wRegOut_1_1[16] , \wRegOut_1_1[15] , 
        \wRegOut_1_1[14] , \wRegOut_1_1[13] , \wRegOut_1_1[12] , 
        \wRegOut_1_1[11] , \wRegOut_1_1[10] , \wRegOut_1_1[9] , 
        \wRegOut_1_1[8] , \wRegOut_1_1[7] , \wRegOut_1_1[6] , \wRegOut_1_1[5] , 
        \wRegOut_1_1[4] , \wRegOut_1_1[3] , \wRegOut_1_1[2] , \wRegOut_1_1[1] , 
        \wRegOut_1_1[0] }), .R_Out({\wRegInTop_1_1[31] , \wRegInTop_1_1[30] , 
        \wRegInTop_1_1[29] , \wRegInTop_1_1[28] , \wRegInTop_1_1[27] , 
        \wRegInTop_1_1[26] , \wRegInTop_1_1[25] , \wRegInTop_1_1[24] , 
        \wRegInTop_1_1[23] , \wRegInTop_1_1[22] , \wRegInTop_1_1[21] , 
        \wRegInTop_1_1[20] , \wRegInTop_1_1[19] , \wRegInTop_1_1[18] , 
        \wRegInTop_1_1[17] , \wRegInTop_1_1[16] , \wRegInTop_1_1[15] , 
        \wRegInTop_1_1[14] , \wRegInTop_1_1[13] , \wRegInTop_1_1[12] , 
        \wRegInTop_1_1[11] , \wRegInTop_1_1[10] , \wRegInTop_1_1[9] , 
        \wRegInTop_1_1[8] , \wRegInTop_1_1[7] , \wRegInTop_1_1[6] , 
        \wRegInTop_1_1[5] , \wRegInTop_1_1[4] , \wRegInTop_1_1[3] , 
        \wRegInTop_1_1[2] , \wRegInTop_1_1[1] , \wRegInTop_1_1[0] }) );
    BHeap_CtrlReg_WIDTH32 BHCR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), 
        .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(\wCtrlOut_1[0] ), 
        .Out(\wCtrlOut_0[0] ), .Enable(\wEnable_0[0] ) );
    BHeap_Control_CWIDTH2_IDWIDTH1_WIDTH32_SCAN1 BHC ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink0[31] , \ScanLink0[30] , \ScanLink0[29] , 
        \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , \ScanLink0[25] , 
        \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , \ScanLink0[21] , 
        \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , \ScanLink0[17] , 
        \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , \ScanLink0[13] , 
        \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , \ScanLink0[9] , 
        \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , \ScanLink0[5] , 
        \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , \ScanLink0[1] , 
        \ScanLink0[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b0), .Id(1'b1), .Go(\wCtrlOut_1[0] ), .Done(\wCtrlOut_0[0] )
         );
endmodule

