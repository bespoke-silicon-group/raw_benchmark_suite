
module BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, 
        n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, 
        n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, n113, 
        n94, n23, n103, n16, n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, 
        n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, 
        n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, 
        n87, n17, n30, n79, n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(B[31]), .Z(n15) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n66), .C(n62), .D(n57), .Z(n65) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U34 ( .A(B[16]), .B(n64), .Z(n67) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n75), .D(n70), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(B[15]), .Z(n66) );
    VMW_INV U101 ( .A(A[6]), .Z(n32) );
    VMW_INV U66 ( .A(B[7]), .Z(n41) );
    VMW_INV U83 ( .A(A[15]), .Z(n69) );
    VMW_INV U98 ( .A(B[13]), .Z(n60) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n69), .C(n67), .D(n65), .Z(n68) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(B[11]), .Z(n54) );
    VMW_INV U74 ( .A(A[3]), .Z(n30) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U40 ( .A(n78), .B(B[20]), .Z(n77) );
    VMW_INV U82 ( .A(B[29]), .Z(n110) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n44) );
    VMW_INV U75 ( .A(B[3]), .Z(n27) );
    VMW_INV U90 ( .A(A[14]), .Z(n58) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n73) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n64) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n107), .D(n102), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_INV U85 ( .A(A[4]), .Z(n25) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_NAND2 U32 ( .A(n64), .B(B[16]), .Z(n63) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n76), .C(n74), .D(n72), .Z(n75) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n76) );
    VMW_INV U95 ( .A(A[1]), .Z(n21) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_INV U79 ( .A(B[19]), .Z(n80) );
    VMW_INV U87 ( .A(A[8]), .Z(n39) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n77), .Z(n85) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n52) );
    VMW_INV U102 ( .A(A[2]), .Z(n18) );
    VMW_INV U80 ( .A(A[10]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n73), .C(n68), .D(n63), .Z(n72) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[18]), .Z(n71) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[25]), .Z(n101) );
    VMW_INV U92 ( .A(A[28]), .Z(n103) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n71), .B(B[18]), .Z(n70) );
    VMW_INV U81 ( .A(B[9]), .Z(n48) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n78), .C(n81), .D(n79), .Z(n82) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(B[25]), .Z(n98) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_INV U88 ( .A(B[21]), .Z(n86) );
    VMW_INV U93 ( .A(A[5]), .Z(n37) );
    VMW_OR2 U38 ( .A(B[18]), .B(n71), .Z(n74) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(B[5]), .Z(n34) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[24]), .Z(n90) );
    VMW_INV U103 ( .A(A[0]), .Z(n20) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_INV U78 ( .A(A[20]), .Z(n78) );
endmodule


module BubbleSort_Node_WIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, 
    AIn, BIn, HiOut, LoOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
output [31:0] LoOut;
input  [31:0] AIn;
input  [31:0] BIn;
output [31:0] HiOut;
input  Clk, Reset, RD, WR;
    wire n159, a58;
    VMW_PULLDOWN U21 ( .Z(n159) );
    VMW_MUX2 U54 ( .A(BIn[9]), .B(AIn[9]), .S(a58), .Z(HiOut[9]) );
    VMW_MUX2 U73 ( .A(BIn[20]), .B(AIn[20]), .S(a58), .Z(HiOut[20]) );
    VMW_MUX2 U22 ( .A(AIn[9]), .B(BIn[9]), .S(a58), .Z(LoOut[9]) );
    VMW_MUX2 U26 ( .A(AIn[5]), .B(BIn[5]), .S(a58), .Z(LoOut[5]) );
    VMW_MUX2 U28 ( .A(AIn[3]), .B(BIn[3]), .S(a58), .Z(LoOut[3]) );
    VMW_MUX2 U33 ( .A(AIn[28]), .B(BIn[28]), .S(a58), .Z(LoOut[28]) );
    VMW_MUX2 U68 ( .A(BIn[25]), .B(AIn[25]), .S(a58), .Z(HiOut[25]) );
    VMW_MUX2 U34 ( .A(AIn[27]), .B(BIn[27]), .S(a58), .Z(LoOut[27]) );
    VMW_MUX2 U41 ( .A(AIn[20]), .B(BIn[20]), .S(a58), .Z(LoOut[20]) );
    VMW_MUX2 U46 ( .A(AIn[16]), .B(BIn[16]), .S(a58), .Z(LoOut[16]) );
    VMW_MUX2 U61 ( .A(BIn[31]), .B(AIn[31]), .S(a58), .Z(HiOut[31]) );
    VMW_MUX2 U84 ( .A(BIn[10]), .B(AIn[10]), .S(a58), .Z(HiOut[10]) );
    VMW_MUX2 U66 ( .A(BIn[27]), .B(AIn[27]), .S(a58), .Z(HiOut[27]) );
    VMW_MUX2 U83 ( .A(BIn[11]), .B(AIn[11]), .S(a58), .Z(HiOut[11]) );
    VMW_MUX2 U48 ( .A(AIn[14]), .B(BIn[14]), .S(a58), .Z(LoOut[14]) );
    VMW_MUX2 U27 ( .A(AIn[4]), .B(BIn[4]), .S(a58), .Z(LoOut[4]) );
    VMW_MUX2 U35 ( .A(AIn[26]), .B(BIn[26]), .S(a58), .Z(LoOut[26]) );
    VMW_MUX2 U53 ( .A(AIn[0]), .B(BIn[0]), .S(a58), .Z(LoOut[0]) );
    VMW_MUX2 U74 ( .A(BIn[1]), .B(AIn[1]), .S(a58), .Z(HiOut[1]) );
    VMW_MUX2 U40 ( .A(AIn[21]), .B(BIn[21]), .S(a58), .Z(LoOut[21]) );
    VMW_MUX2 U82 ( .A(BIn[12]), .B(AIn[12]), .S(a58), .Z(HiOut[12]) );
    VMW_MUX2 U52 ( .A(AIn[10]), .B(BIn[10]), .S(a58), .Z(LoOut[10]) );
    VMW_MUX2 U67 ( .A(BIn[26]), .B(AIn[26]), .S(a58), .Z(HiOut[26]) );
    VMW_MUX2 U75 ( .A(BIn[19]), .B(AIn[19]), .S(a58), .Z(HiOut[19]) );
    VMW_MUX2 U29 ( .A(AIn[31]), .B(BIn[31]), .S(a58), .Z(LoOut[31]) );
    VMW_MUX2 U47 ( .A(AIn[15]), .B(BIn[15]), .S(a58), .Z(LoOut[15]) );
    VMW_MUX2 U49 ( .A(AIn[13]), .B(BIn[13]), .S(a58), .Z(LoOut[13]) );
    VMW_MUX2 U55 ( .A(BIn[8]), .B(AIn[8]), .S(a58), .Z(HiOut[8]) );
    VMW_MUX2 U69 ( .A(BIn[24]), .B(AIn[24]), .S(a58), .Z(HiOut[24]) );
    VMW_MUX2 U72 ( .A(BIn[21]), .B(AIn[21]), .S(a58), .Z(HiOut[21]) );
    VMW_MUX2 U60 ( .A(BIn[3]), .B(AIn[3]), .S(a58), .Z(HiOut[3]) );
    VMW_MUX2 U32 ( .A(AIn[29]), .B(BIn[29]), .S(a58), .Z(LoOut[29]) );
    VMW_MUX2 U85 ( .A(BIn[0]), .B(AIn[0]), .S(a58), .Z(HiOut[0]) );
    VMW_MUX2 U39 ( .A(AIn[22]), .B(BIn[22]), .S(a58), .Z(LoOut[22]) );
    VMW_MUX2 U57 ( .A(BIn[6]), .B(AIn[6]), .S(a58), .Z(HiOut[6]) );
    VMW_MUX2 U70 ( .A(BIn[23]), .B(AIn[23]), .S(a58), .Z(HiOut[23]) );
    VMW_MUX2 U23 ( .A(AIn[8]), .B(BIn[8]), .S(a58), .Z(LoOut[8]) );
    VMW_MUX2 U24 ( .A(AIn[7]), .B(BIn[7]), .S(a58), .Z(LoOut[7]) );
    VMW_MUX2 U25 ( .A(AIn[6]), .B(BIn[6]), .S(a58), .Z(LoOut[6]) );
    VMW_MUX2 U30 ( .A(AIn[30]), .B(BIn[30]), .S(a58), .Z(LoOut[30]) );
    VMW_MUX2 U79 ( .A(BIn[15]), .B(AIn[15]), .S(a58), .Z(HiOut[15]) );
    BubbleSort_Node_WIDTH32_DW01_cmp2_32_0 gt_41 ( .A(BIn), .B(AIn), .LEQ(n159
        ), .TC(n159), .LT_LE(a58) );
    VMW_MUX2 U37 ( .A(AIn[24]), .B(BIn[24]), .S(a58), .Z(LoOut[24]) );
    VMW_MUX2 U42 ( .A(AIn[1]), .B(BIn[1]), .S(a58), .Z(LoOut[1]) );
    VMW_MUX2 U45 ( .A(AIn[17]), .B(BIn[17]), .S(a58), .Z(LoOut[17]) );
    VMW_MUX2 U62 ( .A(BIn[30]), .B(AIn[30]), .S(a58), .Z(HiOut[30]) );
    VMW_MUX2 U65 ( .A(BIn[28]), .B(AIn[28]), .S(a58), .Z(HiOut[28]) );
    VMW_MUX2 U80 ( .A(BIn[14]), .B(AIn[14]), .S(a58), .Z(HiOut[14]) );
    VMW_MUX2 U59 ( .A(BIn[4]), .B(AIn[4]), .S(a58), .Z(HiOut[4]) );
    VMW_MUX2 U36 ( .A(AIn[25]), .B(BIn[25]), .S(a58), .Z(LoOut[25]) );
    VMW_MUX2 U50 ( .A(AIn[12]), .B(BIn[12]), .S(a58), .Z(LoOut[12]) );
    VMW_MUX2 U77 ( .A(BIn[17]), .B(AIn[17]), .S(a58), .Z(HiOut[17]) );
    VMW_MUX2 U58 ( .A(BIn[5]), .B(AIn[5]), .S(a58), .Z(HiOut[5]) );
    VMW_MUX2 U43 ( .A(AIn[19]), .B(BIn[19]), .S(a58), .Z(LoOut[19]) );
    VMW_MUX2 U64 ( .A(BIn[29]), .B(AIn[29]), .S(a58), .Z(HiOut[29]) );
    VMW_MUX2 U81 ( .A(BIn[13]), .B(AIn[13]), .S(a58), .Z(HiOut[13]) );
    VMW_MUX2 U51 ( .A(AIn[11]), .B(BIn[11]), .S(a58), .Z(LoOut[11]) );
    VMW_MUX2 U76 ( .A(BIn[18]), .B(AIn[18]), .S(a58), .Z(HiOut[18]) );
    VMW_MUX2 U31 ( .A(AIn[2]), .B(BIn[2]), .S(a58), .Z(LoOut[2]) );
    VMW_MUX2 U38 ( .A(AIn[23]), .B(BIn[23]), .S(a58), .Z(LoOut[23]) );
    VMW_MUX2 U44 ( .A(AIn[18]), .B(BIn[18]), .S(a58), .Z(LoOut[18]) );
    VMW_MUX2 U56 ( .A(BIn[7]), .B(AIn[7]), .S(a58), .Z(HiOut[7]) );
    VMW_MUX2 U71 ( .A(BIn[22]), .B(AIn[22]), .S(a58), .Z(HiOut[22]) );
    VMW_MUX2 U63 ( .A(BIn[2]), .B(AIn[2]), .S(a58), .Z(HiOut[2]) );
    VMW_MUX2 U78 ( .A(BIn[16]), .B(AIn[16]), .S(a58), .Z(HiOut[16]) );
endmodule


module BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, In, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[31] , \ScanOut[5]1 , \ScanOut[4]1 , n245, n262, n217, n230, 
        n222, n199, n205, n257, n239, \ScanOut[23]1 , \ScanOut[8]1 , n202, 
        n250, n219, n225, n259, n210, n237, \ScanOut[10]1 , \ScanOut[22]1 , 
        \ScanOut[11]1 , n242, \ScanOut[9]1 , n197, n203, n224, n251, n206, 
        \ScanOut[19]1 , n196, n218, \ScanOut[26]1 , \ScanOut[18]1 , 
        \ScanOut[1]1 , \ScanOut[0]1 , n258, n243, \ScanOut[15]1 , n211, n236, 
        n216, n231, \ScanOut[27]1 , n244, \ScanOut[14]1 , n256, n238, n223, 
        n198, n204, n233, n228, n261, n246, n214, \ScanOut[28]1 , n221, 
        \ScanOut[3]1 , \ScanOut[30]1 , \ScanOut[29]1 , \ScanOut[2]1 , n254, 
        \ScanOut[25]1 , \ScanOut[24]1 , \ScanOut[17]1 , n253, n248, 
        \ScanOut[16]1 , n226, n201, n213, n234, n241, n194, n208, 
        \ScanOut[6]1 , n200, n227, n249, \ScanOut[7]1 , n252, n195, n209, n212, 
        n240, n235, n215, n260, n232, n247, \ScanOut[21]1 , n229, 
        \ScanOut[13]1 , \ScanOut[12]1 , n255, \ScanOut[20]1 , n207, n220;
    assign ScanOut[31] = \ScanOut[31] ;
    assign ScanOut[30] = \ScanOut[30]1 ;
    assign ScanOut[29] = \ScanOut[29]1 ;
    assign ScanOut[28] = \ScanOut[28]1 ;
    assign ScanOut[27] = \ScanOut[27]1 ;
    assign ScanOut[26] = \ScanOut[26]1 ;
    assign ScanOut[25] = \ScanOut[25]1 ;
    assign ScanOut[24] = \ScanOut[24]1 ;
    assign ScanOut[23] = \ScanOut[23]1 ;
    assign ScanOut[22] = \ScanOut[22]1 ;
    assign ScanOut[21] = \ScanOut[21]1 ;
    assign ScanOut[20] = \ScanOut[20]1 ;
    assign ScanOut[19] = \ScanOut[19]1 ;
    assign ScanOut[18] = \ScanOut[18]1 ;
    assign ScanOut[17] = \ScanOut[17]1 ;
    assign ScanOut[16] = \ScanOut[16]1 ;
    assign ScanOut[15] = \ScanOut[15]1 ;
    assign ScanOut[14] = \ScanOut[14]1 ;
    assign ScanOut[13] = \ScanOut[13]1 ;
    assign ScanOut[12] = \ScanOut[12]1 ;
    assign ScanOut[11] = \ScanOut[11]1 ;
    assign ScanOut[10] = \ScanOut[10]1 ;
    assign ScanOut[9] = \ScanOut[9]1 ;
    assign ScanOut[8] = \ScanOut[8]1 ;
    assign ScanOut[7] = \ScanOut[7]1 ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[31] = \ScanOut[31] ;
    assign Out[30] = \ScanOut[30]1 ;
    assign Out[29] = \ScanOut[29]1 ;
    assign Out[28] = \ScanOut[28]1 ;
    assign Out[27] = \ScanOut[27]1 ;
    assign Out[26] = \ScanOut[26]1 ;
    assign Out[25] = \ScanOut[25]1 ;
    assign Out[24] = \ScanOut[24]1 ;
    assign Out[23] = \ScanOut[23]1 ;
    assign Out[22] = \ScanOut[22]1 ;
    assign Out[21] = \ScanOut[21]1 ;
    assign Out[20] = \ScanOut[20]1 ;
    assign Out[19] = \ScanOut[19]1 ;
    assign Out[18] = \ScanOut[18]1 ;
    assign Out[17] = \ScanOut[17]1 ;
    assign Out[16] = \ScanOut[16]1 ;
    assign Out[15] = \ScanOut[15]1 ;
    assign Out[14] = \ScanOut[14]1 ;
    assign Out[13] = \ScanOut[13]1 ;
    assign Out[12] = \ScanOut[12]1 ;
    assign Out[11] = \ScanOut[11]1 ;
    assign Out[10] = \ScanOut[10]1 ;
    assign Out[9] = \ScanOut[9]1 ;
    assign Out[8] = \ScanOut[8]1 ;
    assign Out[7] = \ScanOut[7]1 ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U54 ( .A(\ScanOut[25]1 ), .B(n194), .C(n220), .Z(n237) );
    VMW_AO22 U73 ( .A(ScanIn[30]), .B(n230), .C(In[30]), .D(n228), .Z(n225) );
    VMW_AO22 U68 ( .A(ScanIn[6]), .B(n230), .C(In[6]), .D(n228), .Z(n201) );
    VMW_AO22 U96 ( .A(ScanIn[0]), .B(n230), .C(In[0]), .D(n228), .Z(n195) );
    VMW_AO21 U33 ( .A(\ScanOut[4]1 ), .B(n194), .C(n199), .Z(n258) );
    VMW_AO21 U34 ( .A(\ScanOut[5]1 ), .B(n194), .C(n200), .Z(n257) );
    VMW_AO21 U41 ( .A(\ScanOut[12]1 ), .B(n194), .C(n207), .Z(n250) );
    VMW_AO21 U46 ( .A(\ScanOut[17]1 ), .B(n194), .C(n212), .Z(n245) );
    VMW_NOR2 U61 ( .A(Reset), .B(n194), .Z(n227) );
    VMW_AO22 U84 ( .A(ScanIn[20]), .B(n230), .C(In[20]), .D(n228), .Z(n215) );
    VMW_AO22 U66 ( .A(ScanIn[8]), .B(n230), .C(In[8]), .D(n228), .Z(n203) );
    VMW_AO22 U83 ( .A(ScanIn[21]), .B(n230), .C(In[21]), .D(n228), .Z(n216) );
    VMW_AO21 U35 ( .A(\ScanOut[6]1 ), .B(n194), .C(n201), .Z(n256) );
    VMW_AO21 U48 ( .A(\ScanOut[19]1 ), .B(n194), .C(n214), .Z(n243) );
    VMW_AO21 U53 ( .A(\ScanOut[24]1 ), .B(n194), .C(n219), .Z(n238) );
    VMW_AO22 U91 ( .A(ScanIn[14]), .B(n230), .C(In[14]), .D(n228), .Z(n209) );
    VMW_AO22 U74 ( .A(ScanIn[2]), .B(n230), .C(In[2]), .D(n228), .Z(n197) );
    VMW_FD \Out_reg[25]  ( .D(n237), .CP(Clk), .Q(\ScanOut[25]1 ) );
    VMW_FD \Out_reg[16]  ( .D(n246), .CP(Clk), .Q(\ScanOut[16]1 ) );
    VMW_AO21 U29 ( .A(\ScanOut[0]1 ), .B(n194), .C(n195), .Z(n262) );
    VMW_AO21 U40 ( .A(\ScanOut[11]1 ), .B(n194), .C(n206), .Z(n251) );
    VMW_AO22 U82 ( .A(ScanIn[22]), .B(n230), .C(In[22]), .D(n228), .Z(n217) );
    VMW_FD \Out_reg[5]  ( .D(n257), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO21 U47 ( .A(\ScanOut[18]1 ), .B(n194), .C(n213), .Z(n244) );
    VMW_AO21 U49 ( .A(\ScanOut[20]1 ), .B(n194), .C(n215), .Z(n242) );
    VMW_AO21 U52 ( .A(\ScanOut[23]1 ), .B(n194), .C(n218), .Z(n239) );
    VMW_AO22 U67 ( .A(ScanIn[7]), .B(n230), .C(In[7]), .D(n228), .Z(n202) );
    VMW_AO22 U75 ( .A(ScanIn[29]), .B(n230), .C(In[29]), .D(n228), .Z(n224) );
    VMW_FD \Out_reg[12]  ( .D(n250), .CP(Clk), .Q(\ScanOut[12]1 ) );
    VMW_AO22 U90 ( .A(ScanIn[15]), .B(n230), .C(In[15]), .D(n228), .Z(n210) );
    VMW_FD \Out_reg[21]  ( .D(n241), .CP(Clk), .Q(\ScanOut[21]1 ) );
    VMW_FD \Out_reg[31]  ( .D(n231), .CP(Clk), .Q(\ScanOut[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n234), .CP(Clk), .Q(\ScanOut[28]1 ) );
    VMW_FD \Out_reg[8]  ( .D(n254), .CP(Clk), .Q(\ScanOut[8]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n261), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO21 U55 ( .A(\ScanOut[26]1 ), .B(n194), .C(n221), .Z(n236) );
    VMW_AO22 U69 ( .A(ScanIn[5]), .B(n230), .C(In[5]), .D(n228), .Z(n200) );
    VMW_FD \Out_reg[19]  ( .D(n243), .CP(Clk), .Q(\ScanOut[19]1 ) );
    VMW_AO22 U72 ( .A(ScanIn[31]), .B(n230), .C(In[31]), .D(n228), .Z(n226) );
    VMW_INV U97 ( .A(n227), .Z(n229) );
    VMW_FD \Out_reg[3]  ( .D(n259), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[23]  ( .D(n239), .CP(Clk), .Q(\ScanOut[23]1 ) );
    VMW_FD \Out_reg[10]  ( .D(n252), .CP(Clk), .Q(\ScanOut[10]1 ) );
    VMW_AO21 U60 ( .A(\ScanOut[31] ), .B(n194), .C(n226), .Z(n231) );
    VMW_FD \Out_reg[7]  ( .D(n255), .CP(Clk), .Q(\ScanOut[7]1 ) );
    VMW_AO21 U32 ( .A(\ScanOut[3]1 ), .B(n194), .C(n198), .Z(n259) );
    VMW_AO22 U85 ( .A(ScanIn[1]), .B(n230), .C(In[1]), .D(n228), .Z(n196) );
    VMW_FD \Out_reg[27]  ( .D(n235), .CP(Clk), .Q(\ScanOut[27]1 ) );
    VMW_FD \Out_reg[14]  ( .D(n248), .CP(Clk), .Q(\ScanOut[14]1 ) );
    VMW_AO21 U30 ( .A(\ScanOut[1]1 ), .B(n194), .C(n196), .Z(n261) );
    VMW_AO21 U39 ( .A(\ScanOut[10]1 ), .B(n194), .C(n205), .Z(n252) );
    VMW_AO21 U57 ( .A(\ScanOut[28]1 ), .B(n194), .C(n223), .Z(n234) );
    VMW_FD \Out_reg[6]  ( .D(n256), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U70 ( .A(ScanIn[4]), .B(n230), .C(In[4]), .D(n228), .Z(n199) );
    VMW_AO22 U79 ( .A(ScanIn[25]), .B(n230), .C(In[25]), .D(n228), .Z(n220) );
    VMW_AO22 U95 ( .A(ScanIn[10]), .B(n230), .C(In[10]), .D(n228), .Z(n205) );
    VMW_FD \Out_reg[26]  ( .D(n236), .CP(Clk), .Q(\ScanOut[26]1 ) );
    VMW_FD \Out_reg[15]  ( .D(n247), .CP(Clk), .Q(\ScanOut[15]1 ) );
    VMW_FD \Out_reg[18]  ( .D(n244), .CP(Clk), .Q(\ScanOut[18]1 ) );
    VMW_AO21 U31 ( .A(\ScanOut[2]1 ), .B(n194), .C(n197), .Z(n260) );
    VMW_AO21 U36 ( .A(\ScanOut[7]1 ), .B(n194), .C(n202), .Z(n255) );
    VMW_AO21 U37 ( .A(\ScanOut[8]1 ), .B(n194), .C(n203), .Z(n254) );
    VMW_AO21 U42 ( .A(\ScanOut[13]1 ), .B(n194), .C(n208), .Z(n249) );
    VMW_AO21 U45 ( .A(\ScanOut[16]1 ), .B(n194), .C(n211), .Z(n246) );
    VMW_AO22 U87 ( .A(ScanIn[18]), .B(n230), .C(In[18]), .D(n228), .Z(n213) );
    VMW_FD \Out_reg[2]  ( .D(n260), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[11]  ( .D(n251), .CP(Clk), .Q(\ScanOut[11]1 ) );
    VMW_NOR2 U62 ( .A(n229), .B(ScanEnable), .Z(n228) );
    VMW_FD \Out_reg[22]  ( .D(n240), .CP(Clk), .Q(\ScanOut[22]1 ) );
    VMW_AO22 U65 ( .A(ScanIn[9]), .B(n230), .C(In[9]), .D(n228), .Z(n204) );
    VMW_FD \Out_reg[20]  ( .D(n242), .CP(Clk), .Q(\ScanOut[20]1 ) );
    VMW_FD \Out_reg[13]  ( .D(n249), .CP(Clk), .Q(\ScanOut[13]1 ) );
    VMW_AO22 U80 ( .A(ScanIn[24]), .B(n230), .C(In[24]), .D(n228), .Z(n219) );
    VMW_FD \Out_reg[9]  ( .D(n253), .CP(Clk), .Q(\ScanOut[9]1 ) );
    VMW_AO21 U50 ( .A(\ScanOut[21]1 ), .B(n194), .C(n216), .Z(n241) );
    VMW_AO21 U59 ( .A(\ScanOut[30]1 ), .B(n194), .C(n225), .Z(n232) );
    VMW_FD \Out_reg[30]  ( .D(n232), .CP(Clk), .Q(\ScanOut[30]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n262), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_FD \Out_reg[29]  ( .D(n233), .CP(Clk), .Q(\ScanOut[29]1 ) );
    VMW_AO22 U77 ( .A(ScanIn[27]), .B(n230), .C(In[27]), .D(n228), .Z(n222) );
    VMW_AO22 U89 ( .A(ScanIn[16]), .B(n230), .C(In[16]), .D(n228), .Z(n211) );
    VMW_AO22 U92 ( .A(ScanIn[13]), .B(n230), .C(In[13]), .D(n228), .Z(n208) );
    VMW_FD \Out_reg[24]  ( .D(n238), .CP(Clk), .Q(\ScanOut[24]1 ) );
    VMW_FD \Out_reg[17]  ( .D(n245), .CP(Clk), .Q(\ScanOut[17]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n258), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_AO21 U58 ( .A(\ScanOut[29]1 ), .B(n194), .C(n224), .Z(n233) );
    VMW_AO21 U38 ( .A(\ScanOut[9]1 ), .B(n194), .C(n204), .Z(n253) );
    VMW_AO21 U43 ( .A(\ScanOut[14]1 ), .B(n194), .C(n209), .Z(n248) );
    VMW_NOR3 U64 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n194) );
    VMW_AO22 U81 ( .A(ScanIn[23]), .B(n230), .C(In[23]), .D(n228), .Z(n218) );
    VMW_AO21 U51 ( .A(\ScanOut[22]1 ), .B(n194), .C(n217), .Z(n240) );
    VMW_AO22 U76 ( .A(ScanIn[28]), .B(n230), .C(In[28]), .D(n228), .Z(n223) );
    VMW_AO22 U88 ( .A(ScanIn[17]), .B(n230), .C(In[17]), .D(n228), .Z(n212) );
    VMW_AO22 U93 ( .A(ScanIn[12]), .B(n230), .C(In[12]), .D(n228), .Z(n207) );
    VMW_AO21 U44 ( .A(\ScanOut[15]1 ), .B(n194), .C(n210), .Z(n247) );
    VMW_AO21 U56 ( .A(\ScanOut[27]1 ), .B(n194), .C(n222), .Z(n235) );
    VMW_AO22 U94 ( .A(ScanIn[11]), .B(n230), .C(In[11]), .D(n228), .Z(n206) );
    VMW_AO22 U71 ( .A(ScanIn[3]), .B(n230), .C(In[3]), .D(n228), .Z(n198) );
    VMW_AND2 U63 ( .A(ScanEnable), .B(n227), .Z(n230) );
    VMW_AO22 U86 ( .A(ScanIn[19]), .B(n230), .C(In[19]), .D(n228), .Z(n214) );
    VMW_AO22 U78 ( .A(ScanIn[26]), .B(n230), .C(In[26]), .D(n228), .Z(n221) );
endmodule


module BubbleSort_Control_CWIDTH6_IDWIDTH1_WIDTH32_SCAN1_DW01_dec_6_0 ( A, SUM
     );
input  [5:0] A;
output [5:0] SUM;
    wire n5, n7, n9, n6, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[3]), .C(n6), .Z(SUM[3]) );
    VMW_INV U5 ( .A(A[0]), .Z(SUM[0]) );
    VMW_OAI21 U6 ( .A(n7), .B(n8), .C(n5), .Z(SUM[2]) );
    VMW_INV U14 ( .A(n6), .Z(n11) );
    VMW_AND2 U7 ( .A(n6), .B(n10), .Z(n9) );
    VMW_NOR2 U8 ( .A(A[0]), .B(A[1]), .Z(n7) );
    VMW_INV U13 ( .A(A[4]), .Z(n10) );
    VMW_NAND2 U9 ( .A(n7), .B(n8), .Z(n5) );
    VMW_AO22 U12 ( .A(A[4]), .B(n11), .C(n10), .D(n6), .Z(SUM[4]) );
    VMW_INV U15 ( .A(A[2]), .Z(n8) );
    VMW_NOR2 U10 ( .A(n5), .B(A[3]), .Z(n6) );
    VMW_XOR2 U11 ( .A(A[5]), .B(n9), .Z(SUM[5]) );
    VMW_AO21 U4 ( .A(A[0]), .B(A[1]), .C(n7), .Z(SUM[1]) );
endmodule


module BubbleSort_Control_CWIDTH6_IDWIDTH1_WIDTH32_SCAN1 ( Clk, Reset, RD, WR, 
    Addr, DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n330, n317, \count[2] , n362, n345, n339, n357, n322, n325, n350, 
        n319, \count[4] , n342, n365, \count[0] , n359, n356, n337, n318, n351, 
        \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , n324, \count260[3] , 
        \ScanReg[18] , n336, n358, n364, n343, \ScanReg[22] , \ScanReg[11] , 
        \ScanReg[6] , \ScanReg[20] , \ScanReg[13] , \ScanReg[4] , n344, n363, 
        \count260[5] , \ScanReg[29] , n316, \ScanReg[30] , n331, n323, 
        \count260[1] , \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , 
        \ScanReg[9] , n338, n314, n333, \count260[0] , \ScanReg[16] , 
        \ScanReg[25] , \ScanReg[8] , n346, \ScanReg[1] , n361, \ScanReg[7] , 
        n328, \ScanReg[5] , n354, \ScanReg[21] , \ScanReg[12] , \count260[4] , 
        \ScanReg[28] , \ScanReg[31] , n321, \ScanReg[19] , n326, n348, n353, 
        \ScanReg[10] , \ScanReg[23] , n341, \ScanReg[14] , \ScanReg[27] , n313, 
        \ScanReg[3] , n334, \count260[2] , \count[1] , n352, n349, n327, n335, 
        n360, n340, \count[5] , n347, n329, n332, n315, n320, \count[3] , n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U73 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_AOI21 U113 ( .A(n324), .B(n313), .C(Reset), .Z(n317) );
    VMW_INV U134 ( .A(n315), .Z(n316) );
    VMW_AND2 U68 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AND2 U96 ( .A(\ScanReg[16] ), .B(n315), .Z(n337) );
    VMW_AND2 U108 ( .A(n317), .B(n321), .Z(n363) );
    VMW_BUFIZ U141 ( .A(n330), .E(n332), .Z(\arr[10] ) );
    VMW_BUFIZ U166 ( .A(n356), .E(n332), .Z(\arr[22] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AND2 U53 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U61 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U84 ( .A(\ScanReg[7] ), .B(n315), .Z(n351) );
    VMW_BUFIZ U148 ( .A(n338), .E(n332), .Z(\arr[12] ) );
    VMW_BUFIZ U153 ( .A(n343), .E(n332), .Z(\arr[2] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    VMW_FD \count_reg[2]  ( .D(n363), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U66 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U101 ( .A(\ScanReg[10] ), .B(n315), .Z(n330) );
    VMW_AND2 U106 ( .A(n317), .B(n319), .Z(n361) );
    VMW_AO22 U121 ( .A(\count[4] ), .B(n316), .C(\ScanReg[4] ), .D(n315), .Z(
        n333) );
    VMW_OR3 U126 ( .A(\count[3] ), .B(\count[5] ), .C(\count[4] ), .Z(n314) );
    VMW_AND2 U83 ( .A(\ScanReg[26] ), .B(n315), .Z(n353) );
    VMW_BUFIZ U168 ( .A(n358), .E(n332), .Z(\arr[1] ) );
    VMW_FD \count_reg[0]  ( .D(n365), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U91 ( .A(\ScanReg[28] ), .B(n315), .Z(n342) );
    VMW_AND2 U98 ( .A(\ScanReg[14] ), .B(n315), .Z(n335) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(ScanOut[5]), .B(n316), .C(\count260[5] ), .D(n324), .Z(
        n318) );
    VMW_BUFIZ U154 ( .A(n344), .E(n332), .Z(\arr[13] ) );
    VMW_FD \count_reg[4]  ( .D(n361), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n336), .E(n332), .Z(\arr[25] ) );
    VMW_BUFIZ U161 ( .A(n351), .E(n332), .Z(\arr[7] ) );
    VMW_AND2 U74 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_AND2 U114 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AO22 U133 ( .A(ScanOut[0]), .B(n316), .C(\count260[0] ), .D(n324), .Z(
        n323) );
    VMW_AND2 U99 ( .A(\ScanReg[27] ), .B(n315), .Z(n334) );
    VMW_BUFIZ U155 ( .A(n345), .E(n332), .Z(\arr[30] ) );
    VMW_AND2 U52 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U67 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AND2 U82 ( .A(\ScanReg[15] ), .B(n315), .Z(n354) );
    VMW_BUFIZ U169 ( .A(n359), .E(n332), .Z(\arr[8] ) );
    VMW_AND2 U107 ( .A(n317), .B(n320), .Z(n362) );
    VMW_AO22 U120 ( .A(\count[5] ), .B(n316), .C(\ScanReg[5] ), .D(n315), .Z(
        n352) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U55 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U69 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U75 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U115 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AO22 U132 ( .A(ScanOut[1]), .B(n316), .C(\count260[1] ), .D(n324), .Z(
        n322) );
    VMW_AND2 U90 ( .A(\ScanReg[13] ), .B(n315), .Z(n344) );
    VMW_AND2 U109 ( .A(n317), .B(n322), .Z(n364) );
    VMW_AO22 U129 ( .A(ScanOut[4]), .B(n316), .C(\count260[4] ), .D(n324), .Z(
        n319) );
    VMW_BUFIZ U147 ( .A(n337), .E(n332), .Z(\arr[16] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n350), .E(n332), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U97 ( .A(\ScanReg[25] ), .B(n315), .Z(n336) );
    VMW_BUFIZ U140 ( .A(n329), .E(n332), .Z(\arr[23] ) );
    VMW_BUFIZ U167 ( .A(n357), .E(n332), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_AND2 U112 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_XNOR2 U135 ( .A(Addr[0]), .B(ScanId), .Z(n326) );
    BubbleSort_Control_CWIDTH6_IDWIDTH1_WIDTH32_SCAN1_DW01_dec_6_0 sub_202 ( 
        .A({\count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[5] , \count260[4] , \count260[3] , 
        \count260[2] , \count260[1] , \count260[0] }) );
    VMW_AND2 U60 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U85 ( .A(\ScanReg[17] ), .B(n315), .Z(n350) );
    VMW_AND2 U100 ( .A(\ScanReg[9] ), .B(n315), .Z(n331) );
    VMW_NAND2 U127 ( .A(n316), .B(WR), .Z(n324) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n339), .E(n332), .Z(\arr[6] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n342), .E(n332), .Z(\arr[28] ) );
    VMW_NOR4 U51 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n314), 
        .Z(n313) );
    VMW_AND2 U57 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_INV U137 ( .A(n325), .Z(ScanEnable) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U58 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U62 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U70 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AND2 U79 ( .A(\ScanReg[11] ), .B(n315), .Z(n357) );
    VMW_AND2 U95 ( .A(\ScanReg[12] ), .B(n315), .Z(n338) );
    VMW_AND2 U110 ( .A(n317), .B(n323), .Z(n365) );
    VMW_BUFIZ U159 ( .A(n349), .E(n332), .Z(\arr[24] ) );
    VMW_OAI21 U119 ( .A(RD), .B(WR), .C(n326), .Z(n325) );
    VMW_BUFIZ U142 ( .A(n331), .E(n332), .Z(\arr[9] ) );
    VMW_BUFIZ U165 ( .A(n355), .E(n332), .Z(\arr[18] ) );
    VMW_AND2 U87 ( .A(\ScanReg[20] ), .B(n315), .Z(n347) );
    VMW_BUFIZ U150 ( .A(n340), .E(n332), .Z(\arr[31] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(\count[0] ), .B(n316), .C(\ScanReg[0] ), .D(n315), .Z(
        n328) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U65 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U102 ( .A(\ScanReg[23] ), .B(n315), .Z(n329) );
    VMW_AND2 U105 ( .A(n317), .B(n318), .Z(n360) );
    VMW_AND2 U80 ( .A(\ScanReg[22] ), .B(n315), .Z(n356) );
    VMW_AO22 U122 ( .A(\count[3] ), .B(n316), .C(\ScanReg[3] ), .D(n315), .Z(
        n348) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_BUFIZ U139 ( .A(n328), .E(n332), .Z(\arr[0] ) );
    VMW_BUFIZ U157 ( .A(n347), .E(n332), .Z(\arr[20] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AND2 U77 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_AND2 U89 ( .A(\ScanReg[30] ), .B(n315), .Z(n345) );
    VMW_AND2 U92 ( .A(\ScanReg[21] ), .B(n315), .Z(n341) );
    VMW_BUFIZ U145 ( .A(n335), .E(n332), .Z(\arr[14] ) );
    VMW_BUFIZ U162 ( .A(n352), .E(n332), .Z(\arr[5] ) );
    VMW_AND2 U117 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AO22 U130 ( .A(ScanOut[3]), .B(n316), .C(\count260[3] ), .D(n324), .Z(
        n320) );
    VMW_BUFIZ U138 ( .A(n327), .E(n332), .Z(\arr[19] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n360), .CP(Clk), .Q(\count[5] ) );
    VMW_AND2 U64 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AND2 U81 ( .A(\ScanReg[18] ), .B(n315), .Z(n355) );
    VMW_BUFIZ U156 ( .A(n346), .E(n332), .Z(\arr[29] ) );
    VMW_AND2 U104 ( .A(\ScanReg[19] ), .B(n315), .Z(n327) );
    VMW_AND2 U76 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U116 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_AO22 U123 ( .A(\count[2] ), .B(n316), .C(\ScanReg[2] ), .D(n315), .Z(
        n343) );
    VMW_AND2 U56 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U88 ( .A(\ScanReg[29] ), .B(n315), .Z(n346) );
    VMW_AND2 U93 ( .A(\ScanReg[31] ), .B(n315), .Z(n340) );
    VMW_AO22 U131 ( .A(ScanOut[2]), .B(n316), .C(\count260[2] ), .D(n324), .Z(
        n321) );
    VMW_FD \count_reg[1]  ( .D(n364), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[6] ), .B(n315), .Z(n339) );
    VMW_BUFIZ U143 ( .A(n333), .E(n332), .Z(\arr[4] ) );
    VMW_BUFIZ U144 ( .A(n334), .E(n332), .Z(\arr[27] ) );
    VMW_BUFIZ U163 ( .A(n353), .E(n332), .Z(\arr[26] ) );
    VMW_BUFIZ U158 ( .A(n348), .E(n332), .Z(\arr[3] ) );
    VMW_BUFIZ U164 ( .A(n354), .E(n332), .Z(\arr[15] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_FD \count_reg[3]  ( .D(n362), .CP(Clk), .Q(\count[3] ) );
    VMW_INV U136 ( .A(n313), .Z(Enable) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U63 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U71 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_XOR2 U111 ( .A(Addr[0]), .B(Id), .Z(n315) );
    VMW_AO22 U124 ( .A(\count[1] ), .B(n316), .C(\ScanReg[1] ), .D(n315), .Z(
        n358) );
    VMW_AND2 U78 ( .A(\ScanReg[8] ), .B(n315), .Z(n359) );
    VMW_AND2 U86 ( .A(\ScanReg[24] ), .B(n315), .Z(n349) );
    VMW_AO21 U103 ( .A(RD), .B(ScanEnable), .C(n316), .Z(n332) );
    VMW_AND2 U118 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_BUFIZ U151 ( .A(n341), .E(n332), .Z(\arr[21] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wRegInA0[9] , \wAMid11[23] , \wRegInB30[28] , \wAMid27[26] , 
        \wBIn28[21] , \wAIn29[19] , \wRegInB13[19] , \wRegInB30[31] , 
        \wAIn1[3] , \wAIn2[0] , \wBMid9[13] , \wAIn25[6] , \ScanLink51[31] , 
        \ScanLink51[28] , \ScanLink50[8] , \ScanLink24[18] , \wRegInB2[12] , 
        \wRegInA4[17] , \wAMid8[18] , \wBMid9[20] , \wAIn26[5] , 
        \ScanLink0[13] , \wAMid27[15] , \wBIn28[12] , \ScanLink29[3] , 
        \wBIn0[27] , \wBIn0[9] , \wRegInA0[26] , \wRegInA0[15] , \wAIn3[21] , 
        \wAIn3[12] , \wBMid2[9] , \wAMid3[27] , \wAMid3[14] , \wAIn7[10] , 
        \wAMid11[10] , \wBIn24[1] , \wBIn27[2] , \wBMid26[13] , \wRegInB2[21] , 
        \wRegInA4[24] , \ScanLink0[20] , \ScanLink19[22] , \wRegInA6[7] , 
        \wAIn7[23] , \wBMid10[16] , \wRegInA16[2] , \wAIn14[23] , 
        \ScanLink56[6] , \wAIn14[10] , \wBIn15[31] , \wBIn15[28] , 
        \wBMid14[0] , \wBMid17[3] , \wAIn22[26] , \wAIn23[8] , \wRegInA10[21] , 
        \wRegInB18[26] , \wRegInA26[24] , \ScanLink55[5] , \wRegInA5[4] , 
        \wRegInA15[1] , \ScanLink9[6] , \wRegInB18[15] , \ScanLink32[2] , 
        \wAIn22[15] , \wRegInB12[3] , \wBMid10[25] , \wBIn18[5] , \wAMid19[4] , 
        \wBMid26[20] , \wRegInB11[0] , \ScanLink19[11] , \wRegInA10[12] , 
        \ScanLink31[1] , \wRegInA26[17] , \wRegInA14[23] , \wBIn8[1] , 
        \wBIn11[19] , \wRegInA22[26] , \wRegInB28[9] , \ScanLink15[7] , 
        \wAIn26[24] , \wAIn10[21] , \ScanLink16[4] , \wAMid7[16] , 
        \wBMid14[14] , \wAIn19[2] , \wBMid22[11] , \wBMid30[6] , 
        \wRegInA14[10] , \wRegInA22[15] , \wBMid22[22] , \wRegInA31[7] , 
        \wAMid7[25] , \wBMid14[27] , \wAIn10[12] , \wAMid28[28] , \wAIn26[17] , 
        \wAMid28[31] , \wRegInA29[19] , \ScanLink4[11] , \wBMid4[7] , 
        \wAMid26[3] , \wRegInB6[10] , \ScanLink13[9] , \wBMid7[4] , 
        \wAMid25[0] , \wAMid15[21] , \wAMid23[24] , \wRegInB6[23] , 
        \wAIn2[18] , \wBIn5[4] , \wAMid5[0] , \ScanLink4[22] , \wAMid6[3] , 
        \wAMid15[12] , \wAMid23[17] , \wBMid28[4] , \wRegInB17[31] , 
        \wRegInB17[28] , \wBMid7[17] , \wBIn10[20] , \wAIn11[18] , 
        \wRegInB9[0] , \wRegInA29[5] , \ScanLink20[30] , \ScanLink55[19] , 
        \ScanLink20[29] , \wAIn17[4] , \wBIn26[25] , \wAMid29[22] , 
        \wBMid23[31] , \wBMid23[28] , \wAIn14[7] , \wRegInB1[8] , 
        \ScanLink61[9] , \wBIn16[3] , \wBIn4[25] , \wBIn6[7] , \wBMid7[24] , 
        \wBIn10[13] , \wBIn15[0] , \wBIn26[16] , \wAMid29[11] , \wAMid30[7] , 
        \wRegInA15[30] , \wRegInA15[29] , \wAIn9[14] , \ScanLink54[13] , 
        \ScanLink21[23] , \ScanLink18[2] , \wAIn12[9] , \wAMid14[18] , 
        \wBMid25[1] , \wBMid28[17] , \ScanLink62[16] , \ScanLink17[26] , 
        \wRegInB16[22] , \wRegInA24[0] , \ScanLink64[4] , \ScanLink41[27] , 
        \ScanLink34[17] , \wBMid26[2] , \wRegInB4[5] , \wRegInB7[30] , 
        \wRegInB7[6] , \wRegInB20[27] , \wRegInA27[3] , \ScanLink5[28] , 
        \wRegInA28[20] , \ScanLink5[31] , \wRegInB7[29] , \wBIn4[16] , 
        \wAMid8[5] , \wAIn9[27] , \wAMid28[5] , \wRegInB20[14] , \wBMid28[24] , 
        \wRegInB16[11] , \wRegInB20[1] , \ScanLink62[25] , \ScanLink54[20] , 
        \ScanLink41[14] , \ScanLink17[15] , \ScanLink34[24] , \ScanLink21[10] , 
        \wRegInA28[13] , \wBMid9[2] , \wRegInB23[2] , \ScanLink27[5] , 
        \wBIn0[14] , \wAMid9[12] , \wAIn28[20] , \wBIn29[18] , \wRegInB24[25] , 
        \ScanLink39[9] , \wRegInB31[11] , \wRegInB12[20] , \wRegInB19[8] , 
        \ScanLink13[24] , \ScanLink45[25] , \ScanLink30[15] , \ScanLink25[21] , 
        \ScanLink24[6] , \wBIn29[4] , \wRegInB3[18] , \ScanLink50[11] , 
        \ScanLink1[19] , \ScanLink43[1] , \wBMid3[15] , \wAIn6[30] , 
        \wBMid8[19] , \wAMid9[21] , \ScanLink50[22] , \ScanLink40[2] , 
        \ScanLink45[16] , \ScanLink25[12] , \ScanLink13[17] , \wAMid10[30] , 
        \wAIn28[13] , \wRegInB12[13] , \ScanLink30[26] , \wAMid10[29] , 
        \wRegInB31[22] , \wAMid14[1] , \wAIn28[3] , \wRegInB24[16] , 
        \wRegInA11[18] , \wBIn31[6] , \wRegInB8[14] , \wAIn6[29] , 
        \wBIn14[22] , \ScanLink22[8] , \wAMid17[2] , \wBMid19[5] , 
        \wBIn22[27] , \ScanLink58[0] , \wRegInB8[27] , \wBIn0[0] , \wBIn3[3] , 
        \wBMid3[26] , \wBIn14[11] , \wAIn15[30] , \wAIn15[29] , \wAIn30[1] , 
        \wRegInA8[1] , \ScanLink4[3] , \wRegInA18[4] , \ScanLink7[0] , 
        \wBIn22[14] , \wBMid27[19] , \ScanLink18[28] , \ScanLink18[31] , 
        \wAMid14[22] , \wRegInB16[18] , \wRegInB20[8] , \wAMid22[27] , 
        \wBIn10[4] , \wBIn13[7] , \wRegInA1[16] , \wRegInB7[13] , 
        \ScanLink54[30] , \ScanLink54[29] , \ScanLink21[19] , \ScanLink5[12] , 
        \wRegInA0[0] , \wBIn1[24] , \wAIn2[22] , \wAIn2[11] , \wAMid6[15] , 
        \wAIn11[3] , \wAIn12[0] , \wAMid14[11] , \wAMid22[14] , \wBMid25[8] , 
        \wRegInA24[9] , \wRegInA1[25] , \wRegInA28[30] , \wRegInA28[29] , 
        \ScanLink5[21] , \wBMid23[12] , \wRegInB7[20] , \wRegInB26[6] , 
        \wBMid15[17] , \wAMid6[26] , \wBIn10[30] , \wAIn11[22] , \wBIn15[9] , 
        \wAIn27[27] , \wAMid29[18] , \wRegInA15[20] , \wRegInA23[25] , 
        \wRegInB25[5] , \wAIn27[14] , \ScanLink62[3] , \wBIn10[29] , 
        \wAIn11[11] , \wBMid23[6] , \wBMid15[24] , \wAMid2[24] , \wAMid2[17] , 
        \wBIn14[18] , \wBMid20[5] , \wBMid23[21] , \wRegInB1[1] , 
        \wRegInB2[2] , \wRegInA21[4] , \wRegInA22[7] , \wRegInA15[13] , 
        \wRegInA23[16] , \wEnable[0] , \ScanLink61[0] , \wAIn23[25] , 
        \wAIn30[8] , \wRegInA8[8] , \ScanLink58[9] , \wRegInA11[22] , 
        \wRegInA27[27] , \ScanLink45[6] , \wRegInB19[25] , \wAIn15[20] , 
        \ScanLink46[5] , \ScanLink7[9] , \wAIn6[13] , \wBMid11[15] , 
        \wAIn9[2] , \wBMid11[26] , \wAMid14[8] , \wBMid27[10] , 
        \ScanLink18[21] , \wRegInA27[14] , \wBMid27[23] , \wRegInA11[11] , 
        \ScanLink21[2] , \ScanLink18[12] , \wBMid2[25] , \wBMid2[16] , 
        \wAIn6[20] , \wBMid8[23] , \wBMid8[10] , \wAIn15[13] , \wAIn23[16] , 
        \wRegInB19[16] , \ScanLink22[1] , \wRegInB3[11] , \wRegInA5[14] , 
        \ScanLink1[10] , \ScanLink2[4] , \ScanLink43[8] , \wAMid9[31] , 
        \wAMid9[28] , \ScanLink1[7] , \wAMid10[20] , \wAMid26[25] , 
        \wBIn29[22] , \wAMid10[13] , \wAMid12[6] , \wAIn28[29] , 
        \wRegInB3[22] , \wRegInA5[27] , \ScanLink1[23] , \wRegInB12[29] , 
        \wAMid11[5] , \wAMid26[16] , \wAIn28[30] , \wBIn29[11] , 
        \wRegInB31[18] , \wRegInB12[30] , \ScanLink50[18] , \ScanLink39[0] , 
        \ScanLink25[28] , \wRegInB19[1] , \ScanLink25[31] , \wAIn14[19] , 
        \wBIn23[24] , \wBIn15[21] , \wBMid26[30] , \wAIn7[19] , \wBIn21[5] , 
        \wBIn22[6] , \wBMid26[29] , \ScanLink19[18] , \wRegInB9[17] , 
        \wRegInB11[9] , \ScanLink31[8] , \wAIn4[7] , \wBIn15[12] , \wAIn7[4] , 
        \wBMid14[9] , \wAIn20[2] , \wAIn23[1] , \wBIn23[17] , \wRegInA10[31] , 
        \wRegInA10[28] , \wAMid8[11] , \wRegInB9[24] , \wRegInA15[8] , 
        \ScanLink48[3] , \ScanLink24[22] , \wBMid9[30] , \wBMid9[29] , 
        \ScanLink51[12] , \ScanLink44[26] , \ScanLink31[16] , \ScanLink34[5] , 
        \ScanLink12[27] , \wAMid11[19] , \wBIn24[8] , \wAIn29[23] , 
        \wRegInB30[12] , \wRegInB2[31] , \wRegInB2[28] , \wRegInB13[23] , 
        \wRegInB14[4] , \wRegInB17[7] , \wRegInB25[26] , \ScanLink0[30] , 
        \ScanLink0[29] , \wBIn28[28] , \wRegInA10[5] , \ScanLink37[6] , 
        \wBIn1[17] , \wAIn2[9] , \wBIn28[31] , \wRegInB25[15] , \wAIn29[10] , 
        \wRegInB13[10] , \wRegInB30[21] , \ScanLink44[15] , \ScanLink31[25] , 
        \wAMid8[22] , \wBMid11[4] , \ScanLink12[14] , \ScanLink51[21] , 
        \ScanLink50[1] , \wBMid12[7] , \ScanLink24[11] , \wBIn5[26] , 
        \wRegInA3[3] , \ScanLink53[2] , \wRegInA13[6] , \wAMid5[9] , 
        \wAIn8[17] , \wBMid29[14] , \wRegInB17[21] , \wRegInB21[24] , 
        \wRegInA29[23] , \ScanLink63[15] , \ScanLink40[24] , \ScanLink35[14] , 
        \ScanLink16[25] , \wRegInB6[19] , \wRegInB9[9] , \wRegInA29[10] , 
        \ScanLink55[10] , \ScanLink20[20] , \ScanLink4[18] , \wAMid0[4] , 
        \wAIn3[28] , \wAMid3[7] , \wBIn5[15] , \ScanLink13[0] , \wAIn8[24] , 
        \wAMid15[31] , \wAMid15[28] , \wAMid25[9] , \wBMid29[27] , 
        \ScanLink63[26] , \ScanLink55[23] , \ScanLink40[17] , \ScanLink20[13] , 
        \ScanLink10[3] , \ScanLink35[27] , \wRegInB30[2] , \ScanLink16[16] , 
        \wRegInB17[12] , \wRegInA14[19] , \wRegInB21[17] , \wBMid1[3] , 
        \wAIn3[31] , \wBMid2[0] , \wBMid6[14] , \wBIn11[23] , \wBIn27[26] , 
        \wAMid28[21] , \wAIn10[31] , \wAMid20[4] , \wRegInB28[0] , 
        \wAMid28[12] , \wAIn10[28] , \wBIn27[15] , \wAMid2[30] , \wBMid3[11] , 
        \wBMid6[27] , \wBIn8[8] , \wBIn11[10] , \wAMid23[7] , \wBIn14[26] , 
        \wAMid17[6] , \wBIn22[23] , \wBMid22[18] , \wAMid2[29] , \wBMid3[22] , 
        \wBMid11[18] , \wAMid14[5] , \wBIn31[2] , \wRegInB8[10] , 
        \wRegInA27[19] , \wBIn14[15] , \wBIn22[10] , \wAIn23[31] , 
        \wAIn23[28] , \wRegInB19[31] , \wRegInB19[28] , \wAIn30[5] , 
        \wRegInA18[0] , \ScanLink46[8] , \ScanLink7[4] , \wRegInA8[5] , 
        \wBIn0[23] , \wAMid9[16] , \wAMid11[8] , \wBMid19[1] , \wRegInB8[23] , 
        \ScanLink4[7] , \ScanLink58[4] , \ScanLink25[25] , \wAIn28[24] , 
        \wBIn29[0] , \wRegInB31[15] , \ScanLink50[15] , \ScanLink45[21] , 
        \ScanLink30[11] , \ScanLink24[2] , \ScanLink13[20] , \wRegInB12[24] , 
        \wRegInB24[21] , \wBIn0[10] , \wAMid9[25] , \wAMid26[31] , 
        \wAMid26[28] , \wAIn28[7] , \ScanLink27[1] , \wRegInB24[12] , 
        \wAIn28[17] , \wRegInB31[26] , \wRegInB12[17] , \ScanLink50[26] , 
        \ScanLink45[12] , \ScanLink30[22] , \ScanLink13[13] , \ScanLink40[6] , 
        \wRegInA5[19] , \ScanLink25[16] , \wRegInA0[22] , \wRegInA0[11] , 
        \wBIn4[21] , \ScanLink43[5] , \ScanLink2[9] , \wBIn4[12] , \wAMid8[1] , 
        \wAIn9[10] , \wAMid22[19] , \wBMid26[6] , \wRegInA1[31] , 
        \wRegInA1[28] , \wRegInB7[2] , \wRegInA27[7] , \wRegInA28[24] , 
        \wBMid28[13] , \wRegInB4[1] , \wRegInB20[23] , \wRegInB16[26] , 
        \wRegInA24[4] , \ScanLink64[0] , \ScanLink41[23] , \ScanLink34[13] , 
        \ScanLink17[22] , \ScanLink62[12] , \wBMid9[6] , \wBMid25[5] , 
        \ScanLink54[17] , \ScanLink21[27] , \wRegInB23[6] , \wRegInA28[17] , 
        \wBIn5[0] , \wBIn6[3] , \wBMid7[13] , \wAIn9[23] , \wBIn10[9] , 
        \wBMid28[20] , \ScanLink54[24] , \ScanLink41[10] , \ScanLink21[14] , 
        \ScanLink34[20] , \wRegInB16[15] , \wRegInB20[5] , \ScanLink62[21] , 
        \ScanLink17[11] , \wAIn14[3] , \wBMid20[8] , \wAMid28[1] , 
        \wRegInB20[10] , \wBMid15[30] , \wRegInA21[9] , \wBMid15[29] , 
        \wBIn10[24] , \wBIn15[4] , \wAIn17[0] , \wAIn27[19] , \wBIn26[21] , 
        \wAMid29[26] , \wRegInB25[8] , \ScanLink18[6] , \wAMid6[18] , 
        \wBMid7[20] , \wBIn10[17] , \wBIn26[12] , \wAMid30[3] , 
        \wRegInA23[31] , \wRegInA23[28] , \wAMid29[15] , \wBMid4[3] , 
        \wAIn8[30] , \wAMid15[25] , \wBIn16[7] , \wAMid23[20] , \wAIn8[29] , 
        \wBMid7[0] , \wAMid25[4] , \wRegInB6[14] , \wBIn5[18] , \wAMid26[7] , 
        \wAMid5[4] , \wAMid6[7] , \wBMid29[19] , \ScanLink63[18] , 
        \ScanLink16[28] , \ScanLink4[15] , \wRegInB9[4] , \wRegInA29[1] , 
        \ScanLink40[30] , \ScanLink40[29] , \ScanLink35[19] , \ScanLink16[31] , 
        \wRegInB21[29] , \wAMid15[16] , \wAMid23[13] , \wRegInB21[30] , 
        \wBMid28[0] , \ScanLink4[26] , \wAMid0[9] , \wAIn3[25] , \wAIn3[16] , 
        \wAMid7[12] , \wBMid22[15] , \wRegInB6[27] , \wBMid14[10] , 
        \wAMid7[21] , \wBIn8[5] , \wAIn10[25] , \wAIn26[20] , \wBIn27[18] , 
        \ScanLink16[0] , \wAIn10[16] , \wBIn18[1] , \wAMid20[9] , 
        \wRegInA22[22] , \ScanLink15[3] , \wRegInA14[27] , \ScanEnable[0] , 
        \wAIn26[13] , \wBMid14[23] , \wAIn1[7] , \wBMid2[31] , \wAMid3[10] , 
        \wAIn7[9] , \wBMid6[19] , \wBMid22[26] , \wBMid14[4] , \wAIn19[6] , 
        \wBMid30[2] , \wRegInA14[14] , \wRegInA31[3] , \wRegInA22[11] , 
        \wRegInA5[0] , \wRegInB9[30] , \wRegInB9[29] , \wRegInA15[5] , 
        \ScanLink9[2] , \wRegInA10[25] , \wAIn14[27] , \wBMid17[7] , 
        \wAIn22[22] , \wRegInA26[20] , \ScanLink55[1] , \wRegInB18[22] , 
        \ScanLink56[2] , \wAIn7[14] , \wBMid10[12] , \wRegInA16[6] , 
        \wRegInA6[3] , \wBMid2[28] , \wBMid26[17] , \ScanLink19[26] , 
        \wAMid3[23] , \wBMid10[21] , \wAMid19[0] , \wBIn21[8] , 
        \wRegInA10[16] , \wRegInA26[13] , \ScanLink31[5] , \wBMid26[24] , 
        \wRegInB11[4] , \ScanLink19[15] , \wAIn7[27] , \wRegInB12[7] , 
        \wAIn14[14] , \wBIn23[30] , \wAIn22[11] , \wBIn23[29] , 
        \wRegInB18[11] , \ScanLink32[6] , \wAIn26[1] , \ScanLink0[17] , 
        \wRegInA4[13] , \wAIn2[4] , \wRegInB2[16] , \ScanLink31[31] , 
        \ScanLink12[19] , \wBMid9[17] , \wBMid11[9] , \wAIn25[2] , 
        \ScanLink44[18] , \wRegInB25[18] , \ScanLink31[28] , \wBIn1[30] , 
        \wAMid11[27] , \wAMid27[22] , \wRegInA10[8] , \wBIn28[25] , 
        \wRegInB2[25] , \wBIn1[29] , \wAMid11[14] , \wBIn24[5] , \wBIn27[6] , 
        \wRegInA4[20] , \ScanLink0[24] , \wRegInB14[9] , \wRegInA0[18] , 
        \wAMid0[0] , \wBMid6[10] , \wBMid9[24] , \wAMid27[11] , \wBIn28[16] , 
        \ScanLink29[7] , \wBIn11[27] , \wBIn27[22] , \ScanLink34[8] , 
        \wAMid28[25] , \wAMid7[28] , \wBMid1[7] , \wAMid3[3] , \wAMid7[31] , 
        \wBMid6[23] , \wBMid14[19] , \wRegInA22[18] , \wBIn11[14] , 
        \wAMid23[3] , \wAIn26[29] , \wAIn26[30] , \wBMid2[4] , \wBIn18[8] , 
        \wAMid20[0] , \wBIn27[11] , \wAMid28[16] , \ScanLink16[9] , 
        \wBIn5[22] , \wAIn8[13] , \wRegInB28[4] , \wRegInA29[8] , 
        \ScanLink55[14] , \ScanLink20[24] , \wBMid28[9] , \wBMid29[10] , 
        \ScanLink16[21] , \wRegInB17[25] , \ScanLink63[11] , \ScanLink40[20] , 
        \ScanLink35[10] , \wRegInB21[20] , \wRegInA29[27] , \wAIn8[20] , 
        \wBMid7[9] , \wAMid23[30] , \wRegInB21[13] , \wAMid23[29] , 
        \wBMid29[23] , \wRegInB17[16] , \wRegInB30[6] , \ScanLink63[22] , 
        \ScanLink55[27] , \ScanLink40[13] , \ScanLink16[12] , \ScanLink35[23] , 
        \ScanLink20[17] , \ScanLink10[7] , \wBIn1[20] , \wBIn5[11] , 
        \wRegInA4[30] , \wRegInA29[14] , \ScanLink13[4] , \ScanLink37[2] , 
        \wRegInA4[29] , \wRegInB14[0] , \wRegInB17[3] , \wBIn0[19] , 
        \wRegInA0[4] , \wBIn1[13] , \wAMid8[15] , \wAMid27[18] , 
        \wRegInB25[22] , \wAIn29[27] , \wRegInB13[27] , \wRegInB30[16] , 
        \ScanLink44[22] , \ScanLink31[12] , \ScanLink12[23] , \ScanLink34[1] , 
        \ScanLink24[26] , \wBMid12[3] , \wAIn26[8] , \wRegInA3[7] , 
        \wRegInA13[2] , \ScanLink51[16] , \ScanLink53[6] , \wAMid8[26] , 
        \ScanLink51[25] , \ScanLink50[5] , \wBMid11[0] , \ScanLink24[15] , 
        \ScanLink12[10] , \wAIn29[14] , \wRegInB13[14] , \ScanLink44[11] , 
        \ScanLink31[21] , \wRegInB30[25] , \wBMid2[21] , \wBMid2[12] , 
        \wBMid10[31] , \wBMid10[28] , \wAMid19[9] , \wBIn21[1] , 
        \wRegInB9[13] , \wRegInA10[1] , \wRegInB25[11] , \wAIn4[3] , 
        \wAIn7[0] , \wBIn15[25] , \wAIn22[18] , \wBIn22[2] , \wRegInB18[18] , 
        \wBIn23[20] , \wRegInA5[9] , \ScanLink48[7] , \wRegInB9[20] , 
        \wRegInA26[30] , \wRegInA26[29] , \ScanLink55[8] , \wBIn15[16] , 
        \wAIn20[6] , \wAIn23[5] , \wBIn23[13] , \wAMid3[19] , \wBMid8[14] , 
        \wAMid10[24] , \wAMid26[21] , \wBIn29[26] , \ScanLink1[3] , 
        \wRegInB3[15] , \wRegInA5[10] , \ScanLink2[0] , \wAMid2[13] , 
        \wAIn6[17] , \wBMid8[27] , \ScanLink1[14] , \wAMid10[17] , 
        \wAMid11[1] , \wRegInB19[5] , \ScanLink45[28] , \ScanLink30[18] , 
        \ScanLink13[30] , \ScanLink13[29] , \ScanLink45[31] , \wAMid26[12] , 
        \wBIn29[9] , \wBIn29[15] , \wRegInB24[31] , \ScanLink39[4] , 
        \wRegInB24[28] , \wAMid12[2] , \wRegInB3[26] , \wRegInA5[23] , 
        \ScanLink1[27] , \ScanLink27[8] , \wBMid27[14] , \ScanLink18[25] , 
        \wAIn9[6] , \wBMid11[11] , \wAIn15[24] , \wBIn22[19] , \ScanLink46[1] , 
        \wAIn23[21] , \wRegInB19[21] , \wBIn0[31] , \wBIn0[28] , \wBIn0[4] , 
        \wAIn2[26] , \wAIn2[15] , \wAMid2[20] , \wAIn6[24] , \wAIn15[17] , 
        \wBMid19[8] , \wRegInA11[26] , \wRegInA18[9] , \wRegInA27[23] , 
        \ScanLink45[2] , \wAIn23[12] , \wRegInB19[12] , \ScanLink22[5] , 
        \wBMid11[22] , \wBMid3[18] , \wAIn11[26] , \wAIn27[23] , \wBMid27[27] , 
        \wRegInB8[19] , \ScanLink18[16] , \wRegInA11[15] , \ScanLink21[6] , 
        \wRegInA15[24] , \wRegInB25[1] , \wRegInA27[10] , \wRegInA23[21] , 
        \wBIn5[9] , \wAMid6[11] , \wBMid7[30] , \wBMid7[29] , \wBMid15[13] , 
        \wBMid20[1] , \wBMid23[16] , \wRegInB26[2] , \wBMid23[25] , 
        \wRegInB1[5] , \wRegInA15[17] , \wRegInA23[12] , \ScanLink61[4] , 
        \wRegInA21[0] , \wRegInA22[3] , \wRegInB2[6] , \wAMid6[22] , 
        \wBMid15[20] , \wAIn11[15] , \wAIn17[9] , \wBIn26[28] , \wBIn13[3] , 
        \wBMid23[2] , \wBIn26[31] , \wAIn27[10] , \ScanLink62[7] , \wBIn3[7] , 
        \wBMid28[30] , \wRegInA1[12] , \ScanLink5[16] , \wRegInB7[17] , 
        \ScanLink62[31] , \ScanLink41[19] , \wBMid28[29] , \ScanLink62[28] , 
        \ScanLink34[29] , \ScanLink34[30] , \ScanLink17[18] , \wBIn4[31] , 
        \wBIn4[28] , \wBIn10[0] , \wAMid22[23] , \wAIn12[4] , \wAMid14[26] , 
        \wAMid28[8] , \wRegInB20[19] , \wRegInB7[24] , \wAMid8[8] , 
        \wRegInA1[21] , \wAIn9[19] , \wAMid14[15] , \ScanLink5[25] , 
        \wAMid22[10] , \wRegInB4[8] , \wBMid8[16] , \wAIn11[7] , 
        \wRegInB3[17] , \wRegInA5[12] , \ScanLink64[9] , \ScanLink1[16] , 
        \ScanLink30[29] , \ScanLink2[2] , \wAMid10[26] , \wAMid26[23] , 
        \wBIn29[24] , \ScanLink45[19] , \ScanLink30[30] , \ScanLink13[18] , 
        \ScanLink1[1] , \wRegInB24[19] , \wAMid12[0] , \wRegInB3[24] , 
        \wRegInA5[21] , \wBIn0[6] , \wAIn2[24] , \wAIn2[17] , \wAMid2[22] , 
        \wAMid2[11] , \wAIn6[15] , \wAIn9[4] , \wBMid8[25] , \wAMid10[15] , 
        \ScanLink1[25] , \wAMid11[3] , \wAMid26[10] , \wBIn29[17] , 
        \ScanLink39[6] , \ScanLink24[9] , \wAIn15[26] , \wAIn23[23] , 
        \wRegInB8[31] , \wRegInB8[28] , \wRegInB19[7] , \wRegInA11[24] , 
        \wRegInB19[23] , \wRegInA27[21] , \ScanLink45[0] , \ScanLink46[3] , 
        \wBMid11[13] , \wBMid3[30] , \wBMid3[29] , \wBMid27[16] , 
        \ScanLink18[27] , \wAIn6[26] , \wBMid27[25] , \wBIn31[9] , 
        \wRegInA11[17] , \wRegInA27[12] , \ScanLink21[4] , \ScanLink18[14] , 
        \wBMid11[20] , \wAIn15[15] , \wBIn22[28] , \wBIn22[31] , \wAIn23[10] , 
        \wBMid23[14] , \wRegInB19[10] , \ScanLink22[7] , \wRegInB26[0] , 
        \wBIn6[8] , \wAMid6[13] , \wBMid15[11] , \wAIn11[24] , \wBIn26[19] , 
        \wAIn27[21] , \wAMid30[8] , \wRegInA15[26] , \wRegInA23[23] , 
        \wRegInB25[3] , \wAIn11[17] , \wBMid23[0] , \wAIn27[12] , 
        \ScanLink62[5] , \wBIn3[5] , \wAMid6[20] , \wBMid7[18] , \wBMid15[22] , 
        \wAIn14[8] , \wBMid20[3] , \wBMid23[27] , \wRegInA22[1] , 
        \wRegInB1[7] , \wRegInB2[4] , \wRegInA15[15] , \wRegInA21[2] , 
        \ScanLink61[6] , \wAMid14[24] , \wRegInA23[10] , \wAMid22[21] , 
        \wBIn4[19] , \wAIn9[31] , \wAIn9[28] , \wBIn10[2] , \wRegInB7[15] , 
        \wBIn13[1] , \wRegInA1[10] , \ScanLink5[14] , \wRegInA0[30] , 
        \wAMid0[2] , \wAMid3[1] , \wAIn11[5] , \wBMid28[18] , \ScanLink41[31] , 
        \ScanLink41[28] , \ScanLink34[18] , \ScanLink17[30] , \ScanLink62[19] , 
        \ScanLink17[29] , \wAIn12[6] , \wAMid14[17] , \wAMid22[12] , 
        \wRegInB20[31] , \wRegInB20[28] , \wRegInA1[23] , \wRegInB7[9] , 
        \ScanLink5[27] , \wRegInB7[26] , \wBMid30[9] , \wBMid14[28] , 
        \wRegInA31[8] , \wBMid1[5] , \wBMid2[6] , \wBMid6[12] , \wBMid14[31] , 
        \wBIn11[25] , \wAIn26[18] , \wBIn27[20] , \wAMid28[27] , 
        \wRegInA22[30] , \wRegInA22[29] , \ScanLink15[8] , \wAMid20[2] , 
        \wRegInB28[6] , \wBMid6[21] , \wBIn11[16] , \wBIn27[13] , 
        \wAMid28[14] , \wAMid23[1] , \wAMid7[19] , \wRegInA0[29] , 
        \wRegInA0[6] , \wBIn1[22] , \wBIn5[20] , \wBIn5[13] , \wBMid4[8] , 
        \wAIn8[11] , \wAMid23[18] , \wRegInB21[22] , \wRegInA29[25] , 
        \wBMid29[12] , \wRegInB17[27] , \ScanLink63[13] , \ScanLink55[16] , 
        \ScanLink40[22] , \ScanLink16[23] , \ScanLink35[12] , \ScanLink20[26] , 
        \wRegInA29[16] , \ScanLink13[6] , \wAIn8[22] , \ScanLink55[25] , 
        \ScanLink20[15] , \ScanLink10[5] , \wAMid8[17] , \wBMid29[21] , 
        \ScanLink63[20] , \ScanLink16[10] , \wRegInB17[14] , \ScanLink40[11] , 
        \ScanLink35[21] , \wRegInB21[11] , \wRegInB30[4] , \ScanLink51[14] , 
        \wAIn29[25] , \wRegInB13[25] , \ScanLink44[20] , \ScanLink24[24] , 
        \ScanLink12[21] , \ScanLink34[3] , \ScanLink31[10] , \wRegInB14[2] , 
        \wRegInB25[20] , \wRegInB30[14] , \wRegInB17[1] , \ScanLink37[0] , 
        \wAMid27[30] , \wRegInB25[13] , \wAMid27[29] , \wRegInA10[3] , 
        \wRegInA0[20] , \wRegInA0[13] , \wBIn1[11] , \wAMid8[24] , 
        \wBMid11[2] , \wAIn29[16] , \wRegInB13[16] , \wRegInB30[27] , 
        \ScanLink12[12] , \wAIn25[9] , \ScanLink31[23] , \ScanLink50[7] , 
        \ScanLink44[13] , \ScanLink24[17] , \ScanLink51[27] , \wBMid2[23] , 
        \wBMid2[10] , \wBMid12[1] , \wBIn15[27] , \wBIn23[22] , \wRegInA3[5] , 
        \wRegInA4[18] , \wRegInA13[0] , \ScanLink53[4] , \wBIn22[0] , 
        \wAMid3[31] , \wAMid3[28] , \wBMid10[19] , \wBIn21[3] , \wRegInB9[11] , 
        \wRegInA26[18] , \wRegInA6[8] , \wAIn4[1] , \wAIn22[29] , \wAIn23[7] , 
        \wRegInB18[29] , \wAIn7[2] , \wBIn15[14] , \wAIn22[30] , 
        \wRegInB18[30] , \wBIn23[11] , \ScanLink56[9] , \wAIn20[4] , 
        \wAMid26[5] , \wRegInB9[22] , \ScanLink48[5] , \ScanLink9[9] , 
        \ScanLink4[17] , \wBIn5[30] , \wBMid4[1] , \wBMid7[2] , \wAMid25[6] , 
        \wBMid29[28] , \wRegInB6[16] , \ScanLink35[31] , \ScanLink16[19] , 
        \ScanLink63[29] , \wBMid29[31] , \ScanLink35[28] , \ScanLink63[30] , 
        \ScanLink40[18] , \wAMid15[27] , \wAMid23[22] , \wRegInB21[18] , 
        \wRegInB6[25] , \wAIn3[27] , \wAIn3[14] , \wBIn5[29] , \wAMid5[6] , 
        \ScanLink4[24] , \wAMid6[5] , \wAMid15[14] , \wBMid28[2] , 
        \wAMid7[10] , \wAIn8[18] , \wAMid23[11] , \wRegInA29[3] , \wBIn8[7] , 
        \wBIn18[3] , \wRegInB9[6] , \wRegInA14[25] , \wRegInA22[20] , 
        \ScanLink15[1] , \wAIn10[27] , \wAMid23[8] , \wAIn26[22] , 
        \wBMid14[12] , \ScanLink16[2] , \wAMid3[8] , \wBMid6[31] , 
        \wBMid22[17] , \wBMid6[28] , \wAIn19[4] , \wBMid30[0] , 
        \wRegInA22[13] , \wRegInA14[16] , \wRegInA31[1] , \wAMid7[23] , 
        \wBMid22[24] , \wBMid14[21] , \wBMid2[19] , \wAMid3[21] , \wAMid3[12] , 
        \wAIn10[14] , \wBIn27[30] , \wBMid10[10] , \wAIn26[11] , \wBIn27[29] , 
        \wBMid26[15] , \ScanLink19[24] , \wRegInA16[4] , \wAIn4[8] , 
        \wAIn7[16] , \wAIn14[25] , \wRegInA6[1] , \wAIn22[20] , \wBIn23[18] , 
        \ScanLink56[0] , \wRegInB18[20] , \wAIn14[16] , \wBMid14[6] , 
        \wBMid17[5] , \wRegInA10[27] , \wRegInA26[22] , \ScanLink55[3] , 
        \wAIn22[13] , \wRegInA5[2] , \ScanLink9[0] , \wRegInA15[7] , 
        \wRegInB18[13] , \ScanLink32[4] , \wAIn7[25] , \wBMid10[23] , 
        \wBMid26[26] , \wRegInB12[5] , \ScanLink19[17] , \wAMid11[25] , 
        \wAMid19[2] , \wBIn22[9] , \wRegInB9[18] , \wRegInB11[6] , 
        \wRegInA10[14] , \wRegInA26[11] , \ScanLink31[7] , \wAIn1[5] , 
        \wBIn1[18] , \wAIn2[6] , \wAMid27[20] , \wBIn28[27] , \wBMid9[15] , 
        \wBMid12[8] , \wAIn25[0] , \wAIn26[3] , \wRegInB2[14] , \wBMid9[26] , 
        \wRegInA4[11] , \wRegInA13[9] , \ScanLink0[15] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink12[28] , \ScanLink31[19] , \ScanLink12[31] , 
        \wBMid3[13] , \wAMid11[16] , \wBIn24[7] , \wAMid27[13] , \wBIn28[14] , 
        \wRegInB25[30] , \wRegInB25[29] , \ScanLink29[5] , \wBMid11[30] , 
        \wAMid14[7] , \wBIn27[4] , \wRegInB17[8] , \ScanLink0[26] , 
        \wRegInB2[27] , \wRegInA4[22] , \ScanLink37[9] , \wBIn31[0] , 
        \wRegInB8[12] , \wBMid11[29] , \wBIn14[24] , \wAMid17[4] , 
        \wBIn22[21] , \wAIn23[19] , \wRegInB19[19] , \wBMid19[3] , 
        \wRegInB8[21] , \ScanLink58[6] , \wRegInA27[31] , \wBIn0[21] , 
        \wAMid2[18] , \wBMid3[20] , \wBIn14[17] , \wBIn22[12] , \wAIn30[7] , 
        \wRegInA18[2] , \wRegInA27[28] , \ScanLink4[5] , \ScanLink45[9] , 
        \wRegInA8[7] , \ScanLink7[6] , \wRegInA5[28] , \wBIn0[12] , 
        \wAMid9[14] , \wAMid12[9] , \wRegInA5[31] , \ScanLink27[3] , 
        \wAMid26[19] , \wAIn28[26] , \wRegInB31[17] , \wRegInB24[23] , 
        \wRegInB12[26] , \wBIn29[2] , \ScanLink45[23] , \ScanLink30[13] , 
        \ScanLink24[0] , \ScanLink13[22] , \ScanLink50[17] , \ScanLink43[7] , 
        \ScanLink25[27] , \wRegInA0[2] , \wAIn1[8] , \wBIn1[26] , \wBMid2[27] , 
        \wBMid2[14] , \wBIn4[23] , \wAMid8[3] , \wAIn9[12] , \wAMid9[27] , 
        \ScanLink40[4] , \ScanLink1[8] , \ScanLink25[14] , \wBMid25[7] , 
        \wAIn28[15] , \wRegInB31[24] , \ScanLink50[24] , \ScanLink45[10] , 
        \ScanLink30[20] , \ScanLink13[11] , \wAIn28[5] , \wRegInB12[15] , 
        \wRegInB24[10] , \wBMid26[4] , \wBMid28[11] , \ScanLink64[2] , 
        \ScanLink54[15] , \ScanLink41[21] , \ScanLink21[25] , \ScanLink62[10] , 
        \ScanLink34[11] , \wRegInB4[3] , \ScanLink17[20] , \wRegInB7[0] , 
        \wRegInB16[24] , \wRegInB20[21] , \wRegInA24[6] , \wRegInA27[5] , 
        \wRegInA28[26] , \wBIn4[10] , \wAIn9[21] , \wAMid22[31] , 
        \wAMid22[28] , \wAMid28[3] , \wBMid28[22] , \wRegInB16[17] , 
        \wRegInB20[12] , \wRegInB20[7] , \ScanLink62[23] , \ScanLink41[12] , 
        \ScanLink34[22] , \ScanLink17[13] , \ScanLink54[26] , \ScanLink21[16] , 
        \wBIn5[2] , \wAMid6[30] , \wBMid7[11] , \wBIn10[26] , \wBMid9[4] , 
        \wBIn13[8] , \wRegInA1[19] , \wRegInA28[15] , \wAIn17[2] , 
        \wBIn26[23] , \wAMid29[24] , \wRegInB23[4] , \wBMid23[9] , 
        \wRegInA22[8] , \wAMid6[29] , \wAIn14[1] , \wRegInA23[19] , \wBIn6[1] , 
        \wBMid7[22] , \wBIn16[5] , \wBMid15[18] , \wBIn10[15] , \wRegInB26[9] , 
        \wBIn15[6] , \wBIn26[10] , \wAIn27[31] , \wAIn27[28] , \wAMid29[17] , 
        \wAMid30[1] , \wAIn7[31] , \wAIn7[28] , \wBIn21[7] , \wRegInB9[15] , 
        \wRegInA10[19] , \ScanLink18[4] , \wRegInB12[8] , \wBIn22[4] , 
        \wAIn4[5] , \wAIn7[6] , \wBIn15[23] , \wAIn20[0] , \wBIn23[26] , 
        \ScanLink32[9] , \wRegInB9[26] , \ScanLink48[1] , \wAIn14[31] , 
        \wAIn14[28] , \wBIn23[15] , \wBIn15[10] , \wBMid17[8] , \wAIn23[3] , 
        \wBMid26[18] , \ScanLink19[30] , \wRegInA16[9] , \ScanLink19[29] , 
        \wBIn1[15] , \wAMid8[13] , \wBIn27[9] , \wRegInB17[5] , 
        \ScanLink37[4] , \wBIn28[19] , \ScanLink29[8] , \wAIn29[21] , 
        \wRegInB13[21] , \wRegInB14[6] , \wRegInB25[24] , \wRegInB30[10] , 
        \ScanLink51[10] , \ScanLink44[24] , \ScanLink34[7] , \ScanLink31[14] , 
        \ScanLink12[25] , \wRegInB2[19] , \wRegInA3[1] , \ScanLink24[20] , 
        \ScanLink0[18] , \wRegInA13[4] , \ScanLink53[0] , \wBMid12[5] , 
        \wAMid8[20] , \ScanLink50[3] , \ScanLink24[13] , \wBMid9[18] , 
        \ScanLink51[23] , \ScanLink31[27] , \wAMid11[31] , \wAMid11[28] , 
        \wBMid11[6] , \ScanLink44[17] , \ScanLink12[16] , \wAIn29[12] , 
        \wRegInB30[23] , \wRegInA10[7] , \wRegInB13[12] , \wBIn5[24] , 
        \wAMid6[8] , \wAIn8[15] , \wRegInB25[17] , \wAMid15[19] , 
        \wBMid29[16] , \ScanLink55[12] , \ScanLink40[26] , \ScanLink20[22] , 
        \ScanLink35[16] , \ScanLink63[17] , \ScanLink16[27] , \wRegInB17[23] , 
        \wRegInB21[26] , \wRegInB6[31] , \wRegInB6[28] , \wRegInA29[21] , 
        \ScanLink4[30] , \ScanLink4[29] , \wBIn5[17] , \wAIn8[26] , 
        \wBMid29[25] , \wRegInB17[10] , \wRegInB21[15] , \wRegInB30[0] , 
        \ScanLink40[15] , \ScanLink35[25] , \ScanLink16[14] , \ScanLink63[24] , 
        \ScanLink55[21] , \ScanLink20[11] , \ScanLink10[1] , \wAMid26[8] , 
        \ScanLink13[2] , \wBIn0[25] , \wBIn0[2] , \wAMid0[6] , \wBMid6[16] , 
        \wAIn10[19] , \wBIn27[24] , \wRegInA29[12] , \wAMid28[23] , 
        \wBIn11[21] , \wBMid22[30] , \wBMid22[29] , \wBMid1[1] , \wAIn3[19] , 
        \wAMid3[5] , \wAIn19[9] , \wBMid6[25] , \wBIn11[12] , \wAMid23[5] , 
        \wBIn27[17] , \wAMid28[10] , \wBMid2[2] , \wAMid20[6] , 
        \wRegInA14[31] , \wRegInA14[28] , \wBIn13[5] , \wRegInB28[2] , 
        \wAIn2[30] , \wAIn2[20] , \wAIn2[13] , \wBIn3[1] , \wBMid9[9] , 
        \wRegInA28[18] , \ScanLink5[10] , \wRegInA1[14] , \wRegInB23[9] , 
        \wRegInB7[11] , \wAMid6[17] , \wBIn10[18] , \wBIn10[6] , \wAMid22[25] , 
        \wAIn11[1] , \wAIn12[2] , \wAMid14[20] , \wBMid26[9] , \wRegInB7[22] , 
        \wAMid14[13] , \wRegInA1[27] , \wRegInB16[30] , \wRegInB16[29] , 
        \wRegInA27[8] , \ScanLink5[23] , \wAMid22[16] , \ScanLink54[18] , 
        \ScanLink21[28] , \wAIn27[25] , \wRegInA15[22] , \wRegInB25[7] , 
        \ScanLink21[31] , \ScanLink18[9] , \wRegInA23[27] , \wAIn11[20] , 
        \wBIn16[8] , \wBMid15[15] , \wAMid6[24] , \wBMid20[7] , \wBMid23[10] , 
        \wRegInA23[14] , \wRegInB26[4] , \wBMid23[23] , \wRegInB1[3] , 
        \wRegInA15[11] , \wRegInA21[6] , \ScanLink61[2] , \wRegInB2[0] , 
        \wRegInA22[5] , \wBMid15[26] , \wAMid2[26] , \wAMid2[15] , 
        \wAIn11[13] , \wBMid11[17] , \wBMid23[4] , \wAMid29[30] , \wAIn27[16] , 
        \wAMid29[29] , \wBMid27[12] , \ScanLink62[1] , \ScanLink18[23] , 
        \wAIn6[11] , \wAIn9[0] , \wBIn14[30] , \wAIn15[22] , \wAIn23[27] , 
        \wRegInB19[27] , \ScanLink46[7] , \wAIn23[14] , \wRegInA11[20] , 
        \wRegInA27[25] , \ScanLink45[4] , \ScanLink4[8] , \wBIn14[29] , 
        \wRegInB19[14] , \ScanLink22[3] , \wAIn15[11] , \wAMid17[9] , 
        \wAIn6[22] , \wBMid11[24] , \wBMid8[21] , \wBMid8[12] , \wAMid10[22] , 
        \wAIn28[18] , \wBMid27[21] , \ScanLink18[10] , \wRegInA11[13] , 
        \wRegInA27[16] , \ScanLink21[0] , \wRegInB31[30] , \wRegInB12[18] , 
        \wAMid26[27] , \wRegInB31[29] , \wAIn28[8] , \wBIn29[20] , 
        \ScanLink50[30] , \ScanLink50[29] , \ScanLink40[9] , \ScanLink25[19] , 
        \ScanLink1[5] , \wRegInB3[13] , \ScanLink2[6] , \wRegInA5[16] , 
        \wRegInB19[3] , \ScanLink1[12] , \wAMid9[19] , \wAMid10[11] , 
        \wAMid11[7] , \wAMid26[14] , \ScanLink39[2] , \wBIn29[13] , 
        \wAMid12[4] , \wRegInA5[25] , \ScanLink1[21] , \wAIn14[5] , 
        \wRegInB3[20] , \wRegInA15[18] , \wAIn2[29] , \wBIn3[8] , \wBIn4[27] , 
        \wBIn5[6] , \wBIn6[5] , \wBMid7[15] , \wRegInB2[9] , \wBIn10[22] , 
        \ScanLink62[8] , \wBIn15[2] , \wAIn17[6] , \wBIn26[27] , \wAMid29[20] , 
        \ScanLink18[0] , \wBMid7[26] , \wBIn10[11] , \wAIn11[30] , 
        \wAIn11[29] , \wAMid30[5] , \wBIn26[14] , \wAMid29[13] , \wBMid23[19] , 
        \wAMid8[7] , \wBIn16[1] , \wBIn4[14] , \wAIn9[16] , \wAIn11[8] , 
        \wBMid26[0] , \wBMid28[15] , \wRegInB4[7] , \wRegInB7[4] , 
        \wRegInA28[22] , \wRegInB16[20] , \wRegInB20[25] , \wRegInA27[1] , 
        \wRegInA24[2] , \ScanLink64[6] , \ScanLink62[14] , \ScanLink41[25] , 
        \ScanLink17[24] , \ScanLink54[11] , \ScanLink34[15] , \wBMid25[3] , 
        \ScanLink21[21] , \wBMid9[0] , \ScanLink5[19] , \wRegInB7[18] , 
        \wRegInB23[0] , \wRegInA28[11] , \wAIn9[25] , \ScanLink54[22] , 
        \ScanLink21[12] , \wAMid14[30] , \wBMid28[26] , \ScanLink17[17] , 
        \ScanLink62[27] , \ScanLink41[16] , \ScanLink34[26] , \wAMid14[29] , 
        \wRegInB16[13] , \wAMid28[7] , \wRegInB20[3] , \wRegInB20[16] , 
        \wBMid8[31] , \wAMid9[10] , \wBIn29[6] , \ScanLink50[13] , 
        \ScanLink25[23] , \wBMid8[28] , \ScanLink45[27] , \ScanLink13[26] , 
        \ScanLink30[17] , \ScanLink24[4] , \wAMid10[18] , \wAIn28[22] , 
        \wRegInB12[22] , \wRegInB31[13] , \wRegInB3[30] , \wRegInB24[27] , 
        \ScanLink1[31] , \ScanLink1[28] , \wRegInB3[29] , \ScanLink27[7] , 
        \wBIn0[16] , \wAMid9[23] , \wAIn28[11] , \wAIn28[1] , \wBIn29[30] , 
        \wBIn29[29] , \wRegInB24[14] , \wRegInB31[20] , \wRegInB12[11] , 
        \ScanLink45[14] , \ScanLink30[24] , \ScanLink13[15] , \ScanLink40[0] , 
        \ScanLink25[10] , \ScanLink50[20] , \wBMid3[24] , \wBMid3[17] , 
        \wBIn14[20] , \wAIn15[18] , \ScanLink43[3] , \wAMid17[0] , 
        \wBIn22[25] , \wBMid27[28] , \ScanLink18[19] , \wAIn6[18] , \wAIn9[9] , 
        \wAMid14[3] , \wBMid27[31] , \wBIn31[4] , \wRegInB8[16] , 
        \ScanLink21[9] , \wBIn14[13] , \wBIn22[16] , \ScanLink7[2] , 
        \wAIn30[3] , \wRegInA8[3] , \wRegInA11[29] , \wRegInA11[30] , 
        \wRegInA18[6] , \wAIn1[1] , \wBMid19[7] , \ScanLink4[1] , 
        \wRegInA3[8] , \wRegInB8[25] , \ScanLink58[2] , \ScanLink0[11] , 
        \wAIn2[2] , \wBMid9[11] , \wAIn26[7] , \wRegInA4[15] , \wRegInB2[10] , 
        \ScanLink53[9] , \wAIn25[4] , \wAMid8[30] , \wAMid8[29] , 
        \wAMid27[24] , \wBIn28[23] , \wAMid11[21] , \wAMid11[12] , \wBIn27[0] , 
        \wRegInB2[23] , \wRegInA4[26] , \wRegInB13[31] , \wRegInB30[19] , 
        \ScanLink0[22] , \wBIn24[3] , \wAIn29[31] , \wAMid27[17] , 
        \wAIn29[28] , \wRegInB13[28] , \ScanLink29[1] , \wBIn28[10] , 
        \wRegInA0[24] , \wRegInA0[17] , \wBMid1[8] , \wAIn3[10] , \wAMid3[25] , 
        \wAMid3[16] , \wAIn7[12] , \wBMid9[22] , \ScanLink51[19] , 
        \ScanLink24[30] , \ScanLink24[29] , \wAIn14[21] , \wBIn15[19] , 
        \wBMid14[2] , \wAIn20[9] , \wRegInA5[6] , \wRegInA15[3] , 
        \ScanLink48[8] , \ScanLink9[4] , \wBMid17[1] , \wRegInA10[23] , 
        \wRegInA26[26] , \ScanLink55[7] , \wAIn22[24] , \wRegInB18[24] , 
        \ScanLink56[4] , \wBMid10[14] , \wRegInA6[5] , \wRegInA16[0] , 
        \wAIn7[21] , \wAMid19[6] , \wBMid26[11] , \wRegInA10[10] , 
        \wRegInA26[15] , \ScanLink19[20] , \ScanLink31[3] , \wBMid26[22] , 
        \wRegInB11[2] , \ScanLink19[13] , \wRegInB12[1] , \wBMid10[27] , 
        \wAIn14[12] , \wAIn22[17] , \wBMid22[13] , \wRegInB18[17] , 
        \ScanLink32[0] , \wAMid7[14] , \wBMid14[16] , \wAIn10[23] , 
        \wAMid28[19] , \ScanLink16[6] , \wAIn3[23] , \wBIn8[3] , \wAIn10[10] , 
        \wBIn11[31] , \wBIn11[28] , \wBIn18[7] , \wAIn26[26] , \wRegInA22[24] , 
        \ScanLink15[5] , \wRegInA14[21] , \wAIn26[15] , \wBMid4[5] , 
        \wAMid7[27] , \wBMid7[6] , \wBMid14[25] , \wAMid15[23] , \wAIn19[0] , 
        \wBMid22[20] , \wBMid30[4] , \wRegInA14[12] , \wRegInA31[5] , 
        \wRegInA22[17] , \wAMid23[26] , \wRegInB17[19] , \wRegInB30[9] , 
        \wAMid25[2] , \ScanLink55[31] , \ScanLink55[28] , \ScanLink20[18] , 
        \ScanLink10[8] , \wRegInB6[12] , \wAMid26[1] , \wAMid5[2] , 
        \wAMid6[1] , \wAMid23[15] , \wRegInB9[2] , \ScanLink4[13] , 
        \wRegInA29[7] , \wAMid15[10] , \wBMid28[6] , \wRegInA29[31] , 
        \wRegInA29[28] , \ScanLink4[20] , \wAIn1[25] , \wBMid0[31] , 
        \wBMid0[28] , \wBMid0[5] , \wRegInA6[20] , \wRegInB6[21] , 
        \wAMid1[23] , \wAMid1[2] , \wBIn3[30] , \wBIn3[29] , \wBMid3[6] , 
        \wAMid13[14] , \wAMid22[1] , \wRegInB0[25] , \wAMid25[11] , 
        \wRegInA19[30] , \wRegInA19[29] , \ScanLink2[24] , \wAMid30[25] , 
        \wRegInB29[6] , \ScanLink14[8] , \wAMid21[2] , \ScanLink2[17] , 
        \wAMid2[1] , \wAMid13[27] , \wRegInB0[16] , \wRegInA6[13] , 
        \ScanLink46[18] , \ScanLink33[28] , \ScanLink33[31] , \ScanLink10[19] , 
        \wAIn5[27] , \wBIn8[16] , \wAMid25[22] , \wAMid30[16] , \wRegInB31[4] , 
        \wRegInA12[16] , \wRegInB27[18] , \wRegInA30[8] , \wRegInA31[27] , 
        \ScanLink11[5] , \wRegInA24[13] , \wBMid5[8] , \wBMid12[21] , 
        \wBMid24[24] , \ScanLink58[20] , \ScanLink38[24] , \wBIn8[25] , 
        \wAIn16[14] , \wAIn20[11] , \ScanLink12[6] , \wBIn21[30] , 
        \wBIn21[29] , \wAIn16[27] , \wRegInA12[25] , \wRegInA24[20] , 
        \wRegInA31[14] , \ScanLink9[31] , \ScanLink9[28] , \wAMid18[18] , 
        \wAIn20[22] , \ScanLink38[17] , \wBMid24[17] , \wAMid1[10] , 
        \wAIn5[14] , \wBMid12[12] , \ScanLink58[13] , \wBMid4[19] , 
        \wAIn12[16] , \wAIn31[27] , \wBMid13[1] , \wAIn24[13] , 
        \wRegInB28[16] , \ScanLink52[4] , \wBMid20[26] , \wRegInA2[5] , 
        \wRegInA12[0] , \ScanLink49[16] , \wAIn1[16] , \wAMid5[21] , 
        \ScanLink29[12] , \wBMid10[2] , \wBMid16[23] , \wRegInA1[6] , 
        \wRegInA11[3] , \wAIn24[9] , \wRegInA20[11] , \wRegInA16[14] , 
        \ScanLink51[7] , \wAIn5[1] , \wAMid5[12] , \wBMid16[10] , \wAIn6[2] , 
        \wAIn12[25] , \wBMid20[15] , \ScanLink49[25] , \ScanLink29[21] , 
        \wAIn24[20] , \wRegInB16[1] , \wBIn25[18] , \ScanLink36[0] , 
        \wAIn31[14] , \wRegInB28[25] , \wRegInB15[2] , \wRegInA16[27] , 
        \wRegInA20[22] , \ScanLink35[3] , \wAMid17[16] , \wAIn21[4] , 
        \ScanLink61[18] , \ScanLink42[29] , \ScanLink37[19] , \ScanLink14[31] , 
        \ScanLink42[30] , \ScanLink14[28] , \wBIn18[11] , \wAIn19[30] , 
        \wAMid21[13] , \wRegInB23[30] , \ScanLink49[5] , \wAIn19[29] , 
        \wRegInB23[29] , \ScanLink8[9] , \wAIn22[7] , \wRegInB4[27] , 
        \wRegInA7[8] , \ScanLink6[26] , \wAMid17[25] , \wBIn20[3] , 
        \wRegInA2[22] , \ScanLink57[9] , \wAMid21[20] , \wBIn18[22] , 
        \wAMid4[18] , \wBIn7[18] , \wAMid10[3] , \wBIn23[0] , \wRegInA2[11] , 
        \wRegInB4[14] , \wRegInA8[24] , \ScanLink38[6] , \ScanLink6[15] , 
        \wBIn12[17] , \wAMid13[0] , \wBIn31[26] , \wRegInB18[7] , 
        \wRegInA21[31] , \wRegInA21[28] , \ScanLink25[9] , \wBIn24[12] , 
        \wBIn6[21] , \wBIn6[12] , \wBMid5[20] , \wBMid5[13] , \wRegInA8[17] , 
        \ScanLink0[1] , \wBIn12[24] , \wBMid17[30] , \wBMid17[29] , 
        \ScanLink28[18] , \wBIn24[21] , \wAIn25[19] , \wBIn31[15] , 
        \ScanLink3[2] , \wAIn18[10] , \ScanLink60[21] , \ScanLink23[7] , 
        \ScanLink15[11] , \ScanLink56[24] , \ScanLink43[10] , \ScanLink36[20] , 
        \ScanLink23[14] , \ScanLink20[4] , \wBIn19[31] , \wBIn30[9] , 
        \wRegInB22[10] , \wBIn19[28] , \wRegInB14[15] , \wRegInA3[31] , 
        \wRegInA3[28] , \ScanLink47[3] , \wAIn8[4] , \wAIn18[23] , 
        \wRegInB14[26] , \wRegInB22[23] , \wAMid20[19] , \wAMid24[31] , 
        \wRegInB10[17] , \ScanLink60[12] , \ScanLink56[17] , \ScanLink23[27] , 
        \ScanLink44[0] , \ScanLink15[22] , \ScanLink43[23] , \ScanLink36[13] , 
        \wAMid24[28] , \wRegInB0[7] , \wRegInB26[12] , \wRegInA20[2] , 
        \wBIn2[10] , \wAIn15[8] , \wBMid18[27] , \ScanLink60[6] , 
        \ScanLink27[16] , \wBMid21[3] , \ScanLink52[26] , \ScanLink64[23] , 
        \ScanLink11[13] , \ScanLink47[12] , \ScanLink32[22] , \wBMid22[0] , 
        \ScanLink63[5] , \wBMid18[14] , \wRegInB3[4] , \wRegInA7[19] , 
        \wRegInA18[10] , \wRegInA23[1] , \ScanLink64[10] , \ScanLink47[21] , 
        \ScanLink11[20] , \ScanLink32[11] , \wRegInB24[3] , \wRegInB26[21] , 
        \ScanLink52[15] , \ScanLink27[25] , \wAIn0[26] , \wAMid0[30] , 
        \wAMid0[29] , \wBIn2[23] , \wBIn7[8] , \wRegInB10[24] , 
        \wRegInA18[23] , \wRegInB27[0] , \wBMid1[22] , \wAIn10[5] , 
        \wAIn13[6] , \wBMid13[18] , \wBMid30[30] , \ScanLink59[19] , 
        \wBIn20[10] , \wBMid30[29] , \wRegInB6[9] , \wAIn21[28] , \wBIn16[15] , 
        \wAMid19[12] , \wAIn21[31] , \ScanLink8[22] , \wBIn16[26] , 
        \wAMid19[21] , \wBIn20[23] , \wBIn1[6] , \wBIn2[5] , \wBMid1[11] , 
        \wBIn11[2] , \wBIn12[1] , \wAMid4[22] , \wBIn6[31] , \wRegInA25[19] , 
        \ScanLink8[11] , \wBIn6[28] , \wRegInA3[21] , \ScanLink6[6] , 
        \wAMid15[7] , \wAMid16[15] , \wBMid18[3] , \wAMid20[10] , 
        \wRegInB5[24] , \ScanLink59[6] , \ScanLink7[25] , \wAMid16[4] , 
        \wBIn19[12] , \wAIn31[7] , \ScanLink44[9] , \ScanLink5[5] , 
        \wRegInA3[12] , \wRegInB5[17] , \wRegInA9[7] , \wRegInA19[2] , 
        \ScanLink7[16] , \ScanLink36[30] , \ScanLink15[18] , \wAMid16[26] , 
        \ScanLink60[31] , \ScanLink60[28] , \ScanLink43[19] , \ScanLink36[29] , 
        \wAIn18[19] , \wBIn19[21] , \wAMid20[23] , \wBIn30[0] , 
        \wRegInB22[19] , \wAIn29[5] , \wRegInA17[17] , \wRegInA21[12] , 
        \ScanLink41[4] , \ScanLink0[8] , \ScanLink28[11] , \wBMid17[20] , 
        \wAIn0[15] , \wAMid4[11] , \wBMid5[30] , \wAIn13[26] , \wAIn13[15] , 
        \wBMid21[25] , \wAIn25[10] , \ScanLink48[15] , \ScanLink42[7] , 
        \wBIn24[31] , \wBIn24[28] , \wAIn30[24] , \wRegInB29[15] , \wBIn28[2] , 
        \wRegInA17[24] , \wRegInA21[21] , \ScanLink25[0] , \wRegInB29[26] , 
        \wAMid13[9] , \wAIn25[23] , \wAIn30[17] , \ScanLink26[3] , 
        \wBMid21[16] , \wBMid5[29] , \ScanLink48[26] , \wBMid17[13] , 
        \ScanLink28[22] , \wAMid0[20] , \wBMid1[18] , \wBIn12[8] , 
        \wAIn17[17] , \wAMid19[31] , \wAIn21[12] , \wAMid19[28] , 
        \wBMid25[27] , \ScanLink39[27] , \wAMid0[13] , \wAIn4[24] , 
        \wBMid13[22] , \ScanLink59[23] , \wBIn9[15] , \wBMid8[4] , 
        \wBMid30[13] , \wRegInB22[4] , \wBMid13[11] , \wAMid29[3] , 
        \wRegInA13[15] , \wRegInB21[7] , \wRegInA25[10] , \ScanLink8[18] , 
        \wRegInA30[24] , \ScanLink59[10] , \wAIn4[17] , \wBMid30[20] , 
        \wRegInA26[5] , \wRegInB6[0] , \wBIn7[1] , \wBIn9[26] , \wAMid9[3] , 
        \wAIn21[21] , \wBMid25[14] , \ScanLink39[14] , \wBMid27[4] , 
        \wAIn17[24] , \wBIn20[19] , \wBMid24[7] , \wRegInB5[3] , 
        \wRegInA13[26] , \wRegInA25[23] , \wRegInA30[17] , \wRegInA25[6] , 
        \ScanLink64[19] , \ScanLink47[31] , \ScanLink47[28] , \ScanLink11[29] , 
        \ScanLink32[18] , \ScanLink11[30] , \wAMid12[17] , \wBIn14[6] , 
        \wRegInB26[31] , \wRegInB26[28] , \ScanLink19[4] , \wBIn4[2] , 
        \wBIn17[5] , \wAMid24[12] , \ScanLink3[27] , \wAMid12[24] , 
        \wAMid24[21] , \wRegInB1[26] , \wRegInB27[9] , \wRegInA7[23] , 
        \wAIn15[1] , \wAIn16[2] , \wAIn0[5] , \wBMid0[21] , \wAMid1[19] , 
        \wBIn2[19] , \wAMid7[5] , \wBMid22[9] , \wBMid29[2] , \wRegInB1[15] , 
        \wRegInA7[10] , \wRegInA18[19] , \wRegInA23[8] , \ScanLink3[14] , 
        \wBIn17[16] , \wRegInB8[6] , \wRegInA28[3] , \wRegInA24[30] , 
        \ScanLink9[21] , \wRegInA24[29] , \wAMid18[11] , \wBIn21[13] , 
        \wBMid0[12] , \wAMid4[6] , \wBMid6[2] , \wAMid24[6] , \ScanLink9[12] , 
        \wAMid2[8] , \wBIn3[13] , \wBMid5[1] , \wBMid12[31] , \ScanLink58[30] , 
        \wBMid12[28] , \ScanLink58[29] , \wBIn17[25] , \wBIn21[20] , 
        \wAMid27[5] , \wAMid18[22] , \wAIn20[18] , \wRegInA19[13] , 
        \wAIn18[4] , \wBMid19[24] , \ScanLink46[11] , \ScanLink33[21] , 
        \ScanLink26[15] , \ScanLink10[10] , \wRegInA30[1] , \ScanLink53[25] , 
        \wRegInB27[11] , \wBIn3[20] , \wBIn9[7] , \wRegInB11[14] , 
        \wAMid22[8] , \wRegInA6[29] , \wAIn5[8] , \wBIn7[22] , \wBIn7[11] , 
        \wAMid18[2] , \wAIn19[13] , \wBIn19[3] , \wBMid19[17] , \wAMid25[18] , 
        \wRegInA6[30] , \ScanLink17[2] , \wRegInB11[27] , \wRegInA19[20] , 
        \wRegInB27[22] , \ScanLink53[16] , \wAMid21[29] , \wRegInB10[6] , 
        \ScanLink46[22] , \ScanLink26[26] , \ScanLink14[1] , \ScanLink33[12] , 
        \ScanLink10[23] , \wRegInB15[16] , \wAMid21[30] , \wRegInB23[13] , 
        \ScanLink61[22] , \ScanLink57[27] , \ScanLink30[7] , \ScanLink22[17] , 
        \ScanLink42[13] , \ScanLink37[23] , \ScanLink14[12] , \ScanLink33[4] , 
        \wBMid15[6] , \wBIn23[9] , \wRegInA2[18] , \wRegInB13[5] , 
        \ScanLink61[11] , \ScanLink54[3] , \ScanLink42[20] , \ScanLink37[10] , 
        \ScanLink14[21] , \wBIn18[18] , \wAIn19[20] , \wRegInB23[20] , 
        \ScanLink57[14] , \ScanLink22[24] , \ScanLink8[0] , \wRegInA4[2] , 
        \wRegInA7[1] , \wRegInA14[7] , \wRegInB15[25] , \wRegInA17[4] , 
        \wBMid16[5] , \ScanLink57[0] , \wBMid4[23] , \wBIn13[27] , 
        \wBIn13[14] , \wBMid16[19] , \wBIn26[4] , \wRegInB16[8] , 
        \ScanLink29[31] , \wAIn24[30] , \wBIn25[11] , \ScanLink36[9] , 
        \ScanLink29[28] , \wAIn24[29] , \wBIn30[25] , \wBIn25[7] , 
        \wRegInA9[27] , \ScanLink28[5] , \wBIn25[22] , \wBIn30[16] , 
        \wAIn27[3] , \wBIn1[2] , \wBIn2[1] , \wBMid1[26] , \wAIn3[6] , 
        \wBMid4[10] , \wAMid5[31] , \wBMid13[8] , \wAMid5[28] , \wRegInA9[14] , 
        \wRegInA12[9] , \wAIn10[1] , \wAIn24[0] , \wRegInA20[18] , \wAIn13[2] , 
        \wBIn16[11] , \wAMid19[16] , \wBMid27[9] , \ScanLink8[26] , 
        \wAIn17[30] , \wBIn20[14] , \wAIn17[29] , \wRegInA26[8] , 
        \ScanLink39[19] , \wBIn9[18] , \wBMid25[19] , \wRegInA13[18] , 
        \wRegInA30[29] , \ScanLink8[15] , \wRegInA30[30] , \wBIn11[6] , 
        \wBIn2[14] , \wBMid1[15] , \wAIn4[30] , \wAIn4[29] , \wBIn12[5] , 
        \wBMid8[9] , \wRegInB22[9] , \wBIn16[22] , \wAMid19[25] , \wBIn20[27] , 
        \wBMid22[4] , \wRegInB3[0] , \wRegInA18[14] , \wRegInA23[5] , 
        \ScanLink3[19] , \wBMid18[23] , \wBMid21[7] , \wRegInB1[18] , 
        \ScanLink63[1] , \ScanLink47[16] , \ScanLink32[26] , \ScanLink64[27] , 
        \ScanLink11[17] , \ScanLink60[2] , \ScanLink27[12] , \ScanLink52[22] , 
        \wRegInA20[6] , \wBIn2[27] , \wAMid12[30] , \wAMid12[29] , 
        \wRegInB0[3] , \wRegInB26[16] , \wRegInB10[13] , \wBIn17[8] , 
        \wRegInB10[20] , \wRegInA18[27] , \wRegInB27[4] , \ScanLink19[9] , 
        \wAIn0[18] , \wBIn6[25] , \wBIn6[16] , \wAIn18[14] , \wBMid18[10] , 
        \wRegInB24[7] , \wRegInB26[25] , \ScanLink52[11] , \wRegInB14[11] , 
        \ScanLink64[14] , \ScanLink47[25] , \ScanLink27[21] , \ScanLink32[15] , 
        \ScanLink11[24] , \wRegInB22[14] , \ScanLink60[25] , \ScanLink56[20] , 
        \ScanLink23[10] , \ScanLink20[0] , \ScanLink43[14] , \ScanLink36[24] , 
        \ScanLink15[15] , \ScanLink23[3] , \wAIn8[0] , \wAMid16[18] , 
        \wAMid16[9] , \wAIn18[27] , \wRegInB22[27] , \ScanLink60[16] , 
        \ScanLink44[4] , \ScanLink43[27] , \ScanLink36[17] , \ScanLink56[13] , 
        \ScanLink15[26] , \ScanLink5[8] , \ScanLink23[23] , \wRegInB14[22] , 
        \ScanLink7[31] , \ScanLink7[28] , \wBMid5[24] , \wRegInB5[30] , 
        \wRegInB5[29] , \ScanLink47[7] , \wAIn5[5] , \wBMid5[17] , 
        \wAMid10[7] , \wBIn12[13] , \wBIn24[16] , \wAMid13[4] , \wBIn31[22] , 
        \wRegInA17[30] , \wRegInB18[3] , \wRegInA17[29] , \wBIn12[20] , 
        \wRegInA8[20] , \ScanLink38[2] , \wAIn13[18] , \wBIn24[25] , 
        \wBIn31[11] , \ScanLink3[6] , \wAIn30[29] , \wAIn30[30] , 
        \wRegInB29[18] , \wBMid16[8] , \wBMid21[31] , \wBMid21[28] , 
        \ScanLink48[18] , \wAIn29[8] , \wRegInA8[13] , \wRegInA2[26] , 
        \ScanLink41[9] , \ScanLink0[5] , \wAIn6[6] , \wAMid17[12] , 
        \wBIn18[15] , \wAMid21[17] , \wAIn22[3] , \wRegInB4[23] , 
        \wRegInA17[9] , \ScanLink6[22] , \ScanLink49[1] , \wRegInB15[31] , 
        \wRegInB15[28] , \wAIn21[0] , \ScanLink57[19] , \ScanLink22[29] , 
        \wBIn23[4] , \wRegInB13[8] , \ScanLink22[30] , \ScanLink6[11] , 
        \wRegInA2[15] , \wRegInB4[10] , \ScanLink33[9] , \wAIn0[8] , 
        \wAIn1[21] , \wAMid5[25] , \wBMid10[6] , \wAMid17[21] , \wBIn18[26] , 
        \wBIn20[7] , \wAMid21[24] , \wRegInA16[10] , \wRegInA20[15] , 
        \ScanLink51[3] , \wRegInA1[2] , \wRegInA9[19] , \wRegInA11[7] , 
        \ScanLink29[16] , \wBMid16[27] , \wBMid20[22] , \wRegInA2[1] , 
        \wAIn24[17] , \wRegInA12[4] , \ScanLink49[12] , \ScanLink52[0] , 
        \wAIn0[1] , \wAIn1[31] , \wAIn1[12] , \wAMid5[16] , \wAIn12[21] , 
        \wAIn12[12] , \wBMid13[5] , \wAIn31[23] , \wRegInB28[12] , 
        \wRegInB15[6] , \ScanLink28[8] , \wRegInA16[23] , \wRegInA20[26] , 
        \ScanLink35[7] , \wRegInB28[21] , \wBIn13[19] , \wAIn24[24] , 
        \wAIn31[10] , \ScanLink36[4] , \wBIn30[28] , \wBMid16[14] , 
        \wBMid20[11] , \wBIn30[31] , \wRegInB16[5] , \ScanLink49[21] , 
        \wBIn26[9] , \ScanLink29[25] , \wBMid0[1] , \wAMid1[27] , \wAIn16[10] , 
        \wBIn17[31] , \wAMid27[8] , \ScanLink12[2] , \wBIn17[28] , 
        \wAIn20[15] , \wBMid24[20] , \ScanLink38[20] , \wAMid1[14] , 
        \wAIn5[23] , \wBMid12[25] , \ScanLink58[24] , \wBIn8[12] , 
        \wBMid12[16] , \wRegInB31[0] , \wRegInA12[12] , \wRegInA24[17] , 
        \wRegInA31[23] , \ScanLink11[1] , \ScanLink58[17] , \wBMid3[2] , 
        \wAIn5[10] , \wAMid7[8] , \wAIn16[23] , \wAIn20[26] , \wBMid24[13] , 
        \ScanLink38[13] , \wRegInA12[21] , \wRegInA24[24] , \wRegInA31[10] , 
        \wBIn8[21] , \wAMid21[6] , \wRegInB29[2] , \wAMid13[10] , 
        \wAMid30[21] , \wAMid22[5] , \wAMid25[15] , \ScanLink2[20] , 
        \wRegInB0[21] , \wRegInA6[24] , \wAMid1[6] , \wAMid2[5] , 
        \wAMid13[23] , \wAIn18[9] , \wAMid25[26] , \wAMid30[12] , 
        \wRegInB11[19] , \wBMid19[30] , \wBMid19[29] , \ScanLink26[18] , 
        \ScanLink53[28] , \wRegInB0[12] , \wRegInA6[17] , \ScanLink53[31] , 
        \ScanLink2[13] , \wAIn3[2] , \wBMid4[27] , \wAIn12[31] , \wAIn12[28] , 
        \wBIn13[10] , \wBIn25[3] , \wBIn30[21] , \wRegInA9[23] , 
        \ScanLink28[1] , \wRegInB28[28] , \wAIn31[19] , \wRegInB28[31] , 
        \wBMid20[18] , \wBIn25[15] , \wBIn26[0] , \ScanLink49[31] , 
        \ScanLink49[28] , \wAIn24[4] , \wBMid4[14] , \wRegInA2[8] , 
        \wRegInA9[10] , \wRegInA16[19] , \wAIn1[28] , \wBMid0[25] , 
        \wBMid0[8] , \wBIn3[17] , \wBIn7[26] , \wBIn7[15] , \wBIn13[23] , 
        \wBIn25[26] , \wAIn27[7] , \wBIn30[12] , \ScanLink52[9] , 
        \wRegInB13[1] , \ScanLink6[18] , \wBMid16[1] , \wAMid17[31] , 
        \wAMid18[6] , \wAIn19[17] , \wRegInB4[19] , \ScanLink33[0] , 
        \ScanLink61[26] , \ScanLink14[16] , \ScanLink57[23] , \ScanLink42[17] , 
        \ScanLink37[27] , \ScanLink30[3] , \ScanLink22[13] , \wRegInB23[17] , 
        \wAMid17[28] , \wRegInB15[12] , \wRegInB10[2] , \ScanLink57[4] , 
        \wBMid15[2] , \wAIn19[24] , \wRegInA4[6] , \wRegInA7[5] , 
        \wRegInA14[3] , \wRegInB15[21] , \wRegInA17[0] , \wRegInB23[24] , 
        \ScanLink8[4] , \wAIn21[9] , \ScanLink57[10] , \ScanLink49[8] , 
        \ScanLink22[20] , \wAIn18[0] , \wRegInB11[10] , \ScanLink61[15] , 
        \ScanLink54[7] , \ScanLink14[25] , \ScanLink42[24] , \ScanLink37[14] , 
        \wRegInB27[15] , \wRegInA30[5] , \wBMid19[20] , \ScanLink53[21] , 
        \ScanLink26[11] , \ScanLink46[15] , \ScanLink33[25] , \ScanLink10[14] , 
        \wAMid13[19] , \wBIn19[7] , \wBMid19[13] , \wRegInA19[17] , 
        \ScanLink53[12] , \ScanLink46[26] , \ScanLink14[5] , \ScanLink10[27] , 
        \ScanLink33[16] , \wAMid30[31] , \wAMid30[28] , \wRegInB11[23] , 
        \wRegInB27[26] , \ScanLink26[22] , \wRegInA19[24] , \ScanLink17[6] , 
        \ScanLink2[30] , \ScanLink2[29] , \wBIn3[24] , \wAMid4[2] , \wBIn9[3] , 
        \wRegInB0[31] , \wRegInB0[28] , \wBMid0[16] , \wAIn5[19] , \wBMid5[5] , 
        \wAMid7[1] , \wBIn8[31] , \wBIn17[12] , \wAMid18[15] , \wBIn21[17] , 
        \wRegInB8[2] , \wRegInA12[28] , \ScanLink9[25] , \wRegInA12[31] , 
        \wRegInA31[19] , \wRegInA28[7] , \wBIn8[28] , \wBIn17[21] , 
        \wAMid18[26] , \wBMid29[6] , \wAIn16[19] , \wBIn21[24] , \wAMid27[1] , 
        \wBMid24[29] , \ScanLink38[30] , \ScanLink38[29] , \wBIn4[6] , 
        \wBMid6[6] , \wBMid24[30] , \wRegInB31[9] , \ScanLink9[16] , 
        \wBIn17[1] , \wAMid24[2] , \ScanLink11[8] , \wRegInB1[22] , 
        \wRegInA7[27] , \wBIn7[5] , \wAMid12[13] , \wAMid24[16] , 
        \ScanLink19[0] , \ScanLink3[23] , \wRegInB10[30] , \wBIn14[2] , 
        \wRegInB10[29] , \wBMid18[19] , \ScanLink27[31] , \wRegInB1[11] , 
        \wRegInB3[9] , \ScanLink52[18] , \ScanLink27[28] , \ScanLink3[10] , 
        \ScanLink63[8] , \wAMid0[24] , \wBIn2[8] , \wBIn9[11] , \wAMid12[20] , 
        \wAIn15[5] , \wAIn16[6] , \wRegInA7[14] , \wAMid24[25] , 
        \wRegInA13[11] , \wRegInA30[20] , \wRegInB21[3] , \wRegInA25[14] , 
        \wAMid29[7] , \wAIn4[20] , \wBMid8[0] , \wBMid30[17] , \wRegInB22[0] , 
        \wAMid0[17] , \wAIn4[13] , \wBIn9[22] , \wBMid13[26] , 
        \ScanLink59[27] , \wAIn17[13] , \wAIn21[16] , \wBMid25[23] , 
        \ScanLink39[23] , \wAMid9[7] , \wAIn10[8] , \wRegInB5[7] , 
        \wRegInA25[2] , \wRegInA25[27] , \wRegInA30[13] , \wBMid24[3] , 
        \wRegInA13[22] , \wBIn16[18] , \wAIn17[20] , \wBMid27[0] , 
        \wAIn21[25] , \wBMid25[10] , \ScanLink39[10] , \wBMid30[24] , 
        \wRegInB6[4] , \wBMid13[15] , \ScanLink59[14] , \wBIn12[30] , 
        \wBIn12[29] , \wAIn13[11] , \wAIn30[20] , \wRegInA26[1] , 
        \wRegInB29[11] , \wAIn25[14] , \wBIn31[18] , \ScanLink42[3] , 
        \ScanLink48[11] , \wAIn0[22] , \wBMid21[21] , \wAIn0[11] , 
        \wAMid4[26] , \ScanLink28[15] , \wBMid17[24] , \wAIn29[1] , 
        \wRegInA17[13] , \wRegInA21[16] , \ScanLink41[0] , \wBIn4[4] , 
        \wAMid4[15] , \wBMid17[17] , \wBIn7[7] , \wAIn8[9] , \wAIn13[22] , 
        \wBMid21[12] , \ScanLink48[22] , \ScanLink28[26] , \wAIn25[27] , 
        \wAIn30[13] , \ScanLink26[7] , \wRegInB29[22] , \wAMid16[11] , 
        \wBIn19[16] , \wBMid18[7] , \wBIn28[6] , \wAIn31[3] , \wRegInA8[30] , 
        \wRegInA8[29] , \wRegInA17[20] , \wRegInA21[25] , \ScanLink25[4] , 
        \wRegInA9[3] , \wRegInA19[6] , \ScanLink5[1] , \wAMid20[14] , 
        \ScanLink59[2] , \wAMid12[11] , \wAMid15[3] , \wAMid16[22] , 
        \wBIn19[25] , \wAMid20[27] , \wBIn30[4] , \wRegInA3[25] , 
        \wRegInB5[20] , \ScanLink7[21] , \ScanLink6[2] , \wRegInB14[18] , 
        \wAMid16[0] , \wRegInA3[16] , \ScanLink56[30] , \ScanLink56[29] , 
        \ScanLink23[19] , \ScanLink20[9] , \wRegInB5[13] , \ScanLink7[12] , 
        \wBIn14[0] , \wBIn17[3] , \wAMid24[14] , \ScanLink19[2] , 
        \wAMid12[22] , \wAMid24[27] , \wRegInB1[20] , \ScanLink3[21] , 
        \wRegInA7[25] , \wRegInB0[8] , \wAIn15[7] , \wRegInB10[18] , 
        \wBMid18[31] , \ScanLink52[30] , \wBMid18[28] , \ScanLink52[29] , 
        \wRegInA7[16] , \ScanLink60[9] , \ScanLink27[19] , \wAIn0[20] , 
        \wAMid0[26] , \wBIn1[9] , \wAIn16[4] , \wBIn16[30] , \wBIn16[29] , 
        \wAIn17[11] , \wRegInB1[13] , \ScanLink3[12] , \wAIn21[14] , 
        \wAIn4[22] , \wBMid8[2] , \wBMid25[21] , \ScanLink39[21] , 
        \wBMid30[15] , \wRegInB22[2] , \wBMid13[24] , \ScanLink59[25] , 
        \wAMid0[15] , \wAIn4[11] , \wBIn9[13] , \wAMid29[5] , \wRegInA13[13] , 
        \wRegInB21[1] , \wRegInA25[16] , \wRegInA30[22] , \wBMid30[26] , 
        \wRegInB6[6] , \wRegInA26[3] , \wBIn9[20] , \wAMid9[5] , \wAIn13[9] , 
        \wBMid13[17] , \wAIn21[27] , \wBMid25[12] , \ScanLink59[16] , 
        \ScanLink39[12] , \wBMid27[2] , \wAIn17[22] , \wBMid24[1] , 
        \wRegInA30[11] , \wRegInB5[5] , \wRegInA13[20] , \wRegInA25[25] , 
        \wRegInA25[0] , \wAIn29[3] , \wRegInA8[18] , \wRegInA17[11] , 
        \ScanLink41[2] , \wRegInA21[14] , \wAIn0[13] , \wAMid4[24] , 
        \wBMid17[26] , \wBIn12[18] , \wAIn13[20] , \wAIn13[13] , \wBMid21[23] , 
        \ScanLink48[13] , \ScanLink28[17] , \wAIn25[16] , \wAIn30[22] , 
        \ScanLink42[1] , \wRegInB29[13] , \wBIn28[4] , \wRegInB18[8] , 
        \ScanLink38[9] , \wRegInA21[27] , \ScanLink25[6] , \wAIn30[11] , 
        \wRegInA17[22] , \ScanLink26[5] , \wBIn31[30] , \wRegInB29[20] , 
        \wBMid21[10] , \wAIn25[25] , \wBIn31[29] , \ScanLink48[20] , 
        \wAIn0[3] , \wAIn1[19] , \wAMid4[17] , \ScanLink28[24] , \wBMid4[25] , 
        \wAMid15[1] , \wAMid16[13] , \wBMid17[15] , \wAMid20[16] , 
        \wRegInA3[27] , \ScanLink6[0] , \wRegInB5[22] , \ScanLink7[23] , 
        \ScanLink59[0] , \wAMid16[2] , \wBIn19[14] , \wBMid18[5] , \wAIn31[1] , 
        \wRegInA9[1] , \wRegInB14[30] , \wRegInB14[29] , \ScanLink23[31] , 
        \ScanLink5[3] , \wRegInB5[11] , \wRegInA19[4] , \ScanLink23[28] , 
        \ScanLink56[18] , \ScanLink7[10] , \ScanLink23[8] , \wRegInA3[14] , 
        \wAMid16[20] , \wBIn19[27] , \wAMid20[25] , \wBIn30[6] , \wBIn26[2] , 
        \wBIn13[21] , \wBIn13[12] , \wBIn25[17] , \wBIn30[23] , \wBIn25[1] , 
        \wRegInA9[21] , \wRegInA16[31] , \wRegInA16[28] , \ScanLink28[3] , 
        \wBIn30[10] , \wRegInB28[19] , \wAIn3[0] , \wBMid4[16] , \wAIn12[19] , 
        \wAIn31[31] , \wBMid20[30] , \wBMid20[29] , \wBIn25[24] , \wAIn27[5] , 
        \wAIn31[28] , \ScanLink49[19] , \wAIn24[6] , \wRegInA1[9] , 
        \wRegInA9[12] , \ScanLink51[8] , \wAMid18[4] , \wRegInB10[0] , 
        \wRegInB15[10] , \wAIn19[15] , \wRegInB23[15] , \wBMid0[27] , 
        \wBIn3[26] , \wBIn3[15] , \wBIn7[24] , \wBIn7[17] , \ScanLink61[24] , 
        \ScanLink57[21] , \ScanLink30[1] , \ScanLink22[11] , \ScanLink42[15] , 
        \ScanLink14[14] , \ScanLink37[25] , \ScanLink33[2] , \wBMid15[0] , 
        \wRegInB13[3] , \ScanLink61[17] , \ScanLink14[27] , \ScanLink57[12] , 
        \ScanLink54[5] , \ScanLink37[16] , \ScanLink42[26] , \ScanLink22[22] , 
        \wAMid17[19] , \wAIn19[26] , \ScanLink8[6] , \wRegInA4[4] , 
        \wRegInA14[1] , \wRegInB23[26] , \wRegInB15[23] , \wRegInA7[7] , 
        \ScanLink6[29] , \wRegInA17[2] , \ScanLink6[30] , \ScanLink57[6] , 
        \wBMid16[3] , \wAIn22[8] , \wRegInB4[31] , \wRegInB4[28] , 
        \wRegInA19[15] , \ScanLink2[18] , \wBIn9[1] , \wAMid13[31] , 
        \wAIn18[2] , \wBMid19[22] , \wRegInB0[19] , \ScanLink46[17] , 
        \ScanLink10[16] , \ScanLink33[27] , \wRegInB27[17] , \ScanLink53[23] , 
        \ScanLink26[13] , \wRegInA30[7] , \wAMid30[19] , \wRegInB11[12] , 
        \wAMid13[28] , \ScanLink17[4] , \wBMid3[9] , \wBIn19[5] , 
        \wBMid19[11] , \wRegInB11[21] , \wRegInA19[26] , \wRegInB27[24] , 
        \ScanLink26[20] , \ScanLink53[10] , \wRegInB29[9] , \wAMid4[0] , 
        \wAMid7[3] , \wBMid29[4] , \ScanLink46[24] , \ScanLink33[14] , 
        \ScanLink10[25] , \ScanLink14[7] , \wAIn16[31] , \wAIn16[28] , 
        \wBIn17[10] , \wRegInB8[0] , \wRegInA28[5] , \ScanLink9[27] , 
        \wAMid18[17] , \wBIn21[15] , \wBMid24[18] , \wBMid0[14] , \wBMid6[4] , 
        \wAMid24[0] , \ScanLink38[18] , \wBIn8[19] , \wRegInA12[19] , 
        \wRegInA31[31] , \wRegInA31[28] , \ScanLink9[14] , \wAIn5[31] , 
        \wAIn5[28] , \wAIn5[7] , \wAIn6[4] , \wBMid5[7] , \wBIn21[26] , 
        \wAMid27[3] , \ScanLink12[9] , \wBIn17[23] , \wAMid18[24] , 
        \wAIn21[2] , \wBMid15[9] , \wAMid17[10] , \wRegInA14[8] , \wBIn18[17] , 
        \wAMid21[15] , \ScanLink49[3] , \ScanLink6[20] , \wAMid17[23] , 
        \wBIn20[5] , \wAIn22[1] , \wRegInA2[24] , \wRegInB4[21] , 
        \wAMid21[26] , \wRegInB10[9] , \wRegInB15[19] , \wBIn18[24] , 
        \ScanLink57[28] , \wAIn1[23] , \wAMid5[27] , \wAIn12[10] , \wBIn23[6] , 
        \wRegInA2[17] , \ScanLink57[31] , \ScanLink30[8] , \ScanLink22[18] , 
        \wRegInB4[12] , \wRegInB28[10] , \ScanLink6[13] , \wBIn13[31] , 
        \wBMid13[7] , \wAIn31[21] , \wBIn13[28] , \wAIn24[15] , \wBIn30[19] , 
        \ScanLink52[2] , \wBMid16[25] , \wBMid20[20] , \wRegInA2[3] , 
        \wRegInA12[6] , \ScanLink49[10] , \ScanLink29[14] , \wAIn1[10] , 
        \wAIn3[9] , \wBMid10[4] , \wRegInA1[0] , \wRegInA11[5] , 
        \wRegInA20[17] , \wAMid5[14] , \wRegInA16[12] , \ScanLink51[1] , 
        \ScanLink29[27] , \wBMid16[16] , \wBIn1[0] , \wBMid0[3] , \wAMid1[25] , 
        \wBIn8[10] , \wAIn12[23] , \wBMid20[13] , \wRegInB16[7] , \wAIn24[26] , 
        \ScanLink49[23] , \wAMid24[9] , \wBIn25[8] , \wAIn31[12] , 
        \wRegInB28[23] , \wRegInA16[21] , \ScanLink36[6] , \wRegInA20[24] , 
        \ScanLink35[5] , \wRegInA9[31] , \wRegInA9[28] , \wRegInB15[4] , 
        \wRegInA12[10] , \wRegInA24[15] , \wRegInA31[21] , \ScanLink11[3] , 
        \wRegInB31[2] , \wBMid12[27] , \ScanLink58[26] , \wAMid1[16] , 
        \wAMid4[9] , \wAIn5[21] , \wBIn8[23] , \wAIn16[12] , \wAIn20[17] , 
        \wBMid24[22] , \ScanLink38[22] , \ScanLink12[0] , \wAIn16[21] , 
        \wRegInB8[9] , \wRegInA24[26] , \wRegInA12[23] , \wRegInA31[12] , 
        \wBIn17[19] , \wAIn20[24] , \wBMid24[11] , \ScanLink38[11] , 
        \wAIn5[12] , \wBMid12[14] , \ScanLink58[15] , \wAMid1[4] , \wBMid3[0] , 
        \wBIn9[8] , \wAMid22[7] , \wRegInA6[26] , \wRegInB0[23] , 
        \wAMid13[12] , \wAMid25[17] , \ScanLink2[22] , \wAMid30[23] , 
        \wRegInB11[28] , \wRegInB11[31] , \wRegInB29[0] , \wBMid19[18] , 
        \ScanLink53[19] , \ScanLink26[29] , \wAMid21[4] , \ScanLink26[30] , 
        \wBMid1[24] , \wAMid2[7] , \wAMid13[21] , \wAMid30[10] , 
        \wRegInB0[10] , \ScanLink2[11] , \wRegInA6[15] , \wAMid25[24] , 
        \wAIn4[18] , \wBIn9[30] , \wBIn9[29] , \wAIn10[3] , \wAIn13[0] , 
        \wBIn16[13] , \wBIn20[16] , \wAMid19[14] , \wBMid24[8] , 
        \wRegInA13[30] , \wRegInA13[29] , \wRegInA30[18] , \ScanLink8[24] , 
        \wBIn16[20] , \wRegInA25[9] , \wAIn17[18] , \wAMid19[27] , 
        \wBIn20[25] , \wBMid25[31] , \wBIn2[3] , \wBMid1[17] , \wBIn12[7] , 
        \wBIn11[4] , \wBMid25[28] , \ScanLink39[28] , \wRegInB21[8] , 
        \ScanLink39[31] , \wRegInB10[11] , \ScanLink8[17] , \wRegInA20[4] , 
        \wBIn2[16] , \wBMid18[21] , \wRegInB0[1] , \wRegInB26[14] , 
        \wBMid21[5] , \ScanLink64[25] , \ScanLink60[0] , \ScanLink52[20] , 
        \ScanLink27[10] , \ScanLink47[14] , \ScanLink32[24] , \ScanLink63[3] , 
        \ScanLink11[15] , \wBMid18[12] , \wBMid22[6] , \wRegInB3[2] , 
        \wRegInA18[16] , \wRegInA23[7] , \ScanLink64[16] , \ScanLink47[27] , 
        \ScanLink32[17] , \ScanLink11[26] , \ScanLink27[23] , \ScanLink52[13] , 
        \wAIn0[30] , \wAIn0[29] , \wBIn2[25] , \wAMid12[18] , \wRegInB24[5] , 
        \wRegInB26[27] , \wBIn14[9] , \wRegInB10[22] , \wRegInA18[25] , 
        \wRegInB27[6] , \ScanLink3[31] , \ScanLink3[28] , \wBIn6[27] , 
        \wBIn6[14] , \wRegInB1[30] , \wRegInB1[29] , \ScanLink7[19] , 
        \wAMid15[8] , \wRegInB5[18] , \ScanLink43[16] , \ScanLink23[1] , 
        \ScanLink36[26] , \wAMid16[30] , \wAMid16[29] , \wAIn18[16] , 
        \wRegInB22[16] , \ScanLink60[27] , \ScanLink56[22] , \ScanLink15[17] , 
        \ScanLink23[12] , \ScanLink20[2] , \wRegInB14[13] , \ScanLink6[9] , 
        \wBMid5[26] , \wAIn8[2] , \ScanLink47[5] , \wAMid10[5] , \wAIn18[25] , 
        \wRegInB14[20] , \ScanLink59[9] , \wAIn31[8] , \wRegInA9[8] , 
        \wRegInB22[25] , \ScanLink23[21] , \wRegInA8[22] , \ScanLink60[14] , 
        \ScanLink56[11] , \ScanLink44[6] , \ScanLink36[15] , \ScanLink43[25] , 
        \ScanLink15[24] , \ScanLink38[0] , \wBIn12[11] , \wAMid13[6] , 
        \wRegInB18[1] , \wAIn13[30] , \wBIn24[14] , \wBIn31[20] , \wAIn13[29] , 
        \wAIn30[18] , \wRegInB29[30] , \wRegInB29[29] , \wBMid5[15] , 
        \wBMid21[19] , \ScanLink48[29] , \wRegInA8[11] , \wRegInA17[18] , 
        \ScanLink48[30] , \ScanLink0[7] , \wAIn0[24] , \wAIn0[7] , 
        \wBMid0[23] , \wBIn12[22] , \wBIn24[27] , \ScanLink3[4] , \wBIn31[13] , 
        \ScanLink42[8] , \wBMid0[10] , \wAMid1[31] , \wAMid4[4] , \wBMid5[3] , 
        \wAMid7[7] , \wBMid12[19] , \wBIn17[14] , \wAMid18[13] , \wBIn21[11] , 
        \ScanLink58[18] , \wAIn20[30] , \wAIn20[29] , \wRegInB8[4] , 
        \wRegInA28[1] , \ScanLink9[23] , \wBMid29[0] , \wBIn17[27] , 
        \wAMid18[20] , \wBIn21[22] , \wAMid27[7] , \wAMid1[28] , \wAMid1[9] , 
        \wBIn3[11] , \wBMid6[0] , \wAIn18[6] , \wAMid24[4] , \ScanLink9[10] , 
        \wRegInB11[16] , \wRegInA24[18] , \wRegInA30[3] , \wBMid19[26] , 
        \wAMid25[30] , \wAMid25[29] , \wRegInB27[13] , \ScanLink53[27] , 
        \wRegInA6[18] , \ScanLink46[13] , \ScanLink26[17] , \ScanLink33[23] , 
        \ScanLink10[12] , \wRegInA19[11] , \wAIn3[4] , \wBIn3[22] , 
        \wBIn19[1] , \wBMid19[15] , \wAMid21[9] , \ScanLink46[20] , 
        \ScanLink33[10] , \ScanLink14[3] , \ScanLink10[21] , \ScanLink53[14] , 
        \ScanLink26[24] , \wRegInB11[25] , \wRegInB27[20] , \wRegInA19[22] , 
        \wBMid4[21] , \wAMid5[19] , \wAIn6[9] , \wBIn7[20] , \wBIn7[13] , 
        \wBIn9[5] , \ScanLink17[0] , \wRegInB13[7] , \wBMid16[7] , 
        \wBIn18[30] , \wBIn18[29] , \wAMid18[0] , \wBIn20[8] , 
        \ScanLink61[20] , \ScanLink42[11] , \ScanLink33[6] , \ScanLink37[21] , 
        \ScanLink57[25] , \ScanLink14[10] , \ScanLink30[5] , \ScanLink22[15] , 
        \wAIn19[11] , \wRegInB23[11] , \wRegInB10[4] , \wRegInB15[14] , 
        \wAIn19[22] , \wAMid21[18] , \wRegInA2[30] , \wRegInA2[29] , 
        \wRegInA4[0] , \wRegInA7[3] , \wRegInA17[6] , \ScanLink57[2] , 
        \wRegInA14[5] , \wRegInB15[27] , \ScanLink8[2] , \wRegInB23[22] , 
        \wBIn13[16] , \wBMid15[4] , \wBIn25[5] , \ScanLink61[13] , 
        \ScanLink57[16] , \ScanLink22[26] , \ScanLink54[1] , \ScanLink37[12] , 
        \ScanLink42[22] , \ScanLink14[23] , \wRegInA9[25] , \wRegInB15[9] , 
        \wRegInA20[30] , \ScanLink28[7] , \wRegInA20[29] , \ScanLink35[8] , 
        \wBIn25[13] , \wBIn30[27] , \wBIn26[6] , \wBMid10[9] , \wBMid4[12] , 
        \wAIn24[2] , \wRegInA9[16] , \wRegInA11[8] , \wBMid16[31] , 
        \wBMid16[28] , \wBIn25[20] , \wAIn27[1] , \ScanLink29[19] , 
        \wAMid4[20] , \wBIn6[19] , \wBIn13[25] , \wAMid15[5] , \wAMid16[24] , 
        \wAMid16[17] , \wBIn19[10] , \wAIn24[18] , \wBIn30[14] , \wAIn31[5] , 
        \wRegInA9[5] , \wRegInA19[0] , \ScanLink60[19] , \ScanLink43[31] , 
        \ScanLink15[29] , \ScanLink5[7] , \ScanLink43[28] , \ScanLink36[18] , 
        \ScanLink15[30] , \wAIn18[31] , \wAIn18[28] , \wBMid18[1] , 
        \wAMid20[12] , \wRegInB22[28] , \wBIn19[23] , \wAMid20[21] , 
        \wBIn30[2] , \wRegInA3[23] , \wRegInB5[26] , \wRegInB22[31] , 
        \ScanLink59[4] , \ScanLink7[27] , \ScanLink47[8] , \ScanLink6[4] , 
        \wAMid16[6] , \wRegInA3[10] , \wBMid5[18] , \wAIn13[17] , 
        \wRegInB5[15] , \wRegInB29[17] , \ScanLink7[14] , \wBMid21[27] , 
        \wAIn25[12] , \wAIn30[26] , \ScanLink42[5] , \ScanLink3[9] , 
        \ScanLink48[17] , \wBMid17[22] , \ScanLink28[13] , \wAIn0[17] , 
        \wAMid4[13] , \wAIn29[7] , \wRegInA17[15] , \wRegInA21[10] , 
        \ScanLink41[6] , \ScanLink28[20] , \wBMid17[11] , \wAMid0[22] , 
        \wBIn9[17] , \wAMid10[8] , \wAIn13[24] , \wBMid21[14] , \wAIn25[21] , 
        \ScanLink48[24] , \wBIn24[19] , \wAIn30[15] , \wRegInB29[24] , 
        \ScanLink26[1] , \wBIn11[9] , \wBIn28[0] , \wRegInA17[26] , 
        \wRegInA13[17] , \wRegInA21[23] , \ScanLink25[2] , \wRegInB21[5] , 
        \wRegInA25[12] , \wRegInA30[26] , \wAMid29[1] , \wBMid13[20] , 
        \ScanLink59[21] , \wAMid0[11] , \wBMid1[30] , \wAIn4[26] , \wBMid8[6] , 
        \wBMid30[11] , \wRegInB22[6] , \wBIn9[24] , \wAIn17[15] , \wAIn21[10] , 
        \wBMid25[25] , \ScanLink39[25] , \wBIn20[31] , \wBIn20[28] , 
        \wAMid9[1] , \wAIn17[26] , \wBMid24[5] , \wRegInB5[1] , 
        \wRegInA13[24] , \wRegInA25[21] , \wRegInA25[4] , \ScanLink8[29] , 
        \wRegInA30[15] , \ScanLink8[30] , \wAMid19[19] , \wAIn21[23] , 
        \wBMid27[6] , \wBMid1[29] , \wBMid25[16] , \wRegInA26[7] , 
        \ScanLink39[16] , \wBIn2[31] , \wAIn4[15] , \wBMid13[13] , 
        \ScanLink59[12] , \wBMid30[22] , \wRegInB6[2] , \wBIn2[28] , 
        \wBIn4[0] , \wBIn17[7] , \wRegInB1[24] , \wRegInA7[21] , 
        \wRegInA18[28] , \ScanLink3[25] , \wBIn7[3] , \wAMid24[10] , 
        \wRegInA18[31] , \wRegInB24[8] , \ScanLink19[6] , \wAMid12[15] , 
        \wBIn14[4] , \wAIn16[0] , \wRegInB1[17] , \ScanLink3[16] , 
        \wRegInA7[12] , \wAMid12[26] , \wAIn15[3] , \wBMid21[8] , 
        \ScanLink64[28] , \ScanLink64[31] , \ScanLink32[30] , \ScanLink11[18] , 
        \ScanLink47[19] , \ScanLink32[29] , \wRegInB26[19] , \wRegInA20[9] , 
        \wAMid4[30] , \wAMid4[29] , \wBMid5[22] , \wAMid24[23] , \wAMid10[1] , 
        \wBIn12[15] , \wBMid17[18] , \ScanLink28[29] , \wBIn24[10] , 
        \ScanLink28[30] , \wAIn25[28] , \ScanLink26[8] , \wBIn31[24] , 
        \wAMid13[2] , \wAIn25[31] , \wRegInB18[5] , \wBIn12[26] , \wBIn28[9] , 
        \wBIn31[17] , \wRegInA8[26] , \ScanLink38[4] , \ScanLink3[0] , 
        \wBIn24[23] , \wBIn6[23] , \wBIn6[10] , \wBMid5[11] , \wAIn18[12] , 
        \wRegInA8[15] , \wRegInB14[17] , \wRegInA21[19] , \ScanLink0[3] , 
        \wRegInB22[12] , \wAMid20[31] , \wAMid20[28] , \wRegInA3[19] , 
        \ScanLink60[23] , \ScanLink56[26] , \ScanLink23[16] , \ScanLink20[6] , 
        \ScanLink43[12] , \ScanLink15[13] , \ScanLink36[22] , \ScanLink23[5] , 
        \wAIn8[6] , \wAIn18[21] , \wRegInA19[9] , \ScanLink60[10] , 
        \ScanLink15[20] , \ScanLink44[2] , \ScanLink36[11] , \ScanLink43[21] , 
        \ScanLink23[25] , \ScanLink56[15] , \wBIn19[19] , \wRegInB14[24] , 
        \wRegInB22[21] , \wBMid18[8] , \ScanLink47[1] , \wAIn16[9] , 
        \wRegInB3[6] , \wRegInA23[3] , \wRegInA18[12] , \wBIn2[12] , 
        \wBMid18[25] , \wBMid21[1] , \wBMid22[2] , \ScanLink64[21] , 
        \ScanLink63[7] , \ScanLink52[24] , \ScanLink47[10] , \ScanLink11[11] , 
        \ScanLink32[20] , \wRegInB0[5] , \wRegInB26[10] , \ScanLink60[4] , 
        \ScanLink27[14] , \wRegInA20[0] , \wBIn2[21] , \wRegInA7[31] , 
        \wRegInB10[15] , \wBIn4[9] , \wRegInA7[28] , \wRegInA18[21] , 
        \wAMid24[19] , \wRegInB10[26] , \wRegInB27[2] , \wRegInB24[1] , 
        \wRegInB26[23] , \wAMid0[18] , \wAMid9[8] , \wAIn10[7] , \wBMid18[16] , 
        \ScanLink52[17] , \ScanLink27[27] , \wRegInB5[8] , \ScanLink64[12] , 
        \ScanLink11[22] , \ScanLink47[23] , \ScanLink32[13] , \ScanLink8[20] , 
        \wAIn13[4] , \wRegInA25[31] , \wRegInA25[28] , \wBIn16[17] , 
        \wAMid19[10] , \wBIn20[12] , \wAIn1[27] , \wBIn1[4] , \wBIn2[7] , 
        \wBMid1[20] , \wBIn11[0] , \ScanLink8[13] , \wAMid29[8] , \wBMid0[19] , 
        \wBMid0[7] , \wBMid1[13] , \wBIn12[3] , \wBMid3[4] , \wBMid13[30] , 
        \wBMid13[29] , \wBMid30[18] , \ScanLink59[28] , \wBIn16[24] , 
        \wAMid19[23] , \wBIn20[21] , \ScanLink59[31] , \wAIn21[19] , 
        \wBIn19[8] , \wAMid21[0] , \wRegInB29[4] , \ScanLink46[29] , 
        \ScanLink33[19] , \ScanLink10[31] , \ScanLink10[28] , \wAMid13[16] , 
        \ScanLink46[30] , \wAMid22[3] , \wAMid25[13] , \wAMid30[27] , 
        \wRegInB0[27] , \wRegInB27[30] , \wRegInB27[29] , \ScanLink2[26] , 
        \wAMid1[0] , \wAMid2[3] , \wAMid13[25] , \wAMid25[20] , \wRegInA6[22] , 
        \ScanLink17[9] , \wBIn3[18] , \wAMid30[14] , \wRegInA6[11] , 
        \wRegInB0[14] , \wRegInA19[18] , \wAIn16[16] , \ScanLink2[15] , 
        \wAMid18[30] , \wAMid18[29] , \wAIn20[13] , \ScanLink12[4] , 
        \wAMid1[21] , \wAIn5[25] , \wBMid24[26] , \ScanLink38[26] , 
        \wBMid12[23] , \ScanLink58[22] , \wAMid1[12] , \wAIn5[16] , 
        \wBMid6[9] , \wBIn8[14] , \wRegInB31[6] , \wRegInA24[11] , 
        \wRegInA31[25] , \ScanLink11[7] , \wRegInA12[14] , \ScanLink9[19] , 
        \wBIn8[27] , \wBMid12[10] , \ScanLink58[11] , \wAIn16[25] , 
        \wAIn20[20] , \wBMid24[15] , \ScanLink38[15] , \wBIn21[18] , 
        \wBMid29[9] , \wRegInA12[27] , \wRegInA28[8] , \wRegInA31[16] , 
        \wRegInA24[22] , \wBMid10[0] , \wRegInA16[16] , \ScanLink51[5] , 
        \wRegInA1[4] , \wRegInA20[13] , \wRegInA11[1] , \wAIn1[14] , 
        \wBMid4[31] , \wBMid4[28] , \wAMid5[23] , \wBMid16[21] , \wAIn12[27] , 
        \wAIn12[14] , \wBMid13[3] , \wBMid20[24] , \wRegInA2[7] , 
        \wRegInA12[2] , \ScanLink29[10] , \ScanLink49[14] , \wAIn24[11] , 
        \wBIn25[30] , \wBIn25[29] , \wAIn27[8] , \ScanLink52[6] , \wAIn31[25] , 
        \wRegInB28[14] , \wAIn31[16] , \wRegInB15[0] , \wRegInA16[25] , 
        \wRegInA20[20] , \ScanLink35[1] , \ScanLink36[2] , \wAIn24[22] , 
        \wRegInB28[27] , \wRegInB16[3] , \ScanLink49[27] , \wBMid20[17] , 
        \wAIn5[3] , \wAMid5[10] , \ScanLink29[23] , \wBIn7[30] , \wBIn7[29] , 
        \wBMid16[12] , \wRegInA2[20] , \wAIn22[5] , \wRegInB4[25] , \wAIn6[0] , 
        \wAMid17[14] , \wBIn18[13] , \wAMid21[11] , \ScanLink6[24] , 
        \ScanLink49[7] , \wRegInA4[9] , \ScanLink54[8] , \wAIn21[6] , 
        \wBIn23[2] , \ScanLink6[17] , \wRegInA2[13] , \wRegInB4[16] , 
        \wAIn0[25] , \wAIn0[6] , \wBMid0[22] , \wAMid1[8] , \wBIn3[10] , 
        \wAMid17[27] , \wBIn18[20] , \ScanLink61[30] , \ScanLink61[29] , 
        \ScanLink42[18] , \ScanLink37[28] , \ScanLink37[31] , \ScanLink14[19] , 
        \wAMid18[9] , \wBIn20[1] , \wAMid21[22] , \wRegInB23[18] , 
        \wAIn19[18] , \wRegInA6[19] , \wRegInA19[10] , \wBIn3[23] , \wBIn9[4] , 
        \wAIn18[7] , \wAMid25[31] , \wRegInB27[12] , \wBMid19[27] , 
        \wAMid25[28] , \wRegInA30[2] , \wRegInB11[17] , \ScanLink46[12] , 
        \ScanLink10[13] , \ScanLink33[22] , \wRegInA19[23] , \ScanLink53[26] , 
        \ScanLink26[16] , \ScanLink17[1] , \wAMid4[5] , \wAMid7[6] , 
        \wBIn19[0] , \ScanLink26[25] , \wBMid19[14] , \wAMid21[8] , 
        \ScanLink53[15] , \wBMid29[1] , \wRegInB8[5] , \wRegInB11[24] , 
        \ScanLink46[21] , \ScanLink33[11] , \ScanLink10[20] , \ScanLink14[2] , 
        \wRegInB27[21] , \wRegInA28[0] , \ScanLink9[22] , \wBMid12[18] , 
        \ScanLink58[19] , \wBMid0[11] , \wBMid5[2] , \wBMid6[1] , \wBIn17[15] , 
        \wAIn20[28] , \wAMid18[12] , \wAIn20[31] , \wBIn21[10] , \wAMid24[5] , 
        \wRegInA24[19] , \wBIn21[23] , \wAMid27[6] , \ScanLink9[11] , 
        \wBIn17[26] , \wAMid18[21] , \wAMid1[30] , \wAMid1[29] , \wBMid4[20] , 
        \wBIn13[17] , \wBIn25[12] , \wBIn30[26] , \wBMid4[13] , \wAMid5[18] , 
        \wBMid16[30] , \wBMid16[29] , \wBIn25[4] , \wBIn26[7] , \wRegInA9[24] , 
        \wRegInB15[8] , \ScanLink28[6] , \wRegInA20[31] , \wRegInA20[28] , 
        \ScanLink35[9] , \ScanLink29[18] , \wBIn13[24] , \wAIn24[19] , 
        \wBIn30[15] , \wAIn3[5] , \wAIn24[3] , \wBIn25[21] , \wAIn27[0] , 
        \wAIn6[8] , \wBIn7[12] , \wBMid10[8] , \wBIn18[31] , \wRegInA9[17] , 
        \wRegInA11[9] , \wRegInB15[15] , \ScanLink61[21] , \ScanLink57[24] , 
        \ScanLink30[4] , \ScanLink22[14] , \ScanLink42[10] , \ScanLink14[11] , 
        \ScanLink37[20] , \wBIn18[28] , \wRegInB10[5] , \wAMid18[1] , 
        \wAIn19[10] , \wRegInB23[10] , \wBIn20[9] , \wRegInB13[6] , 
        \ScanLink33[7] , \wBMid15[5] , \wAIn19[23] , \wAMid21[19] , 
        \wRegInB23[23] , \ScanLink8[3] , \wRegInA4[1] , \wRegInA14[4] , 
        \wRegInB15[26] , \ScanLink61[12] , \ScanLink14[22] , \ScanLink57[17] , 
        \ScanLink54[0] , \ScanLink42[23] , \ScanLink37[13] , \ScanLink22[27] , 
        \wBIn7[21] , \wRegInA2[31] , \ScanLink57[3] , \wAIn13[16] , 
        \wBMid16[6] , \wRegInA2[28] , \wAIn25[13] , \wAIn29[6] , \wRegInA7[2] , 
        \wRegInA17[7] , \wRegInA17[14] , \ScanLink41[7] , \wRegInA21[11] , 
        \ScanLink3[8] , \wAIn30[27] , \ScanLink42[4] , \wRegInB29[16] , 
        \wAIn0[16] , \wAMid4[21] , \wBMid17[23] , \wBMid5[19] , 
        \ScanLink48[16] , \ScanLink28[12] , \wAMid10[9] , \wBMid21[26] , 
        \wBIn28[1] , \wRegInA21[22] , \ScanLink25[3] , \wBMid21[15] , 
        \wRegInA17[27] , \ScanLink48[25] , \wBIn2[30] , \wBIn2[29] , 
        \wAMid4[12] , \ScanLink28[21] , \wBIn6[18] , \wAIn13[25] , 
        \wBMid17[10] , \wBIn24[18] , \wAIn30[14] , \ScanLink26[0] , 
        \wAMid16[16] , \wAIn18[30] , \wAIn25[20] , \wRegInB29[25] , 
        \wAIn31[4] , \wRegInA3[22] , \ScanLink7[26] , \ScanLink6[5] , 
        \wRegInB5[27] , \ScanLink47[9] , \wRegInA9[4] , \ScanLink60[18] , 
        \ScanLink43[30] , \ScanLink43[29] , \ScanLink36[19] , \ScanLink15[31] , 
        \ScanLink15[28] , \ScanLink5[6] , \wRegInA19[1] , \wAIn18[29] , 
        \wAMid20[13] , \wRegInB22[30] , \ScanLink59[5] , \wRegInB22[29] , 
        \wAMid16[7] , \wBIn19[11] , \wBMid18[0] , \wRegInB5[14] , 
        \wRegInA3[11] , \wBIn7[2] , \wAMid12[14] , \wAMid15[4] , \wAMid16[25] , 
        \ScanLink7[15] , \wBIn19[22] , \wAMid20[20] , \wBIn30[3] , \wBIn14[5] , 
        \wAMid24[11] , \wRegInB1[25] , \wRegInB24[9] , \ScanLink19[7] , 
        \wRegInA7[20] , \wBIn4[1] , \wRegInA18[30] , \wAIn15[2] , \wBIn17[6] , 
        \wRegInA18[29] , \ScanLink3[24] , \ScanLink64[30] , \wBMid21[9] , 
        \ScanLink64[29] , \ScanLink47[18] , \ScanLink32[28] , \ScanLink32[31] , 
        \ScanLink11[19] , \wAMid24[22] , \wRegInA20[8] , \wAMid12[27] , 
        \wRegInB26[18] , \wRegInA7[13] , \ScanLink3[17] , \wAMid0[23] , 
        \wAIn4[27] , \wBMid8[7] , \wAIn16[1] , \wBMid25[24] , \wRegInB1[16] , 
        \ScanLink39[24] , \wBMid30[10] , \wRegInB22[7] , \wBMid13[21] , 
        \ScanLink59[20] , \wAMid0[19] , \wAMid0[10] , \wAIn4[14] , \wBIn9[16] , 
        \wAIn17[14] , \wBIn20[30] , \wBIn20[29] , \wAIn21[11] , \wAMid29[0] , 
        \wRegInA13[16] , \wRegInA25[13] , \wRegInA30[27] , \wAMid9[0] , 
        \wBIn11[8] , \wAIn17[27] , \wAMid19[18] , \wRegInB21[4] , \wAIn21[22] , 
        \wBMid27[7] , \wBMid30[23] , \wRegInB6[3] , \wRegInA26[6] , 
        \wBMid1[31] , \wBMid1[28] , \wBMid13[12] , \ScanLink59[13] , 
        \ScanLink39[17] , \wBMid1[21] , \wAMid4[31] , \wBIn6[22] , \wBIn6[11] , 
        \wBIn9[25] , \wBMid25[17] , \wRegInB5[0] , \wRegInA25[5] , 
        \wBMid24[4] , \wRegInA30[14] , \ScanLink8[31] , \ScanLink8[28] , 
        \wRegInA3[18] , \wRegInA13[25] , \wRegInA25[20] , \wAIn8[7] , 
        \wAIn18[13] , \wAMid20[30] , \wAMid20[29] , \ScanLink23[4] , 
        \wRegInB22[13] , \wRegInB14[16] , \ScanLink60[22] , \ScanLink43[13] , 
        \ScanLink36[23] , \ScanLink56[27] , \ScanLink15[12] , \ScanLink23[17] , 
        \ScanLink20[7] , \wBMid5[23] , \wAMid10[0] , \wAIn18[20] , 
        \wBIn19[18] , \wRegInA19[8] , \ScanLink47[0] , \ScanLink60[11] , 
        \ScanLink56[14] , \ScanLink23[24] , \ScanLink44[3] , \ScanLink43[20] , 
        \ScanLink36[10] , \ScanLink15[21] , \wBMid18[9] , \wRegInB14[25] , 
        \wBIn28[8] , \wRegInB22[20] , \wBMid17[19] , \wRegInA8[27] , 
        \wRegInB18[4] , \ScanLink38[5] , \ScanLink28[31] , \ScanLink28[28] , 
        \wBMid5[10] , \wBIn12[27] , \wBIn12[14] , \wAMid13[3] , \wAIn25[30] , 
        \wBIn24[22] , \wBIn24[11] , \wAIn25[29] , \wBIn31[25] , \wRegInA8[14] , 
        \ScanLink26[9] , \wRegInA21[18] , \ScanLink0[2] , \ScanLink3[1] , 
        \wBIn31[16] , \wAMid4[28] , \wAMid9[9] , \wBIn20[13] , \wAIn13[5] , 
        \wBIn16[16] , \wAMid19[11] , \wBIn1[5] , \wBMid1[12] , \wAIn10[6] , 
        \wRegInB5[9] , \wRegInA25[30] , \wRegInA25[29] , \wBIn12[2] , 
        \wBMid13[31] , \wBMid30[19] , \ScanLink8[21] , \ScanLink59[30] , 
        \wBMid13[28] , \ScanLink59[29] , \wBIn2[6] , \wBIn16[25] , 
        \wAMid19[22] , \wBIn20[20] , \wAIn21[18] , \wAMid29[9] , 
        \ScanLink8[12] , \wBIn11[1] , \wBMid18[24] , \wBMid21[0] , 
        \ScanLink64[20] , \ScanLink60[5] , \ScanLink52[25] , \ScanLink47[11] , 
        \ScanLink27[15] , \ScanLink32[21] , \ScanLink11[10] , \wRegInB10[14] , 
        \wBIn2[13] , \wRegInB0[4] , \wRegInA20[1] , \wRegInB3[7] , 
        \wRegInA18[13] , \wRegInB26[11] , \wRegInA23[2] , \ScanLink63[6] , 
        \wBMid22[3] , \wAIn16[8] , \wAMid24[18] , \wBMid0[18] , \wAMid1[20] , 
        \wBIn2[20] , \wBMid18[17] , \wRegInB10[27] , \wRegInB24[0] , 
        \wRegInB26[22] , \ScanLink64[13] , \ScanLink47[22] , \ScanLink32[12] , 
        \ScanLink11[23] , \ScanLink27[26] , \ScanLink52[16] , \wBIn4[8] , 
        \wRegInA7[30] , \wRegInA7[29] , \wRegInB27[3] , \wBMid6[8] , 
        \wBIn8[15] , \wRegInB31[7] , \wRegInA18[20] , \wRegInA12[15] , 
        \wBMid12[22] , \wAIn16[17] , \wAMid18[31] , \wRegInA24[10] , 
        \wRegInA31[24] , \ScanLink9[18] , \ScanLink11[6] , \wAMid18[28] , 
        \wAIn20[12] , \ScanLink12[5] , \ScanLink58[23] , \wAIn5[24] , 
        \wBMid24[27] , \ScanLink38[27] , \wBMid0[6] , \wAMid1[13] , 
        \wBIn8[26] , \wRegInA12[26] , \wRegInA24[23] , \wRegInA28[9] , 
        \wRegInA31[17] , \wBMid24[14] , \wBMid29[8] , \ScanLink38[14] , 
        \wAIn5[17] , \wBMid12[11] , \ScanLink58[10] , \wAIn16[24] , 
        \wAIn20[21] , \wBIn21[19] , \ScanLink17[8] , \ScanLink2[27] , 
        \wAMid1[1] , \wBIn3[19] , \wBMid3[5] , \wAMid22[2] , \wRegInA6[23] , 
        \wRegInB0[26] , \ScanLink10[29] , \wAMid13[17] , \wBIn19[9] , 
        \wRegInB29[5] , \ScanLink46[31] , \ScanLink46[28] , \ScanLink33[18] , 
        \ScanLink10[30] , \wAMid21[1] , \wAMid25[12] , \wRegInB27[28] , 
        \wAMid30[26] , \wRegInB27[31] , \wRegInB0[15] , \wRegInA6[10] , 
        \wRegInA19[19] , \wAMid2[2] , \wAMid30[15] , \ScanLink2[14] , 
        \wAIn5[2] , \wAIn6[1] , \wAMid13[24] , \wAMid17[15] , \wAMid25[21] , 
        \wBIn18[12] , \wRegInA4[8] , \wAIn21[7] , \wAMid21[10] , 
        \ScanLink49[6] , \ScanLink54[9] , \wBIn7[31] , \wAIn22[4] , 
        \wRegInB4[24] , \wBIn7[28] , \wRegInA2[21] , \ScanLink61[31] , 
        \ScanLink61[28] , \ScanLink6[25] , \ScanLink37[30] , \ScanLink14[18] , 
        \ScanLink42[19] , \ScanLink37[29] , \wAMid0[27] , \wAIn1[26] , 
        \wAMid5[22] , \wBMid16[20] , \wAMid17[26] , \wAMid18[8] , 
        \wRegInB23[19] , \wAIn19[19] , \wBIn20[0] , \wAMid21[23] , 
        \wBIn18[21] , \wBMid20[25] , \wBIn23[3] , \wRegInA2[12] , 
        \ScanLink6[16] , \wRegInB4[17] , \wRegInA2[6] , \wRegInA12[3] , 
        \ScanLink49[15] , \ScanLink29[11] , \wAIn1[15] , \wAMid5[11] , 
        \wBMid10[1] , \wAIn12[15] , \wRegInB28[15] , \wBMid13[2] , 
        \wAIn24[10] , \wBIn25[31] , \wBIn25[28] , \wAIn27[9] , \wAIn31[24] , 
        \wRegInA20[12] , \ScanLink52[7] , \wAIn12[26] , \wAIn24[23] , 
        \wRegInA1[5] , \wRegInA11[0] , \wRegInA16[17] , \ScanLink51[4] , 
        \wAIn31[17] , \wRegInB28[26] , \ScanLink36[3] , \ScanLink29[22] , 
        \wBMid16[13] , \wBMid4[30] , \wRegInB16[2] , \wBMid4[29] , 
        \wBMid20[16] , \wBIn9[12] , \wAMid29[4] , \wRegInB15[1] , 
        \ScanLink49[26] , \wRegInA16[24] , \wRegInA20[21] , \ScanLink35[0] , 
        \wRegInB21[0] , \wBMid13[25] , \wBIn16[31] , \wRegInA13[12] , 
        \wRegInA25[17] , \wRegInA30[23] , \wBIn16[28] , \wAIn21[15] , 
        \wAIn17[10] , \ScanLink59[24] , \wAMid0[14] , \wBIn1[8] , \wAIn4[23] , 
        \wBMid8[3] , \wBMid30[14] , \wRegInB22[3] , \wBMid25[20] , 
        \ScanLink39[20] , \wBIn9[21] , \wBMid24[0] , \wRegInA13[21] , 
        \wRegInA25[24] , \wRegInA30[10] , \wBMid25[13] , \wRegInB5[4] , 
        \wRegInA25[1] , \wRegInA26[2] , \ScanLink39[13] , \wAIn4[10] , 
        \wBMid13[16] , \ScanLink59[17] , \wBIn4[5] , \wAMid9[4] , \wAIn17[23] , 
        \wBMid30[27] , \wRegInB6[7] , \wAIn13[8] , \wAIn21[26] , \wBMid27[3] , 
        \ScanLink3[20] , \wBIn7[6] , \wBIn14[1] , \wBIn17[2] , \wAMid24[15] , 
        \wRegInB1[21] , \wRegInA7[24] , \ScanLink19[3] , \wAMid12[10] , 
        \wAIn16[5] , \wRegInB1[12] , \wRegInA7[17] , \wAIn0[21] , \wAMid4[25] , 
        \wAMid12[23] , \wRegInB10[19] , \ScanLink3[13] , \wAIn15[6] , 
        \wBMid18[30] , \wBMid18[29] , \wAMid24[26] , \wRegInB0[9] , 
        \ScanLink60[8] , \ScanLink52[28] , \ScanLink27[18] , \ScanLink52[31] , 
        \wAMid15[0] , \wAMid16[12] , \wBIn19[15] , \wRegInB14[28] , 
        \wBMid18[4] , \wAMid20[17] , \wRegInB14[31] , \wAIn31[0] , 
        \wRegInA19[5] , \ScanLink59[1] , \ScanLink23[29] , \wRegInA3[26] , 
        \wRegInB5[23] , \wRegInA9[0] , \ScanLink56[19] , \ScanLink23[30] , 
        \ScanLink5[2] , \ScanLink6[1] , \ScanLink7[22] , \wAMid16[21] , 
        \wBIn19[26] , \wAMid20[24] , \wBIn30[7] , \wAMid16[3] , 
        \ScanLink7[11] , \wBMid17[27] , \wBMid21[22] , \wRegInA3[15] , 
        \wRegInB5[10] , \ScanLink23[9] , \ScanLink48[12] , \ScanLink28[16] , 
        \wAIn0[12] , \wAMid4[16] , \wBIn12[19] , \wAIn13[12] , \wRegInB29[12] , 
        \wAIn25[24] , \wAIn25[17] , \wAIn30[23] , \wAIn29[2] , \wRegInA17[10] , 
        \wRegInA21[15] , \ScanLink42[0] , \ScanLink41[3] , \wBIn31[28] , 
        \wRegInA8[19] , \wBIn31[31] , \wAIn13[21] , \wAIn30[10] , 
        \wRegInB29[21] , \ScanLink28[25] , \ScanLink26[4] , \wBMid17[14] , 
        \wBIn7[16] , \wBMid21[11] , \wBIn28[5] , \wRegInA17[23] , 
        \ScanLink48[21] , \ScanLink38[8] , \wRegInB18[9] , \wRegInA21[26] , 
        \ScanLink25[7] , \wAMid18[5] , \wRegInB13[2] , \ScanLink33[3] , 
        \wAIn19[14] , \wRegInB23[14] , \wRegInB10[1] , \wRegInB15[11] , 
        \ScanLink61[25] , \ScanLink42[14] , \ScanLink37[24] , \ScanLink14[15] , 
        \wAIn0[2] , \wAIn1[18] , \wBIn7[25] , \wBMid16[2] , \wAIn22[9] , 
        \wRegInA7[6] , \wRegInA17[3] , \ScanLink57[20] , \ScanLink30[0] , 
        \ScanLink22[10] , \ScanLink6[31] , \ScanLink6[28] , \wRegInB4[29] , 
        \wRegInB4[30] , \wBMid15[1] , \ScanLink57[7] , \wAMid17[18] , 
        \ScanLink61[16] , \ScanLink57[13] , \ScanLink22[23] , \ScanLink54[4] , 
        \ScanLink42[27] , \ScanLink37[17] , \ScanLink14[26] , \wAIn19[27] , 
        \wRegInA4[5] , \wRegInA14[0] , \wRegInB15[22] , \wBIn25[0] , 
        \wRegInA16[30] , \wRegInB23[27] , \ScanLink8[7] , \wRegInA16[29] , 
        \wRegInA9[20] , \ScanLink28[2] , \wAIn3[1] , \wBMid4[24] , \wBIn26[3] , 
        \wBIn13[13] , \wBIn25[16] , \wBIn30[22] , \wRegInA1[8] , 
        \wRegInA9[13] , \wAIn12[18] , \wAIn24[7] , \wBIn25[25] , \wAIn27[4] , 
        \ScanLink51[9] , \wAIn31[29] , \wAIn31[30] , \wRegInB28[18] , 
        \wAIn1[22] , \wBMid0[26] , \wBMid4[17] , \wBIn13[20] , \wBMid20[31] , 
        \wBIn30[11] , \ScanLink49[18] , \wAIn16[30] , \wBIn21[14] , 
        \wBMid20[28] , \wAIn16[29] , \wBIn17[11] , \wAMid18[16] , 
        \ScanLink38[19] , \wBMid0[15] , \wAMid4[1] , \wAIn5[30] , \wAIn5[29] , 
        \wAMid7[2] , \wBMid24[19] , \wBMid29[5] , \wRegInB8[1] , 
        \wRegInA28[4] , \ScanLink9[26] , \wAIn3[8] , \wBIn3[27] , \wBIn3[14] , 
        \wBMid5[6] , \wBMid6[5] , \wBIn17[22] , \wAMid18[25] , \wBIn21[27] , 
        \ScanLink12[8] , \wAMid27[2] , \wRegInA12[18] , \wRegInA31[30] , 
        \wRegInA31[29] , \wBIn8[18] , \wAMid24[1] , \ScanLink9[15] , 
        \wAMid13[30] , \wAMid13[29] , \wBMid19[23] , \ScanLink53[22] , 
        \ScanLink46[16] , \ScanLink26[12] , \ScanLink33[26] , \ScanLink10[17] , 
        \wAMid30[18] , \wRegInB11[13] , \wAIn18[3] , \wRegInB0[18] , 
        \wRegInA19[14] , \wRegInB27[16] , \wRegInA30[6] , \ScanLink2[19] , 
        \wBMid3[8] , \wRegInB11[20] , \wRegInB27[25] , \ScanLink46[25] , 
        \ScanLink33[15] , \ScanLink14[6] , \wBIn19[4] , \wRegInB29[8] , 
        \ScanLink10[24] , \ScanLink26[21] , \wBMid19[10] , \ScanLink53[11] , 
        \wBIn9[0] , \ScanLink17[5] , \wRegInA1[1] , \wRegInA19[27] , 
        \wRegInA11[4] , \wRegInA16[13] , \ScanLink51[0] , \wBMid10[5] , 
        \wAIn12[11] , \wBIn13[30] , \wBIn13[29] , \wRegInA20[16] , 
        \wAIn24[14] , \wBMid13[6] , \wBIn30[18] , \wAIn31[20] , 
        \ScanLink52[3] , \wRegInB28[11] , \wAIn1[11] , \wAMid5[26] , 
        \wBMid16[24] , \wBMid20[21] , \wRegInA12[7] , \ScanLink49[11] , 
        \ScanLink29[15] , \wBMid20[12] , \wBIn25[9] , \wRegInA2[2] , 
        \wRegInA9[30] , \wRegInA9[29] , \wRegInB15[5] , \wRegInA16[20] , 
        \wRegInA20[25] , \ScanLink35[4] , \wRegInB16[6] , \ScanLink49[22] , 
        \wAIn5[6] , \wAMid5[15] , \ScanLink29[26] , \wAIn12[22] , 
        \wBMid16[17] , \wAIn31[13] , \ScanLink36[7] , \wAIn22[0] , 
        \wAIn24[27] , \wRegInB28[22] , \wRegInA2[25] , \ScanLink6[21] , 
        \wRegInB4[20] , \wAIn6[5] , \wBMid15[8] , \wAMid17[22] , \wAMid17[11] , 
        \wBIn18[16] , \wAIn21[3] , \wAMid21[14] , \ScanLink49[2] , 
        \wBIn18[25] , \wBIn23[7] , \wRegInA2[16] , \wRegInB4[13] , 
        \wRegInA14[9] , \ScanLink6[12] , \wRegInB10[8] , \wBIn20[4] , 
        \wAMid21[27] , \wRegInB15[18] , \ScanLink57[30] , \ScanLink57[29] , 
        \wBMid0[2] , \wBMid3[1] , \wAMid13[13] , \ScanLink30[9] , 
        \ScanLink22[19] , \wBMid19[19] , \wAMid21[5] , \wAMid25[16] , 
        \wAMid30[22] , \wRegInB11[30] , \wRegInB11[29] , \ScanLink26[31] , 
        \ScanLink26[28] , \ScanLink53[18] , \wBIn9[9] , \wRegInB29[1] , 
        \wAMid22[6] , \wRegInB0[22] , \wAMid1[24] , \wAMid1[5] , \wAMid2[6] , 
        \wAMid25[25] , \wRegInA6[27] , \ScanLink2[23] , \wAMid13[20] , 
        \wAMid30[11] , \wAIn5[20] , \wBMid24[23] , \wRegInB0[11] , 
        \wRegInA6[14] , \ScanLink2[10] , \ScanLink38[23] , \wBMid12[26] , 
        \ScanLink58[27] , \wAMid1[17] , \wAIn5[13] , \wBIn8[11] , \wAIn16[13] , 
        \wAIn20[16] , \wAMid24[8] , \ScanLink12[1] , \wRegInA12[11] , 
        \wRegInA24[14] , \wRegInA31[20] , \ScanLink11[2] , \wAIn16[20] , 
        \wBIn17[18] , \wRegInB31[3] , \wAIn20[25] , \wBIn2[17] , \wAMid4[8] , 
        \wBMid12[15] , \ScanLink58[14] , \wBMid24[10] , \ScanLink38[10] , 
        \wBIn8[22] , \wRegInB8[8] , \wRegInA31[13] , \wRegInA12[22] , 
        \wRegInA24[27] , \wBMid22[7] , \wRegInB0[0] , \wRegInB3[3] , 
        \wRegInA23[6] , \ScanLink63[2] , \wRegInA18[17] , \wRegInB26[15] , 
        \wBIn2[24] , \wBMid18[20] , \wBMid21[4] , \wRegInB10[10] , 
        \wRegInA20[5] , \ScanLink64[24] , \ScanLink11[14] , \ScanLink52[21] , 
        \ScanLink47[15] , \ScanLink32[25] , \wRegInB1[31] , \wRegInA18[24] , 
        \ScanLink60[1] , \ScanLink27[11] , \ScanLink3[29] , \wRegInB27[7] , 
        \ScanLink3[30] , \wRegInB1[28] , \wAMid12[19] , \wBIn14[8] , 
        \wBMid18[13] , \ScanLink52[12] , \ScanLink27[22] , \wRegInB10[23] , 
        \ScanLink64[17] , \ScanLink11[27] , \ScanLink47[26] , \ScanLink32[16] , 
        \wRegInB24[4] , \wRegInB26[26] , \wAIn0[31] , \wBIn1[1] , \wBIn2[2] , 
        \wBMid1[25] , \wAIn4[19] , \wBIn9[31] , \wAIn10[2] , \wBMid24[9] , 
        \ScanLink8[25] , \wRegInA13[28] , \wRegInA13[31] , \wRegInA25[8] , 
        \wRegInA30[19] , \wBIn9[28] , \wAIn13[1] , \wBIn16[12] , \wAMid19[15] , 
        \wBIn20[17] , \wBMid1[16] , \wBIn11[5] , \wBIn12[6] , \wBIn16[21] , 
        \wAIn17[19] , \wRegInB21[9] , \ScanLink8[16] , \wAMid19[26] , 
        \wBIn20[24] , \wBMid25[30] , \wBMid25[29] , \ScanLink39[30] , 
        \ScanLink39[29] , \wBMid5[27] , \wBIn12[10] , \wAIn13[31] , 
        \wAIn13[28] , \wRegInB29[28] , \wBIn24[15] , \wAIn30[19] , 
        \wBIn31[21] , \wRegInB29[31] , \wAMid13[7] , \wBMid21[18] , 
        \ScanLink48[31] , \wAMid10[4] , \wRegInA8[23] , \ScanLink48[28] , 
        \ScanLink38[1] , \wRegInB18[0] , \wAIn0[28] , \wBIn6[26] , \wBIn6[15] , 
        \wBMid5[14] , \wBIn12[23] , \wBIn31[12] , \ScanLink42[9] , 
        \ScanLink3[5] , \wAMid15[9] , \wBIn24[26] , \wRegInA8[10] , 
        \wRegInA17[19] , \ScanLink0[6] , \ScanLink60[26] , \ScanLink56[23] , 
        \ScanLink23[13] , \ScanLink20[3] , \wAMid16[31] , \wRegInB14[12] , 
        \ScanLink43[17] , \ScanLink15[16] , \ScanLink36[27] , \wAMid16[28] , 
        \wAIn18[17] , \wRegInB22[17] , \wRegInB5[19] , \ScanLink7[18] , 
        \ScanLink23[0] , \wAIn18[24] , \wAIn31[9] , \wRegInB14[21] , 
        \wRegInB22[24] , \ScanLink59[8] , \ScanLink60[15] , \ScanLink15[25] , 
        \ScanLink44[7] , \ScanLink43[24] , \ScanLink36[14] , \wRegInA9[9] , 
        \ScanLink56[10] , \ScanLink23[20] , \ScanLink47[4] , \ScanLink6[8] , 
        \wAIn8[3] , \wAMid12[31] , \wBMid18[22] , \ScanLink60[3] , 
        \ScanLink27[13] , \wBMid21[6] , \ScanLink52[23] , \ScanLink11[16] , 
        \ScanLink64[26] , \ScanLink47[17] , \ScanLink32[27] , \wAMid12[28] , 
        \wRegInB10[12] , \wRegInB0[2] , \wRegInB26[17] , \wBIn2[15] , 
        \wBMid22[5] , \wRegInB1[19] , \wRegInB3[1] , \wRegInA18[15] , 
        \wRegInA20[7] , \ScanLink3[18] , \wRegInA23[4] , \ScanLink63[0] , 
        \wRegInB24[6] , \wRegInB26[24] , \wAIn0[19] , \wBIn1[3] , \wBIn2[26] , 
        \wBMid18[11] , \wRegInB10[21] , \ScanLink19[8] , \ScanLink64[15] , 
        \ScanLink47[24] , \ScanLink11[25] , \ScanLink32[14] , \ScanLink52[10] , 
        \ScanLink27[20] , \wBMid1[27] , \wAIn13[3] , \wAIn17[31] , 
        \wAIn17[28] , \wBIn17[9] , \wRegInA18[26] , \wRegInB27[5] , 
        \wBIn20[15] , \wBIn16[10] , \wBMid27[8] , \wAMid19[17] , \wBMid25[18] , 
        \wBMid1[14] , \wAIn4[31] , \wAIn10[0] , \wRegInA26[9] , 
        \ScanLink39[18] , \ScanLink8[27] , \wAIn4[28] , \wBMid8[8] , 
        \wRegInB22[8] , \wBIn12[4] , \wBIn2[0] , \wBIn16[23] , \wAMid19[24] , 
        \wBIn20[26] , \wRegInA13[19] , \ScanLink8[14] , \wRegInA30[31] , 
        \wRegInA30[28] , \wBIn9[19] , \wBIn11[7] , \wAMid10[6] , 
        \wRegInA17[28] , \wRegInA8[21] , \wRegInA17[31] , \wRegInB18[2] , 
        \ScanLink38[3] , \wAIn0[9] , \wAIn1[20] , \wBIn6[24] , \wBIn6[17] , 
        \wBMid5[25] , \wBMid5[16] , \wBIn12[21] , \wBIn12[12] , \wAMid13[5] , 
        \wBIn31[23] , \wAIn13[19] , \wBIn24[17] , \wAIn29[9] , \wRegInA8[12] , 
        \ScanLink41[8] , \ScanLink0[4] , \wBIn24[24] , \wAIn30[31] , 
        \wRegInB29[19] , \wAIn30[28] , \wBIn31[10] , \wBMid21[29] , 
        \ScanLink3[7] , \wBMid21[30] , \ScanLink48[19] , \wAIn8[1] , 
        \wAMid16[8] , \wAIn18[15] , \ScanLink23[2] , \wRegInB14[10] , 
        \wRegInB22[15] , \ScanLink60[24] , \ScanLink15[14] , \ScanLink56[21] , 
        \ScanLink43[15] , \ScanLink36[25] , \ScanLink23[11] , \ScanLink20[1] , 
        \wRegInB5[31] , \ScanLink7[30] , \ScanLink7[29] , \wRegInB5[28] , 
        \ScanLink47[6] , \wAMid16[19] , \wRegInB14[23] , \ScanLink60[17] , 
        \ScanLink56[12] , \ScanLink23[22] , \ScanLink44[5] , \ScanLink43[26] , 
        \ScanLink15[27] , \ScanLink5[9] , \ScanLink36[16] , \wAIn18[26] , 
        \wRegInB22[26] , \wBMid20[23] , \wRegInA12[5] , \ScanLink49[13] , 
        \wRegInA2[0] , \wAMid5[24] , \ScanLink29[17] , \wAIn12[13] , 
        \wBMid16[26] , \wAIn31[22] , \wBMid13[4] , \wAIn1[13] , \wBMid10[7] , 
        \wAIn24[16] , \wRegInB28[13] , \ScanLink52[1] , \wAIn12[20] , 
        \wBIn13[18] , \wRegInA1[3] , \wRegInA9[18] , \wRegInA16[11] , 
        \wRegInA20[14] , \ScanLink51[2] , \wRegInA11[6] , \wAIn24[25] , 
        \wBIn30[30] , \wBIn30[29] , \wAIn31[11] , \ScanLink36[5] , 
        \wRegInB28[20] , \wAIn5[4] , \wAMid5[17] , \wBMid16[15] , \wBIn26[8] , 
        \wAIn6[7] , \wAMid17[13] , \wBMid20[10] , \ScanLink49[20] , 
        \ScanLink29[24] , \wRegInB15[30] , \wRegInB15[7] , \wRegInB16[4] , 
        \wRegInA16[22] , \ScanLink28[9] , \wRegInA20[27] , \ScanLink35[6] , 
        \wBIn18[14] , \wAMid21[16] , \wRegInB15[29] , \ScanLink49[0] , 
        \wAIn21[1] , \ScanLink57[18] , \ScanLink22[31] , \ScanLink22[28] , 
        \wAIn22[2] , \wRegInB4[22] , \wBMid16[9] , \wRegInA2[27] , 
        \wRegInA17[8] , \ScanLink6[23] , \wAIn0[0] , \wAIn1[30] , \wAIn1[29] , 
        \wBMid0[0] , \wAMid17[20] , \wBIn20[6] , \wAMid21[25] , \wBIn18[27] , 
        \wBIn23[5] , \wRegInA2[14] , \wRegInB13[9] , \ScanLink6[10] , 
        \wRegInB4[11] , \ScanLink33[8] , \wRegInA6[25] , \ScanLink2[21] , 
        \wAMid1[26] , \wAMid1[7] , \wBMid3[3] , \wAMid22[4] , \wRegInB0[20] , 
        \wAMid13[11] , \wAMid21[7] , \wRegInB29[3] , \wAMid25[14] , 
        \wAMid30[20] , \wRegInB0[13] , \wRegInA6[16] , \ScanLink2[12] , 
        \wAMid2[4] , \wAIn5[22] , \wBIn8[13] , \wAMid13[22] , \wAIn18[8] , 
        \wAMid25[27] , \wAMid30[13] , \wRegInB11[18] , \wBMid19[31] , 
        \ScanLink53[30] , \wBMid19[28] , \ScanLink53[29] , \ScanLink26[19] , 
        \wRegInB31[1] , \wAIn16[11] , \wBIn17[30] , \wBIn17[29] , 
        \wRegInA12[13] , \wRegInA31[22] , \ScanLink11[0] , \wRegInA24[16] , 
        \wAIn20[14] , \ScanLink12[3] , \wAMid27[9] , \wAMid1[15] , \wAIn5[11] , 
        \wAMid7[9] , \wBMid12[24] , \wBMid24[21] , \ScanLink58[25] , 
        \ScanLink38[21] , \wRegInA12[20] , \wRegInA24[25] , \wRegInA31[11] , 
        \wBIn8[20] , \wBMid24[12] , \ScanLink38[12] , \wBMid12[17] , 
        \ScanLink58[16] , \wBMid4[26] , \wBIn7[27] , \wBIn7[14] , \wAIn16[22] , 
        \wAMid17[30] , \wAMid17[29] , \wAIn20[27] , \ScanLink61[27] , 
        \ScanLink57[22] , \ScanLink30[2] , \ScanLink22[12] , \ScanLink42[16] , 
        \ScanLink37[26] , \ScanLink14[17] , \wRegInB10[3] , \wAMid18[7] , 
        \wAIn19[16] , \wRegInB15[13] , \wRegInB23[16] , \wRegInB4[18] , 
        \wRegInB13[0] , \ScanLink6[19] , \ScanLink33[1] , \wBMid15[3] , 
        \wAIn19[25] , \wRegInB23[25] , \ScanLink49[9] , \wRegInA4[7] , 
        \ScanLink8[5] , \wRegInA14[2] , \wRegInB15[20] , \ScanLink61[14] , 
        \ScanLink54[6] , \ScanLink42[25] , \ScanLink37[15] , \ScanLink14[24] , 
        \wAIn21[8] , \ScanLink57[11] , \ScanLink22[21] , \wAIn12[30] , 
        \wBMid16[0] , \ScanLink57[5] , \wBIn25[14] , \wAIn31[18] , 
        \wRegInA7[4] , \wRegInA17[1] , \wRegInB28[30] , \wAIn12[29] , 
        \wRegInB28[29] , \wBIn13[11] , \wBIn30[20] , \ScanLink49[29] , 
        \wBMid20[19] , \ScanLink49[30] , \wBIn25[2] , \wBIn26[1] , 
        \wRegInA9[22] , \ScanLink28[0] , \wBMid4[15] , \wBIn13[22] , 
        \wRegInA2[9] , \wBIn25[27] , \wBIn30[13] , \ScanLink52[8] , 
        \wAIn27[6] , \wAMid0[25] , \wBMid0[24] , \wAIn3[3] , \wRegInA16[18] , 
        \wAIn5[18] , \wAMid7[0] , \wAIn24[5] , \wBMid29[7] , \wRegInB8[3] , 
        \wRegInA9[11] , \wRegInA12[30] , \wRegInA31[18] , \wRegInA12[29] , 
        \wRegInA28[6] , \ScanLink9[24] , \wBIn8[30] , \wBIn8[29] , 
        \wBMid0[17] , \wAMid4[3] , \wBMid5[4] , \wBMid6[7] , \wBIn17[13] , 
        \wAMid18[14] , \wBIn21[16] , \wAMid24[3] , \wRegInB31[8] , 
        \ScanLink11[9] , \ScanLink9[17] , \wAIn16[18] , \wBIn21[25] , 
        \wBIn17[20] , \wAMid27[0] , \wAMid18[27] , \wBMid0[9] , \wBIn3[25] , 
        \wBIn3[16] , \wBMid24[31] , \ScanLink38[28] , \wBMid24[28] , 
        \ScanLink38[31] , \wBIn9[2] , \wAIn18[1] , \wRegInA19[16] , 
        \wBMid19[21] , \wRegInB11[11] , \wRegInB27[14] , \wRegInA30[4] , 
        \ScanLink46[14] , \ScanLink33[24] , \ScanLink26[10] , \ScanLink10[15] , 
        \wRegInA19[25] , \ScanLink53[20] , \ScanLink2[31] , \ScanLink2[28] , 
        \wRegInB0[30] , \wRegInB0[29] , \wAMid13[18] , \wBIn19[6] , 
        \ScanLink17[7] , \wBMid19[12] , \wAMid30[30] , \ScanLink53[13] , 
        \ScanLink46[27] , \ScanLink26[23] , \ScanLink33[17] , \ScanLink14[4] , 
        \ScanLink10[26] , \wBMid25[22] , \wAMid30[29] , \wRegInB11[22] , 
        \wRegInB27[27] , \ScanLink39[22] , \wBIn2[9] , \wAIn4[21] , 
        \wBMid13[27] , \ScanLink59[26] , \wBMid8[1] , \wAIn17[12] , 
        \wBMid30[16] , \wRegInB22[1] , \wAIn21[17] , \wRegInA13[10] , 
        \wRegInA25[15] , \wRegInA30[21] , \wAMid0[16] , \wBIn9[10] , 
        \wAMid9[6] , \wBIn16[19] , \wAIn21[24] , \wAMid29[6] , \wRegInB21[2] , 
        \wBMid27[1] , \wBMid13[14] , \wAIn17[21] , \ScanLink59[15] , 
        \wAIn4[12] , \wBMid30[25] , \wRegInA26[0] , \wRegInB6[5] , \wBIn4[7] , 
        \wBIn7[4] , \wBIn9[23] , \wBMid25[11] , \wRegInB5[6] , 
        \ScanLink39[11] , \wRegInA25[3] , \wAIn10[9] , \wBMid24[2] , 
        \wRegInA13[23] , \wRegInA30[12] , \wBIn14[3] , \wRegInB10[28] , 
        \wRegInA25[26] , \wAMid12[12] , \wRegInB10[31] , \wBMid18[18] , 
        \wAMid24[17] , \ScanLink19[1] , \ScanLink52[19] , \wRegInB1[23] , 
        \ScanLink27[30] , \ScanLink27[29] , \wRegInA7[26] , \ScanLink3[22] , 
        \wAMid12[21] , \wAIn15[4] , \wBIn17[0] , \wAMid24[24] , \wAIn16[7] , 
        \wRegInB3[8] , \ScanLink3[11] , \wAIn0[23] , \wAMid4[27] , \wAIn8[8] , 
        \wRegInB1[10] , \wRegInA7[15] , \ScanLink63[9] , \wBIn12[31] , 
        \wAMid15[2] , \wAMid16[23] , \wAMid16[10] , \wBMid18[6] , 
        \wAMid20[15] , \wAIn31[2] , \wRegInA3[24] , \ScanLink7[20] , 
        \wRegInB5[21] , \ScanLink6[3] , \wRegInA19[7] , \ScanLink5[0] , 
        \wRegInA9[2] , \ScanLink59[3] , \wAMid16[1] , \wBIn19[17] , 
        \wRegInA3[17] , \wRegInB5[12] , \wRegInB14[19] , \ScanLink7[13] , 
        \wBIn19[24] , \wAMid20[26] , \wBIn30[5] , \ScanLink56[31] , 
        \ScanLink56[28] , \ScanLink23[18] , \ScanLink20[8] , \wAIn29[0] , 
        \wBIn31[19] , \wRegInA17[12] , \wRegInA21[17] , \ScanLink41[1] , 
        \ScanLink42[2] , \wBIn12[28] , \wAIn25[15] , \wAIn13[10] , 
        \wAIn30[21] , \wRegInB29[10] , \ScanLink28[14] , \wBMid17[25] , 
        \wAIn0[10] , \wAMid4[14] , \wBMid17[16] , \wBMid21[20] , \wBMid21[13] , 
        \wBIn28[7] , \wRegInA17[21] , \wRegInA21[24] , \ScanLink48[10] , 
        \ScanLink25[5] , \wRegInA8[31] , \wRegInA8[28] , \ScanLink48[23] , 
        \ScanLink28[27] , \wBMid0[30] , \wAMid1[22] , \wAIn13[23] , 
        \wRegInB29[23] , \wAIn25[26] , \wAIn30[12] , \ScanLink26[6] , 
        \wBMid24[25] , \ScanLink38[25] , \wAMid1[11] , \wAIn5[26] , 
        \wBMid12[20] , \ScanLink58[21] , \wBMid5[9] , \wAIn16[15] , 
        \wAIn20[10] , \wBIn21[31] , \wBIn21[28] , \ScanLink12[7] , \wBIn8[17] , 
        \wRegInA12[17] , \wRegInA24[12] , \wRegInA31[26] , \ScanLink11[4] , 
        \wBMid12[13] , \wAIn16[26] , \wAMid18[19] , \wAIn20[23] , 
        \wRegInB31[5] , \ScanLink58[12] , \wAIn5[15] , \wBMid24[16] , 
        \wBMid0[29] , \wBMid0[4] , \wBIn3[31] , \wBMid3[7] , \wBIn8[24] , 
        \ScanLink38[16] , \wAMid13[15] , \wAMid30[24] , \wRegInA12[24] , 
        \wRegInA24[21] , \wRegInA31[15] , \ScanLink9[29] , \ScanLink9[30] , 
        \wAMid21[3] , \wAMid25[10] , \wAMid22[0] , \wRegInB29[7] , 
        \ScanLink14[9] , \wRegInB0[24] , \wBIn3[28] , \wRegInA6[21] , 
        \wAMid1[3] , \wAMid2[0] , \wAMid25[23] , \wRegInA19[31] , 
        \wRegInA19[28] , \ScanLink2[25] , \wRegInB27[19] , \ScanLink46[19] , 
        \ScanLink33[30] , \ScanLink10[18] , \ScanLink33[29] , \wAMid30[17] , 
        \wRegInA30[9] , \wAMid13[26] , \ScanLink2[16] , \wAIn5[0] , 
        \wRegInB0[17] , \wRegInA6[12] , \wRegInA2[23] , \wRegInA7[9] , 
        \ScanLink57[8] , \ScanLink6[27] , \wAIn6[3] , \wAIn21[5] , \wAIn22[6] , 
        \wRegInB4[26] , \ScanLink61[19] , \ScanLink42[31] , \ScanLink42[28] , 
        \ScanLink14[29] , \ScanLink37[18] , \ScanLink14[30] , \wBIn7[19] , 
        \wAMid17[17] , \wBIn18[10] , \wAIn19[31] , \wAIn19[28] , 
        \wRegInB23[28] , \wRegInB23[31] , \ScanLink49[4] , \ScanLink8[8] , 
        \wAMid21[12] , \wRegInB4[15] , \wAMid17[24] , \wBIn18[23] , 
        \wBIn23[1] , \wRegInA2[10] , \ScanLink6[14] , \wBIn20[2] , 
        \wAMid21[21] , \wAMid0[31] , \wAIn1[24] , \wAMid5[20] , \wBMid10[3] , 
        \wAIn24[8] , \wRegInA1[7] , \wRegInA11[2] , \wRegInA16[15] , 
        \ScanLink51[6] , \wRegInA20[10] , \wAIn12[17] , \wBMid13[0] , 
        \wAIn24[12] , \ScanLink52[5] , \wAIn31[26] , \wRegInB28[17] , 
        \ScanLink29[13] , \wBMid16[22] , \wAIn1[17] , \wBMid4[18] , 
        \wBMid20[27] , \wRegInA2[4] , \wAMid5[13] , \wBMid16[11] , 
        \wBMid20[14] , \wRegInA12[1] , \wRegInB15[3] , \wRegInA16[26] , 
        \wRegInA20[23] , \ScanLink49[17] , \ScanLink35[2] , \wRegInB16[0] , 
        \ScanLink49[24] , \ScanLink29[20] , \wBIn1[7] , \wBIn2[4] , 
        \wBMid1[23] , \wAMid4[19] , \wBIn6[20] , \wBIn6[13] , \wAIn12[24] , 
        \wRegInB28[24] , \wAIn18[11] , \wBIn19[30] , \wBIn19[29] , 
        \wAIn24[21] , \wBIn25[19] , \ScanLink36[1] , \wAIn31[15] , 
        \ScanLink60[20] , \ScanLink56[25] , \ScanLink23[15] , \ScanLink20[5] , 
        \ScanLink43[11] , \ScanLink36[21] , \ScanLink15[10] , \wBIn30[8] , 
        \wRegInB14[14] , \wRegInB22[11] , \ScanLink23[6] , \wAIn18[22] , 
        \wAMid20[18] , \wRegInB22[22] , \wRegInA3[29] , \wRegInB14[27] , 
        \ScanLink60[13] , \ScanLink44[1] , \ScanLink43[22] , \ScanLink36[12] , 
        \ScanLink56[16] , \ScanLink15[23] , \ScanLink23[26] , \wBMid5[21] , 
        \wAIn8[5] , \wRegInA3[30] , \ScanLink47[2] , \wBIn12[16] , 
        \wBIn24[13] , \wAMid13[1] , \wBIn31[27] , \wBMid5[12] , \wAMid10[2] , 
        \wRegInA8[25] , \wRegInB18[6] , \wRegInA21[30] , \ScanLink38[7] , 
        \wRegInA21[29] , \ScanLink25[8] , \wBMid17[31] , \wBMid17[28] , 
        \ScanLink28[19] , \wAIn10[4] , \wBIn12[25] , \wBIn24[20] , 
        \wAIn25[18] , \ScanLink3[3] , \wBIn31[14] , \wRegInA8[16] , 
        \ScanLink0[0] , \wBMid13[19] , \wBMid30[31] , \wBMid30[28] , 
        \ScanLink8[23] , \wRegInB6[8] , \ScanLink59[18] , \wAIn13[7] , 
        \wBIn16[14] , \wAMid19[13] , \wAIn21[30] , \wBIn20[11] , \wAIn21[29] , 
        \wBMid1[10] , \wBIn11[3] , \wBIn16[27] , \wAMid19[20] , \wBIn20[22] , 
        \wRegInA25[18] , \ScanLink8[10] , \wBIn12[0] , \wAMid0[28] , 
        \wBIn2[11] , \wBMid22[1] , \wAMid24[29] , \wRegInB3[5] , 
        \wRegInA7[18] , \ScanLink63[4] , \wRegInA18[11] , \wRegInA23[0] , 
        \wBIn2[22] , \wAIn15[9] , \wAMid24[30] , \wRegInA20[3] , \wRegInB0[6] , 
        \wRegInB10[16] , \wRegInB26[13] , \ScanLink32[23] , \wBMid18[26] , 
        \wBMid21[2] , \ScanLink47[13] , \ScanLink11[12] , \ScanLink64[22] , 
        \ScanLink60[7] , \ScanLink52[27] , \ScanLink27[17] , \wRegInA18[22] , 
        \wRegInB27[1] , \wBIn7[9] , \wBMid18[15] , \ScanLink52[14] , 
        \wRegInB10[25] , \ScanLink64[11] , \ScanLink47[20] , \ScanLink27[24] , 
        \ScanLink32[10] , \ScanLink11[21] , \wAIn0[27] , \wBMid21[24] , 
        \wRegInB24[2] , \wRegInB26[20] , \ScanLink48[14] , \wAIn0[14] , 
        \wAMid4[23] , \ScanLink28[10] , \wAIn13[27] , \wAIn13[14] , 
        \wBMid17[21] , \wBIn24[30] , \wBIn24[29] , \wAIn30[25] , \wAMid13[8] , 
        \wAIn25[11] , \wRegInB29[14] , \ScanLink42[6] , \wAIn29[4] , 
        \wRegInA17[16] , \wRegInA21[13] , \ScanLink41[5] , \ScanLink0[9] , 
        \wAIn25[22] , \wAIn30[16] , \ScanLink26[2] , \wRegInB29[27] , 
        \wBIn4[3] , \wAMid4[10] , \wBMid17[12] , \wBIn6[30] , \wBIn6[29] , 
        \wBMid5[31] , \wBMid5[28] , \ScanLink48[27] , \ScanLink28[23] , 
        \wBMid21[17] , \wAMid16[14] , \wBIn19[13] , \wBMid18[2] , \wBIn28[3] , 
        \wRegInA17[25] , \wRegInA21[20] , \ScanLink25[1] , \wAMid20[11] , 
        \ScanLink59[7] , \wAIn31[6] , \wRegInA9[6] , \wRegInA19[3] , 
        \wRegInA3[20] , \wRegInB5[25] , \ScanLink44[8] , \ScanLink5[4] , 
        \ScanLink6[7] , \wAMid15[6] , \ScanLink60[30] , \ScanLink43[18] , 
        \ScanLink36[28] , \ScanLink7[24] , \ScanLink60[29] , \ScanLink36[31] , 
        \ScanLink15[19] , \wAMid16[27] , \wAIn18[18] , \wAMid20[22] , 
        \wBIn30[1] , \wBIn19[20] , \wRegInB22[18] , \wAMid16[5] , 
        \wRegInA3[13] , \ScanLink7[17] , \wRegInB5[16] , \wRegInB27[8] , 
        \wBIn17[4] , \wRegInB1[27] , \wRegInA7[22] , \ScanLink3[26] , 
        \ScanLink64[18] , \ScanLink47[29] , \ScanLink32[19] , \ScanLink11[31] , 
        \ScanLink47[30] , \ScanLink11[28] , \wBIn2[18] , \wBIn7[0] , 
        \wAMid12[16] , \wAMid24[13] , \wRegInB26[30] , \ScanLink19[5] , 
        \wRegInB26[29] , \wBIn14[7] , \wRegInB1[14] , \wBMid22[8] , \wAIn0[4] , 
        \wAMid0[21] , \wAIn4[25] , \wBIn9[14] , \wAMid12[25] , \wAIn16[3] , 
        \wRegInA7[11] , \wRegInA18[18] , \ScanLink3[15] , \wRegInA23[9] , 
        \wAIn15[0] , \wAMid24[20] , \wRegInB21[6] , \wAIn17[16] , 
        \wAMid19[30] , \wAMid19[29] , \wAMid29[2] , \wRegInA13[14] , 
        \wRegInA30[25] , \ScanLink8[19] , \wRegInA25[11] , \wAIn21[13] , 
        \wBMid8[5] , \wBMid30[12] , \wRegInB22[5] , \wAMid0[12] , \wBMid1[19] , 
        \wBIn12[9] , \wBMid13[23] , \ScanLink59[22] , \wAIn4[16] , \wBIn9[27] , 
        \wBMid24[6] , \wBMid25[26] , \ScanLink39[26] , \wRegInA13[27] , 
        \wRegInA25[22] , \wRegInA30[16] , \wBMid25[15] , \wRegInB5[2] , 
        \wRegInA25[7] , \ScanLink39[15] , \wBMid30[21] , \wRegInB6[1] , 
        \wBMid13[10] , \ScanLink59[11] , \wBMid0[20] , \wAMid2[9] , 
        \wAMid9[2] , \wBIn20[18] , \wRegInA26[4] , \wAIn17[25] , \wBMid19[25] , 
        \wAIn21[20] , \wBMid27[5] , \ScanLink53[24] , \ScanLink26[14] , 
        \wRegInB11[15] , \ScanLink46[10] , \ScanLink33[20] , \ScanLink10[11] , 
        \wBIn3[21] , \wBIn3[12] , \wAIn18[5] , \wRegInB27[10] , 
        \wRegInA19[12] , \wRegInA30[0] , \wBIn19[2] , \wAMid25[19] , 
        \wRegInB27[23] , \wRegInB11[26] , \ScanLink46[23] , \ScanLink10[22] , 
        \ScanLink33[13] , \ScanLink14[0] , \wBMid19[16] , \ScanLink53[17] , 
        \wRegInA6[31] , \ScanLink26[27] , \wRegInA6[28] , \ScanLink17[3] , 
        \wAMid4[7] , \wBIn9[6] , \wAMid22[9] , \wBIn17[17] , \wAMid18[10] , 
        \wBIn21[12] , \wRegInA19[21] , \wBMid0[13] , \wAMid1[18] , \wAMid7[4] , 
        \wBMid12[30] , \wBMid12[29] , \wBMid29[3] , \wRegInB8[7] , 
        \wRegInA24[31] , \wRegInA24[28] , \ScanLink9[20] , \wRegInA28[2] , 
        \ScanLink58[28] , \ScanLink58[31] , \wAIn3[7] , \wBMid4[22] , 
        \wBMid5[0] , \wBIn17[24] , \wAMid18[23] , \wAIn20[19] , \wBMid6[3] , 
        \wBIn21[21] , \wAMid27[4] , \ScanLink9[13] , \wBMid16[18] , 
        \wAMid24[7] , \wBIn25[6] , \wBIn26[5] , \wRegInA9[26] , 
        \ScanLink28[4] , \wRegInB16[9] , \ScanLink29[30] , \ScanLink29[29] , 
        \wBIn13[15] , \wAIn24[28] , \wBIn30[24] , \wAIn24[31] , \wAIn24[1] , 
        \wBIn25[10] , \ScanLink36[8] , \wRegInA9[15] , \wRegInA20[19] , 
        \wBMid13[9] , \wRegInA0[3] , \wBIn1[27] , \wAIn5[9] , \wBMid4[11] , 
        \wBIn13[26] , \wBIn25[23] , \wAIn27[2] , \wBIn30[17] , \wAMid5[30] , 
        \wAMid5[29] , \wRegInA12[8] , \wBIn7[10] , \wAMid18[3] , \wAIn19[12] , 
        \wAMid21[31] , \wBIn23[8] , \wRegInA2[19] , \ScanLink33[5] , 
        \wRegInB13[4] , \wRegInB23[12] , \wAMid21[28] , \wRegInA7[0] , 
        \wRegInB10[7] , \wRegInB15[17] , \ScanLink61[23] , \ScanLink14[13] , 
        \ScanLink57[26] , \ScanLink42[12] , \ScanLink37[22] , \ScanLink30[6] , 
        \ScanLink22[16] , \wRegInA17[5] , \wBIn7[23] , \wBMid16[4] , 
        \ScanLink57[1] , \wAMid8[12] , \wBMid15[7] , \ScanLink57[15] , 
        \ScanLink22[25] , \wBIn18[19] , \wRegInA4[3] , \wRegInA14[6] , 
        \wRegInB15[24] , \ScanLink61[10] , \ScanLink54[2] , \ScanLink42[21] , 
        \ScanLink14[20] , \ScanLink37[11] , \wAIn19[21] , \wRegInB23[21] , 
        \wBIn28[18] , \wAIn29[20] , \wRegInB13[20] , \ScanLink8[1] , 
        \wRegInB14[7] , \wRegInB25[25] , \wRegInB30[11] , \ScanLink29[9] , 
        \ScanLink51[11] , \ScanLink44[25] , \ScanLink34[6] , \ScanLink24[21] , 
        \ScanLink12[24] , \ScanLink37[5] , \ScanLink31[15] , \wAMid8[21] , 
        \wBMid9[19] , \wBMid11[7] , \wBIn27[8] , \wRegInB17[4] , 
        \ScanLink12[17] , \ScanLink44[16] , \ScanLink31[26] , \ScanLink24[12] , 
        \wRegInB25[16] , \ScanLink51[22] , \ScanLink50[2] , \wAMid0[7] , 
        \wAIn1[9] , \wAMid11[30] , \wRegInA10[6] , \wAMid11[29] , \wAIn29[13] , 
        \wRegInB13[13] , \wRegInA3[0] , \wRegInA13[5] , \wRegInB30[22] , 
        \ScanLink0[19] , \wBIn1[14] , \wBMid2[26] , \wBMid2[15] , \wBMid12[4] , 
        \wBIn22[5] , \wRegInB2[18] , \ScanLink53[1] , \wAIn4[4] , \wAIn7[30] , 
        \wAIn7[29] , \wBIn15[22] , \wBIn23[27] , \wRegInB12[9] , 
        \ScanLink32[8] , \wBMid17[9] , \wBIn21[6] , \wRegInA10[18] , 
        \wAIn23[2] , \wRegInB9[14] , \wAIn14[30] , \wAIn14[29] , \wBIn15[11] , 
        \wBIn23[14] , \wBMid26[19] , \wRegInA16[8] , \ScanLink19[28] , 
        \wAMid3[4] , \wAIn7[7] , \wRegInB9[27] , \ScanLink19[31] , 
        \ScanLink48[0] , \wAIn20[1] , \wAIn10[18] , \wBIn11[20] , \wAIn19[8] , 
        \wBIn27[25] , \wAMid28[22] , \wBMid1[0] , \wAIn3[18] , \wBMid2[3] , 
        \wBMid6[17] , \wBMid22[28] , \wBMid22[31] , \wRegInB28[3] , 
        \wBMid6[24] , \wAMid20[7] , \wRegInA14[29] , \wRegInA14[30] , 
        \wBIn5[25] , \wBIn11[13] , \wBIn27[16] , \wAMid28[11] , \wAMid23[4] , 
        \wRegInA29[20] , \ScanLink4[31] , \ScanLink4[28] , \wAMid6[9] , 
        \wAIn8[14] , \wBMid29[17] , \wRegInB6[30] , \wRegInB6[29] , 
        \ScanLink63[16] , \ScanLink55[13] , \ScanLink40[27] , \ScanLink16[26] , 
        \ScanLink35[17] , \ScanLink20[23] , \wAMid15[18] , \wRegInB17[22] , 
        \wRegInB21[27] , \ScanLink13[3] , \wBIn0[3] , \wAIn2[21] , \wAIn2[12] , 
        \wBIn5[16] , \wAIn8[27] , \wAMid26[9] , \wRegInB17[11] , 
        \wRegInA29[13] , \wRegInB21[14] , \wRegInB30[1] , \ScanLink55[20] , 
        \ScanLink20[10] , \ScanLink10[0] , \wBIn10[19] , \wAIn11[21] , 
        \wBMid29[24] , \ScanLink63[25] , \ScanLink16[15] , \ScanLink40[14] , 
        \ScanLink35[24] , \wBMid23[11] , \wAIn27[24] , \wRegInB26[5] , 
        \wAMid6[16] , \wBIn16[9] , \wBMid15[14] , \wRegInA15[23] , 
        \wRegInA23[26] , \wRegInB25[6] , \ScanLink18[8] , \wBIn3[0] , 
        \wAMid6[25] , \wBIn10[7] , \wAIn11[12] , \wBMid15[27] , \wBMid23[22] , 
        \wRegInB2[1] , \wRegInA22[4] , \wBMid23[5] , \wAIn27[17] , 
        \wAMid29[28] , \ScanLink62[0] , \wAMid29[31] , \wAMid14[21] , 
        \wBMid20[6] , \wRegInA15[10] , \ScanLink61[3] , \wRegInB1[2] , 
        \wRegInA23[15] , \wRegInA21[7] , \wAMid22[24] , \wBMid9[8] , 
        \wRegInB23[8] , \ScanLink5[11] , \wAIn2[31] , \wAIn2[28] , 
        \wAMid2[27] , \wAMid2[14] , \wAIn6[10] , \wAIn9[1] , \wBMid8[20] , 
        \wBMid8[13] , \wAMid10[23] , \wAIn11[0] , \wBIn13[4] , \wAMid14[12] , 
        \wAMid22[17] , \wRegInA1[15] , \wRegInB7[10] , \wRegInA28[19] , 
        \wRegInB16[31] , \wRegInB16[28] , \ScanLink54[19] , \ScanLink21[30] , 
        \wAIn12[3] , \wRegInA1[26] , \ScanLink21[29] , \wRegInB7[23] , 
        \wAMid26[26] , \wBMid26[8] , \wBIn29[21] , \wRegInB3[12] , 
        \wRegInA5[17] , \wRegInA27[9] , \ScanLink5[22] , \ScanLink2[7] , 
        \ScanLink1[13] , \wAIn28[9] , \wAIn28[19] , \wRegInB31[28] , 
        \wRegInB31[31] , \wRegInB12[19] , \wAMid9[18] , \wAMid11[6] , 
        \wAMid12[5] , \wRegInB3[21] , \ScanLink50[31] , \ScanLink50[28] , 
        \ScanLink40[8] , \ScanLink25[18] , \ScanLink1[4] , \ScanLink1[20] , 
        \wRegInA5[24] , \wAMid10[10] , \wRegInB19[2] , \wAMid26[15] , 
        \wBIn29[12] , \ScanLink39[3] , \wRegInA11[21] , \wRegInA27[24] , 
        \ScanLink45[5] , \ScanLink4[9] , \wBMid11[16] , \wAIn6[23] , 
        \wBIn14[31] , \wBIn14[28] , \wAIn15[23] , \wAIn23[26] , \wBMid27[13] , 
        \wRegInB19[26] , \ScanLink18[22] , \ScanLink46[6] , \wAIn15[10] , 
        \wRegInA11[12] , \wRegInA27[17] , \ScanLink21[1] , \wAMid17[8] , 
        \wAIn23[15] , \wBMid27[20] , \wRegInB19[15] , \ScanLink22[2] , 
        \ScanLink18[11] , \wBIn3[9] , \wBIn4[26] , \wAMid8[6] , \wAIn9[17] , 
        \wBMid11[25] , \wBMid25[2] , \wRegInB4[6] , \wRegInB16[21] , 
        \wRegInB20[24] , \wRegInA24[3] , \wAIn11[9] , \ScanLink54[10] , 
        \ScanLink21[20] , \wBMid26[1] , \wBMid28[14] , \ScanLink64[7] , 
        \ScanLink62[15] , \ScanLink41[24] , \ScanLink34[14] , \ScanLink17[25] , 
        \wAIn9[24] , \wBMid28[27] , \wRegInB7[5] , \wRegInA27[0] , 
        \wRegInA28[23] , \ScanLink62[26] , \ScanLink41[17] , \ScanLink34[27] , 
        \ScanLink17[16] , \ScanLink54[23] , \ScanLink21[13] , \wBIn4[15] , 
        \wBMid9[1] , \wAMid14[31] , \wAMid14[28] , \wAMid28[6] , 
        \wRegInB20[17] , \wRegInB20[2] , \wRegInB16[12] , \wRegInB23[1] , 
        \wRegInA28[10] , \ScanLink5[18] , \wBMid7[14] , \wRegInB7[19] , 
        \wRegInB2[8] , \wBMid3[16] , \wBIn5[7] , \wBIn10[23] , \wAIn17[7] , 
        \wBIn26[26] , \wAMid29[21] , \wBIn10[10] , \wAIn14[4] , 
        \ScanLink62[9] , \wRegInA15[19] , \wAIn11[31] , \wAIn11[28] , 
        \wBIn26[15] , \wAMid29[12] , \wBIn16[0] , \wBIn6[4] , \wBMid7[27] , 
        \wBMid23[18] , \wBIn14[21] , \wAMid14[2] , \wBIn15[3] , \wAMid30[4] , 
        \ScanLink18[1] , \wBIn31[5] , \wRegInB8[17] , \ScanLink21[8] , 
        \wAIn15[19] , \wBIn22[24] , \wAMid17[1] , \wBMid27[30] , \wBMid27[29] , 
        \ScanLink18[18] , \ScanLink4[0] , \wBIn0[24] , \wBMid3[25] , 
        \wBMid19[6] , \wAIn30[2] , \wRegInA11[31] , \wRegInA8[2] , 
        \wRegInA11[28] , \wRegInA18[7] , \wRegInB8[24] , \ScanLink58[3] , 
        \wAIn6[19] , \wAIn9[8] , \wBIn14[12] , \wBIn22[17] , \ScanLink7[3] , 
        \ScanLink1[30] , \ScanLink1[29] , \wBIn0[17] , \wBMid8[30] , 
        \wBMid8[29] , \wRegInB3[31] , \wRegInB3[28] , \ScanLink27[6] , 
        \ScanLink45[26] , \ScanLink24[5] , \ScanLink30[16] , \wAMid9[11] , 
        \wBIn29[7] , \ScanLink50[12] , \ScanLink13[27] , \wAMid10[19] , 
        \wRegInB31[12] , \wRegInB24[26] , \ScanLink25[22] , \wAIn28[23] , 
        \wRegInB12[23] , \ScanLink43[2] , \wAIn2[3] , \wAMid3[24] , 
        \wAMid3[17] , \wAMid9[22] , \wAIn28[10] , \wRegInB31[21] , \wAIn28[0] , 
        \wBIn29[28] , \wRegInB12[10] , \wBIn29[31] , \wRegInB24[15] , 
        \ScanLink25[11] , \wBMid10[15] , \wAIn14[20] , \ScanLink50[21] , 
        \ScanLink40[1] , \ScanLink45[15] , \ScanLink30[25] , \ScanLink13[14] , 
        \wBIn15[18] , \wBMid17[0] , \wAIn22[25] , \wRegInB18[25] , 
        \ScanLink56[5] , \wBMid26[10] , \ScanLink19[21] , \wRegInA16[1] , 
        \wAIn7[13] , \wBMid14[3] , \wRegInA5[7] , \wRegInA6[4] , 
        \ScanLink48[9] , \ScanLink9[5] , \wRegInA10[22] , \wRegInA15[2] , 
        \wRegInA26[27] , \ScanLink55[6] , \wAIn20[8] , \wAIn7[20] , 
        \wBMid10[26] , \wAMid8[31] , \wAMid8[28] , \wAIn14[13] , \wAIn22[16] , 
        \wBMid26[23] , \wRegInB12[0] , \ScanLink19[12] , \wRegInB18[16] , 
        \ScanLink32[1] , \wAMid19[7] , \wRegInA10[11] , \wRegInB11[3] , 
        \wRegInA26[14] , \ScanLink31[2] , \wBMid9[10] , \wAMid11[20] , 
        \wAIn25[5] , \wAIn1[0] , \wAIn26[6] , \wAMid27[25] , \wBIn28[22] , 
        \wRegInB2[11] , \wRegInA3[9] , \ScanLink0[10] , \ScanLink53[8] , 
        \wRegInA4[14] , \wBIn0[30] , \wRegInA0[25] , \wRegInA0[16] , 
        \wBMid9[23] , \wAMid11[13] , \wBIn24[2] , \wAMid27[16] , \wBIn28[11] , 
        \ScanLink29[0] , \wAIn29[30] , \wAIn29[29] , \wRegInB13[29] , 
        \wRegInB13[30] , \wRegInB30[18] , \wAMid26[0] , \wBIn27[1] , 
        \wRegInB2[22] , \wRegInA4[27] , \ScanLink51[18] , \ScanLink24[31] , 
        \ScanLink24[28] , \ScanLink0[23] , \wBMid4[4] , \wAMid5[3] , 
        \wBMid7[7] , \wAMid15[22] , \wAMid23[27] , \wRegInB6[13] , 
        \ScanLink4[12] , \wRegInB17[18] , \wAMid25[3] , \wRegInB30[8] , 
        \ScanLink55[30] , \ScanLink55[29] , \ScanLink20[19] , \ScanLink10[9] , 
        \wRegInA29[30] , \wRegInA29[29] , \ScanLink4[21] , \wRegInB6[20] , 
        \wBMid1[9] , \wAIn3[11] , \wAMid6[0] , \wAMid15[11] , \wBMid28[7] , 
        \wRegInB9[3] , \wRegInA29[6] , \wAMid7[15] , \wBMid14[17] , 
        \wBIn18[6] , \wAMid23[14] , \wRegInA14[20] , \wRegInA22[25] , 
        \ScanLink15[4] , \wBIn8[2] , \wBMid22[12] , \wAIn26[27] , \wAMid2[23] , 
        \wAMid2[10] , \wAIn3[22] , \wAMid7[26] , \wAIn10[22] , \wAIn10[11] , 
        \wAIn19[1] , \wAMid28[18] , \ScanLink16[7] , \wRegInA31[4] , 
        \wBMid30[5] , \wRegInA22[16] , \wRegInA14[13] , \wBIn11[30] , 
        \wAIn26[14] , \wBIn11[29] , \wBMid22[21] , \wBMid14[24] , \wBMid3[31] , 
        \wAIn15[27] , \wAIn23[22] , \wRegInB19[22] , \ScanLink46[2] , 
        \wBMid27[17] , \ScanLink18[26] , \wBMid3[28] , \wBMid11[12] , 
        \wAIn6[14] , \wAIn9[5] , \wRegInB8[30] , \wRegInB8[29] , 
        \wRegInA11[25] , \wRegInA27[20] , \ScanLink45[1] , \wAIn6[27] , 
        \wBMid11[21] , \wBMid8[24] , \wBMid8[17] , \wAIn15[14] , \wBIn22[30] , 
        \wAIn23[11] , \wBMid27[24] , \ScanLink18[15] , \wRegInB19[11] , 
        \ScanLink22[6] , \wBIn22[29] , \wBIn31[8] , \wRegInA11[16] , 
        \wRegInA27[13] , \ScanLink21[5] , \ScanLink30[31] , \ScanLink1[0] , 
        \ScanLink13[19] , \wAMid10[27] , \ScanLink45[18] , \ScanLink30[28] , 
        \wAMid10[14] , \wAMid26[22] , \wRegInB24[18] , \wAMid26[11] , 
        \wBIn29[25] , \wRegInB3[16] , \ScanLink2[3] , \ScanLink1[17] , 
        \wRegInA5[13] , \ScanLink39[7] , \wBIn29[16] , \wRegInB19[6] , 
        \ScanLink24[8] , \wAMid11[2] , \wBIn0[29] , \wRegInA5[20] , \wBIn0[7] , 
        \wBIn4[18] , \wAMid12[1] , \wRegInB3[25] , \ScanLink1[24] , 
        \wRegInA1[11] , \wRegInB7[14] , \wRegInA0[31] , \wRegInA0[28] , 
        \wAIn2[25] , \wAIn2[16] , \wBIn3[4] , \wBIn10[3] , \wBIn13[0] , 
        \ScanLink5[15] , \wBIn6[9] , \wAIn9[30] , \wAMid14[25] , \wAMid22[20] , 
        \wAIn9[29] , \wAIn11[4] , \wAIn12[7] , \wRegInB7[27] , \wRegInB7[8] , 
        \ScanLink5[26] , \wRegInA1[22] , \wAMid14[16] , \wBMid28[19] , 
        \ScanLink62[18] , \ScanLink41[30] , \ScanLink41[29] , \ScanLink17[28] , 
        \ScanLink34[19] , \ScanLink17[31] , \wAMid22[13] , \wRegInB20[30] , 
        \wRegInB20[29] , \wAMid30[9] , \wRegInA15[27] , \wRegInA23[22] , 
        \wAMid6[12] , \wBMid15[10] , \wRegInB25[2] , \wAMid6[21] , 
        \wBMid7[19] , \wAIn11[25] , \wBMid23[15] , \wAIn27[20] , 
        \wRegInB26[1] , \wAIn11[16] , \wAIn14[9] , \wBIn26[18] , \wRegInB1[6] , 
        \wRegInA21[3] , \wRegInA23[11] , \wBMid20[2] , \wRegInA15[14] , 
        \ScanLink61[7] , \wBMid23[26] , \wBMid23[1] , \wAIn27[13] , 
        \wRegInB2[5] , \ScanLink62[4] , \wRegInA22[0] , \wBMid15[23] , 
        \wAIn8[10] , \wAMid23[19] , \wRegInB17[26] , \wRegInB21[23] , 
        \wBMid29[13] , \ScanLink55[17] , \ScanLink40[23] , \ScanLink20[27] , 
        \ScanLink35[13] , \ScanLink63[12] , \ScanLink16[22] , \wBIn5[21] , 
        \wBIn5[12] , \wAIn8[23] , \wBMid29[20] , \wRegInA29[24] , 
        \ScanLink40[10] , \ScanLink35[20] , \ScanLink16[11] , \ScanLink63[21] , 
        \wRegInB17[15] , \wRegInB21[10] , \ScanLink55[24] , \ScanLink20[14] , 
        \ScanLink10[4] , \wRegInB30[5] , \wRegInA29[17] , \ScanLink13[7] , 
        \wAMid0[3] , \wBMid4[9] , \wBMid6[13] , \wBIn1[23] , \wBMid1[4] , 
        \wAMid3[0] , \wBIn11[24] , \wBMid14[30] , \wBMid14[29] , \wBIn27[21] , 
        \wAMid28[26] , \wAIn26[19] , \wBMid30[8] , \wRegInA31[9] , 
        \wBIn11[17] , \wAMid23[0] , \wBIn27[12] , \wAMid28[15] , \wBMid2[22] , 
        \wBMid2[11] , \wBMid2[7] , \wBMid6[20] , \wAMid7[18] , \wAMid20[3] , 
        \wRegInA22[31] , \wRegInB28[7] , \wAMid3[30] , \wBIn15[26] , 
        \wBIn21[2] , \wRegInB9[10] , \wRegInA22[28] , \ScanLink15[9] , 
        \wRegInA26[19] , \wBIn23[23] , \wAMid3[29] , \wBIn22[1] , \wAIn7[3] , 
        \wAIn20[5] , \wRegInB9[23] , \ScanLink48[4] , \ScanLink9[8] , 
        \wAIn4[0] , \wBMid10[18] , \wRegInA6[9] , \wBIn23[10] , 
        \ScanLink56[8] , \wRegInB18[31] , \wBIn15[15] , \wAIn22[31] , 
        \wAIn22[28] , \wRegInB18[28] , \wAIn23[6] , \wRegInB17[0] , 
        \wBIn1[10] , \wAMid8[16] , \ScanLink51[15] , \ScanLink44[21] , 
        \ScanLink37[1] , \ScanLink34[2] , \ScanLink31[11] , \ScanLink12[20] , 
        \wAIn29[24] , \wRegInB13[24] , \wRegInB14[3] , \wRegInB25[21] , 
        \ScanLink24[25] , \wRegInB30[15] , \ScanLink53[5] , \wBMid12[0] , 
        \wAMid27[28] , \wAIn29[17] , \wRegInA3[4] , \wRegInA4[19] , 
        \wRegInA13[1] , \wRegInB30[26] , \wRegInB13[17] , \wRegInA10[2] , 
        \wAMid27[31] , \wRegInA0[21] , \wRegInA0[12] , \wRegInA0[7] , 
        \wRegInB25[12] , \wAIn3[26] , \wAIn3[15] , \wBMid6[30] , \wBMid6[29] , 
        \wBIn8[6] , \wAMid8[25] , \ScanLink24[16] , \wAIn10[26] , \wBMid11[3] , 
        \wAIn25[8] , \ScanLink51[26] , \ScanLink50[6] , \ScanLink44[12] , 
        \ScanLink31[22] , \ScanLink16[3] , \ScanLink12[13] , \wAMid23[9] , 
        \wAIn26[23] , \wBMid22[16] , \wAMid7[11] , \wBMid14[13] , \wBIn18[2] , 
        \wRegInA22[21] , \ScanLink15[0] , \wRegInA14[24] , \wAMid3[9] , 
        \wAMid7[22] , \wAIn10[15] , \wBMid14[20] , \wBMid22[25] , \wAIn26[10] , 
        \wBIn27[28] , \wBIn27[31] , \wBMid30[1] , \wRegInA14[17] , 
        \wRegInA22[12] , \wBMid4[0] , \wBMid7[3] , \wAIn19[5] , \wRegInA31[0] , 
        \wAMid15[26] , \wAMid25[7] , \wBMid29[30] , \ScanLink63[31] , 
        \ScanLink35[29] , \ScanLink40[19] , \ScanLink35[30] , \ScanLink16[18] , 
        \wBMid29[29] , \ScanLink63[28] , \wAMid23[23] , \wRegInB6[17] , 
        \wRegInB21[19] , \ScanLink4[16] , \wAMid26[4] , \wAMid6[4] , 
        \wAMid23[10] , \wAIn8[19] , \wAMid15[15] , \wBMid28[3] , \wRegInB9[7] , 
        \wRegInA29[2] , \wAIn1[4] , \wBIn5[31] , \wBIn5[28] , \wAMid5[7] , 
        \wRegInB6[24] , \ScanLink4[25] , \wBIn1[19] , \wBMid12[9] , 
        \wAIn26[2] , \wRegInA4[10] , \wAMid27[21] , \wRegInB2[15] , 
        \wRegInA13[8] , \ScanLink0[14] , \wBIn28[26] , \wAIn2[7] , 
        \wBMid9[14] , \wAMid11[24] , \wAIn25[1] , \wBMid9[27] , \wBIn27[5] , 
        \wRegInB2[26] , \wRegInB17[9] , \ScanLink0[27] , \wRegInA4[23] , 
        \ScanLink44[28] , \ScanLink37[8] , \ScanLink12[30] , \wAMid11[17] , 
        \ScanLink44[31] , \ScanLink31[18] , \ScanLink12[29] , \wBIn24[6] , 
        \wAMid27[12] , \wRegInB25[31] , \ScanLink29[4] , \wBIn28[15] , 
        \wRegInB25[28] , \wBIn0[20] , \wBMid2[18] , \wAMid3[13] , \wAIn7[17] , 
        \wBMid14[7] , \wRegInA5[3] , \wRegInA10[26] , \wRegInA15[6] , 
        \wRegInA26[23] , \ScanLink55[2] , \ScanLink9[1] , \wBMid10[11] , 
        \wRegInA6[0] , \wRegInA16[5] , \wAIn4[9] , \wBMid17[4] , \wBMid26[14] , 
        \ScanLink19[25] , \wAIn14[24] , \wAIn22[21] , \wRegInB18[21] , 
        \wBIn23[19] , \ScanLink56[1] , \wAIn14[17] , \wAMid19[3] , 
        \wRegInB9[19] , \wRegInA10[15] , \wRegInB11[7] , \wRegInA26[10] , 
        \ScanLink31[6] , \wAIn22[12] , \wRegInB18[12] , \ScanLink32[5] , 
        \wAMid3[20] , \wAIn7[24] , \wBIn22[8] , \wBMid26[27] , 
        \ScanLink19[16] , \wRegInB12[4] , \wAMid9[15] , \wBMid10[22] , 
        \wAMid26[18] , \wAIn28[27] , \wRegInB12[27] , \wRegInB31[16] , 
        \wRegInB24[22] , \wBIn29[3] , \ScanLink50[16] , \wAMid12[8] , 
        \ScanLink45[22] , \ScanLink25[26] , \ScanLink24[1] , \ScanLink13[23] , 
        \ScanLink30[12] , \wRegInA5[30] , \ScanLink27[2] , \wRegInA5[29] , 
        \wBIn0[13] , \wAMid9[26] , \ScanLink45[11] , \ScanLink30[21] , 
        \ScanLink13[10] , \ScanLink25[15] , \wAIn28[14] , \wAIn28[4] , 
        \wRegInB24[11] , \ScanLink50[25] , \ScanLink40[5] , \ScanLink1[9] , 
        \wRegInB31[25] , \wRegInB12[14] , \wAMid2[19] , \wBMid3[12] , 
        \ScanLink43[6] , \wBMid11[31] , \wBMid11[28] , \wBIn14[25] , 
        \wAMid17[5] , \wBIn22[20] , \wAIn23[18] , \wRegInB19[18] , 
        \wBIn14[16] , \wAMid14[6] , \wBIn31[1] , \wRegInB8[13] , \wBIn22[13] , 
        \ScanLink7[7] , \wBMid3[21] , \wBMid19[2] , \wAIn30[6] , \wRegInA8[6] , 
        \wRegInB8[20] , \ScanLink58[7] , \wRegInA18[3] , \wRegInA27[30] , 
        \wRegInA27[29] , \ScanLink45[8] , \ScanLink4[4] , \wBIn0[22] , 
        \wBIn4[22] , \wBIn5[3] , \wBIn6[0] , \wAMid6[31] , \wAMid6[28] , 
        \wBIn10[27] , \wAIn14[0] , \wRegInA23[18] , \wAIn17[3] , \wBMid23[8] , 
        \wBIn26[22] , \wAMid29[25] , \wBMid7[10] , \wAMid30[0] , 
        \wRegInA22[9] , \ScanLink18[5] , \wBMid7[23] , \wBIn15[7] , 
        \wRegInB26[8] , \wBIn16[4] , \wBMid15[19] , \wAMid8[2] , \wBIn10[14] , 
        \wBIn26[11] , \wAIn27[30] , \wAIn27[29] , \wAMid29[16] , \wRegInB7[1] , 
        \wRegInA28[27] , \wRegInA27[4] , \wBIn4[11] , \wAIn9[13] , 
        \wBMid25[6] , \wBMid26[5] , \wBMid28[10] , \ScanLink64[3] , 
        \ScanLink62[11] , \ScanLink17[21] , \ScanLink54[14] , \ScanLink41[20] , 
        \ScanLink34[10] , \ScanLink21[24] , \wRegInB4[2] , \wRegInB16[25] , 
        \wRegInB20[20] , \wRegInA24[7] , \wAIn9[20] , \wBMid9[5] , 
        \wRegInA1[18] , \wRegInB23[5] , \wBIn13[9] , \wAMid22[30] , 
        \wRegInB16[16] , \wRegInA28[14] , \wRegInB20[6] , \wAMid22[29] , 
        \wAMid28[2] , \wRegInB20[13] , \ScanLink54[27] , \ScanLink21[17] , 
        \wBMid28[23] , \ScanLink17[12] , \ScanLink62[22] , \ScanLink41[13] , 
        \ScanLink34[23] , \ScanLink27[0] , \wBIn0[11] , \wAMid9[17] , 
        \ScanLink45[20] , \ScanLink30[10] , \ScanLink13[21] , \ScanLink24[3] , 
        \ScanLink25[24] , \wAMid11[9] , \wBIn29[1] , \ScanLink50[14] , 
        \wAIn28[25] , \wRegInB24[20] , \wRegInB31[14] , \wRegInB12[25] , 
        \wRegInA5[18] , \ScanLink43[4] , \ScanLink2[8] , \wAMid2[31] , 
        \wAMid2[28] , \wAMid9[24] , \wAMid26[30] , \wAIn28[16] , 
        \wRegInB12[16] , \wRegInB31[27] , \wRegInB24[13] , \wAMid26[29] , 
        \wAIn28[6] , \ScanLink50[27] , \wBIn14[27] , \wAMid14[4] , \wBIn31[3] , 
        \wRegInB8[11] , \ScanLink45[13] , \ScanLink40[7] , \ScanLink25[17] , 
        \ScanLink13[12] , \ScanLink30[23] , \wRegInA27[18] , \wAMid17[7] , 
        \wBIn22[22] , \wBMid3[10] , \ScanLink4[6] , \wRegInA0[23] , 
        \wRegInA0[10] , \wAMid0[8] , \wAIn3[17] , \wBIn4[20] , \wBMid3[23] , 
        \wBMid19[0] , \wAIn30[4] , \wRegInA8[4] , \wRegInA18[1] , 
        \ScanLink58[5] , \wRegInB8[22] , \wBIn5[1] , \wAMid6[19] , 
        \wBMid7[12] , \wBMid11[19] , \wBIn14[14] , \wBIn22[11] , 
        \ScanLink7[5] , \wAIn23[30] , \wAIn23[29] , \ScanLink46[9] , 
        \wRegInB19[29] , \wRegInB19[30] , \wBIn10[25] , \wBMid15[31] , 
        \wBMid15[28] , \wAIn17[1] , \wBIn26[20] , \wAMid29[27] , \wAIn27[18] , 
        \wBIn10[16] , \wAIn14[2] , \wBMid20[9] , \wRegInA21[8] , \wBIn26[13] , 
        \wAMid29[14] , \wBIn16[6] , \wBIn6[2] , \wBMid7[21] , \wAIn9[11] , 
        \wBIn15[5] , \wAMid22[18] , \wAMid30[2] , \wRegInB25[9] , 
        \ScanLink18[7] , \wRegInB4[0] , \wRegInB16[27] , \wRegInA23[30] , 
        \wRegInA23[29] , \wRegInA24[5] , \wRegInB20[22] , \ScanLink54[16] , 
        \ScanLink21[26] , \wBMid25[4] , \wBMid26[7] , \wBMid28[12] , 
        \ScanLink62[13] , \ScanLink17[23] , \ScanLink64[1] , \ScanLink34[12] , 
        \ScanLink41[22] , \wRegInA1[30] , \wBIn4[13] , \wAMid8[0] , 
        \wRegInA1[29] , \wAIn9[22] , \wBMid28[21] , \wRegInB7[3] , 
        \wRegInA27[6] , \wRegInA28[25] , \ScanLink62[20] , \ScanLink54[25] , 
        \ScanLink41[11] , \ScanLink17[10] , \ScanLink34[21] , \ScanLink21[15] , 
        \wBIn10[8] , \wAMid28[0] , \wRegInB20[11] , \wBMid9[7] , 
        \wRegInB16[14] , \wRegInB20[4] , \wRegInB23[7] , \wRegInA28[16] , 
        \wBIn18[0] , \wAMid20[8] , \wRegInA14[26] , \wRegInA22[23] , 
        \ScanLink15[2] , \wBMid6[18] , \wAMid7[13] , \wBIn8[4] , \wBMid14[11] , 
        \wBMid22[14] , \wAIn26[21] , \wAIn10[24] , \wBIn27[19] , 
        \ScanLink16[1] , \wAIn10[17] , \wAIn19[7] , \wRegInA31[2] , 
        \wBMid30[3] , \wRegInA14[15] , \wRegInA22[10] , \wAIn26[12] , 
        \wBMid22[27] , \wAIn3[24] , \wAMid7[20] , \wBMid14[22] , \wBIn5[19] , 
        \wAMid26[6] , \wBMid4[2] , \wRegInB6[15] , \wAMid5[5] , \wAIn8[31] , 
        \wAIn8[28] , \wBMid7[1] , \wAMid15[24] , \wAMid23[21] , 
        \ScanLink4[14] , \wAMid25[5] , \ScanLink4[27] , \wRegInB6[26] , 
        \wAIn2[5] , \wAMid6[6] , \wAMid15[17] , \wBMid29[18] , \wRegInB9[5] , 
        \wRegInA29[0] , \ScanLink40[28] , \ScanLink35[18] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink63[19] , \ScanLink40[31] , \wAMid23[12] , 
        \wBMid28[1] , \wRegInB21[31] , \wBMid9[16] , \wAIn25[3] , 
        \wRegInB21[28] , \ScanLink44[19] , \ScanLink31[29] , \wBMid11[8] , 
        \ScanLink12[18] , \wAMid11[26] , \ScanLink31[30] , \wAMid27[23] , 
        \wBIn28[24] , \wRegInA10[9] , \wAIn1[6] , \wRegInB2[17] , 
        \wRegInB25[19] , \ScanLink0[16] , \wRegInA4[12] , \wAIn26[0] , 
        \wAMid27[10] , \wBIn28[17] , \wRegInB14[8] , \ScanLink29[6] , 
        \wRegInA0[19] , \wBIn1[31] , \wBIn1[28] , \wBMid9[25] , \wAMid11[15] , 
        \wBIn24[4] , \ScanLink34[9] , \wRegInA4[21] , \wBMid2[30] , 
        \wBMid2[29] , \wAIn14[26] , \wBIn27[7] , \wRegInB2[24] , 
        \ScanLink56[3] , \ScanLink0[25] , \wBMid17[6] , \wAIn22[23] , 
        \wRegInB18[23] , \wAMid3[22] , \wAMid3[11] , \wAIn7[15] , 
        \wBMid26[16] , \ScanLink19[27] , \wRegInA6[2] , \wAIn7[26] , 
        \wAIn7[8] , \wBMid10[13] , \wRegInA16[7] , \wRegInA5[1] , 
        \wRegInB9[28] , \wRegInA15[4] , \ScanLink9[3] , \wRegInB9[31] , 
        \wRegInA26[21] , \ScanLink55[0] , \wBMid14[5] , \wRegInA10[24] , 
        \wRegInB12[6] , \wBMid10[20] , \wBIn5[23] , \wAIn14[15] , \wAIn22[10] , 
        \wBMid26[25] , \wRegInB18[10] , \ScanLink19[14] , \ScanLink32[7] , 
        \wBIn23[28] , \wAMid19[1] , \wBIn23[31] , \wRegInA10[17] , 
        \ScanLink31[4] , \wRegInB11[5] , \wRegInA26[12] , \wBIn21[9] , 
        \wRegInA29[26] , \wAIn8[12] , \wBMid29[11] , \ScanLink63[10] , 
        \ScanLink40[21] , \ScanLink35[11] , \ScanLink16[20] , \wBMid28[8] , 
        \wRegInB21[21] , \wRegInA29[9] , \ScanLink20[25] , \ScanLink55[15] , 
        \wRegInB17[24] , \ScanLink13[5] , \wAMid0[1] , \wAMid3[2] , 
        \wBIn5[10] , \wAIn8[21] , \wBMid7[8] , \wAMid23[31] , \wAMid23[28] , 
        \wRegInB17[17] , \wRegInA29[15] , \wRegInB30[7] , \wRegInB21[12] , 
        \wBMid29[22] , \ScanLink63[23] , \ScanLink55[26] , \ScanLink40[12] , 
        \ScanLink20[16] , \ScanLink10[6] , \ScanLink35[22] , \ScanLink16[13] , 
        \wAMid7[30] , \wBIn11[26] , \wRegInA22[19] , \wBIn27[23] , 
        \wAMid28[24] , \wBMid1[6] , \wBMid2[5] , \wBMid6[11] , \wAMid7[29] , 
        \wRegInB28[5] , \wBMid6[22] , \wBIn18[9] , \wAMid20[1] , \wBMid14[18] , 
        \wBIn27[10] , \wAMid28[17] , \ScanLink16[8] , \wBMid2[20] , 
        \wBMid2[13] , \wBIn11[15] , \wAMid23[2] , \wAIn26[31] , \wAIn26[28] , 
        \wAMid3[18] , \wAIn4[2] , \wBMid10[30] , \wBIn22[3] , \wBMid10[29] , 
        \wBIn15[24] , \wBIn23[21] , \wBIn15[17] , \wAMid19[8] , \wAIn22[19] , 
        \wRegInB18[19] , \wBIn21[0] , \wRegInB9[12] , \wAIn23[4] , 
        \wBIn23[12] , \wAIn7[1] , \wAIn20[7] , \wRegInA5[8] , \wRegInB9[21] , 
        \ScanLink48[6] , \wAMid27[19] , \wAIn29[26] , \wRegInA26[31] , 
        \wRegInA26[28] , \ScanLink55[9] , \wRegInB30[17] , \wRegInB13[26] , 
        \wRegInB14[1] , \wRegInB25[23] , \wRegInA0[5] , \wBIn1[21] , 
        \wAMid8[14] , \ScanLink24[27] , \ScanLink51[17] , \ScanLink44[23] , 
        \ScanLink34[0] , \ScanLink31[13] , \ScanLink12[22] , \wAMid8[27] , 
        \wBMid11[1] , \wRegInA4[31] , \wRegInA4[28] , \ScanLink37[3] , 
        \wRegInB17[2] , \ScanLink44[10] , \ScanLink31[20] , \ScanLink51[24] , 
        \ScanLink12[11] , \wRegInA10[0] , \ScanLink50[4] , \ScanLink24[14] , 
        \wRegInB25[10] , \wBIn1[12] , \wBMid12[2] , \wAIn29[15] , 
        \wRegInB13[15] , \wRegInB30[24] , \wRegInA3[6] , \wRegInA13[3] , 
        \wAIn26[9] , \wRegInA11[27] , \ScanLink53[7] , \wRegInA18[8] , 
        \wRegInA27[22] , \ScanLink45[3] , \wBIn0[18] , \wAMid2[21] , 
        \wAMid2[12] , \wBMid19[9] , \wBMid3[19] , \wAIn6[16] , \wBMid11[10] , 
        \wAIn9[7] , \wAIn15[25] , \wAIn23[20] , \wBMid27[15] , 
        \ScanLink18[24] , \wRegInB19[20] , \wAIn15[16] , \wBIn22[18] , 
        \wRegInB8[18] , \ScanLink46[0] , \wRegInA11[14] , \wRegInA27[11] , 
        \ScanLink21[7] , \wAIn23[13] , \wRegInB19[13] , \ScanLink22[4] , 
        \wBMid27[26] , \ScanLink18[17] , \wBMid11[23] , \wAIn6[25] , 
        \wRegInA5[11] , \wBIn0[5] , \wBIn3[6] , \wBMid8[26] , \wBMid8[15] , 
        \wAMid10[25] , \wAMid26[20] , \wBIn29[27] , \wRegInB3[14] , 
        \ScanLink2[1] , \ScanLink1[15] , \wAMid11[0] , \wAMid12[3] , 
        \ScanLink1[26] , \ScanLink1[2] , \wBIn29[8] , \wRegInB3[27] , 
        \wRegInA5[22] , \ScanLink27[9] , \wRegInB19[4] , \ScanLink45[30] , 
        \ScanLink13[28] , \ScanLink30[19] , \wBIn10[1] , \wAMid10[16] , 
        \ScanLink45[29] , \ScanLink13[31] , \wAMid14[27] , \wAMid26[13] , 
        \wBIn29[14] , \wRegInB24[29] , \wBMid28[31] , \wBMid28[28] , 
        \wRegInB24[30] , \ScanLink39[5] , \ScanLink62[29] , \ScanLink41[18] , 
        \ScanLink34[31] , \ScanLink17[19] , \ScanLink62[30] , \ScanLink34[28] , 
        \wAMid28[9] , \wRegInB20[18] , \wAMid22[22] , \ScanLink5[17] , 
        \wAIn1[2] , \wAIn2[27] , \wAIn2[14] , \wBIn4[30] , \wAIn9[18] , 
        \wAIn11[6] , \wBIn13[2] , \wAMid14[14] , \wAMid22[11] , \wRegInA1[13] , 
        \wRegInB7[16] , \wRegInB4[9] , \ScanLink64[8] , \wBIn4[29] , 
        \wBIn5[8] , \wAMid6[10] , \wBMid7[31] , \wAMid8[9] , \wAIn11[27] , 
        \wAIn12[5] , \wRegInA1[20] , \wRegInB7[25] , \ScanLink5[24] , 
        \wAIn27[22] , \wBMid7[28] , \wBMid23[17] , \wRegInB26[3] , 
        \wBMid15[12] , \wAMid6[23] , \wBMid15[21] , \wRegInA15[25] , 
        \wRegInA23[20] , \wRegInB25[0] , \wAMid3[26] , \wAMid3[15] , 
        \wAIn11[14] , \wBMid23[24] , \wRegInB2[7] , \wBMid23[3] , \wBIn26[30] , 
        \wAIn27[11] , \wRegInA22[2] , \ScanLink62[6] , \wBMid14[1] , 
        \wAIn17[8] , \wBMid20[0] , \wBIn26[29] , \wRegInA15[16] , 
        \wRegInA23[13] , \ScanLink61[5] , \wRegInB1[4] , \wRegInA21[1] , 
        \wRegInA5[5] , \wRegInA10[20] , \wRegInA26[25] , \ScanLink55[4] , 
        \wRegInA15[0] , \ScanLink9[7] , \wAIn7[11] , \wBMid10[17] , 
        \wRegInA16[3] , \wRegInA6[6] , \wBMid10[24] , \wAIn14[22] , 
        \wBMid17[2] , \wAIn22[27] , \wBMid26[12] , \ScanLink19[23] , 
        \wAIn23[9] , \wRegInB18[27] , \wAIn14[11] , \wAMid19[5] , 
        \ScanLink56[7] , \wRegInA10[13] , \wRegInB11[1] , \wRegInA26[16] , 
        \ScanLink31[0] , \wBIn15[30] , \wAIn22[14] , \wRegInB18[14] , 
        \ScanLink32[3] , \wBIn15[29] , \wBMid26[21] , \ScanLink19[10] , 
        \wAIn7[22] , \wRegInB12[2] , \wAIn26[4] , \wRegInA4[16] , 
        \wRegInB2[13] , \ScanLink0[12] , \wRegInA0[8] , \wAIn2[1] , 
        \wAMid11[22] , \wAMid27[27] , \wBIn28[20] , \wAIn29[18] , 
        \wRegInB13[18] , \wRegInB30[30] , \wRegInB30[29] , \wAMid8[19] , 
        \wBMid9[12] , \wAIn25[7] , \wBIn27[3] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink50[9] , \ScanLink24[19] , \ScanLink0[21] , 
        \wRegInB2[20] , \wRegInA4[25] , \wBMid9[21] , \wAMid11[11] , 
        \wBIn24[0] , \wBIn0[8] , \wRegInA0[27] , \wRegInA0[14] , \wBMid4[6] , 
        \wBMid7[5] , \wAMid27[14] , \wBIn28[13] , \ScanLink29[2] , 
        \wAMid15[20] , \wAMid25[1] , \wAMid23[25] , \wRegInA29[18] , 
        \ScanLink4[10] , \wRegInB6[11] , \ScanLink13[8] , \wAMid6[2] , 
        \wAMid26[2] , \wAMid15[13] , \wAMid23[16] , \wRegInB17[29] , 
        \wBMid28[5] , \wRegInB17[30] , \wRegInB9[1] , \wRegInA29[4] , 
        \ScanLink20[28] , \ScanLink55[18] , \ScanLink20[31] , \wAIn3[20] , 
        \wAIn3[13] , \wAMid5[1] , \wRegInB6[22] , \wAMid7[17] , \wBIn8[0] , 
        \wAIn10[20] , \ScanLink4[23] , \wAIn26[25] , \ScanLink16[5] , 
        \wBIn11[18] , \wBMid22[10] , \wBMid14[15] , \wBMid2[8] , 
        \wRegInA22[27] , \wRegInB28[8] , \ScanLink15[6] , \wAMid7[24] , 
        \wBMid14[26] , \wBIn18[4] , \wRegInA14[22] , \wBIn4[24] , \wAIn10[13] , 
        \wBMid22[23] , \wAIn26[16] , \wAMid28[30] , \wAIn19[3] , \wAMid28[29] , 
        \wBMid30[7] , \wRegInA14[11] , \wRegInA22[14] , \wRegInA31[6] , 
        \wRegInB7[7] , \wRegInA27[2] , \wRegInA28[21] , \ScanLink5[30] , 
        \ScanLink5[29] , \wBIn4[17] , \wAMid8[4] , \wAIn9[15] , \wAIn12[8] , 
        \wBMid26[3] , \wRegInB7[31] , \wRegInB7[28] , \wBMid28[16] , 
        \ScanLink64[5] , \ScanLink34[16] , \ScanLink41[26] , \ScanLink17[27] , 
        \ScanLink62[17] , \wAMid14[19] , \wBMid25[0] , \wRegInB4[4] , 
        \wRegInB20[26] , \ScanLink54[12] , \ScanLink21[22] , \wRegInB16[23] , 
        \wRegInA24[1] , \wBMid9[3] , \wRegInB23[3] , \wRegInA28[12] , 
        \wAIn2[19] , \wBIn6[6] , \wBMid7[16] , \wAIn9[26] , \wAMid28[4] , 
        \wRegInB16[10] , \wRegInB20[0] , \wRegInB20[15] , \wBIn10[21] , 
        \wAIn14[6] , \wBMid28[25] , \ScanLink54[21] , \ScanLink41[15] , 
        \ScanLink21[11] , \ScanLink34[25] , \wRegInB1[9] , \ScanLink62[24] , 
        \ScanLink17[14] , \ScanLink61[8] , \wAIn11[19] , \wAIn17[5] , 
        \wBIn26[24] , \wAMid29[23] , \wBMid23[30] , \wBMid23[29] , 
        \wAMid30[6] , \wRegInA15[31] , \wRegInA15[28] , \ScanLink18[3] , 
        \wBMid7[25] , \wBIn15[1] , \wBMid3[27] , \wBMid3[14] , \wBIn5[5] , 
        \wBIn16[2] , \wBIn10[12] , \wBIn26[17] , \wAMid29[10] , \wAIn6[31] , 
        \wAIn6[28] , \wBIn14[23] , \wAMid17[3] , \wBIn22[26] , \wBIn14[10] , 
        \wAMid14[0] , \ScanLink22[9] , \wBIn31[7] , \wRegInA11[19] , 
        \wRegInB8[15] , \wAIn15[31] , \wAIn15[28] , \wBIn22[15] , 
        \ScanLink18[30] , \ScanLink7[1] , \wBMid19[4] , \wBMid27[18] , 
        \ScanLink18[29] , \wRegInB8[26] , \wAIn30[0] , \ScanLink58[1] , 
        \wRegInA8[0] , \wRegInA18[5] , \ScanLink4[2] , \wBIn0[26] , 
        \wAMid9[13] , \wAIn28[21] , \wRegInB31[10] , \wBIn29[19] , 
        \wRegInB12[21] , \wRegInB24[24] , \ScanLink39[8] , \ScanLink25[20] , 
        \wBIn29[5] , \ScanLink50[10] , \wRegInB19[9] , \ScanLink45[24] , 
        \ScanLink30[14] , \ScanLink24[7] , \ScanLink13[25] , \wBIn0[15] , 
        \wBMid8[18] , \ScanLink45[17] , \ScanLink27[4] , \ScanLink30[27] , 
        \wAMid9[20] , \ScanLink50[23] , \ScanLink13[16] , \wAMid10[31] , 
        \wAMid10[28] , \wAIn28[2] , \ScanLink40[3] , \ScanLink25[13] , 
        \wRegInB31[23] , \wRegInB24[17] , \wRegInB12[12] , \wAIn28[12] , 
        \ScanLink1[18] , \wBIn0[1] , \wAIn2[23] , \wAIn2[10] , \wBIn15[8] , 
        \wRegInB3[19] , \wRegInA15[21] , \ScanLink43[0] , \wRegInA23[24] , 
        \wRegInB25[4] , \wAMid6[14] , \wBIn10[31] , \wBIn10[28] , \wAIn11[23] , 
        \wBMid15[16] , \wBMid23[13] , \wRegInB26[7] , \wAIn27[26] , 
        \wAMid29[19] , \wAIn11[10] , \wBMid20[4] , \wRegInB1[0] , 
        \wRegInA21[5] , \wRegInA15[12] , \wRegInA23[17] , \ScanLink61[1] , 
        \wBMid23[7] , \ScanLink62[2] , \wBMid23[20] , \wAIn27[15] , 
        \wRegInB2[3] , \wRegInA22[6] , \wAMid6[27] , \wBMid15[25] , 
        \wRegInA1[17] , \wRegInB7[12] , \wRegInA0[1] , \wBIn1[25] , 
        \wAMid2[25] , \wAMid2[16] , \wBIn3[2] , \wBIn10[5] , \wBIn13[6] , 
        \ScanLink5[13] , \wAIn6[12] , \wBMid8[22] , \wBMid8[11] , \wAMid9[30] , 
        \wAIn11[2] , \wAIn12[1] , \wAMid14[23] , \wAMid22[26] , \wRegInB20[9] , 
        \wRegInB16[19] , \wRegInA28[31] , \ScanLink54[31] , \ScanLink54[28] , 
        \ScanLink21[18] , \ScanLink5[20] , \wRegInA28[28] , \wBMid25[9] , 
        \wRegInA1[24] , \wRegInB7[21] , \wAMid14[10] , \wAMid22[15] , 
        \wRegInA24[8] , \ScanLink1[6] , \wAMid9[29] , \wAMid10[21] , 
        \wAMid10[12] , \wAMid26[24] , \wAMid26[17] , \wBIn29[23] , 
        \wRegInB3[10] , \ScanLink1[11] , \wRegInA5[15] , \ScanLink43[9] , 
        \ScanLink2[5] , \wAIn28[31] , \wBIn29[10] , \ScanLink39[1] , 
        \wAIn28[28] , \wRegInB31[19] , \wRegInB12[31] , \wRegInB12[28] , 
        \wAMid11[4] , \wRegInB19[0] , \ScanLink25[30] , \wAMid12[7] , 
        \wRegInB3[23] , \wRegInA5[26] , \ScanLink50[19] , \ScanLink25[29] , 
        \wBIn14[19] , \wAIn15[21] , \ScanLink46[4] , \ScanLink1[22] , 
        \ScanLink7[8] , \wAIn23[24] , \wBMid27[11] , \wRegInB19[24] , 
        \ScanLink18[20] , \wAIn9[3] , \wAIn6[21] , \wBMid11[14] , \wAIn30[9] , 
        \wRegInA27[26] , \ScanLink58[8] , \ScanLink45[7] , \wRegInA8[9] , 
        \wRegInA11[23] , \wBMid11[27] , \wAMid14[9] , \wAIn15[12] , 
        \wAIn23[17] , \wBMid27[22] , \wRegInB19[17] , \ScanLink18[13] , 
        \ScanLink22[0] , \wRegInA11[10] , \ScanLink21[3] , \wRegInB17[6] , 
        \wRegInA27[15] , \ScanLink37[7] , \ScanLink0[31] , \ScanLink0[28] , 
        \wBIn1[16] , \wAMid8[10] , \wBMid9[31] , \wRegInB2[30] , 
        \wRegInB2[29] , \ScanLink12[26] , \wBMid9[28] , \ScanLink31[17] , 
        \ScanLink44[27] , \ScanLink34[4] , \ScanLink24[23] , \wAMid11[18] , 
        \wBIn24[9] , \wAIn29[22] , \wRegInB14[5] , \ScanLink51[13] , 
        \wRegInB25[27] , \wRegInB13[22] , \wBMid12[6] , \wRegInB30[13] , 
        \ScanLink53[3] , \wAIn29[11] , \wRegInA3[2] , \wRegInA13[7] , 
        \wRegInB13[11] , \wRegInB25[14] , \wRegInB30[20] , \wAMid0[5] , 
        \wAIn2[8] , \wAMid8[23] , \wBIn28[30] , \wBIn28[29] , \wRegInA10[4] , 
        \ScanLink51[20] , \wBMid11[5] , \ScanLink50[0] , \ScanLink24[10] , 
        \wAIn3[30] , \wBMid2[24] , \wBMid2[17] , \wAIn14[18] , \wBIn15[20] , 
        \wBIn21[4] , \wRegInB9[16] , \wRegInB11[8] , \ScanLink44[14] , 
        \ScanLink12[15] , \ScanLink31[24] , \ScanLink31[9] , \wBIn23[25] , 
        \wBMid26[31] , \wBMid26[28] , \ScanLink19[19] , \wAIn7[5] , 
        \wBIn22[7] , \wBMid14[8] , \wRegInA10[29] , \wAIn20[3] , 
        \wRegInB9[25] , \wRegInA10[30] , \wRegInA15[9] , \ScanLink48[2] , 
        \wAIn4[6] , \wAIn7[18] , \wBIn15[13] , \wAIn23[0] , \wBIn23[16] , 
        \wBMid6[15] , \wBMid1[2] , \wAIn3[29] , \wAMid3[6] , \wBIn11[22] , 
        \wBIn27[27] , \wAMid28[20] , \wRegInA14[18] , \wBIn8[9] , \wBIn11[11] , 
        \wAMid23[6] , \wBMid2[1] , \wBMid6[26] , \wAIn10[30] , \wAIn10[29] , 
        \wBIn27[14] , \wBMid22[19] , \wAMid28[13] , \wAMid20[5] , 
        \wRegInB28[1] , \wBIn5[27] , \wAIn8[16] , \wRegInB9[8] , 
        \wRegInB17[20] , \wRegInB21[25] , \ScanLink55[11] , \ScanLink20[21] , 
        \wBMid29[15] , \ScanLink16[24] , \ScanLink63[14] , \ScanLink40[25] , 
        \ScanLink35[15] , \wBIn5[14] , \wAMid5[8] , \wRegInA29[22] , 
        \wAIn8[25] , \wAMid25[8] , \wBMid29[26] , \ScanLink63[27] , 
        \ScanLink55[22] , \ScanLink40[16] , \ScanLink16[17] , \ScanLink35[26] , 
        \ScanLink20[12] , \ScanLink10[2] , \wAMid15[30] , \wRegInB17[13] , 
        \wRegInB21[16] , \wAMid15[29] , \wRegInB30[3] , \wRegInA29[11] , 
        \ScanLink4[19] , \wRegInB6[18] , \ScanLink13[1] ;
    BubbleSort_Node_WIDTH32 BSN1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn0[31] , 
        \wAIn0[30] , \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , \wAIn0[26] , 
        \wAIn0[25] , \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , \wAIn0[21] , 
        \wAIn0[20] , \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , \wAIn0[16] , 
        \wAIn0[15] , \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , \wAIn0[11] , 
        \wAIn0[10] , \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , \wAIn0[6] , 
        \wAIn0[5] , \wAIn0[4] , \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , \wAIn0[0] 
        }), .BIn({\wBIn0[31] , \wBIn0[30] , \wBIn0[29] , \wBIn0[28] , 
        \wBIn0[27] , \wBIn0[26] , \wBIn0[25] , \wBIn0[24] , \wBIn0[23] , 
        \wBIn0[22] , \wBIn0[21] , \wBIn0[20] , \wBIn0[19] , \wBIn0[18] , 
        \wBIn0[17] , \wBIn0[16] , \wBIn0[15] , \wBIn0[14] , \wBIn0[13] , 
        \wBIn0[12] , \wBIn0[11] , \wBIn0[10] , \wBIn0[9] , \wBIn0[8] , 
        \wBIn0[7] , \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , \wBIn0[3] , \wBIn0[2] , 
        \wBIn0[1] , \wBIn0[0] }), .HiOut({\wRegInA0[31] , \wRegInA0[30] , 
        \wRegInA0[29] , \wRegInA0[28] , \wRegInA0[27] , \wRegInA0[26] , 
        \wRegInA0[25] , \wRegInA0[24] , \wRegInA0[23] , \wRegInA0[22] , 
        \wRegInA0[21] , \wRegInA0[20] , \wRegInA0[19] , \wRegInA0[18] , 
        \wRegInA0[17] , \wRegInA0[16] , \wRegInA0[15] , \wRegInA0[14] , 
        \wRegInA0[13] , \wRegInA0[12] , \wRegInA0[11] , \wRegInA0[10] , 
        \wRegInA0[9] , \wRegInA0[8] , \wRegInA0[7] , \wRegInA0[6] , 
        \wRegInA0[5] , \wRegInA0[4] , \wRegInA0[3] , \wRegInA0[2] , 
        \wRegInA0[1] , \wRegInA0[0] }), .LoOut({\wAMid0[31] , \wAMid0[30] , 
        \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , \wAMid0[25] , 
        \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , \wAMid0[20] , 
        \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , \wAMid0[15] , 
        \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , \wAMid0[10] , 
        \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , \wAMid0[5] , 
        \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , \wAMid0[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn2[31] , 
        \wAIn2[30] , \wAIn2[29] , \wAIn2[28] , \wAIn2[27] , \wAIn2[26] , 
        \wAIn2[25] , \wAIn2[24] , \wAIn2[23] , \wAIn2[22] , \wAIn2[21] , 
        \wAIn2[20] , \wAIn2[19] , \wAIn2[18] , \wAIn2[17] , \wAIn2[16] , 
        \wAIn2[15] , \wAIn2[14] , \wAIn2[13] , \wAIn2[12] , \wAIn2[11] , 
        \wAIn2[10] , \wAIn2[9] , \wAIn2[8] , \wAIn2[7] , \wAIn2[6] , 
        \wAIn2[5] , \wAIn2[4] , \wAIn2[3] , \wAIn2[2] , \wAIn2[1] , \wAIn2[0] 
        }), .BIn({\wBIn2[31] , \wBIn2[30] , \wBIn2[29] , \wBIn2[28] , 
        \wBIn2[27] , \wBIn2[26] , \wBIn2[25] , \wBIn2[24] , \wBIn2[23] , 
        \wBIn2[22] , \wBIn2[21] , \wBIn2[20] , \wBIn2[19] , \wBIn2[18] , 
        \wBIn2[17] , \wBIn2[16] , \wBIn2[15] , \wBIn2[14] , \wBIn2[13] , 
        \wBIn2[12] , \wBIn2[11] , \wBIn2[10] , \wBIn2[9] , \wBIn2[8] , 
        \wBIn2[7] , \wBIn2[6] , \wBIn2[5] , \wBIn2[4] , \wBIn2[3] , \wBIn2[2] , 
        \wBIn2[1] , \wBIn2[0] }), .HiOut({\wBMid1[31] , \wBMid1[30] , 
        \wBMid1[29] , \wBMid1[28] , \wBMid1[27] , \wBMid1[26] , \wBMid1[25] , 
        \wBMid1[24] , \wBMid1[23] , \wBMid1[22] , \wBMid1[21] , \wBMid1[20] , 
        \wBMid1[19] , \wBMid1[18] , \wBMid1[17] , \wBMid1[16] , \wBMid1[15] , 
        \wBMid1[14] , \wBMid1[13] , \wBMid1[12] , \wBMid1[11] , \wBMid1[10] , 
        \wBMid1[9] , \wBMid1[8] , \wBMid1[7] , \wBMid1[6] , \wBMid1[5] , 
        \wBMid1[4] , \wBMid1[3] , \wBMid1[2] , \wBMid1[1] , \wBMid1[0] }), 
        .LoOut({\wAMid2[31] , \wAMid2[30] , \wAMid2[29] , \wAMid2[28] , 
        \wAMid2[27] , \wAMid2[26] , \wAMid2[25] , \wAMid2[24] , \wAMid2[23] , 
        \wAMid2[22] , \wAMid2[21] , \wAMid2[20] , \wAMid2[19] , \wAMid2[18] , 
        \wAMid2[17] , \wAMid2[16] , \wAMid2[15] , \wAMid2[14] , \wAMid2[13] , 
        \wAMid2[12] , \wAMid2[11] , \wAMid2[10] , \wAMid2[9] , \wAMid2[8] , 
        \wAMid2[7] , \wAMid2[6] , \wAMid2[5] , \wAMid2[4] , \wAMid2[3] , 
        \wAMid2[2] , \wAMid2[1] , \wAMid2[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn3[31] , 
        \wAIn3[30] , \wAIn3[29] , \wAIn3[28] , \wAIn3[27] , \wAIn3[26] , 
        \wAIn3[25] , \wAIn3[24] , \wAIn3[23] , \wAIn3[22] , \wAIn3[21] , 
        \wAIn3[20] , \wAIn3[19] , \wAIn3[18] , \wAIn3[17] , \wAIn3[16] , 
        \wAIn3[15] , \wAIn3[14] , \wAIn3[13] , \wAIn3[12] , \wAIn3[11] , 
        \wAIn3[10] , \wAIn3[9] , \wAIn3[8] , \wAIn3[7] , \wAIn3[6] , 
        \wAIn3[5] , \wAIn3[4] , \wAIn3[3] , \wAIn3[2] , \wAIn3[1] , \wAIn3[0] 
        }), .BIn({\wBIn3[31] , \wBIn3[30] , \wBIn3[29] , \wBIn3[28] , 
        \wBIn3[27] , \wBIn3[26] , \wBIn3[25] , \wBIn3[24] , \wBIn3[23] , 
        \wBIn3[22] , \wBIn3[21] , \wBIn3[20] , \wBIn3[19] , \wBIn3[18] , 
        \wBIn3[17] , \wBIn3[16] , \wBIn3[15] , \wBIn3[14] , \wBIn3[13] , 
        \wBIn3[12] , \wBIn3[11] , \wBIn3[10] , \wBIn3[9] , \wBIn3[8] , 
        \wBIn3[7] , \wBIn3[6] , \wBIn3[5] , \wBIn3[4] , \wBIn3[3] , \wBIn3[2] , 
        \wBIn3[1] , \wBIn3[0] }), .HiOut({\wBMid2[31] , \wBMid2[30] , 
        \wBMid2[29] , \wBMid2[28] , \wBMid2[27] , \wBMid2[26] , \wBMid2[25] , 
        \wBMid2[24] , \wBMid2[23] , \wBMid2[22] , \wBMid2[21] , \wBMid2[20] , 
        \wBMid2[19] , \wBMid2[18] , \wBMid2[17] , \wBMid2[16] , \wBMid2[15] , 
        \wBMid2[14] , \wBMid2[13] , \wBMid2[12] , \wBMid2[11] , \wBMid2[10] , 
        \wBMid2[9] , \wBMid2[8] , \wBMid2[7] , \wBMid2[6] , \wBMid2[5] , 
        \wBMid2[4] , \wBMid2[3] , \wBMid2[2] , \wBMid2[1] , \wBMid2[0] }), 
        .LoOut({\wAMid3[31] , \wAMid3[30] , \wAMid3[29] , \wAMid3[28] , 
        \wAMid3[27] , \wAMid3[26] , \wAMid3[25] , \wAMid3[24] , \wAMid3[23] , 
        \wAMid3[22] , \wAMid3[21] , \wAMid3[20] , \wAMid3[19] , \wAMid3[18] , 
        \wAMid3[17] , \wAMid3[16] , \wAMid3[15] , \wAMid3[14] , \wAMid3[13] , 
        \wAMid3[12] , \wAMid3[11] , \wAMid3[10] , \wAMid3[9] , \wAMid3[8] , 
        \wAMid3[7] , \wAMid3[6] , \wAMid3[5] , \wAMid3[4] , \wAMid3[3] , 
        \wAMid3[2] , \wAMid3[1] , \wAMid3[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn4[31] , 
        \wAIn4[30] , \wAIn4[29] , \wAIn4[28] , \wAIn4[27] , \wAIn4[26] , 
        \wAIn4[25] , \wAIn4[24] , \wAIn4[23] , \wAIn4[22] , \wAIn4[21] , 
        \wAIn4[20] , \wAIn4[19] , \wAIn4[18] , \wAIn4[17] , \wAIn4[16] , 
        \wAIn4[15] , \wAIn4[14] , \wAIn4[13] , \wAIn4[12] , \wAIn4[11] , 
        \wAIn4[10] , \wAIn4[9] , \wAIn4[8] , \wAIn4[7] , \wAIn4[6] , 
        \wAIn4[5] , \wAIn4[4] , \wAIn4[3] , \wAIn4[2] , \wAIn4[1] , \wAIn4[0] 
        }), .BIn({\wBIn4[31] , \wBIn4[30] , \wBIn4[29] , \wBIn4[28] , 
        \wBIn4[27] , \wBIn4[26] , \wBIn4[25] , \wBIn4[24] , \wBIn4[23] , 
        \wBIn4[22] , \wBIn4[21] , \wBIn4[20] , \wBIn4[19] , \wBIn4[18] , 
        \wBIn4[17] , \wBIn4[16] , \wBIn4[15] , \wBIn4[14] , \wBIn4[13] , 
        \wBIn4[12] , \wBIn4[11] , \wBIn4[10] , \wBIn4[9] , \wBIn4[8] , 
        \wBIn4[7] , \wBIn4[6] , \wBIn4[5] , \wBIn4[4] , \wBIn4[3] , \wBIn4[2] , 
        \wBIn4[1] , \wBIn4[0] }), .HiOut({\wBMid3[31] , \wBMid3[30] , 
        \wBMid3[29] , \wBMid3[28] , \wBMid3[27] , \wBMid3[26] , \wBMid3[25] , 
        \wBMid3[24] , \wBMid3[23] , \wBMid3[22] , \wBMid3[21] , \wBMid3[20] , 
        \wBMid3[19] , \wBMid3[18] , \wBMid3[17] , \wBMid3[16] , \wBMid3[15] , 
        \wBMid3[14] , \wBMid3[13] , \wBMid3[12] , \wBMid3[11] , \wBMid3[10] , 
        \wBMid3[9] , \wBMid3[8] , \wBMid3[7] , \wBMid3[6] , \wBMid3[5] , 
        \wBMid3[4] , \wBMid3[3] , \wBMid3[2] , \wBMid3[1] , \wBMid3[0] }), 
        .LoOut({\wAMid4[31] , \wAMid4[30] , \wAMid4[29] , \wAMid4[28] , 
        \wAMid4[27] , \wAMid4[26] , \wAMid4[25] , \wAMid4[24] , \wAMid4[23] , 
        \wAMid4[22] , \wAMid4[21] , \wAMid4[20] , \wAMid4[19] , \wAMid4[18] , 
        \wAMid4[17] , \wAMid4[16] , \wAMid4[15] , \wAMid4[14] , \wAMid4[13] , 
        \wAMid4[12] , \wAMid4[11] , \wAMid4[10] , \wAMid4[9] , \wAMid4[8] , 
        \wAMid4[7] , \wAMid4[6] , \wAMid4[5] , \wAMid4[4] , \wAMid4[3] , 
        \wAMid4[2] , \wAMid4[1] , \wAMid4[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn12[31] , \wAIn12[30] , \wAIn12[29] , \wAIn12[28] , \wAIn12[27] , 
        \wAIn12[26] , \wAIn12[25] , \wAIn12[24] , \wAIn12[23] , \wAIn12[22] , 
        \wAIn12[21] , \wAIn12[20] , \wAIn12[19] , \wAIn12[18] , \wAIn12[17] , 
        \wAIn12[16] , \wAIn12[15] , \wAIn12[14] , \wAIn12[13] , \wAIn12[12] , 
        \wAIn12[11] , \wAIn12[10] , \wAIn12[9] , \wAIn12[8] , \wAIn12[7] , 
        \wAIn12[6] , \wAIn12[5] , \wAIn12[4] , \wAIn12[3] , \wAIn12[2] , 
        \wAIn12[1] , \wAIn12[0] }), .BIn({\wBIn12[31] , \wBIn12[30] , 
        \wBIn12[29] , \wBIn12[28] , \wBIn12[27] , \wBIn12[26] , \wBIn12[25] , 
        \wBIn12[24] , \wBIn12[23] , \wBIn12[22] , \wBIn12[21] , \wBIn12[20] , 
        \wBIn12[19] , \wBIn12[18] , \wBIn12[17] , \wBIn12[16] , \wBIn12[15] , 
        \wBIn12[14] , \wBIn12[13] , \wBIn12[12] , \wBIn12[11] , \wBIn12[10] , 
        \wBIn12[9] , \wBIn12[8] , \wBIn12[7] , \wBIn12[6] , \wBIn12[5] , 
        \wBIn12[4] , \wBIn12[3] , \wBIn12[2] , \wBIn12[1] , \wBIn12[0] }), 
        .HiOut({\wBMid11[31] , \wBMid11[30] , \wBMid11[29] , \wBMid11[28] , 
        \wBMid11[27] , \wBMid11[26] , \wBMid11[25] , \wBMid11[24] , 
        \wBMid11[23] , \wBMid11[22] , \wBMid11[21] , \wBMid11[20] , 
        \wBMid11[19] , \wBMid11[18] , \wBMid11[17] , \wBMid11[16] , 
        \wBMid11[15] , \wBMid11[14] , \wBMid11[13] , \wBMid11[12] , 
        \wBMid11[11] , \wBMid11[10] , \wBMid11[9] , \wBMid11[8] , \wBMid11[7] , 
        \wBMid11[6] , \wBMid11[5] , \wBMid11[4] , \wBMid11[3] , \wBMid11[2] , 
        \wBMid11[1] , \wBMid11[0] }), .LoOut({\wAMid12[31] , \wAMid12[30] , 
        \wAMid12[29] , \wAMid12[28] , \wAMid12[27] , \wAMid12[26] , 
        \wAMid12[25] , \wAMid12[24] , \wAMid12[23] , \wAMid12[22] , 
        \wAMid12[21] , \wAMid12[20] , \wAMid12[19] , \wAMid12[18] , 
        \wAMid12[17] , \wAMid12[16] , \wAMid12[15] , \wAMid12[14] , 
        \wAMid12[13] , \wAMid12[12] , \wAMid12[11] , \wAMid12[10] , 
        \wAMid12[9] , \wAMid12[8] , \wAMid12[7] , \wAMid12[6] , \wAMid12[5] , 
        \wAMid12[4] , \wAMid12[3] , \wAMid12[2] , \wAMid12[1] , \wAMid12[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid8[31] , 
        \wAMid8[30] , \wAMid8[29] , \wAMid8[28] , \wAMid8[27] , \wAMid8[26] , 
        \wAMid8[25] , \wAMid8[24] , \wAMid8[23] , \wAMid8[22] , \wAMid8[21] , 
        \wAMid8[20] , \wAMid8[19] , \wAMid8[18] , \wAMid8[17] , \wAMid8[16] , 
        \wAMid8[15] , \wAMid8[14] , \wAMid8[13] , \wAMid8[12] , \wAMid8[11] , 
        \wAMid8[10] , \wAMid8[9] , \wAMid8[8] , \wAMid8[7] , \wAMid8[6] , 
        \wAMid8[5] , \wAMid8[4] , \wAMid8[3] , \wAMid8[2] , \wAMid8[1] , 
        \wAMid8[0] }), .BIn({\wBMid8[31] , \wBMid8[30] , \wBMid8[29] , 
        \wBMid8[28] , \wBMid8[27] , \wBMid8[26] , \wBMid8[25] , \wBMid8[24] , 
        \wBMid8[23] , \wBMid8[22] , \wBMid8[21] , \wBMid8[20] , \wBMid8[19] , 
        \wBMid8[18] , \wBMid8[17] , \wBMid8[16] , \wBMid8[15] , \wBMid8[14] , 
        \wBMid8[13] , \wBMid8[12] , \wBMid8[11] , \wBMid8[10] , \wBMid8[9] , 
        \wBMid8[8] , \wBMid8[7] , \wBMid8[6] , \wBMid8[5] , \wBMid8[4] , 
        \wBMid8[3] , \wBMid8[2] , \wBMid8[1] , \wBMid8[0] }), .HiOut({
        \wRegInB8[31] , \wRegInB8[30] , \wRegInB8[29] , \wRegInB8[28] , 
        \wRegInB8[27] , \wRegInB8[26] , \wRegInB8[25] , \wRegInB8[24] , 
        \wRegInB8[23] , \wRegInB8[22] , \wRegInB8[21] , \wRegInB8[20] , 
        \wRegInB8[19] , \wRegInB8[18] , \wRegInB8[17] , \wRegInB8[16] , 
        \wRegInB8[15] , \wRegInB8[14] , \wRegInB8[13] , \wRegInB8[12] , 
        \wRegInB8[11] , \wRegInB8[10] , \wRegInB8[9] , \wRegInB8[8] , 
        \wRegInB8[7] , \wRegInB8[6] , \wRegInB8[5] , \wRegInB8[4] , 
        \wRegInB8[3] , \wRegInB8[2] , \wRegInB8[1] , \wRegInB8[0] }), .LoOut({
        \wRegInA9[31] , \wRegInA9[30] , \wRegInA9[29] , \wRegInA9[28] , 
        \wRegInA9[27] , \wRegInA9[26] , \wRegInA9[25] , \wRegInA9[24] , 
        \wRegInA9[23] , \wRegInA9[22] , \wRegInA9[21] , \wRegInA9[20] , 
        \wRegInA9[19] , \wRegInA9[18] , \wRegInA9[17] , \wRegInA9[16] , 
        \wRegInA9[15] , \wRegInA9[14] , \wRegInA9[13] , \wRegInA9[12] , 
        \wRegInA9[11] , \wRegInA9[10] , \wRegInA9[9] , \wRegInA9[8] , 
        \wRegInA9[7] , \wRegInA9[6] , \wRegInA9[5] , \wRegInA9[4] , 
        \wRegInA9[3] , \wRegInA9[2] , \wRegInA9[1] , \wRegInA9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_32 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink33[31] , \ScanLink33[30] , \ScanLink33[29] , 
        \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , \ScanLink33[25] , 
        \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , \ScanLink33[21] , 
        \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , \ScanLink33[17] , 
        \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , \ScanLink33[13] , 
        \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , \ScanLink33[9] , 
        \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , \ScanLink33[5] , 
        \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , \ScanLink33[1] , 
        \ScanLink33[0] }), .ScanOut({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB15[31] , \wRegInB15[30] , 
        \wRegInB15[29] , \wRegInB15[28] , \wRegInB15[27] , \wRegInB15[26] , 
        \wRegInB15[25] , \wRegInB15[24] , \wRegInB15[23] , \wRegInB15[22] , 
        \wRegInB15[21] , \wRegInB15[20] , \wRegInB15[19] , \wRegInB15[18] , 
        \wRegInB15[17] , \wRegInB15[16] , \wRegInB15[15] , \wRegInB15[14] , 
        \wRegInB15[13] , \wRegInB15[12] , \wRegInB15[11] , \wRegInB15[10] , 
        \wRegInB15[9] , \wRegInB15[8] , \wRegInB15[7] , \wRegInB15[6] , 
        \wRegInB15[5] , \wRegInB15[4] , \wRegInB15[3] , \wRegInB15[2] , 
        \wRegInB15[1] , \wRegInB15[0] }), .Out({\wBIn15[31] , \wBIn15[30] , 
        \wBIn15[29] , \wBIn15[28] , \wBIn15[27] , \wBIn15[26] , \wBIn15[25] , 
        \wBIn15[24] , \wBIn15[23] , \wBIn15[22] , \wBIn15[21] , \wBIn15[20] , 
        \wBIn15[19] , \wBIn15[18] , \wBIn15[17] , \wBIn15[16] , \wBIn15[15] , 
        \wBIn15[14] , \wBIn15[13] , \wBIn15[12] , \wBIn15[11] , \wBIn15[10] , 
        \wBIn15[9] , \wBIn15[8] , \wBIn15[7] , \wBIn15[6] , \wBIn15[5] , 
        \wBIn15[4] , \wBIn15[3] , \wBIn15[2] , \wBIn15[1] , \wBIn15[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_15 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[31] , \ScanLink16[30] , \ScanLink16[29] , 
        \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , \ScanLink16[25] , 
        \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , \ScanLink16[21] , 
        \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , \ScanLink16[17] , 
        \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , \ScanLink16[13] , 
        \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , \ScanLink16[9] , 
        \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA24[31] , \wRegInA24[30] , 
        \wRegInA24[29] , \wRegInA24[28] , \wRegInA24[27] , \wRegInA24[26] , 
        \wRegInA24[25] , \wRegInA24[24] , \wRegInA24[23] , \wRegInA24[22] , 
        \wRegInA24[21] , \wRegInA24[20] , \wRegInA24[19] , \wRegInA24[18] , 
        \wRegInA24[17] , \wRegInA24[16] , \wRegInA24[15] , \wRegInA24[14] , 
        \wRegInA24[13] , \wRegInA24[12] , \wRegInA24[11] , \wRegInA24[10] , 
        \wRegInA24[9] , \wRegInA24[8] , \wRegInA24[7] , \wRegInA24[6] , 
        \wRegInA24[5] , \wRegInA24[4] , \wRegInA24[3] , \wRegInA24[2] , 
        \wRegInA24[1] , \wRegInA24[0] }), .Out({\wAIn24[31] , \wAIn24[30] , 
        \wAIn24[29] , \wAIn24[28] , \wAIn24[27] , \wAIn24[26] , \wAIn24[25] , 
        \wAIn24[24] , \wAIn24[23] , \wAIn24[22] , \wAIn24[21] , \wAIn24[20] , 
        \wAIn24[19] , \wAIn24[18] , \wAIn24[17] , \wAIn24[16] , \wAIn24[15] , 
        \wAIn24[14] , \wAIn24[13] , \wAIn24[12] , \wAIn24[11] , \wAIn24[10] , 
        \wAIn24[9] , \wAIn24[8] , \wAIn24[7] , \wAIn24[6] , \wAIn24[5] , 
        \wAIn24[4] , \wAIn24[3] , \wAIn24[2] , \wAIn24[1] , \wAIn24[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_29 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink30[31] , \ScanLink30[30] , \ScanLink30[29] , 
        \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , \ScanLink30[25] , 
        \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , \ScanLink30[21] , 
        \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , \ScanLink30[17] , 
        \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , \ScanLink30[13] , 
        \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , \ScanLink30[9] , 
        \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , \ScanLink30[5] , 
        \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , \ScanLink30[1] , 
        \ScanLink30[0] }), .ScanOut({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA17[31] , \wRegInA17[30] , 
        \wRegInA17[29] , \wRegInA17[28] , \wRegInA17[27] , \wRegInA17[26] , 
        \wRegInA17[25] , \wRegInA17[24] , \wRegInA17[23] , \wRegInA17[22] , 
        \wRegInA17[21] , \wRegInA17[20] , \wRegInA17[19] , \wRegInA17[18] , 
        \wRegInA17[17] , \wRegInA17[16] , \wRegInA17[15] , \wRegInA17[14] , 
        \wRegInA17[13] , \wRegInA17[12] , \wRegInA17[11] , \wRegInA17[10] , 
        \wRegInA17[9] , \wRegInA17[8] , \wRegInA17[7] , \wRegInA17[6] , 
        \wRegInA17[5] , \wRegInA17[4] , \wRegInA17[3] , \wRegInA17[2] , 
        \wRegInA17[1] , \wRegInA17[0] }), .Out({\wAIn17[31] , \wAIn17[30] , 
        \wAIn17[29] , \wAIn17[28] , \wAIn17[27] , \wAIn17[26] , \wAIn17[25] , 
        \wAIn17[24] , \wAIn17[23] , \wAIn17[22] , \wAIn17[21] , \wAIn17[20] , 
        \wAIn17[19] , \wAIn17[18] , \wAIn17[17] , \wAIn17[16] , \wAIn17[15] , 
        \wAIn17[14] , \wAIn17[13] , \wAIn17[12] , \wAIn17[11] , \wAIn17[10] , 
        \wAIn17[9] , \wAIn17[8] , \wAIn17[7] , \wAIn17[6] , \wAIn17[5] , 
        \wAIn17[4] , \wAIn17[3] , \wAIn17[2] , \wAIn17[1] , \wAIn17[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_60 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink61[31] , \ScanLink61[30] , \ScanLink61[29] , 
        \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , \ScanLink61[25] , 
        \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , \ScanLink61[21] , 
        \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , \ScanLink61[17] , 
        \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , \ScanLink61[13] , 
        \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , \ScanLink61[9] , 
        \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , \ScanLink61[5] , 
        \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , \ScanLink61[1] , 
        \ScanLink61[0] }), .ScanOut({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB1[31] , \wRegInB1[30] , 
        \wRegInB1[29] , \wRegInB1[28] , \wRegInB1[27] , \wRegInB1[26] , 
        \wRegInB1[25] , \wRegInB1[24] , \wRegInB1[23] , \wRegInB1[22] , 
        \wRegInB1[21] , \wRegInB1[20] , \wRegInB1[19] , \wRegInB1[18] , 
        \wRegInB1[17] , \wRegInB1[16] , \wRegInB1[15] , \wRegInB1[14] , 
        \wRegInB1[13] , \wRegInB1[12] , \wRegInB1[11] , \wRegInB1[10] , 
        \wRegInB1[9] , \wRegInB1[8] , \wRegInB1[7] , \wRegInB1[6] , 
        \wRegInB1[5] , \wRegInB1[4] , \wRegInB1[3] , \wRegInB1[2] , 
        \wRegInB1[1] , \wRegInB1[0] }), .Out({\wBIn1[31] , \wBIn1[30] , 
        \wBIn1[29] , \wBIn1[28] , \wBIn1[27] , \wBIn1[26] , \wBIn1[25] , 
        \wBIn1[24] , \wBIn1[23] , \wBIn1[22] , \wBIn1[21] , \wBIn1[20] , 
        \wBIn1[19] , \wBIn1[18] , \wBIn1[17] , \wBIn1[16] , \wBIn1[15] , 
        \wBIn1[14] , \wBIn1[13] , \wBIn1[12] , \wBIn1[11] , \wBIn1[10] , 
        \wBIn1[9] , \wBIn1[8] , \wBIn1[7] , \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , 
        \wBIn1[3] , \wBIn1[2] , \wBIn1[1] , \wBIn1[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_4 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[31] , \ScanLink5[30] , \ScanLink5[29] , 
        \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , \ScanLink5[25] , 
        \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , \ScanLink5[21] , 
        \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , \ScanLink5[17] , 
        \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , \ScanLink5[13] , 
        \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , \ScanLink5[9] , 
        \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB29[31] , \wRegInB29[30] , 
        \wRegInB29[29] , \wRegInB29[28] , \wRegInB29[27] , \wRegInB29[26] , 
        \wRegInB29[25] , \wRegInB29[24] , \wRegInB29[23] , \wRegInB29[22] , 
        \wRegInB29[21] , \wRegInB29[20] , \wRegInB29[19] , \wRegInB29[18] , 
        \wRegInB29[17] , \wRegInB29[16] , \wRegInB29[15] , \wRegInB29[14] , 
        \wRegInB29[13] , \wRegInB29[12] , \wRegInB29[11] , \wRegInB29[10] , 
        \wRegInB29[9] , \wRegInB29[8] , \wRegInB29[7] , \wRegInB29[6] , 
        \wRegInB29[5] , \wRegInB29[4] , \wRegInB29[3] , \wRegInB29[2] , 
        \wRegInB29[1] , \wRegInB29[0] }), .Out({\wBIn29[31] , \wBIn29[30] , 
        \wBIn29[29] , \wBIn29[28] , \wBIn29[27] , \wBIn29[26] , \wBIn29[25] , 
        \wBIn29[24] , \wBIn29[23] , \wBIn29[22] , \wBIn29[21] , \wBIn29[20] , 
        \wBIn29[19] , \wBIn29[18] , \wBIn29[17] , \wBIn29[16] , \wBIn29[15] , 
        \wBIn29[14] , \wBIn29[13] , \wBIn29[12] , \wBIn29[11] , \wBIn29[10] , 
        \wBIn29[9] , \wBIn29[8] , \wBIn29[7] , \wBIn29[6] , \wBIn29[5] , 
        \wBIn29[4] , \wBIn29[3] , \wBIn29[2] , \wBIn29[1] , \wBIn29[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn15[31] , \wAIn15[30] , \wAIn15[29] , \wAIn15[28] , \wAIn15[27] , 
        \wAIn15[26] , \wAIn15[25] , \wAIn15[24] , \wAIn15[23] , \wAIn15[22] , 
        \wAIn15[21] , \wAIn15[20] , \wAIn15[19] , \wAIn15[18] , \wAIn15[17] , 
        \wAIn15[16] , \wAIn15[15] , \wAIn15[14] , \wAIn15[13] , \wAIn15[12] , 
        \wAIn15[11] , \wAIn15[10] , \wAIn15[9] , \wAIn15[8] , \wAIn15[7] , 
        \wAIn15[6] , \wAIn15[5] , \wAIn15[4] , \wAIn15[3] , \wAIn15[2] , 
        \wAIn15[1] , \wAIn15[0] }), .BIn({\wBIn15[31] , \wBIn15[30] , 
        \wBIn15[29] , \wBIn15[28] , \wBIn15[27] , \wBIn15[26] , \wBIn15[25] , 
        \wBIn15[24] , \wBIn15[23] , \wBIn15[22] , \wBIn15[21] , \wBIn15[20] , 
        \wBIn15[19] , \wBIn15[18] , \wBIn15[17] , \wBIn15[16] , \wBIn15[15] , 
        \wBIn15[14] , \wBIn15[13] , \wBIn15[12] , \wBIn15[11] , \wBIn15[10] , 
        \wBIn15[9] , \wBIn15[8] , \wBIn15[7] , \wBIn15[6] , \wBIn15[5] , 
        \wBIn15[4] , \wBIn15[3] , \wBIn15[2] , \wBIn15[1] , \wBIn15[0] }), 
        .HiOut({\wBMid14[31] , \wBMid14[30] , \wBMid14[29] , \wBMid14[28] , 
        \wBMid14[27] , \wBMid14[26] , \wBMid14[25] , \wBMid14[24] , 
        \wBMid14[23] , \wBMid14[22] , \wBMid14[21] , \wBMid14[20] , 
        \wBMid14[19] , \wBMid14[18] , \wBMid14[17] , \wBMid14[16] , 
        \wBMid14[15] , \wBMid14[14] , \wBMid14[13] , \wBMid14[12] , 
        \wBMid14[11] , \wBMid14[10] , \wBMid14[9] , \wBMid14[8] , \wBMid14[7] , 
        \wBMid14[6] , \wBMid14[5] , \wBMid14[4] , \wBMid14[3] , \wBMid14[2] , 
        \wBMid14[1] , \wBMid14[0] }), .LoOut({\wAMid15[31] , \wAMid15[30] , 
        \wAMid15[29] , \wAMid15[28] , \wAMid15[27] , \wAMid15[26] , 
        \wAMid15[25] , \wAMid15[24] , \wAMid15[23] , \wAMid15[22] , 
        \wAMid15[21] , \wAMid15[20] , \wAMid15[19] , \wAMid15[18] , 
        \wAMid15[17] , \wAMid15[16] , \wAMid15[15] , \wAMid15[14] , 
        \wAMid15[13] , \wAMid15[12] , \wAMid15[11] , \wAMid15[10] , 
        \wAMid15[9] , \wAMid15[8] , \wAMid15[7] , \wAMid15[6] , \wAMid15[5] , 
        \wAMid15[4] , \wAMid15[3] , \wAMid15[2] , \wAMid15[1] , \wAMid15[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn20[31] , \wAIn20[30] , \wAIn20[29] , \wAIn20[28] , \wAIn20[27] , 
        \wAIn20[26] , \wAIn20[25] , \wAIn20[24] , \wAIn20[23] , \wAIn20[22] , 
        \wAIn20[21] , \wAIn20[20] , \wAIn20[19] , \wAIn20[18] , \wAIn20[17] , 
        \wAIn20[16] , \wAIn20[15] , \wAIn20[14] , \wAIn20[13] , \wAIn20[12] , 
        \wAIn20[11] , \wAIn20[10] , \wAIn20[9] , \wAIn20[8] , \wAIn20[7] , 
        \wAIn20[6] , \wAIn20[5] , \wAIn20[4] , \wAIn20[3] , \wAIn20[2] , 
        \wAIn20[1] , \wAIn20[0] }), .BIn({\wBIn20[31] , \wBIn20[30] , 
        \wBIn20[29] , \wBIn20[28] , \wBIn20[27] , \wBIn20[26] , \wBIn20[25] , 
        \wBIn20[24] , \wBIn20[23] , \wBIn20[22] , \wBIn20[21] , \wBIn20[20] , 
        \wBIn20[19] , \wBIn20[18] , \wBIn20[17] , \wBIn20[16] , \wBIn20[15] , 
        \wBIn20[14] , \wBIn20[13] , \wBIn20[12] , \wBIn20[11] , \wBIn20[10] , 
        \wBIn20[9] , \wBIn20[8] , \wBIn20[7] , \wBIn20[6] , \wBIn20[5] , 
        \wBIn20[4] , \wBIn20[3] , \wBIn20[2] , \wBIn20[1] , \wBIn20[0] }), 
        .HiOut({\wBMid19[31] , \wBMid19[30] , \wBMid19[29] , \wBMid19[28] , 
        \wBMid19[27] , \wBMid19[26] , \wBMid19[25] , \wBMid19[24] , 
        \wBMid19[23] , \wBMid19[22] , \wBMid19[21] , \wBMid19[20] , 
        \wBMid19[19] , \wBMid19[18] , \wBMid19[17] , \wBMid19[16] , 
        \wBMid19[15] , \wBMid19[14] , \wBMid19[13] , \wBMid19[12] , 
        \wBMid19[11] , \wBMid19[10] , \wBMid19[9] , \wBMid19[8] , \wBMid19[7] , 
        \wBMid19[6] , \wBMid19[5] , \wBMid19[4] , \wBMid19[3] , \wBMid19[2] , 
        \wBMid19[1] , \wBMid19[0] }), .LoOut({\wAMid20[31] , \wAMid20[30] , 
        \wAMid20[29] , \wAMid20[28] , \wAMid20[27] , \wAMid20[26] , 
        \wAMid20[25] , \wAMid20[24] , \wAMid20[23] , \wAMid20[22] , 
        \wAMid20[21] , \wAMid20[20] , \wAMid20[19] , \wAMid20[18] , 
        \wAMid20[17] , \wAMid20[16] , \wAMid20[15] , \wAMid20[14] , 
        \wAMid20[13] , \wAMid20[12] , \wAMid20[11] , \wAMid20[10] , 
        \wAMid20[9] , \wAMid20[8] , \wAMid20[7] , \wAMid20[6] , \wAMid20[5] , 
        \wAMid20[4] , \wAMid20[3] , \wAMid20[2] , \wAMid20[1] , \wAMid20[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn27[31] , \wAIn27[30] , \wAIn27[29] , \wAIn27[28] , \wAIn27[27] , 
        \wAIn27[26] , \wAIn27[25] , \wAIn27[24] , \wAIn27[23] , \wAIn27[22] , 
        \wAIn27[21] , \wAIn27[20] , \wAIn27[19] , \wAIn27[18] , \wAIn27[17] , 
        \wAIn27[16] , \wAIn27[15] , \wAIn27[14] , \wAIn27[13] , \wAIn27[12] , 
        \wAIn27[11] , \wAIn27[10] , \wAIn27[9] , \wAIn27[8] , \wAIn27[7] , 
        \wAIn27[6] , \wAIn27[5] , \wAIn27[4] , \wAIn27[3] , \wAIn27[2] , 
        \wAIn27[1] , \wAIn27[0] }), .BIn({\wBIn27[31] , \wBIn27[30] , 
        \wBIn27[29] , \wBIn27[28] , \wBIn27[27] , \wBIn27[26] , \wBIn27[25] , 
        \wBIn27[24] , \wBIn27[23] , \wBIn27[22] , \wBIn27[21] , \wBIn27[20] , 
        \wBIn27[19] , \wBIn27[18] , \wBIn27[17] , \wBIn27[16] , \wBIn27[15] , 
        \wBIn27[14] , \wBIn27[13] , \wBIn27[12] , \wBIn27[11] , \wBIn27[10] , 
        \wBIn27[9] , \wBIn27[8] , \wBIn27[7] , \wBIn27[6] , \wBIn27[5] , 
        \wBIn27[4] , \wBIn27[3] , \wBIn27[2] , \wBIn27[1] , \wBIn27[0] }), 
        .HiOut({\wBMid26[31] , \wBMid26[30] , \wBMid26[29] , \wBMid26[28] , 
        \wBMid26[27] , \wBMid26[26] , \wBMid26[25] , \wBMid26[24] , 
        \wBMid26[23] , \wBMid26[22] , \wBMid26[21] , \wBMid26[20] , 
        \wBMid26[19] , \wBMid26[18] , \wBMid26[17] , \wBMid26[16] , 
        \wBMid26[15] , \wBMid26[14] , \wBMid26[13] , \wBMid26[12] , 
        \wBMid26[11] , \wBMid26[10] , \wBMid26[9] , \wBMid26[8] , \wBMid26[7] , 
        \wBMid26[6] , \wBMid26[5] , \wBMid26[4] , \wBMid26[3] , \wBMid26[2] , 
        \wBMid26[1] , \wBMid26[0] }), .LoOut({\wAMid27[31] , \wAMid27[30] , 
        \wAMid27[29] , \wAMid27[28] , \wAMid27[27] , \wAMid27[26] , 
        \wAMid27[25] , \wAMid27[24] , \wAMid27[23] , \wAMid27[22] , 
        \wAMid27[21] , \wAMid27[20] , \wAMid27[19] , \wAMid27[18] , 
        \wAMid27[17] , \wAMid27[16] , \wAMid27[15] , \wAMid27[14] , 
        \wAMid27[13] , \wAMid27[12] , \wAMid27[11] , \wAMid27[10] , 
        \wAMid27[9] , \wAMid27[8] , \wAMid27[7] , \wAMid27[6] , \wAMid27[5] , 
        \wAMid27[4] , \wAMid27[3] , \wAMid27[2] , \wAMid27[1] , \wAMid27[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid22[31] , \wAMid22[30] , \wAMid22[29] , \wAMid22[28] , 
        \wAMid22[27] , \wAMid22[26] , \wAMid22[25] , \wAMid22[24] , 
        \wAMid22[23] , \wAMid22[22] , \wAMid22[21] , \wAMid22[20] , 
        \wAMid22[19] , \wAMid22[18] , \wAMid22[17] , \wAMid22[16] , 
        \wAMid22[15] , \wAMid22[14] , \wAMid22[13] , \wAMid22[12] , 
        \wAMid22[11] , \wAMid22[10] , \wAMid22[9] , \wAMid22[8] , \wAMid22[7] , 
        \wAMid22[6] , \wAMid22[5] , \wAMid22[4] , \wAMid22[3] , \wAMid22[2] , 
        \wAMid22[1] , \wAMid22[0] }), .BIn({\wBMid22[31] , \wBMid22[30] , 
        \wBMid22[29] , \wBMid22[28] , \wBMid22[27] , \wBMid22[26] , 
        \wBMid22[25] , \wBMid22[24] , \wBMid22[23] , \wBMid22[22] , 
        \wBMid22[21] , \wBMid22[20] , \wBMid22[19] , \wBMid22[18] , 
        \wBMid22[17] , \wBMid22[16] , \wBMid22[15] , \wBMid22[14] , 
        \wBMid22[13] , \wBMid22[12] , \wBMid22[11] , \wBMid22[10] , 
        \wBMid22[9] , \wBMid22[8] , \wBMid22[7] , \wBMid22[6] , \wBMid22[5] , 
        \wBMid22[4] , \wBMid22[3] , \wBMid22[2] , \wBMid22[1] , \wBMid22[0] }), 
        .HiOut({\wRegInB22[31] , \wRegInB22[30] , \wRegInB22[29] , 
        \wRegInB22[28] , \wRegInB22[27] , \wRegInB22[26] , \wRegInB22[25] , 
        \wRegInB22[24] , \wRegInB22[23] , \wRegInB22[22] , \wRegInB22[21] , 
        \wRegInB22[20] , \wRegInB22[19] , \wRegInB22[18] , \wRegInB22[17] , 
        \wRegInB22[16] , \wRegInB22[15] , \wRegInB22[14] , \wRegInB22[13] , 
        \wRegInB22[12] , \wRegInB22[11] , \wRegInB22[10] , \wRegInB22[9] , 
        \wRegInB22[8] , \wRegInB22[7] , \wRegInB22[6] , \wRegInB22[5] , 
        \wRegInB22[4] , \wRegInB22[3] , \wRegInB22[2] , \wRegInB22[1] , 
        \wRegInB22[0] }), .LoOut({\wRegInA23[31] , \wRegInA23[30] , 
        \wRegInA23[29] , \wRegInA23[28] , \wRegInA23[27] , \wRegInA23[26] , 
        \wRegInA23[25] , \wRegInA23[24] , \wRegInA23[23] , \wRegInA23[22] , 
        \wRegInA23[21] , \wRegInA23[20] , \wRegInA23[19] , \wRegInA23[18] , 
        \wRegInA23[17] , \wRegInA23[16] , \wRegInA23[15] , \wRegInA23[14] , 
        \wRegInA23[13] , \wRegInA23[12] , \wRegInA23[11] , \wRegInA23[10] , 
        \wRegInA23[9] , \wRegInA23[8] , \wRegInA23[7] , \wRegInA23[6] , 
        \wRegInA23[5] , \wRegInA23[4] , \wRegInA23[3] , \wRegInA23[2] , 
        \wRegInA23[1] , \wRegInA23[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_47 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink48[31] , \ScanLink48[30] , \ScanLink48[29] , 
        \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , \ScanLink48[25] , 
        \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , \ScanLink48[21] , 
        \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , \ScanLink48[17] , 
        \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , \ScanLink48[13] , 
        \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , \ScanLink48[9] , 
        \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , \ScanLink48[5] , 
        \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , \ScanLink48[1] , 
        \ScanLink48[0] }), .ScanOut({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA8[31] , \wRegInA8[30] , 
        \wRegInA8[29] , \wRegInA8[28] , \wRegInA8[27] , \wRegInA8[26] , 
        \wRegInA8[25] , \wRegInA8[24] , \wRegInA8[23] , \wRegInA8[22] , 
        \wRegInA8[21] , \wRegInA8[20] , \wRegInA8[19] , \wRegInA8[18] , 
        \wRegInA8[17] , \wRegInA8[16] , \wRegInA8[15] , \wRegInA8[14] , 
        \wRegInA8[13] , \wRegInA8[12] , \wRegInA8[11] , \wRegInA8[10] , 
        \wRegInA8[9] , \wRegInA8[8] , \wRegInA8[7] , \wRegInA8[6] , 
        \wRegInA8[5] , \wRegInA8[4] , \wRegInA8[3] , \wRegInA8[2] , 
        \wRegInA8[1] , \wRegInA8[0] }), .Out({\wAIn8[31] , \wAIn8[30] , 
        \wAIn8[29] , \wAIn8[28] , \wAIn8[27] , \wAIn8[26] , \wAIn8[25] , 
        \wAIn8[24] , \wAIn8[23] , \wAIn8[22] , \wAIn8[21] , \wAIn8[20] , 
        \wAIn8[19] , \wAIn8[18] , \wAIn8[17] , \wAIn8[16] , \wAIn8[15] , 
        \wAIn8[14] , \wAIn8[13] , \wAIn8[12] , \wAIn8[11] , \wAIn8[10] , 
        \wAIn8[9] , \wAIn8[8] , \wAIn8[7] , \wAIn8[6] , \wAIn8[5] , \wAIn8[4] , 
        \wAIn8[3] , \wAIn8[2] , \wAIn8[1] , \wAIn8[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid1[31] , 
        \wAMid1[30] , \wAMid1[29] , \wAMid1[28] , \wAMid1[27] , \wAMid1[26] , 
        \wAMid1[25] , \wAMid1[24] , \wAMid1[23] , \wAMid1[22] , \wAMid1[21] , 
        \wAMid1[20] , \wAMid1[19] , \wAMid1[18] , \wAMid1[17] , \wAMid1[16] , 
        \wAMid1[15] , \wAMid1[14] , \wAMid1[13] , \wAMid1[12] , \wAMid1[11] , 
        \wAMid1[10] , \wAMid1[9] , \wAMid1[8] , \wAMid1[7] , \wAMid1[6] , 
        \wAMid1[5] , \wAMid1[4] , \wAMid1[3] , \wAMid1[2] , \wAMid1[1] , 
        \wAMid1[0] }), .BIn({\wBMid1[31] , \wBMid1[30] , \wBMid1[29] , 
        \wBMid1[28] , \wBMid1[27] , \wBMid1[26] , \wBMid1[25] , \wBMid1[24] , 
        \wBMid1[23] , \wBMid1[22] , \wBMid1[21] , \wBMid1[20] , \wBMid1[19] , 
        \wBMid1[18] , \wBMid1[17] , \wBMid1[16] , \wBMid1[15] , \wBMid1[14] , 
        \wBMid1[13] , \wBMid1[12] , \wBMid1[11] , \wBMid1[10] , \wBMid1[9] , 
        \wBMid1[8] , \wBMid1[7] , \wBMid1[6] , \wBMid1[5] , \wBMid1[4] , 
        \wBMid1[3] , \wBMid1[2] , \wBMid1[1] , \wBMid1[0] }), .HiOut({
        \wRegInB1[31] , \wRegInB1[30] , \wRegInB1[29] , \wRegInB1[28] , 
        \wRegInB1[27] , \wRegInB1[26] , \wRegInB1[25] , \wRegInB1[24] , 
        \wRegInB1[23] , \wRegInB1[22] , \wRegInB1[21] , \wRegInB1[20] , 
        \wRegInB1[19] , \wRegInB1[18] , \wRegInB1[17] , \wRegInB1[16] , 
        \wRegInB1[15] , \wRegInB1[14] , \wRegInB1[13] , \wRegInB1[12] , 
        \wRegInB1[11] , \wRegInB1[10] , \wRegInB1[9] , \wRegInB1[8] , 
        \wRegInB1[7] , \wRegInB1[6] , \wRegInB1[5] , \wRegInB1[4] , 
        \wRegInB1[3] , \wRegInB1[2] , \wRegInB1[1] , \wRegInB1[0] }), .LoOut({
        \wRegInA2[31] , \wRegInA2[30] , \wRegInA2[29] , \wRegInA2[28] , 
        \wRegInA2[27] , \wRegInA2[26] , \wRegInA2[25] , \wRegInA2[24] , 
        \wRegInA2[23] , \wRegInA2[22] , \wRegInA2[21] , \wRegInA2[20] , 
        \wRegInA2[19] , \wRegInA2[18] , \wRegInA2[17] , \wRegInA2[16] , 
        \wRegInA2[15] , \wRegInA2[14] , \wRegInA2[13] , \wRegInA2[12] , 
        \wRegInA2[11] , \wRegInA2[10] , \wRegInA2[9] , \wRegInA2[8] , 
        \wRegInA2[7] , \wRegInA2[6] , \wRegInA2[5] , \wRegInA2[4] , 
        \wRegInA2[3] , \wRegInA2[2] , \wRegInA2[1] , \wRegInA2[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid17[31] , \wAMid17[30] , \wAMid17[29] , \wAMid17[28] , 
        \wAMid17[27] , \wAMid17[26] , \wAMid17[25] , \wAMid17[24] , 
        \wAMid17[23] , \wAMid17[22] , \wAMid17[21] , \wAMid17[20] , 
        \wAMid17[19] , \wAMid17[18] , \wAMid17[17] , \wAMid17[16] , 
        \wAMid17[15] , \wAMid17[14] , \wAMid17[13] , \wAMid17[12] , 
        \wAMid17[11] , \wAMid17[10] , \wAMid17[9] , \wAMid17[8] , \wAMid17[7] , 
        \wAMid17[6] , \wAMid17[5] , \wAMid17[4] , \wAMid17[3] , \wAMid17[2] , 
        \wAMid17[1] , \wAMid17[0] }), .BIn({\wBMid17[31] , \wBMid17[30] , 
        \wBMid17[29] , \wBMid17[28] , \wBMid17[27] , \wBMid17[26] , 
        \wBMid17[25] , \wBMid17[24] , \wBMid17[23] , \wBMid17[22] , 
        \wBMid17[21] , \wBMid17[20] , \wBMid17[19] , \wBMid17[18] , 
        \wBMid17[17] , \wBMid17[16] , \wBMid17[15] , \wBMid17[14] , 
        \wBMid17[13] , \wBMid17[12] , \wBMid17[11] , \wBMid17[10] , 
        \wBMid17[9] , \wBMid17[8] , \wBMid17[7] , \wBMid17[6] , \wBMid17[5] , 
        \wBMid17[4] , \wBMid17[3] , \wBMid17[2] , \wBMid17[1] , \wBMid17[0] }), 
        .HiOut({\wRegInB17[31] , \wRegInB17[30] , \wRegInB17[29] , 
        \wRegInB17[28] , \wRegInB17[27] , \wRegInB17[26] , \wRegInB17[25] , 
        \wRegInB17[24] , \wRegInB17[23] , \wRegInB17[22] , \wRegInB17[21] , 
        \wRegInB17[20] , \wRegInB17[19] , \wRegInB17[18] , \wRegInB17[17] , 
        \wRegInB17[16] , \wRegInB17[15] , \wRegInB17[14] , \wRegInB17[13] , 
        \wRegInB17[12] , \wRegInB17[11] , \wRegInB17[10] , \wRegInB17[9] , 
        \wRegInB17[8] , \wRegInB17[7] , \wRegInB17[6] , \wRegInB17[5] , 
        \wRegInB17[4] , \wRegInB17[3] , \wRegInB17[2] , \wRegInB17[1] , 
        \wRegInB17[0] }), .LoOut({\wRegInA18[31] , \wRegInA18[30] , 
        \wRegInA18[29] , \wRegInA18[28] , \wRegInA18[27] , \wRegInA18[26] , 
        \wRegInA18[25] , \wRegInA18[24] , \wRegInA18[23] , \wRegInA18[22] , 
        \wRegInA18[21] , \wRegInA18[20] , \wRegInA18[19] , \wRegInA18[18] , 
        \wRegInA18[17] , \wRegInA18[16] , \wRegInA18[15] , \wRegInA18[14] , 
        \wRegInA18[13] , \wRegInA18[12] , \wRegInA18[11] , \wRegInA18[10] , 
        \wRegInA18[9] , \wRegInA18[8] , \wRegInA18[7] , \wRegInA18[6] , 
        \wRegInA18[5] , \wRegInA18[4] , \wRegInA18[3] , \wRegInA18[2] , 
        \wRegInA18[1] , \wRegInA18[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid30[31] , \wAMid30[30] , \wAMid30[29] , \wAMid30[28] , 
        \wAMid30[27] , \wAMid30[26] , \wAMid30[25] , \wAMid30[24] , 
        \wAMid30[23] , \wAMid30[22] , \wAMid30[21] , \wAMid30[20] , 
        \wAMid30[19] , \wAMid30[18] , \wAMid30[17] , \wAMid30[16] , 
        \wAMid30[15] , \wAMid30[14] , \wAMid30[13] , \wAMid30[12] , 
        \wAMid30[11] , \wAMid30[10] , \wAMid30[9] , \wAMid30[8] , \wAMid30[7] , 
        \wAMid30[6] , \wAMid30[5] , \wAMid30[4] , \wAMid30[3] , \wAMid30[2] , 
        \wAMid30[1] , \wAMid30[0] }), .BIn({\wBMid30[31] , \wBMid30[30] , 
        \wBMid30[29] , \wBMid30[28] , \wBMid30[27] , \wBMid30[26] , 
        \wBMid30[25] , \wBMid30[24] , \wBMid30[23] , \wBMid30[22] , 
        \wBMid30[21] , \wBMid30[20] , \wBMid30[19] , \wBMid30[18] , 
        \wBMid30[17] , \wBMid30[16] , \wBMid30[15] , \wBMid30[14] , 
        \wBMid30[13] , \wBMid30[12] , \wBMid30[11] , \wBMid30[10] , 
        \wBMid30[9] , \wBMid30[8] , \wBMid30[7] , \wBMid30[6] , \wBMid30[5] , 
        \wBMid30[4] , \wBMid30[3] , \wBMid30[2] , \wBMid30[1] , \wBMid30[0] }), 
        .HiOut({\wRegInB30[31] , \wRegInB30[30] , \wRegInB30[29] , 
        \wRegInB30[28] , \wRegInB30[27] , \wRegInB30[26] , \wRegInB30[25] , 
        \wRegInB30[24] , \wRegInB30[23] , \wRegInB30[22] , \wRegInB30[21] , 
        \wRegInB30[20] , \wRegInB30[19] , \wRegInB30[18] , \wRegInB30[17] , 
        \wRegInB30[16] , \wRegInB30[15] , \wRegInB30[14] , \wRegInB30[13] , 
        \wRegInB30[12] , \wRegInB30[11] , \wRegInB30[10] , \wRegInB30[9] , 
        \wRegInB30[8] , \wRegInB30[7] , \wRegInB30[6] , \wRegInB30[5] , 
        \wRegInB30[4] , \wRegInB30[3] , \wRegInB30[2] , \wRegInB30[1] , 
        \wRegInB30[0] }), .LoOut({\wRegInA31[31] , \wRegInA31[30] , 
        \wRegInA31[29] , \wRegInA31[28] , \wRegInA31[27] , \wRegInA31[26] , 
        \wRegInA31[25] , \wRegInA31[24] , \wRegInA31[23] , \wRegInA31[22] , 
        \wRegInA31[21] , \wRegInA31[20] , \wRegInA31[19] , \wRegInA31[18] , 
        \wRegInA31[17] , \wRegInA31[16] , \wRegInA31[15] , \wRegInA31[14] , 
        \wRegInA31[13] , \wRegInA31[12] , \wRegInA31[11] , \wRegInA31[10] , 
        \wRegInA31[9] , \wRegInA31[8] , \wRegInA31[7] , \wRegInA31[6] , 
        \wRegInA31[5] , \wRegInA31[4] , \wRegInA31[3] , \wRegInA31[2] , 
        \wRegInA31[1] , \wRegInA31[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_55 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink56[31] , \ScanLink56[30] , \ScanLink56[29] , 
        \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , \ScanLink56[25] , 
        \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , \ScanLink56[21] , 
        \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , \ScanLink56[17] , 
        \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , \ScanLink56[13] , 
        \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , \ScanLink56[9] , 
        \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , \ScanLink56[5] , 
        \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , \ScanLink56[1] , 
        \ScanLink56[0] }), .ScanOut({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA4[31] , \wRegInA4[30] , 
        \wRegInA4[29] , \wRegInA4[28] , \wRegInA4[27] , \wRegInA4[26] , 
        \wRegInA4[25] , \wRegInA4[24] , \wRegInA4[23] , \wRegInA4[22] , 
        \wRegInA4[21] , \wRegInA4[20] , \wRegInA4[19] , \wRegInA4[18] , 
        \wRegInA4[17] , \wRegInA4[16] , \wRegInA4[15] , \wRegInA4[14] , 
        \wRegInA4[13] , \wRegInA4[12] , \wRegInA4[11] , \wRegInA4[10] , 
        \wRegInA4[9] , \wRegInA4[8] , \wRegInA4[7] , \wRegInA4[6] , 
        \wRegInA4[5] , \wRegInA4[4] , \wRegInA4[3] , \wRegInA4[2] , 
        \wRegInA4[1] , \wRegInA4[0] }), .Out({\wAIn4[31] , \wAIn4[30] , 
        \wAIn4[29] , \wAIn4[28] , \wAIn4[27] , \wAIn4[26] , \wAIn4[25] , 
        \wAIn4[24] , \wAIn4[23] , \wAIn4[22] , \wAIn4[21] , \wAIn4[20] , 
        \wAIn4[19] , \wAIn4[18] , \wAIn4[17] , \wAIn4[16] , \wAIn4[15] , 
        \wAIn4[14] , \wAIn4[13] , \wAIn4[12] , \wAIn4[11] , \wAIn4[10] , 
        \wAIn4[9] , \wAIn4[8] , \wAIn4[7] , \wAIn4[6] , \wAIn4[5] , \wAIn4[4] , 
        \wAIn4[3] , \wAIn4[2] , \wAIn4[1] , \wAIn4[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_20 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink21[31] , \ScanLink21[30] , \ScanLink21[29] , 
        \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , \ScanLink21[25] , 
        \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , \ScanLink21[21] , 
        \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , \ScanLink21[17] , 
        \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , \ScanLink21[13] , 
        \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , \ScanLink21[9] , 
        \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , \ScanLink21[5] , 
        \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , \ScanLink21[1] , 
        \ScanLink21[0] }), .ScanOut({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB21[31] , \wRegInB21[30] , 
        \wRegInB21[29] , \wRegInB21[28] , \wRegInB21[27] , \wRegInB21[26] , 
        \wRegInB21[25] , \wRegInB21[24] , \wRegInB21[23] , \wRegInB21[22] , 
        \wRegInB21[21] , \wRegInB21[20] , \wRegInB21[19] , \wRegInB21[18] , 
        \wRegInB21[17] , \wRegInB21[16] , \wRegInB21[15] , \wRegInB21[14] , 
        \wRegInB21[13] , \wRegInB21[12] , \wRegInB21[11] , \wRegInB21[10] , 
        \wRegInB21[9] , \wRegInB21[8] , \wRegInB21[7] , \wRegInB21[6] , 
        \wRegInB21[5] , \wRegInB21[4] , \wRegInB21[3] , \wRegInB21[2] , 
        \wRegInB21[1] , \wRegInB21[0] }), .Out({\wBIn21[31] , \wBIn21[30] , 
        \wBIn21[29] , \wBIn21[28] , \wBIn21[27] , \wBIn21[26] , \wBIn21[25] , 
        \wBIn21[24] , \wBIn21[23] , \wBIn21[22] , \wBIn21[21] , \wBIn21[20] , 
        \wBIn21[19] , \wBIn21[18] , \wBIn21[17] , \wBIn21[16] , \wBIn21[15] , 
        \wBIn21[14] , \wBIn21[13] , \wBIn21[12] , \wBIn21[11] , \wBIn21[10] , 
        \wBIn21[9] , \wBIn21[8] , \wBIn21[7] , \wBIn21[6] , \wBIn21[5] , 
        \wBIn21[4] , \wBIn21[3] , \wBIn21[2] , \wBIn21[1] , \wBIn21[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid6[31] , 
        \wAMid6[30] , \wAMid6[29] , \wAMid6[28] , \wAMid6[27] , \wAMid6[26] , 
        \wAMid6[25] , \wAMid6[24] , \wAMid6[23] , \wAMid6[22] , \wAMid6[21] , 
        \wAMid6[20] , \wAMid6[19] , \wAMid6[18] , \wAMid6[17] , \wAMid6[16] , 
        \wAMid6[15] , \wAMid6[14] , \wAMid6[13] , \wAMid6[12] , \wAMid6[11] , 
        \wAMid6[10] , \wAMid6[9] , \wAMid6[8] , \wAMid6[7] , \wAMid6[6] , 
        \wAMid6[5] , \wAMid6[4] , \wAMid6[3] , \wAMid6[2] , \wAMid6[1] , 
        \wAMid6[0] }), .BIn({\wBMid6[31] , \wBMid6[30] , \wBMid6[29] , 
        \wBMid6[28] , \wBMid6[27] , \wBMid6[26] , \wBMid6[25] , \wBMid6[24] , 
        \wBMid6[23] , \wBMid6[22] , \wBMid6[21] , \wBMid6[20] , \wBMid6[19] , 
        \wBMid6[18] , \wBMid6[17] , \wBMid6[16] , \wBMid6[15] , \wBMid6[14] , 
        \wBMid6[13] , \wBMid6[12] , \wBMid6[11] , \wBMid6[10] , \wBMid6[9] , 
        \wBMid6[8] , \wBMid6[7] , \wBMid6[6] , \wBMid6[5] , \wBMid6[4] , 
        \wBMid6[3] , \wBMid6[2] , \wBMid6[1] , \wBMid6[0] }), .HiOut({
        \wRegInB6[31] , \wRegInB6[30] , \wRegInB6[29] , \wRegInB6[28] , 
        \wRegInB6[27] , \wRegInB6[26] , \wRegInB6[25] , \wRegInB6[24] , 
        \wRegInB6[23] , \wRegInB6[22] , \wRegInB6[21] , \wRegInB6[20] , 
        \wRegInB6[19] , \wRegInB6[18] , \wRegInB6[17] , \wRegInB6[16] , 
        \wRegInB6[15] , \wRegInB6[14] , \wRegInB6[13] , \wRegInB6[12] , 
        \wRegInB6[11] , \wRegInB6[10] , \wRegInB6[9] , \wRegInB6[8] , 
        \wRegInB6[7] , \wRegInB6[6] , \wRegInB6[5] , \wRegInB6[4] , 
        \wRegInB6[3] , \wRegInB6[2] , \wRegInB6[1] , \wRegInB6[0] }), .LoOut({
        \wRegInA7[31] , \wRegInA7[30] , \wRegInA7[29] , \wRegInA7[28] , 
        \wRegInA7[27] , \wRegInA7[26] , \wRegInA7[25] , \wRegInA7[24] , 
        \wRegInA7[23] , \wRegInA7[22] , \wRegInA7[21] , \wRegInA7[20] , 
        \wRegInA7[19] , \wRegInA7[18] , \wRegInA7[17] , \wRegInA7[16] , 
        \wRegInA7[15] , \wRegInA7[14] , \wRegInA7[13] , \wRegInA7[12] , 
        \wRegInA7[11] , \wRegInA7[10] , \wRegInA7[9] , \wRegInA7[8] , 
        \wRegInA7[7] , \wRegInA7[6] , \wRegInA7[5] , \wRegInA7[4] , 
        \wRegInA7[3] , \wRegInA7[2] , \wRegInA7[1] , \wRegInA7[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid10[31] , \wAMid10[30] , \wAMid10[29] , \wAMid10[28] , 
        \wAMid10[27] , \wAMid10[26] , \wAMid10[25] , \wAMid10[24] , 
        \wAMid10[23] , \wAMid10[22] , \wAMid10[21] , \wAMid10[20] , 
        \wAMid10[19] , \wAMid10[18] , \wAMid10[17] , \wAMid10[16] , 
        \wAMid10[15] , \wAMid10[14] , \wAMid10[13] , \wAMid10[12] , 
        \wAMid10[11] , \wAMid10[10] , \wAMid10[9] , \wAMid10[8] , \wAMid10[7] , 
        \wAMid10[6] , \wAMid10[5] , \wAMid10[4] , \wAMid10[3] , \wAMid10[2] , 
        \wAMid10[1] , \wAMid10[0] }), .BIn({\wBMid10[31] , \wBMid10[30] , 
        \wBMid10[29] , \wBMid10[28] , \wBMid10[27] , \wBMid10[26] , 
        \wBMid10[25] , \wBMid10[24] , \wBMid10[23] , \wBMid10[22] , 
        \wBMid10[21] , \wBMid10[20] , \wBMid10[19] , \wBMid10[18] , 
        \wBMid10[17] , \wBMid10[16] , \wBMid10[15] , \wBMid10[14] , 
        \wBMid10[13] , \wBMid10[12] , \wBMid10[11] , \wBMid10[10] , 
        \wBMid10[9] , \wBMid10[8] , \wBMid10[7] , \wBMid10[6] , \wBMid10[5] , 
        \wBMid10[4] , \wBMid10[3] , \wBMid10[2] , \wBMid10[1] , \wBMid10[0] }), 
        .HiOut({\wRegInB10[31] , \wRegInB10[30] , \wRegInB10[29] , 
        \wRegInB10[28] , \wRegInB10[27] , \wRegInB10[26] , \wRegInB10[25] , 
        \wRegInB10[24] , \wRegInB10[23] , \wRegInB10[22] , \wRegInB10[21] , 
        \wRegInB10[20] , \wRegInB10[19] , \wRegInB10[18] , \wRegInB10[17] , 
        \wRegInB10[16] , \wRegInB10[15] , \wRegInB10[14] , \wRegInB10[13] , 
        \wRegInB10[12] , \wRegInB10[11] , \wRegInB10[10] , \wRegInB10[9] , 
        \wRegInB10[8] , \wRegInB10[7] , \wRegInB10[6] , \wRegInB10[5] , 
        \wRegInB10[4] , \wRegInB10[3] , \wRegInB10[2] , \wRegInB10[1] , 
        \wRegInB10[0] }), .LoOut({\wRegInA11[31] , \wRegInA11[30] , 
        \wRegInA11[29] , \wRegInA11[28] , \wRegInA11[27] , \wRegInA11[26] , 
        \wRegInA11[25] , \wRegInA11[24] , \wRegInA11[23] , \wRegInA11[22] , 
        \wRegInA11[21] , \wRegInA11[20] , \wRegInA11[19] , \wRegInA11[18] , 
        \wRegInA11[17] , \wRegInA11[16] , \wRegInA11[15] , \wRegInA11[14] , 
        \wRegInA11[13] , \wRegInA11[12] , \wRegInA11[11] , \wRegInA11[10] , 
        \wRegInA11[9] , \wRegInA11[8] , \wRegInA11[7] , \wRegInA11[6] , 
        \wRegInA11[5] , \wRegInA11[4] , \wRegInA11[3] , \wRegInA11[2] , 
        \wRegInA11[1] , \wRegInA11[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_52 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink53[31] , \ScanLink53[30] , \ScanLink53[29] , 
        \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , \ScanLink53[25] , 
        \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , \ScanLink53[21] , 
        \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , \ScanLink53[17] , 
        \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , \ScanLink53[13] , 
        \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , \ScanLink53[9] , 
        \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , \ScanLink53[5] , 
        \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , \ScanLink53[1] , 
        \ScanLink53[0] }), .ScanOut({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB5[31] , \wRegInB5[30] , 
        \wRegInB5[29] , \wRegInB5[28] , \wRegInB5[27] , \wRegInB5[26] , 
        \wRegInB5[25] , \wRegInB5[24] , \wRegInB5[23] , \wRegInB5[22] , 
        \wRegInB5[21] , \wRegInB5[20] , \wRegInB5[19] , \wRegInB5[18] , 
        \wRegInB5[17] , \wRegInB5[16] , \wRegInB5[15] , \wRegInB5[14] , 
        \wRegInB5[13] , \wRegInB5[12] , \wRegInB5[11] , \wRegInB5[10] , 
        \wRegInB5[9] , \wRegInB5[8] , \wRegInB5[7] , \wRegInB5[6] , 
        \wRegInB5[5] , \wRegInB5[4] , \wRegInB5[3] , \wRegInB5[2] , 
        \wRegInB5[1] , \wRegInB5[0] }), .Out({\wBIn5[31] , \wBIn5[30] , 
        \wBIn5[29] , \wBIn5[28] , \wBIn5[27] , \wBIn5[26] , \wBIn5[25] , 
        \wBIn5[24] , \wBIn5[23] , \wBIn5[22] , \wBIn5[21] , \wBIn5[20] , 
        \wBIn5[19] , \wBIn5[18] , \wBIn5[17] , \wBIn5[16] , \wBIn5[15] , 
        \wBIn5[14] , \wBIn5[13] , \wBIn5[12] , \wBIn5[11] , \wBIn5[10] , 
        \wBIn5[9] , \wBIn5[8] , \wBIn5[7] , \wBIn5[6] , \wBIn5[5] , \wBIn5[4] , 
        \wBIn5[3] , \wBIn5[2] , \wBIn5[1] , \wBIn5[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_49 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink50[31] , \ScanLink50[30] , \ScanLink50[29] , 
        \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , \ScanLink50[25] , 
        \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , \ScanLink50[21] , 
        \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , \ScanLink50[17] , 
        \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , \ScanLink50[13] , 
        \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , \ScanLink50[9] , 
        \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , \ScanLink50[5] , 
        \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , \ScanLink50[1] , 
        \ScanLink50[0] }), .ScanOut({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA7[31] , \wRegInA7[30] , 
        \wRegInA7[29] , \wRegInA7[28] , \wRegInA7[27] , \wRegInA7[26] , 
        \wRegInA7[25] , \wRegInA7[24] , \wRegInA7[23] , \wRegInA7[22] , 
        \wRegInA7[21] , \wRegInA7[20] , \wRegInA7[19] , \wRegInA7[18] , 
        \wRegInA7[17] , \wRegInA7[16] , \wRegInA7[15] , \wRegInA7[14] , 
        \wRegInA7[13] , \wRegInA7[12] , \wRegInA7[11] , \wRegInA7[10] , 
        \wRegInA7[9] , \wRegInA7[8] , \wRegInA7[7] , \wRegInA7[6] , 
        \wRegInA7[5] , \wRegInA7[4] , \wRegInA7[3] , \wRegInA7[2] , 
        \wRegInA7[1] , \wRegInA7[0] }), .Out({\wAIn7[31] , \wAIn7[30] , 
        \wAIn7[29] , \wAIn7[28] , \wAIn7[27] , \wAIn7[26] , \wAIn7[25] , 
        \wAIn7[24] , \wAIn7[23] , \wAIn7[22] , \wAIn7[21] , \wAIn7[20] , 
        \wAIn7[19] , \wAIn7[18] , \wAIn7[17] , \wAIn7[16] , \wAIn7[15] , 
        \wAIn7[14] , \wAIn7[13] , \wAIn7[12] , \wAIn7[11] , \wAIn7[10] , 
        \wAIn7[9] , \wAIn7[8] , \wAIn7[7] , \wAIn7[6] , \wAIn7[5] , \wAIn7[4] , 
        \wAIn7[3] , \wAIn7[2] , \wAIn7[1] , \wAIn7[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_27 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink28[31] , \ScanLink28[30] , \ScanLink28[29] , 
        \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , \ScanLink28[25] , 
        \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , \ScanLink28[21] , 
        \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , \ScanLink28[17] , 
        \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , \ScanLink28[13] , 
        \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , \ScanLink28[9] , 
        \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , \ScanLink28[5] , 
        \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , \ScanLink28[1] , 
        \ScanLink28[0] }), .ScanOut({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA18[31] , \wRegInA18[30] , 
        \wRegInA18[29] , \wRegInA18[28] , \wRegInA18[27] , \wRegInA18[26] , 
        \wRegInA18[25] , \wRegInA18[24] , \wRegInA18[23] , \wRegInA18[22] , 
        \wRegInA18[21] , \wRegInA18[20] , \wRegInA18[19] , \wRegInA18[18] , 
        \wRegInA18[17] , \wRegInA18[16] , \wRegInA18[15] , \wRegInA18[14] , 
        \wRegInA18[13] , \wRegInA18[12] , \wRegInA18[11] , \wRegInA18[10] , 
        \wRegInA18[9] , \wRegInA18[8] , \wRegInA18[7] , \wRegInA18[6] , 
        \wRegInA18[5] , \wRegInA18[4] , \wRegInA18[3] , \wRegInA18[2] , 
        \wRegInA18[1] , \wRegInA18[0] }), .Out({\wAIn18[31] , \wAIn18[30] , 
        \wAIn18[29] , \wAIn18[28] , \wAIn18[27] , \wAIn18[26] , \wAIn18[25] , 
        \wAIn18[24] , \wAIn18[23] , \wAIn18[22] , \wAIn18[21] , \wAIn18[20] , 
        \wAIn18[19] , \wAIn18[18] , \wAIn18[17] , \wAIn18[16] , \wAIn18[15] , 
        \wAIn18[14] , \wAIn18[13] , \wAIn18[12] , \wAIn18[11] , \wAIn18[10] , 
        \wAIn18[9] , \wAIn18[8] , \wAIn18[7] , \wAIn18[6] , \wAIn18[5] , 
        \wAIn18[4] , \wAIn18[3] , \wAIn18[2] , \wAIn18[1] , \wAIn18[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid25[31] , \wAMid25[30] , \wAMid25[29] , \wAMid25[28] , 
        \wAMid25[27] , \wAMid25[26] , \wAMid25[25] , \wAMid25[24] , 
        \wAMid25[23] , \wAMid25[22] , \wAMid25[21] , \wAMid25[20] , 
        \wAMid25[19] , \wAMid25[18] , \wAMid25[17] , \wAMid25[16] , 
        \wAMid25[15] , \wAMid25[14] , \wAMid25[13] , \wAMid25[12] , 
        \wAMid25[11] , \wAMid25[10] , \wAMid25[9] , \wAMid25[8] , \wAMid25[7] , 
        \wAMid25[6] , \wAMid25[5] , \wAMid25[4] , \wAMid25[3] , \wAMid25[2] , 
        \wAMid25[1] , \wAMid25[0] }), .BIn({\wBMid25[31] , \wBMid25[30] , 
        \wBMid25[29] , \wBMid25[28] , \wBMid25[27] , \wBMid25[26] , 
        \wBMid25[25] , \wBMid25[24] , \wBMid25[23] , \wBMid25[22] , 
        \wBMid25[21] , \wBMid25[20] , \wBMid25[19] , \wBMid25[18] , 
        \wBMid25[17] , \wBMid25[16] , \wBMid25[15] , \wBMid25[14] , 
        \wBMid25[13] , \wBMid25[12] , \wBMid25[11] , \wBMid25[10] , 
        \wBMid25[9] , \wBMid25[8] , \wBMid25[7] , \wBMid25[6] , \wBMid25[5] , 
        \wBMid25[4] , \wBMid25[3] , \wBMid25[2] , \wBMid25[1] , \wBMid25[0] }), 
        .HiOut({\wRegInB25[31] , \wRegInB25[30] , \wRegInB25[29] , 
        \wRegInB25[28] , \wRegInB25[27] , \wRegInB25[26] , \wRegInB25[25] , 
        \wRegInB25[24] , \wRegInB25[23] , \wRegInB25[22] , \wRegInB25[21] , 
        \wRegInB25[20] , \wRegInB25[19] , \wRegInB25[18] , \wRegInB25[17] , 
        \wRegInB25[16] , \wRegInB25[15] , \wRegInB25[14] , \wRegInB25[13] , 
        \wRegInB25[12] , \wRegInB25[11] , \wRegInB25[10] , \wRegInB25[9] , 
        \wRegInB25[8] , \wRegInB25[7] , \wRegInB25[6] , \wRegInB25[5] , 
        \wRegInB25[4] , \wRegInB25[3] , \wRegInB25[2] , \wRegInB25[1] , 
        \wRegInB25[0] }), .LoOut({\wRegInA26[31] , \wRegInA26[30] , 
        \wRegInA26[29] , \wRegInA26[28] , \wRegInA26[27] , \wRegInA26[26] , 
        \wRegInA26[25] , \wRegInA26[24] , \wRegInA26[23] , \wRegInA26[22] , 
        \wRegInA26[21] , \wRegInA26[20] , \wRegInA26[19] , \wRegInA26[18] , 
        \wRegInA26[17] , \wRegInA26[16] , \wRegInA26[15] , \wRegInA26[14] , 
        \wRegInA26[13] , \wRegInA26[12] , \wRegInA26[11] , \wRegInA26[10] , 
        \wRegInA26[9] , \wRegInA26[8] , \wRegInA26[7] , \wRegInA26[6] , 
        \wRegInA26[5] , \wRegInA26[4] , \wRegInA26[3] , \wRegInA26[2] , 
        \wRegInA26[1] , \wRegInA26[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_40 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink41[31] , \ScanLink41[30] , \ScanLink41[29] , 
        \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , \ScanLink41[25] , 
        \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , \ScanLink41[21] , 
        \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , \ScanLink41[17] , 
        \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , \ScanLink41[13] , 
        \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , \ScanLink41[9] , 
        \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , \ScanLink41[5] , 
        \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , \ScanLink41[1] , 
        \ScanLink41[0] }), .ScanOut({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB11[31] , \wRegInB11[30] , 
        \wRegInB11[29] , \wRegInB11[28] , \wRegInB11[27] , \wRegInB11[26] , 
        \wRegInB11[25] , \wRegInB11[24] , \wRegInB11[23] , \wRegInB11[22] , 
        \wRegInB11[21] , \wRegInB11[20] , \wRegInB11[19] , \wRegInB11[18] , 
        \wRegInB11[17] , \wRegInB11[16] , \wRegInB11[15] , \wRegInB11[14] , 
        \wRegInB11[13] , \wRegInB11[12] , \wRegInB11[11] , \wRegInB11[10] , 
        \wRegInB11[9] , \wRegInB11[8] , \wRegInB11[7] , \wRegInB11[6] , 
        \wRegInB11[5] , \wRegInB11[4] , \wRegInB11[3] , \wRegInB11[2] , 
        \wRegInB11[1] , \wRegInB11[0] }), .Out({\wBIn11[31] , \wBIn11[30] , 
        \wBIn11[29] , \wBIn11[28] , \wBIn11[27] , \wBIn11[26] , \wBIn11[25] , 
        \wBIn11[24] , \wBIn11[23] , \wBIn11[22] , \wBIn11[21] , \wBIn11[20] , 
        \wBIn11[19] , \wBIn11[18] , \wBIn11[17] , \wBIn11[16] , \wBIn11[15] , 
        \wBIn11[14] , \wBIn11[13] , \wBIn11[12] , \wBIn11[11] , \wBIn11[10] , 
        \wBIn11[9] , \wBIn11[8] , \wBIn11[7] , \wBIn11[6] , \wBIn11[5] , 
        \wBIn11[4] , \wBIn11[3] , \wBIn11[2] , \wBIn11[1] , \wBIn11[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn29[31] , \wAIn29[30] , \wAIn29[29] , \wAIn29[28] , \wAIn29[27] , 
        \wAIn29[26] , \wAIn29[25] , \wAIn29[24] , \wAIn29[23] , \wAIn29[22] , 
        \wAIn29[21] , \wAIn29[20] , \wAIn29[19] , \wAIn29[18] , \wAIn29[17] , 
        \wAIn29[16] , \wAIn29[15] , \wAIn29[14] , \wAIn29[13] , \wAIn29[12] , 
        \wAIn29[11] , \wAIn29[10] , \wAIn29[9] , \wAIn29[8] , \wAIn29[7] , 
        \wAIn29[6] , \wAIn29[5] , \wAIn29[4] , \wAIn29[3] , \wAIn29[2] , 
        \wAIn29[1] , \wAIn29[0] }), .BIn({\wBIn29[31] , \wBIn29[30] , 
        \wBIn29[29] , \wBIn29[28] , \wBIn29[27] , \wBIn29[26] , \wBIn29[25] , 
        \wBIn29[24] , \wBIn29[23] , \wBIn29[22] , \wBIn29[21] , \wBIn29[20] , 
        \wBIn29[19] , \wBIn29[18] , \wBIn29[17] , \wBIn29[16] , \wBIn29[15] , 
        \wBIn29[14] , \wBIn29[13] , \wBIn29[12] , \wBIn29[11] , \wBIn29[10] , 
        \wBIn29[9] , \wBIn29[8] , \wBIn29[7] , \wBIn29[6] , \wBIn29[5] , 
        \wBIn29[4] , \wBIn29[3] , \wBIn29[2] , \wBIn29[1] , \wBIn29[0] }), 
        .HiOut({\wBMid28[31] , \wBMid28[30] , \wBMid28[29] , \wBMid28[28] , 
        \wBMid28[27] , \wBMid28[26] , \wBMid28[25] , \wBMid28[24] , 
        \wBMid28[23] , \wBMid28[22] , \wBMid28[21] , \wBMid28[20] , 
        \wBMid28[19] , \wBMid28[18] , \wBMid28[17] , \wBMid28[16] , 
        \wBMid28[15] , \wBMid28[14] , \wBMid28[13] , \wBMid28[12] , 
        \wBMid28[11] , \wBMid28[10] , \wBMid28[9] , \wBMid28[8] , \wBMid28[7] , 
        \wBMid28[6] , \wBMid28[5] , \wBMid28[4] , \wBMid28[3] , \wBMid28[2] , 
        \wBMid28[1] , \wBMid28[0] }), .LoOut({\wAMid29[31] , \wAMid29[30] , 
        \wAMid29[29] , \wAMid29[28] , \wAMid29[27] , \wAMid29[26] , 
        \wAMid29[25] , \wAMid29[24] , \wAMid29[23] , \wAMid29[22] , 
        \wAMid29[21] , \wAMid29[20] , \wAMid29[19] , \wAMid29[18] , 
        \wAMid29[17] , \wAMid29[16] , \wAMid29[15] , \wAMid29[14] , 
        \wAMid29[13] , \wAMid29[12] , \wAMid29[11] , \wAMid29[10] , 
        \wAMid29[9] , \wAMid29[8] , \wAMid29[7] , \wAMid29[6] , \wAMid29[5] , 
        \wAMid29[4] , \wAMid29[3] , \wAMid29[2] , \wAMid29[1] , \wAMid29[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_35 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink36[31] , \ScanLink36[30] , \ScanLink36[29] , 
        \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , \ScanLink36[25] , 
        \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , \ScanLink36[21] , 
        \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , \ScanLink36[17] , 
        \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , \ScanLink36[13] , 
        \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , \ScanLink36[9] , 
        \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , \ScanLink36[5] , 
        \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , \ScanLink36[1] , 
        \ScanLink36[0] }), .ScanOut({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA14[31] , \wRegInA14[30] , 
        \wRegInA14[29] , \wRegInA14[28] , \wRegInA14[27] , \wRegInA14[26] , 
        \wRegInA14[25] , \wRegInA14[24] , \wRegInA14[23] , \wRegInA14[22] , 
        \wRegInA14[21] , \wRegInA14[20] , \wRegInA14[19] , \wRegInA14[18] , 
        \wRegInA14[17] , \wRegInA14[16] , \wRegInA14[15] , \wRegInA14[14] , 
        \wRegInA14[13] , \wRegInA14[12] , \wRegInA14[11] , \wRegInA14[10] , 
        \wRegInA14[9] , \wRegInA14[8] , \wRegInA14[7] , \wRegInA14[6] , 
        \wRegInA14[5] , \wRegInA14[4] , \wRegInA14[3] , \wRegInA14[2] , 
        \wRegInA14[1] , \wRegInA14[0] }), .Out({\wAIn14[31] , \wAIn14[30] , 
        \wAIn14[29] , \wAIn14[28] , \wAIn14[27] , \wAIn14[26] , \wAIn14[25] , 
        \wAIn14[24] , \wAIn14[23] , \wAIn14[22] , \wAIn14[21] , \wAIn14[20] , 
        \wAIn14[19] , \wAIn14[18] , \wAIn14[17] , \wAIn14[16] , \wAIn14[15] , 
        \wAIn14[14] , \wAIn14[13] , \wAIn14[12] , \wAIn14[11] , \wAIn14[10] , 
        \wAIn14[9] , \wAIn14[8] , \wAIn14[7] , \wAIn14[6] , \wAIn14[5] , 
        \wAIn14[4] , \wAIn14[3] , \wAIn14[2] , \wAIn14[1] , \wAIn14[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_3 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[31] , \ScanLink4[30] , \ScanLink4[29] , 
        \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , \ScanLink4[25] , 
        \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , \ScanLink4[21] , 
        \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , \ScanLink4[17] , 
        \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , \ScanLink4[13] , 
        \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , \ScanLink4[9] , 
        \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA30[31] , \wRegInA30[30] , 
        \wRegInA30[29] , \wRegInA30[28] , \wRegInA30[27] , \wRegInA30[26] , 
        \wRegInA30[25] , \wRegInA30[24] , \wRegInA30[23] , \wRegInA30[22] , 
        \wRegInA30[21] , \wRegInA30[20] , \wRegInA30[19] , \wRegInA30[18] , 
        \wRegInA30[17] , \wRegInA30[16] , \wRegInA30[15] , \wRegInA30[14] , 
        \wRegInA30[13] , \wRegInA30[12] , \wRegInA30[11] , \wRegInA30[10] , 
        \wRegInA30[9] , \wRegInA30[8] , \wRegInA30[7] , \wRegInA30[6] , 
        \wRegInA30[5] , \wRegInA30[4] , \wRegInA30[3] , \wRegInA30[2] , 
        \wRegInA30[1] , \wRegInA30[0] }), .Out({\wAIn30[31] , \wAIn30[30] , 
        \wAIn30[29] , \wAIn30[28] , \wAIn30[27] , \wAIn30[26] , \wAIn30[25] , 
        \wAIn30[24] , \wAIn30[23] , \wAIn30[22] , \wAIn30[21] , \wAIn30[20] , 
        \wAIn30[19] , \wAIn30[18] , \wAIn30[17] , \wAIn30[16] , \wAIn30[15] , 
        \wAIn30[14] , \wAIn30[13] , \wAIn30[12] , \wAIn30[11] , \wAIn30[10] , 
        \wAIn30[9] , \wAIn30[8] , \wAIn30[7] , \wAIn30[6] , \wAIn30[5] , 
        \wAIn30[4] , \wAIn30[3] , \wAIn30[2] , \wAIn30[1] , \wAIn30[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_12 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[31] , \ScanLink13[30] , \ScanLink13[29] , 
        \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , \ScanLink13[25] , 
        \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , \ScanLink13[21] , 
        \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , \ScanLink13[17] , 
        \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , \ScanLink13[13] , 
        \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , \ScanLink13[9] , 
        \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB25[31] , \wRegInB25[30] , 
        \wRegInB25[29] , \wRegInB25[28] , \wRegInB25[27] , \wRegInB25[26] , 
        \wRegInB25[25] , \wRegInB25[24] , \wRegInB25[23] , \wRegInB25[22] , 
        \wRegInB25[21] , \wRegInB25[20] , \wRegInB25[19] , \wRegInB25[18] , 
        \wRegInB25[17] , \wRegInB25[16] , \wRegInB25[15] , \wRegInB25[14] , 
        \wRegInB25[13] , \wRegInB25[12] , \wRegInB25[11] , \wRegInB25[10] , 
        \wRegInB25[9] , \wRegInB25[8] , \wRegInB25[7] , \wRegInB25[6] , 
        \wRegInB25[5] , \wRegInB25[4] , \wRegInB25[3] , \wRegInB25[2] , 
        \wRegInB25[1] , \wRegInB25[0] }), .Out({\wBIn25[31] , \wBIn25[30] , 
        \wBIn25[29] , \wBIn25[28] , \wBIn25[27] , \wBIn25[26] , \wBIn25[25] , 
        \wBIn25[24] , \wBIn25[23] , \wBIn25[22] , \wBIn25[21] , \wBIn25[20] , 
        \wBIn25[19] , \wBIn25[18] , \wBIn25[17] , \wBIn25[16] , \wBIn25[15] , 
        \wBIn25[14] , \wBIn25[13] , \wBIn25[12] , \wBIn25[11] , \wBIn25[10] , 
        \wBIn25[9] , \wBIn25[8] , \wBIn25[7] , \wBIn25[6] , \wBIn25[5] , 
        \wBIn25[4] , \wBIn25[3] , \wBIn25[2] , \wBIn25[1] , \wBIn25[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid19[31] , \wAMid19[30] , \wAMid19[29] , \wAMid19[28] , 
        \wAMid19[27] , \wAMid19[26] , \wAMid19[25] , \wAMid19[24] , 
        \wAMid19[23] , \wAMid19[22] , \wAMid19[21] , \wAMid19[20] , 
        \wAMid19[19] , \wAMid19[18] , \wAMid19[17] , \wAMid19[16] , 
        \wAMid19[15] , \wAMid19[14] , \wAMid19[13] , \wAMid19[12] , 
        \wAMid19[11] , \wAMid19[10] , \wAMid19[9] , \wAMid19[8] , \wAMid19[7] , 
        \wAMid19[6] , \wAMid19[5] , \wAMid19[4] , \wAMid19[3] , \wAMid19[2] , 
        \wAMid19[1] , \wAMid19[0] }), .BIn({\wBMid19[31] , \wBMid19[30] , 
        \wBMid19[29] , \wBMid19[28] , \wBMid19[27] , \wBMid19[26] , 
        \wBMid19[25] , \wBMid19[24] , \wBMid19[23] , \wBMid19[22] , 
        \wBMid19[21] , \wBMid19[20] , \wBMid19[19] , \wBMid19[18] , 
        \wBMid19[17] , \wBMid19[16] , \wBMid19[15] , \wBMid19[14] , 
        \wBMid19[13] , \wBMid19[12] , \wBMid19[11] , \wBMid19[10] , 
        \wBMid19[9] , \wBMid19[8] , \wBMid19[7] , \wBMid19[6] , \wBMid19[5] , 
        \wBMid19[4] , \wBMid19[3] , \wBMid19[2] , \wBMid19[1] , \wBMid19[0] }), 
        .HiOut({\wRegInB19[31] , \wRegInB19[30] , \wRegInB19[29] , 
        \wRegInB19[28] , \wRegInB19[27] , \wRegInB19[26] , \wRegInB19[25] , 
        \wRegInB19[24] , \wRegInB19[23] , \wRegInB19[22] , \wRegInB19[21] , 
        \wRegInB19[20] , \wRegInB19[19] , \wRegInB19[18] , \wRegInB19[17] , 
        \wRegInB19[16] , \wRegInB19[15] , \wRegInB19[14] , \wRegInB19[13] , 
        \wRegInB19[12] , \wRegInB19[11] , \wRegInB19[10] , \wRegInB19[9] , 
        \wRegInB19[8] , \wRegInB19[7] , \wRegInB19[6] , \wRegInB19[5] , 
        \wRegInB19[4] , \wRegInB19[3] , \wRegInB19[2] , \wRegInB19[1] , 
        \wRegInB19[0] }), .LoOut({\wRegInA20[31] , \wRegInA20[30] , 
        \wRegInA20[29] , \wRegInA20[28] , \wRegInA20[27] , \wRegInA20[26] , 
        \wRegInA20[25] , \wRegInA20[24] , \wRegInA20[23] , \wRegInA20[22] , 
        \wRegInA20[21] , \wRegInA20[20] , \wRegInA20[19] , \wRegInA20[18] , 
        \wRegInA20[17] , \wRegInA20[16] , \wRegInA20[15] , \wRegInA20[14] , 
        \wRegInA20[13] , \wRegInA20[12] , \wRegInA20[11] , \wRegInA20[10] , 
        \wRegInA20[9] , \wRegInA20[8] , \wRegInA20[7] , \wRegInA20[6] , 
        \wRegInA20[5] , \wRegInA20[4] , \wRegInA20[3] , \wRegInA20[2] , 
        \wRegInA20[1] , \wRegInA20[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn21[31] , \wAIn21[30] , \wAIn21[29] , \wAIn21[28] , \wAIn21[27] , 
        \wAIn21[26] , \wAIn21[25] , \wAIn21[24] , \wAIn21[23] , \wAIn21[22] , 
        \wAIn21[21] , \wAIn21[20] , \wAIn21[19] , \wAIn21[18] , \wAIn21[17] , 
        \wAIn21[16] , \wAIn21[15] , \wAIn21[14] , \wAIn21[13] , \wAIn21[12] , 
        \wAIn21[11] , \wAIn21[10] , \wAIn21[9] , \wAIn21[8] , \wAIn21[7] , 
        \wAIn21[6] , \wAIn21[5] , \wAIn21[4] , \wAIn21[3] , \wAIn21[2] , 
        \wAIn21[1] , \wAIn21[0] }), .BIn({\wBIn21[31] , \wBIn21[30] , 
        \wBIn21[29] , \wBIn21[28] , \wBIn21[27] , \wBIn21[26] , \wBIn21[25] , 
        \wBIn21[24] , \wBIn21[23] , \wBIn21[22] , \wBIn21[21] , \wBIn21[20] , 
        \wBIn21[19] , \wBIn21[18] , \wBIn21[17] , \wBIn21[16] , \wBIn21[15] , 
        \wBIn21[14] , \wBIn21[13] , \wBIn21[12] , \wBIn21[11] , \wBIn21[10] , 
        \wBIn21[9] , \wBIn21[8] , \wBIn21[7] , \wBIn21[6] , \wBIn21[5] , 
        \wBIn21[4] , \wBIn21[3] , \wBIn21[2] , \wBIn21[1] , \wBIn21[0] }), 
        .HiOut({\wBMid20[31] , \wBMid20[30] , \wBMid20[29] , \wBMid20[28] , 
        \wBMid20[27] , \wBMid20[26] , \wBMid20[25] , \wBMid20[24] , 
        \wBMid20[23] , \wBMid20[22] , \wBMid20[21] , \wBMid20[20] , 
        \wBMid20[19] , \wBMid20[18] , \wBMid20[17] , \wBMid20[16] , 
        \wBMid20[15] , \wBMid20[14] , \wBMid20[13] , \wBMid20[12] , 
        \wBMid20[11] , \wBMid20[10] , \wBMid20[9] , \wBMid20[8] , \wBMid20[7] , 
        \wBMid20[6] , \wBMid20[5] , \wBMid20[4] , \wBMid20[3] , \wBMid20[2] , 
        \wBMid20[1] , \wBMid20[0] }), .LoOut({\wAMid21[31] , \wAMid21[30] , 
        \wAMid21[29] , \wAMid21[28] , \wAMid21[27] , \wAMid21[26] , 
        \wAMid21[25] , \wAMid21[24] , \wAMid21[23] , \wAMid21[22] , 
        \wAMid21[21] , \wAMid21[20] , \wAMid21[19] , \wAMid21[18] , 
        \wAMid21[17] , \wAMid21[16] , \wAMid21[15] , \wAMid21[14] , 
        \wAMid21[13] , \wAMid21[12] , \wAMid21[11] , \wAMid21[10] , 
        \wAMid21[9] , \wAMid21[8] , \wAMid21[7] , \wAMid21[6] , \wAMid21[5] , 
        \wAMid21[4] , \wAMid21[3] , \wAMid21[2] , \wAMid21[1] , \wAMid21[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_53 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink54[31] , \ScanLink54[30] , \ScanLink54[29] , 
        \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , \ScanLink54[25] , 
        \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , \ScanLink54[21] , 
        \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , \ScanLink54[17] , 
        \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , \ScanLink54[13] , 
        \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , \ScanLink54[9] , 
        \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , \ScanLink54[5] , 
        \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , \ScanLink54[1] , 
        \ScanLink54[0] }), .ScanOut({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA5[31] , \wRegInA5[30] , 
        \wRegInA5[29] , \wRegInA5[28] , \wRegInA5[27] , \wRegInA5[26] , 
        \wRegInA5[25] , \wRegInA5[24] , \wRegInA5[23] , \wRegInA5[22] , 
        \wRegInA5[21] , \wRegInA5[20] , \wRegInA5[19] , \wRegInA5[18] , 
        \wRegInA5[17] , \wRegInA5[16] , \wRegInA5[15] , \wRegInA5[14] , 
        \wRegInA5[13] , \wRegInA5[12] , \wRegInA5[11] , \wRegInA5[10] , 
        \wRegInA5[9] , \wRegInA5[8] , \wRegInA5[7] , \wRegInA5[6] , 
        \wRegInA5[5] , \wRegInA5[4] , \wRegInA5[3] , \wRegInA5[2] , 
        \wRegInA5[1] , \wRegInA5[0] }), .Out({\wAIn5[31] , \wAIn5[30] , 
        \wAIn5[29] , \wAIn5[28] , \wAIn5[27] , \wAIn5[26] , \wAIn5[25] , 
        \wAIn5[24] , \wAIn5[23] , \wAIn5[22] , \wAIn5[21] , \wAIn5[20] , 
        \wAIn5[19] , \wAIn5[18] , \wAIn5[17] , \wAIn5[16] , \wAIn5[15] , 
        \wAIn5[14] , \wAIn5[13] , \wAIn5[12] , \wAIn5[11] , \wAIn5[10] , 
        \wAIn5[9] , \wAIn5[8] , \wAIn5[7] , \wAIn5[6] , \wAIn5[5] , \wAIn5[4] , 
        \wAIn5[3] , \wAIn5[2] , \wAIn5[1] , \wAIn5[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn28[31] , \wAIn28[30] , \wAIn28[29] , \wAIn28[28] , \wAIn28[27] , 
        \wAIn28[26] , \wAIn28[25] , \wAIn28[24] , \wAIn28[23] , \wAIn28[22] , 
        \wAIn28[21] , \wAIn28[20] , \wAIn28[19] , \wAIn28[18] , \wAIn28[17] , 
        \wAIn28[16] , \wAIn28[15] , \wAIn28[14] , \wAIn28[13] , \wAIn28[12] , 
        \wAIn28[11] , \wAIn28[10] , \wAIn28[9] , \wAIn28[8] , \wAIn28[7] , 
        \wAIn28[6] , \wAIn28[5] , \wAIn28[4] , \wAIn28[3] , \wAIn28[2] , 
        \wAIn28[1] , \wAIn28[0] }), .BIn({\wBIn28[31] , \wBIn28[30] , 
        \wBIn28[29] , \wBIn28[28] , \wBIn28[27] , \wBIn28[26] , \wBIn28[25] , 
        \wBIn28[24] , \wBIn28[23] , \wBIn28[22] , \wBIn28[21] , \wBIn28[20] , 
        \wBIn28[19] , \wBIn28[18] , \wBIn28[17] , \wBIn28[16] , \wBIn28[15] , 
        \wBIn28[14] , \wBIn28[13] , \wBIn28[12] , \wBIn28[11] , \wBIn28[10] , 
        \wBIn28[9] , \wBIn28[8] , \wBIn28[7] , \wBIn28[6] , \wBIn28[5] , 
        \wBIn28[4] , \wBIn28[3] , \wBIn28[2] , \wBIn28[1] , \wBIn28[0] }), 
        .HiOut({\wBMid27[31] , \wBMid27[30] , \wBMid27[29] , \wBMid27[28] , 
        \wBMid27[27] , \wBMid27[26] , \wBMid27[25] , \wBMid27[24] , 
        \wBMid27[23] , \wBMid27[22] , \wBMid27[21] , \wBMid27[20] , 
        \wBMid27[19] , \wBMid27[18] , \wBMid27[17] , \wBMid27[16] , 
        \wBMid27[15] , \wBMid27[14] , \wBMid27[13] , \wBMid27[12] , 
        \wBMid27[11] , \wBMid27[10] , \wBMid27[9] , \wBMid27[8] , \wBMid27[7] , 
        \wBMid27[6] , \wBMid27[5] , \wBMid27[4] , \wBMid27[3] , \wBMid27[2] , 
        \wBMid27[1] , \wBMid27[0] }), .LoOut({\wAMid28[31] , \wAMid28[30] , 
        \wAMid28[29] , \wAMid28[28] , \wAMid28[27] , \wAMid28[26] , 
        \wAMid28[25] , \wAMid28[24] , \wAMid28[23] , \wAMid28[22] , 
        \wAMid28[21] , \wAMid28[20] , \wAMid28[19] , \wAMid28[18] , 
        \wAMid28[17] , \wAMid28[16] , \wAMid28[15] , \wAMid28[14] , 
        \wAMid28[13] , \wAMid28[12] , \wAMid28[11] , \wAMid28[10] , 
        \wAMid28[9] , \wAMid28[8] , \wAMid28[7] , \wAMid28[6] , \wAMid28[5] , 
        \wAMid28[4] , \wAMid28[3] , \wAMid28[2] , \wAMid28[1] , \wAMid28[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid7[31] , 
        \wAMid7[30] , \wAMid7[29] , \wAMid7[28] , \wAMid7[27] , \wAMid7[26] , 
        \wAMid7[25] , \wAMid7[24] , \wAMid7[23] , \wAMid7[22] , \wAMid7[21] , 
        \wAMid7[20] , \wAMid7[19] , \wAMid7[18] , \wAMid7[17] , \wAMid7[16] , 
        \wAMid7[15] , \wAMid7[14] , \wAMid7[13] , \wAMid7[12] , \wAMid7[11] , 
        \wAMid7[10] , \wAMid7[9] , \wAMid7[8] , \wAMid7[7] , \wAMid7[6] , 
        \wAMid7[5] , \wAMid7[4] , \wAMid7[3] , \wAMid7[2] , \wAMid7[1] , 
        \wAMid7[0] }), .BIn({\wBMid7[31] , \wBMid7[30] , \wBMid7[29] , 
        \wBMid7[28] , \wBMid7[27] , \wBMid7[26] , \wBMid7[25] , \wBMid7[24] , 
        \wBMid7[23] , \wBMid7[22] , \wBMid7[21] , \wBMid7[20] , \wBMid7[19] , 
        \wBMid7[18] , \wBMid7[17] , \wBMid7[16] , \wBMid7[15] , \wBMid7[14] , 
        \wBMid7[13] , \wBMid7[12] , \wBMid7[11] , \wBMid7[10] , \wBMid7[9] , 
        \wBMid7[8] , \wBMid7[7] , \wBMid7[6] , \wBMid7[5] , \wBMid7[4] , 
        \wBMid7[3] , \wBMid7[2] , \wBMid7[1] , \wBMid7[0] }), .HiOut({
        \wRegInB7[31] , \wRegInB7[30] , \wRegInB7[29] , \wRegInB7[28] , 
        \wRegInB7[27] , \wRegInB7[26] , \wRegInB7[25] , \wRegInB7[24] , 
        \wRegInB7[23] , \wRegInB7[22] , \wRegInB7[21] , \wRegInB7[20] , 
        \wRegInB7[19] , \wRegInB7[18] , \wRegInB7[17] , \wRegInB7[16] , 
        \wRegInB7[15] , \wRegInB7[14] , \wRegInB7[13] , \wRegInB7[12] , 
        \wRegInB7[11] , \wRegInB7[10] , \wRegInB7[9] , \wRegInB7[8] , 
        \wRegInB7[7] , \wRegInB7[6] , \wRegInB7[5] , \wRegInB7[4] , 
        \wRegInB7[3] , \wRegInB7[2] , \wRegInB7[1] , \wRegInB7[0] }), .LoOut({
        \wRegInA8[31] , \wRegInA8[30] , \wRegInA8[29] , \wRegInA8[28] , 
        \wRegInA8[27] , \wRegInA8[26] , \wRegInA8[25] , \wRegInA8[24] , 
        \wRegInA8[23] , \wRegInA8[22] , \wRegInA8[21] , \wRegInA8[20] , 
        \wRegInA8[19] , \wRegInA8[18] , \wRegInA8[17] , \wRegInA8[16] , 
        \wRegInA8[15] , \wRegInA8[14] , \wRegInA8[13] , \wRegInA8[12] , 
        \wRegInA8[11] , \wRegInA8[10] , \wRegInA8[9] , \wRegInA8[8] , 
        \wRegInA8[7] , \wRegInA8[6] , \wRegInA8[5] , \wRegInA8[4] , 
        \wRegInA8[3] , \wRegInA8[2] , \wRegInA8[1] , \wRegInA8[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid11[31] , \wAMid11[30] , \wAMid11[29] , \wAMid11[28] , 
        \wAMid11[27] , \wAMid11[26] , \wAMid11[25] , \wAMid11[24] , 
        \wAMid11[23] , \wAMid11[22] , \wAMid11[21] , \wAMid11[20] , 
        \wAMid11[19] , \wAMid11[18] , \wAMid11[17] , \wAMid11[16] , 
        \wAMid11[15] , \wAMid11[14] , \wAMid11[13] , \wAMid11[12] , 
        \wAMid11[11] , \wAMid11[10] , \wAMid11[9] , \wAMid11[8] , \wAMid11[7] , 
        \wAMid11[6] , \wAMid11[5] , \wAMid11[4] , \wAMid11[3] , \wAMid11[2] , 
        \wAMid11[1] , \wAMid11[0] }), .BIn({\wBMid11[31] , \wBMid11[30] , 
        \wBMid11[29] , \wBMid11[28] , \wBMid11[27] , \wBMid11[26] , 
        \wBMid11[25] , \wBMid11[24] , \wBMid11[23] , \wBMid11[22] , 
        \wBMid11[21] , \wBMid11[20] , \wBMid11[19] , \wBMid11[18] , 
        \wBMid11[17] , \wBMid11[16] , \wBMid11[15] , \wBMid11[14] , 
        \wBMid11[13] , \wBMid11[12] , \wBMid11[11] , \wBMid11[10] , 
        \wBMid11[9] , \wBMid11[8] , \wBMid11[7] , \wBMid11[6] , \wBMid11[5] , 
        \wBMid11[4] , \wBMid11[3] , \wBMid11[2] , \wBMid11[1] , \wBMid11[0] }), 
        .HiOut({\wRegInB11[31] , \wRegInB11[30] , \wRegInB11[29] , 
        \wRegInB11[28] , \wRegInB11[27] , \wRegInB11[26] , \wRegInB11[25] , 
        \wRegInB11[24] , \wRegInB11[23] , \wRegInB11[22] , \wRegInB11[21] , 
        \wRegInB11[20] , \wRegInB11[19] , \wRegInB11[18] , \wRegInB11[17] , 
        \wRegInB11[16] , \wRegInB11[15] , \wRegInB11[14] , \wRegInB11[13] , 
        \wRegInB11[12] , \wRegInB11[11] , \wRegInB11[10] , \wRegInB11[9] , 
        \wRegInB11[8] , \wRegInB11[7] , \wRegInB11[6] , \wRegInB11[5] , 
        \wRegInB11[4] , \wRegInB11[3] , \wRegInB11[2] , \wRegInB11[1] , 
        \wRegInB11[0] }), .LoOut({\wRegInA12[31] , \wRegInA12[30] , 
        \wRegInA12[29] , \wRegInA12[28] , \wRegInA12[27] , \wRegInA12[26] , 
        \wRegInA12[25] , \wRegInA12[24] , \wRegInA12[23] , \wRegInA12[22] , 
        \wRegInA12[21] , \wRegInA12[20] , \wRegInA12[19] , \wRegInA12[18] , 
        \wRegInA12[17] , \wRegInA12[16] , \wRegInA12[15] , \wRegInA12[14] , 
        \wRegInA12[13] , \wRegInA12[12] , \wRegInA12[11] , \wRegInA12[10] , 
        \wRegInA12[9] , \wRegInA12[8] , \wRegInA12[7] , \wRegInA12[6] , 
        \wRegInA12[5] , \wRegInA12[4] , \wRegInA12[3] , \wRegInA12[2] , 
        \wRegInA12[1] , \wRegInA12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_26 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink27[31] , \ScanLink27[30] , \ScanLink27[29] , 
        \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , \ScanLink27[25] , 
        \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , \ScanLink27[21] , 
        \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , \ScanLink27[17] , 
        \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , \ScanLink27[13] , 
        \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , \ScanLink27[9] , 
        \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , \ScanLink27[5] , 
        \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , \ScanLink27[1] , 
        \ScanLink27[0] }), .ScanOut({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB18[31] , \wRegInB18[30] , 
        \wRegInB18[29] , \wRegInB18[28] , \wRegInB18[27] , \wRegInB18[26] , 
        \wRegInB18[25] , \wRegInB18[24] , \wRegInB18[23] , \wRegInB18[22] , 
        \wRegInB18[21] , \wRegInB18[20] , \wRegInB18[19] , \wRegInB18[18] , 
        \wRegInB18[17] , \wRegInB18[16] , \wRegInB18[15] , \wRegInB18[14] , 
        \wRegInB18[13] , \wRegInB18[12] , \wRegInB18[11] , \wRegInB18[10] , 
        \wRegInB18[9] , \wRegInB18[8] , \wRegInB18[7] , \wRegInB18[6] , 
        \wRegInB18[5] , \wRegInB18[4] , \wRegInB18[3] , \wRegInB18[2] , 
        \wRegInB18[1] , \wRegInB18[0] }), .Out({\wBIn18[31] , \wBIn18[30] , 
        \wBIn18[29] , \wBIn18[28] , \wBIn18[27] , \wBIn18[26] , \wBIn18[25] , 
        \wBIn18[24] , \wBIn18[23] , \wBIn18[22] , \wBIn18[21] , \wBIn18[20] , 
        \wBIn18[19] , \wBIn18[18] , \wBIn18[17] , \wBIn18[16] , \wBIn18[15] , 
        \wBIn18[14] , \wBIn18[13] , \wBIn18[12] , \wBIn18[11] , \wBIn18[10] , 
        \wBIn18[9] , \wBIn18[8] , \wBIn18[7] , \wBIn18[6] , \wBIn18[5] , 
        \wBIn18[4] , \wBIn18[3] , \wBIn18[2] , \wBIn18[1] , \wBIn18[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid18[31] , \wAMid18[30] , \wAMid18[29] , \wAMid18[28] , 
        \wAMid18[27] , \wAMid18[26] , \wAMid18[25] , \wAMid18[24] , 
        \wAMid18[23] , \wAMid18[22] , \wAMid18[21] , \wAMid18[20] , 
        \wAMid18[19] , \wAMid18[18] , \wAMid18[17] , \wAMid18[16] , 
        \wAMid18[15] , \wAMid18[14] , \wAMid18[13] , \wAMid18[12] , 
        \wAMid18[11] , \wAMid18[10] , \wAMid18[9] , \wAMid18[8] , \wAMid18[7] , 
        \wAMid18[6] , \wAMid18[5] , \wAMid18[4] , \wAMid18[3] , \wAMid18[2] , 
        \wAMid18[1] , \wAMid18[0] }), .BIn({\wBMid18[31] , \wBMid18[30] , 
        \wBMid18[29] , \wBMid18[28] , \wBMid18[27] , \wBMid18[26] , 
        \wBMid18[25] , \wBMid18[24] , \wBMid18[23] , \wBMid18[22] , 
        \wBMid18[21] , \wBMid18[20] , \wBMid18[19] , \wBMid18[18] , 
        \wBMid18[17] , \wBMid18[16] , \wBMid18[15] , \wBMid18[14] , 
        \wBMid18[13] , \wBMid18[12] , \wBMid18[11] , \wBMid18[10] , 
        \wBMid18[9] , \wBMid18[8] , \wBMid18[7] , \wBMid18[6] , \wBMid18[5] , 
        \wBMid18[4] , \wBMid18[3] , \wBMid18[2] , \wBMid18[1] , \wBMid18[0] }), 
        .HiOut({\wRegInB18[31] , \wRegInB18[30] , \wRegInB18[29] , 
        \wRegInB18[28] , \wRegInB18[27] , \wRegInB18[26] , \wRegInB18[25] , 
        \wRegInB18[24] , \wRegInB18[23] , \wRegInB18[22] , \wRegInB18[21] , 
        \wRegInB18[20] , \wRegInB18[19] , \wRegInB18[18] , \wRegInB18[17] , 
        \wRegInB18[16] , \wRegInB18[15] , \wRegInB18[14] , \wRegInB18[13] , 
        \wRegInB18[12] , \wRegInB18[11] , \wRegInB18[10] , \wRegInB18[9] , 
        \wRegInB18[8] , \wRegInB18[7] , \wRegInB18[6] , \wRegInB18[5] , 
        \wRegInB18[4] , \wRegInB18[3] , \wRegInB18[2] , \wRegInB18[1] , 
        \wRegInB18[0] }), .LoOut({\wRegInA19[31] , \wRegInA19[30] , 
        \wRegInA19[29] , \wRegInA19[28] , \wRegInA19[27] , \wRegInA19[26] , 
        \wRegInA19[25] , \wRegInA19[24] , \wRegInA19[23] , \wRegInA19[22] , 
        \wRegInA19[21] , \wRegInA19[20] , \wRegInA19[19] , \wRegInA19[18] , 
        \wRegInA19[17] , \wRegInA19[16] , \wRegInA19[15] , \wRegInA19[14] , 
        \wRegInA19[13] , \wRegInA19[12] , \wRegInA19[11] , \wRegInA19[10] , 
        \wRegInA19[9] , \wRegInA19[8] , \wRegInA19[7] , \wRegInA19[6] , 
        \wRegInA19[5] , \wRegInA19[4] , \wRegInA19[3] , \wRegInA19[2] , 
        \wRegInA19[1] , \wRegInA19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_48 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink49[31] , \ScanLink49[30] , \ScanLink49[29] , 
        \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , \ScanLink49[25] , 
        \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , \ScanLink49[21] , 
        \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , \ScanLink49[17] , 
        \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , \ScanLink49[13] , 
        \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , \ScanLink49[9] , 
        \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , \ScanLink49[5] , 
        \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , \ScanLink49[1] , 
        \ScanLink49[0] }), .ScanOut({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB7[31] , \wRegInB7[30] , 
        \wRegInB7[29] , \wRegInB7[28] , \wRegInB7[27] , \wRegInB7[26] , 
        \wRegInB7[25] , \wRegInB7[24] , \wRegInB7[23] , \wRegInB7[22] , 
        \wRegInB7[21] , \wRegInB7[20] , \wRegInB7[19] , \wRegInB7[18] , 
        \wRegInB7[17] , \wRegInB7[16] , \wRegInB7[15] , \wRegInB7[14] , 
        \wRegInB7[13] , \wRegInB7[12] , \wRegInB7[11] , \wRegInB7[10] , 
        \wRegInB7[9] , \wRegInB7[8] , \wRegInB7[7] , \wRegInB7[6] , 
        \wRegInB7[5] , \wRegInB7[4] , \wRegInB7[3] , \wRegInB7[2] , 
        \wRegInB7[1] , \wRegInB7[0] }), .Out({\wBIn7[31] , \wBIn7[30] , 
        \wBIn7[29] , \wBIn7[28] , \wBIn7[27] , \wBIn7[26] , \wBIn7[25] , 
        \wBIn7[24] , \wBIn7[23] , \wBIn7[22] , \wBIn7[21] , \wBIn7[20] , 
        \wBIn7[19] , \wBIn7[18] , \wBIn7[17] , \wBIn7[16] , \wBIn7[15] , 
        \wBIn7[14] , \wBIn7[13] , \wBIn7[12] , \wBIn7[11] , \wBIn7[10] , 
        \wBIn7[9] , \wBIn7[8] , \wBIn7[7] , \wBIn7[6] , \wBIn7[5] , \wBIn7[4] , 
        \wBIn7[3] , \wBIn7[2] , \wBIn7[1] , \wBIn7[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn5[31] , 
        \wAIn5[30] , \wAIn5[29] , \wAIn5[28] , \wAIn5[27] , \wAIn5[26] , 
        \wAIn5[25] , \wAIn5[24] , \wAIn5[23] , \wAIn5[22] , \wAIn5[21] , 
        \wAIn5[20] , \wAIn5[19] , \wAIn5[18] , \wAIn5[17] , \wAIn5[16] , 
        \wAIn5[15] , \wAIn5[14] , \wAIn5[13] , \wAIn5[12] , \wAIn5[11] , 
        \wAIn5[10] , \wAIn5[9] , \wAIn5[8] , \wAIn5[7] , \wAIn5[6] , 
        \wAIn5[5] , \wAIn5[4] , \wAIn5[3] , \wAIn5[2] , \wAIn5[1] , \wAIn5[0] 
        }), .BIn({\wBIn5[31] , \wBIn5[30] , \wBIn5[29] , \wBIn5[28] , 
        \wBIn5[27] , \wBIn5[26] , \wBIn5[25] , \wBIn5[24] , \wBIn5[23] , 
        \wBIn5[22] , \wBIn5[21] , \wBIn5[20] , \wBIn5[19] , \wBIn5[18] , 
        \wBIn5[17] , \wBIn5[16] , \wBIn5[15] , \wBIn5[14] , \wBIn5[13] , 
        \wBIn5[12] , \wBIn5[11] , \wBIn5[10] , \wBIn5[9] , \wBIn5[8] , 
        \wBIn5[7] , \wBIn5[6] , \wBIn5[5] , \wBIn5[4] , \wBIn5[3] , \wBIn5[2] , 
        \wBIn5[1] , \wBIn5[0] }), .HiOut({\wBMid4[31] , \wBMid4[30] , 
        \wBMid4[29] , \wBMid4[28] , \wBMid4[27] , \wBMid4[26] , \wBMid4[25] , 
        \wBMid4[24] , \wBMid4[23] , \wBMid4[22] , \wBMid4[21] , \wBMid4[20] , 
        \wBMid4[19] , \wBMid4[18] , \wBMid4[17] , \wBMid4[16] , \wBMid4[15] , 
        \wBMid4[14] , \wBMid4[13] , \wBMid4[12] , \wBMid4[11] , \wBMid4[10] , 
        \wBMid4[9] , \wBMid4[8] , \wBMid4[7] , \wBMid4[6] , \wBMid4[5] , 
        \wBMid4[4] , \wBMid4[3] , \wBMid4[2] , \wBMid4[1] , \wBMid4[0] }), 
        .LoOut({\wAMid5[31] , \wAMid5[30] , \wAMid5[29] , \wAMid5[28] , 
        \wAMid5[27] , \wAMid5[26] , \wAMid5[25] , \wAMid5[24] , \wAMid5[23] , 
        \wAMid5[22] , \wAMid5[21] , \wAMid5[20] , \wAMid5[19] , \wAMid5[18] , 
        \wAMid5[17] , \wAMid5[16] , \wAMid5[15] , \wAMid5[14] , \wAMid5[13] , 
        \wAMid5[12] , \wAMid5[11] , \wAMid5[10] , \wAMid5[9] , \wAMid5[8] , 
        \wAMid5[7] , \wAMid5[6] , \wAMid5[5] , \wAMid5[4] , \wAMid5[3] , 
        \wAMid5[2] , \wAMid5[1] , \wAMid5[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn13[31] , \wAIn13[30] , \wAIn13[29] , \wAIn13[28] , \wAIn13[27] , 
        \wAIn13[26] , \wAIn13[25] , \wAIn13[24] , \wAIn13[23] , \wAIn13[22] , 
        \wAIn13[21] , \wAIn13[20] , \wAIn13[19] , \wAIn13[18] , \wAIn13[17] , 
        \wAIn13[16] , \wAIn13[15] , \wAIn13[14] , \wAIn13[13] , \wAIn13[12] , 
        \wAIn13[11] , \wAIn13[10] , \wAIn13[9] , \wAIn13[8] , \wAIn13[7] , 
        \wAIn13[6] , \wAIn13[5] , \wAIn13[4] , \wAIn13[3] , \wAIn13[2] , 
        \wAIn13[1] , \wAIn13[0] }), .BIn({\wBIn13[31] , \wBIn13[30] , 
        \wBIn13[29] , \wBIn13[28] , \wBIn13[27] , \wBIn13[26] , \wBIn13[25] , 
        \wBIn13[24] , \wBIn13[23] , \wBIn13[22] , \wBIn13[21] , \wBIn13[20] , 
        \wBIn13[19] , \wBIn13[18] , \wBIn13[17] , \wBIn13[16] , \wBIn13[15] , 
        \wBIn13[14] , \wBIn13[13] , \wBIn13[12] , \wBIn13[11] , \wBIn13[10] , 
        \wBIn13[9] , \wBIn13[8] , \wBIn13[7] , \wBIn13[6] , \wBIn13[5] , 
        \wBIn13[4] , \wBIn13[3] , \wBIn13[2] , \wBIn13[1] , \wBIn13[0] }), 
        .HiOut({\wBMid12[31] , \wBMid12[30] , \wBMid12[29] , \wBMid12[28] , 
        \wBMid12[27] , \wBMid12[26] , \wBMid12[25] , \wBMid12[24] , 
        \wBMid12[23] , \wBMid12[22] , \wBMid12[21] , \wBMid12[20] , 
        \wBMid12[19] , \wBMid12[18] , \wBMid12[17] , \wBMid12[16] , 
        \wBMid12[15] , \wBMid12[14] , \wBMid12[13] , \wBMid12[12] , 
        \wBMid12[11] , \wBMid12[10] , \wBMid12[9] , \wBMid12[8] , \wBMid12[7] , 
        \wBMid12[6] , \wBMid12[5] , \wBMid12[4] , \wBMid12[3] , \wBMid12[2] , 
        \wBMid12[1] , \wBMid12[0] }), .LoOut({\wAMid13[31] , \wAMid13[30] , 
        \wAMid13[29] , \wAMid13[28] , \wAMid13[27] , \wAMid13[26] , 
        \wAMid13[25] , \wAMid13[24] , \wAMid13[23] , \wAMid13[22] , 
        \wAMid13[21] , \wAMid13[20] , \wAMid13[19] , \wAMid13[18] , 
        \wAMid13[17] , \wAMid13[16] , \wAMid13[15] , \wAMid13[14] , 
        \wAMid13[13] , \wAMid13[12] , \wAMid13[11] , \wAMid13[10] , 
        \wAMid13[9] , \wAMid13[8] , \wAMid13[7] , \wAMid13[6] , \wAMid13[5] , 
        \wAMid13[4] , \wAMid13[3] , \wAMid13[2] , \wAMid13[1] , \wAMid13[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn14[31] , \wAIn14[30] , \wAIn14[29] , \wAIn14[28] , \wAIn14[27] , 
        \wAIn14[26] , \wAIn14[25] , \wAIn14[24] , \wAIn14[23] , \wAIn14[22] , 
        \wAIn14[21] , \wAIn14[20] , \wAIn14[19] , \wAIn14[18] , \wAIn14[17] , 
        \wAIn14[16] , \wAIn14[15] , \wAIn14[14] , \wAIn14[13] , \wAIn14[12] , 
        \wAIn14[11] , \wAIn14[10] , \wAIn14[9] , \wAIn14[8] , \wAIn14[7] , 
        \wAIn14[6] , \wAIn14[5] , \wAIn14[4] , \wAIn14[3] , \wAIn14[2] , 
        \wAIn14[1] , \wAIn14[0] }), .BIn({\wBIn14[31] , \wBIn14[30] , 
        \wBIn14[29] , \wBIn14[28] , \wBIn14[27] , \wBIn14[26] , \wBIn14[25] , 
        \wBIn14[24] , \wBIn14[23] , \wBIn14[22] , \wBIn14[21] , \wBIn14[20] , 
        \wBIn14[19] , \wBIn14[18] , \wBIn14[17] , \wBIn14[16] , \wBIn14[15] , 
        \wBIn14[14] , \wBIn14[13] , \wBIn14[12] , \wBIn14[11] , \wBIn14[10] , 
        \wBIn14[9] , \wBIn14[8] , \wBIn14[7] , \wBIn14[6] , \wBIn14[5] , 
        \wBIn14[4] , \wBIn14[3] , \wBIn14[2] , \wBIn14[1] , \wBIn14[0] }), 
        .HiOut({\wBMid13[31] , \wBMid13[30] , \wBMid13[29] , \wBMid13[28] , 
        \wBMid13[27] , \wBMid13[26] , \wBMid13[25] , \wBMid13[24] , 
        \wBMid13[23] , \wBMid13[22] , \wBMid13[21] , \wBMid13[20] , 
        \wBMid13[19] , \wBMid13[18] , \wBMid13[17] , \wBMid13[16] , 
        \wBMid13[15] , \wBMid13[14] , \wBMid13[13] , \wBMid13[12] , 
        \wBMid13[11] , \wBMid13[10] , \wBMid13[9] , \wBMid13[8] , \wBMid13[7] , 
        \wBMid13[6] , \wBMid13[5] , \wBMid13[4] , \wBMid13[3] , \wBMid13[2] , 
        \wBMid13[1] , \wBMid13[0] }), .LoOut({\wAMid14[31] , \wAMid14[30] , 
        \wAMid14[29] , \wAMid14[28] , \wAMid14[27] , \wAMid14[26] , 
        \wAMid14[25] , \wAMid14[24] , \wAMid14[23] , \wAMid14[22] , 
        \wAMid14[21] , \wAMid14[20] , \wAMid14[19] , \wAMid14[18] , 
        \wAMid14[17] , \wAMid14[16] , \wAMid14[15] , \wAMid14[14] , 
        \wAMid14[13] , \wAMid14[12] , \wAMid14[11] , \wAMid14[10] , 
        \wAMid14[9] , \wAMid14[8] , \wAMid14[7] , \wAMid14[6] , \wAMid14[5] , 
        \wAMid14[4] , \wAMid14[3] , \wAMid14[2] , \wAMid14[1] , \wAMid14[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_34 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink35[31] , \ScanLink35[30] , \ScanLink35[29] , 
        \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , \ScanLink35[25] , 
        \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , \ScanLink35[21] , 
        \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , \ScanLink35[17] , 
        \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , \ScanLink35[13] , 
        \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , \ScanLink35[9] , 
        \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , \ScanLink35[5] , 
        \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , \ScanLink35[1] , 
        \ScanLink35[0] }), .ScanOut({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB14[31] , \wRegInB14[30] , 
        \wRegInB14[29] , \wRegInB14[28] , \wRegInB14[27] , \wRegInB14[26] , 
        \wRegInB14[25] , \wRegInB14[24] , \wRegInB14[23] , \wRegInB14[22] , 
        \wRegInB14[21] , \wRegInB14[20] , \wRegInB14[19] , \wRegInB14[18] , 
        \wRegInB14[17] , \wRegInB14[16] , \wRegInB14[15] , \wRegInB14[14] , 
        \wRegInB14[13] , \wRegInB14[12] , \wRegInB14[11] , \wRegInB14[10] , 
        \wRegInB14[9] , \wRegInB14[8] , \wRegInB14[7] , \wRegInB14[6] , 
        \wRegInB14[5] , \wRegInB14[4] , \wRegInB14[3] , \wRegInB14[2] , 
        \wRegInB14[1] , \wRegInB14[0] }), .Out({\wBIn14[31] , \wBIn14[30] , 
        \wBIn14[29] , \wBIn14[28] , \wBIn14[27] , \wBIn14[26] , \wBIn14[25] , 
        \wBIn14[24] , \wBIn14[23] , \wBIn14[22] , \wBIn14[21] , \wBIn14[20] , 
        \wBIn14[19] , \wBIn14[18] , \wBIn14[17] , \wBIn14[16] , \wBIn14[15] , 
        \wBIn14[14] , \wBIn14[13] , \wBIn14[12] , \wBIn14[11] , \wBIn14[10] , 
        \wBIn14[9] , \wBIn14[8] , \wBIn14[7] , \wBIn14[6] , \wBIn14[5] , 
        \wBIn14[4] , \wBIn14[3] , \wBIn14[2] , \wBIn14[1] , \wBIn14[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_13 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[31] , \ScanLink14[30] , \ScanLink14[29] , 
        \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , \ScanLink14[25] , 
        \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , \ScanLink14[21] , 
        \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , \ScanLink14[17] , 
        \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , \ScanLink14[13] , 
        \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , \ScanLink14[9] , 
        \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA25[31] , \wRegInA25[30] , 
        \wRegInA25[29] , \wRegInA25[28] , \wRegInA25[27] , \wRegInA25[26] , 
        \wRegInA25[25] , \wRegInA25[24] , \wRegInA25[23] , \wRegInA25[22] , 
        \wRegInA25[21] , \wRegInA25[20] , \wRegInA25[19] , \wRegInA25[18] , 
        \wRegInA25[17] , \wRegInA25[16] , \wRegInA25[15] , \wRegInA25[14] , 
        \wRegInA25[13] , \wRegInA25[12] , \wRegInA25[11] , \wRegInA25[10] , 
        \wRegInA25[9] , \wRegInA25[8] , \wRegInA25[7] , \wRegInA25[6] , 
        \wRegInA25[5] , \wRegInA25[4] , \wRegInA25[3] , \wRegInA25[2] , 
        \wRegInA25[1] , \wRegInA25[0] }), .Out({\wAIn25[31] , \wAIn25[30] , 
        \wAIn25[29] , \wAIn25[28] , \wAIn25[27] , \wAIn25[26] , \wAIn25[25] , 
        \wAIn25[24] , \wAIn25[23] , \wAIn25[22] , \wAIn25[21] , \wAIn25[20] , 
        \wAIn25[19] , \wAIn25[18] , \wAIn25[17] , \wAIn25[16] , \wAIn25[15] , 
        \wAIn25[14] , \wAIn25[13] , \wAIn25[12] , \wAIn25[11] , \wAIn25[10] , 
        \wAIn25[9] , \wAIn25[8] , \wAIn25[7] , \wAIn25[6] , \wAIn25[5] , 
        \wAIn25[4] , \wAIn25[3] , \wAIn25[2] , \wAIn25[1] , \wAIn25[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid9[31] , 
        \wAMid9[30] , \wAMid9[29] , \wAMid9[28] , \wAMid9[27] , \wAMid9[26] , 
        \wAMid9[25] , \wAMid9[24] , \wAMid9[23] , \wAMid9[22] , \wAMid9[21] , 
        \wAMid9[20] , \wAMid9[19] , \wAMid9[18] , \wAMid9[17] , \wAMid9[16] , 
        \wAMid9[15] , \wAMid9[14] , \wAMid9[13] , \wAMid9[12] , \wAMid9[11] , 
        \wAMid9[10] , \wAMid9[9] , \wAMid9[8] , \wAMid9[7] , \wAMid9[6] , 
        \wAMid9[5] , \wAMid9[4] , \wAMid9[3] , \wAMid9[2] , \wAMid9[1] , 
        \wAMid9[0] }), .BIn({\wBMid9[31] , \wBMid9[30] , \wBMid9[29] , 
        \wBMid9[28] , \wBMid9[27] , \wBMid9[26] , \wBMid9[25] , \wBMid9[24] , 
        \wBMid9[23] , \wBMid9[22] , \wBMid9[21] , \wBMid9[20] , \wBMid9[19] , 
        \wBMid9[18] , \wBMid9[17] , \wBMid9[16] , \wBMid9[15] , \wBMid9[14] , 
        \wBMid9[13] , \wBMid9[12] , \wBMid9[11] , \wBMid9[10] , \wBMid9[9] , 
        \wBMid9[8] , \wBMid9[7] , \wBMid9[6] , \wBMid9[5] , \wBMid9[4] , 
        \wBMid9[3] , \wBMid9[2] , \wBMid9[1] , \wBMid9[0] }), .HiOut({
        \wRegInB9[31] , \wRegInB9[30] , \wRegInB9[29] , \wRegInB9[28] , 
        \wRegInB9[27] , \wRegInB9[26] , \wRegInB9[25] , \wRegInB9[24] , 
        \wRegInB9[23] , \wRegInB9[22] , \wRegInB9[21] , \wRegInB9[20] , 
        \wRegInB9[19] , \wRegInB9[18] , \wRegInB9[17] , \wRegInB9[16] , 
        \wRegInB9[15] , \wRegInB9[14] , \wRegInB9[13] , \wRegInB9[12] , 
        \wRegInB9[11] , \wRegInB9[10] , \wRegInB9[9] , \wRegInB9[8] , 
        \wRegInB9[7] , \wRegInB9[6] , \wRegInB9[5] , \wRegInB9[4] , 
        \wRegInB9[3] , \wRegInB9[2] , \wRegInB9[1] , \wRegInB9[0] }), .LoOut({
        \wRegInA10[31] , \wRegInA10[30] , \wRegInA10[29] , \wRegInA10[28] , 
        \wRegInA10[27] , \wRegInA10[26] , \wRegInA10[25] , \wRegInA10[24] , 
        \wRegInA10[23] , \wRegInA10[22] , \wRegInA10[21] , \wRegInA10[20] , 
        \wRegInA10[19] , \wRegInA10[18] , \wRegInA10[17] , \wRegInA10[16] , 
        \wRegInA10[15] , \wRegInA10[14] , \wRegInA10[13] , \wRegInA10[12] , 
        \wRegInA10[11] , \wRegInA10[10] , \wRegInA10[9] , \wRegInA10[8] , 
        \wRegInA10[7] , \wRegInA10[6] , \wRegInA10[5] , \wRegInA10[4] , 
        \wRegInA10[3] , \wRegInA10[2] , \wRegInA10[1] , \wRegInA10[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid24[31] , \wAMid24[30] , \wAMid24[29] , \wAMid24[28] , 
        \wAMid24[27] , \wAMid24[26] , \wAMid24[25] , \wAMid24[24] , 
        \wAMid24[23] , \wAMid24[22] , \wAMid24[21] , \wAMid24[20] , 
        \wAMid24[19] , \wAMid24[18] , \wAMid24[17] , \wAMid24[16] , 
        \wAMid24[15] , \wAMid24[14] , \wAMid24[13] , \wAMid24[12] , 
        \wAMid24[11] , \wAMid24[10] , \wAMid24[9] , \wAMid24[8] , \wAMid24[7] , 
        \wAMid24[6] , \wAMid24[5] , \wAMid24[4] , \wAMid24[3] , \wAMid24[2] , 
        \wAMid24[1] , \wAMid24[0] }), .BIn({\wBMid24[31] , \wBMid24[30] , 
        \wBMid24[29] , \wBMid24[28] , \wBMid24[27] , \wBMid24[26] , 
        \wBMid24[25] , \wBMid24[24] , \wBMid24[23] , \wBMid24[22] , 
        \wBMid24[21] , \wBMid24[20] , \wBMid24[19] , \wBMid24[18] , 
        \wBMid24[17] , \wBMid24[16] , \wBMid24[15] , \wBMid24[14] , 
        \wBMid24[13] , \wBMid24[12] , \wBMid24[11] , \wBMid24[10] , 
        \wBMid24[9] , \wBMid24[8] , \wBMid24[7] , \wBMid24[6] , \wBMid24[5] , 
        \wBMid24[4] , \wBMid24[3] , \wBMid24[2] , \wBMid24[1] , \wBMid24[0] }), 
        .HiOut({\wRegInB24[31] , \wRegInB24[30] , \wRegInB24[29] , 
        \wRegInB24[28] , \wRegInB24[27] , \wRegInB24[26] , \wRegInB24[25] , 
        \wRegInB24[24] , \wRegInB24[23] , \wRegInB24[22] , \wRegInB24[21] , 
        \wRegInB24[20] , \wRegInB24[19] , \wRegInB24[18] , \wRegInB24[17] , 
        \wRegInB24[16] , \wRegInB24[15] , \wRegInB24[14] , \wRegInB24[13] , 
        \wRegInB24[12] , \wRegInB24[11] , \wRegInB24[10] , \wRegInB24[9] , 
        \wRegInB24[8] , \wRegInB24[7] , \wRegInB24[6] , \wRegInB24[5] , 
        \wRegInB24[4] , \wRegInB24[3] , \wRegInB24[2] , \wRegInB24[1] , 
        \wRegInB24[0] }), .LoOut({\wRegInA25[31] , \wRegInA25[30] , 
        \wRegInA25[29] , \wRegInA25[28] , \wRegInA25[27] , \wRegInA25[26] , 
        \wRegInA25[25] , \wRegInA25[24] , \wRegInA25[23] , \wRegInA25[22] , 
        \wRegInA25[21] , \wRegInA25[20] , \wRegInA25[19] , \wRegInA25[18] , 
        \wRegInA25[17] , \wRegInA25[16] , \wRegInA25[15] , \wRegInA25[14] , 
        \wRegInA25[13] , \wRegInA25[12] , \wRegInA25[11] , \wRegInA25[10] , 
        \wRegInA25[9] , \wRegInA25[8] , \wRegInA25[7] , \wRegInA25[6] , 
        \wRegInA25[5] , \wRegInA25[4] , \wRegInA25[3] , \wRegInA25[2] , 
        \wRegInA25[1] , \wRegInA25[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_41 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink42[31] , \ScanLink42[30] , \ScanLink42[29] , 
        \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , \ScanLink42[25] , 
        \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , \ScanLink42[21] , 
        \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , \ScanLink42[17] , 
        \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , \ScanLink42[13] , 
        \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , \ScanLink42[9] , 
        \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , \ScanLink42[5] , 
        \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , \ScanLink42[1] , 
        \ScanLink42[0] }), .ScanOut({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA11[31] , \wRegInA11[30] , 
        \wRegInA11[29] , \wRegInA11[28] , \wRegInA11[27] , \wRegInA11[26] , 
        \wRegInA11[25] , \wRegInA11[24] , \wRegInA11[23] , \wRegInA11[22] , 
        \wRegInA11[21] , \wRegInA11[20] , \wRegInA11[19] , \wRegInA11[18] , 
        \wRegInA11[17] , \wRegInA11[16] , \wRegInA11[15] , \wRegInA11[14] , 
        \wRegInA11[13] , \wRegInA11[12] , \wRegInA11[11] , \wRegInA11[10] , 
        \wRegInA11[9] , \wRegInA11[8] , \wRegInA11[7] , \wRegInA11[6] , 
        \wRegInA11[5] , \wRegInA11[4] , \wRegInA11[3] , \wRegInA11[2] , 
        \wRegInA11[1] , \wRegInA11[0] }), .Out({\wAIn11[31] , \wAIn11[30] , 
        \wAIn11[29] , \wAIn11[28] , \wAIn11[27] , \wAIn11[26] , \wAIn11[25] , 
        \wAIn11[24] , \wAIn11[23] , \wAIn11[22] , \wAIn11[21] , \wAIn11[20] , 
        \wAIn11[19] , \wAIn11[18] , \wAIn11[17] , \wAIn11[16] , \wAIn11[15] , 
        \wAIn11[14] , \wAIn11[13] , \wAIn11[12] , \wAIn11[11] , \wAIn11[10] , 
        \wAIn11[9] , \wAIn11[8] , \wAIn11[7] , \wAIn11[6] , \wAIn11[5] , 
        \wAIn11[4] , \wAIn11[3] , \wAIn11[2] , \wAIn11[1] , \wAIn11[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_2 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[31] , \ScanLink3[30] , \ScanLink3[29] , 
        \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , \ScanLink3[25] , 
        \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , \ScanLink3[21] , 
        \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , \ScanLink3[17] , 
        \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , \ScanLink3[13] , 
        \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , \ScanLink3[9] , 
        \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB30[31] , \wRegInB30[30] , 
        \wRegInB30[29] , \wRegInB30[28] , \wRegInB30[27] , \wRegInB30[26] , 
        \wRegInB30[25] , \wRegInB30[24] , \wRegInB30[23] , \wRegInB30[22] , 
        \wRegInB30[21] , \wRegInB30[20] , \wRegInB30[19] , \wRegInB30[18] , 
        \wRegInB30[17] , \wRegInB30[16] , \wRegInB30[15] , \wRegInB30[14] , 
        \wRegInB30[13] , \wRegInB30[12] , \wRegInB30[11] , \wRegInB30[10] , 
        \wRegInB30[9] , \wRegInB30[8] , \wRegInB30[7] , \wRegInB30[6] , 
        \wRegInB30[5] , \wRegInB30[4] , \wRegInB30[3] , \wRegInB30[2] , 
        \wRegInB30[1] , \wRegInB30[0] }), .Out({\wBIn30[31] , \wBIn30[30] , 
        \wBIn30[29] , \wBIn30[28] , \wBIn30[27] , \wBIn30[26] , \wBIn30[25] , 
        \wBIn30[24] , \wBIn30[23] , \wBIn30[22] , \wBIn30[21] , \wBIn30[20] , 
        \wBIn30[19] , \wBIn30[18] , \wBIn30[17] , \wBIn30[16] , \wBIn30[15] , 
        \wBIn30[14] , \wBIn30[13] , \wBIn30[12] , \wBIn30[11] , \wBIn30[10] , 
        \wBIn30[9] , \wBIn30[8] , \wBIn30[7] , \wBIn30[6] , \wBIn30[5] , 
        \wBIn30[4] , \wBIn30[3] , \wBIn30[2] , \wBIn30[1] , \wBIn30[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid23[31] , \wAMid23[30] , \wAMid23[29] , \wAMid23[28] , 
        \wAMid23[27] , \wAMid23[26] , \wAMid23[25] , \wAMid23[24] , 
        \wAMid23[23] , \wAMid23[22] , \wAMid23[21] , \wAMid23[20] , 
        \wAMid23[19] , \wAMid23[18] , \wAMid23[17] , \wAMid23[16] , 
        \wAMid23[15] , \wAMid23[14] , \wAMid23[13] , \wAMid23[12] , 
        \wAMid23[11] , \wAMid23[10] , \wAMid23[9] , \wAMid23[8] , \wAMid23[7] , 
        \wAMid23[6] , \wAMid23[5] , \wAMid23[4] , \wAMid23[3] , \wAMid23[2] , 
        \wAMid23[1] , \wAMid23[0] }), .BIn({\wBMid23[31] , \wBMid23[30] , 
        \wBMid23[29] , \wBMid23[28] , \wBMid23[27] , \wBMid23[26] , 
        \wBMid23[25] , \wBMid23[24] , \wBMid23[23] , \wBMid23[22] , 
        \wBMid23[21] , \wBMid23[20] , \wBMid23[19] , \wBMid23[18] , 
        \wBMid23[17] , \wBMid23[16] , \wBMid23[15] , \wBMid23[14] , 
        \wBMid23[13] , \wBMid23[12] , \wBMid23[11] , \wBMid23[10] , 
        \wBMid23[9] , \wBMid23[8] , \wBMid23[7] , \wBMid23[6] , \wBMid23[5] , 
        \wBMid23[4] , \wBMid23[3] , \wBMid23[2] , \wBMid23[1] , \wBMid23[0] }), 
        .HiOut({\wRegInB23[31] , \wRegInB23[30] , \wRegInB23[29] , 
        \wRegInB23[28] , \wRegInB23[27] , \wRegInB23[26] , \wRegInB23[25] , 
        \wRegInB23[24] , \wRegInB23[23] , \wRegInB23[22] , \wRegInB23[21] , 
        \wRegInB23[20] , \wRegInB23[19] , \wRegInB23[18] , \wRegInB23[17] , 
        \wRegInB23[16] , \wRegInB23[15] , \wRegInB23[14] , \wRegInB23[13] , 
        \wRegInB23[12] , \wRegInB23[11] , \wRegInB23[10] , \wRegInB23[9] , 
        \wRegInB23[8] , \wRegInB23[7] , \wRegInB23[6] , \wRegInB23[5] , 
        \wRegInB23[4] , \wRegInB23[3] , \wRegInB23[2] , \wRegInB23[1] , 
        \wRegInB23[0] }), .LoOut({\wRegInA24[31] , \wRegInA24[30] , 
        \wRegInA24[29] , \wRegInA24[28] , \wRegInA24[27] , \wRegInA24[26] , 
        \wRegInA24[25] , \wRegInA24[24] , \wRegInA24[23] , \wRegInA24[22] , 
        \wRegInA24[21] , \wRegInA24[20] , \wRegInA24[19] , \wRegInA24[18] , 
        \wRegInA24[17] , \wRegInA24[16] , \wRegInA24[15] , \wRegInA24[14] , 
        \wRegInA24[13] , \wRegInA24[12] , \wRegInA24[11] , \wRegInA24[10] , 
        \wRegInA24[9] , \wRegInA24[8] , \wRegInA24[7] , \wRegInA24[6] , 
        \wRegInA24[5] , \wRegInA24[4] , \wRegInA24[3] , \wRegInA24[2] , 
        \wRegInA24[1] , \wRegInA24[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_61 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink62[31] , \ScanLink62[30] , \ScanLink62[29] , 
        \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , \ScanLink62[25] , 
        \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , \ScanLink62[21] , 
        \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , \ScanLink62[17] , 
        \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , \ScanLink62[13] , 
        \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , \ScanLink62[9] , 
        \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , \ScanLink62[5] , 
        \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , \ScanLink62[1] , 
        \ScanLink62[0] }), .ScanOut({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA1[31] , \wRegInA1[30] , 
        \wRegInA1[29] , \wRegInA1[28] , \wRegInA1[27] , \wRegInA1[26] , 
        \wRegInA1[25] , \wRegInA1[24] , \wRegInA1[23] , \wRegInA1[22] , 
        \wRegInA1[21] , \wRegInA1[20] , \wRegInA1[19] , \wRegInA1[18] , 
        \wRegInA1[17] , \wRegInA1[16] , \wRegInA1[15] , \wRegInA1[14] , 
        \wRegInA1[13] , \wRegInA1[12] , \wRegInA1[11] , \wRegInA1[10] , 
        \wRegInA1[9] , \wRegInA1[8] , \wRegInA1[7] , \wRegInA1[6] , 
        \wRegInA1[5] , \wRegInA1[4] , \wRegInA1[3] , \wRegInA1[2] , 
        \wRegInA1[1] , \wRegInA1[0] }), .Out({\wAIn1[31] , \wAIn1[30] , 
        \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , \wAIn1[26] , \wAIn1[25] , 
        \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , \wAIn1[21] , \wAIn1[20] , 
        \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , \wAIn1[16] , \wAIn1[15] , 
        \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , \wAIn1[11] , \wAIn1[10] , 
        \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , \wAIn1[6] , \wAIn1[5] , \wAIn1[4] , 
        \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , \wAIn1[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_5 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[31] , \ScanLink6[30] , \ScanLink6[29] , 
        \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , \ScanLink6[25] , 
        \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , \ScanLink6[21] , 
        \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , \ScanLink6[17] , 
        \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , \ScanLink6[13] , 
        \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , \ScanLink6[9] , 
        \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA29[31] , \wRegInA29[30] , 
        \wRegInA29[29] , \wRegInA29[28] , \wRegInA29[27] , \wRegInA29[26] , 
        \wRegInA29[25] , \wRegInA29[24] , \wRegInA29[23] , \wRegInA29[22] , 
        \wRegInA29[21] , \wRegInA29[20] , \wRegInA29[19] , \wRegInA29[18] , 
        \wRegInA29[17] , \wRegInA29[16] , \wRegInA29[15] , \wRegInA29[14] , 
        \wRegInA29[13] , \wRegInA29[12] , \wRegInA29[11] , \wRegInA29[10] , 
        \wRegInA29[9] , \wRegInA29[8] , \wRegInA29[7] , \wRegInA29[6] , 
        \wRegInA29[5] , \wRegInA29[4] , \wRegInA29[3] , \wRegInA29[2] , 
        \wRegInA29[1] , \wRegInA29[0] }), .Out({\wAIn29[31] , \wAIn29[30] , 
        \wAIn29[29] , \wAIn29[28] , \wAIn29[27] , \wAIn29[26] , \wAIn29[25] , 
        \wAIn29[24] , \wAIn29[23] , \wAIn29[22] , \wAIn29[21] , \wAIn29[20] , 
        \wAIn29[19] , \wAIn29[18] , \wAIn29[17] , \wAIn29[16] , \wAIn29[15] , 
        \wAIn29[14] , \wAIn29[13] , \wAIn29[12] , \wAIn29[11] , \wAIn29[10] , 
        \wAIn29[9] , \wAIn29[8] , \wAIn29[7] , \wAIn29[6] , \wAIn29[5] , 
        \wAIn29[4] , \wAIn29[3] , \wAIn29[2] , \wAIn29[1] , \wAIn29[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_46 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink47[31] , \ScanLink47[30] , \ScanLink47[29] , 
        \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , \ScanLink47[25] , 
        \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , \ScanLink47[21] , 
        \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , \ScanLink47[17] , 
        \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , \ScanLink47[13] , 
        \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , \ScanLink47[9] , 
        \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , \ScanLink47[5] , 
        \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , \ScanLink47[1] , 
        \ScanLink47[0] }), .ScanOut({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB8[31] , \wRegInB8[30] , 
        \wRegInB8[29] , \wRegInB8[28] , \wRegInB8[27] , \wRegInB8[26] , 
        \wRegInB8[25] , \wRegInB8[24] , \wRegInB8[23] , \wRegInB8[22] , 
        \wRegInB8[21] , \wRegInB8[20] , \wRegInB8[19] , \wRegInB8[18] , 
        \wRegInB8[17] , \wRegInB8[16] , \wRegInB8[15] , \wRegInB8[14] , 
        \wRegInB8[13] , \wRegInB8[12] , \wRegInB8[11] , \wRegInB8[10] , 
        \wRegInB8[9] , \wRegInB8[8] , \wRegInB8[7] , \wRegInB8[6] , 
        \wRegInB8[5] , \wRegInB8[4] , \wRegInB8[3] , \wRegInB8[2] , 
        \wRegInB8[1] , \wRegInB8[0] }), .Out({\wBIn8[31] , \wBIn8[30] , 
        \wBIn8[29] , \wBIn8[28] , \wBIn8[27] , \wBIn8[26] , \wBIn8[25] , 
        \wBIn8[24] , \wBIn8[23] , \wBIn8[22] , \wBIn8[21] , \wBIn8[20] , 
        \wBIn8[19] , \wBIn8[18] , \wBIn8[17] , \wBIn8[16] , \wBIn8[15] , 
        \wBIn8[14] , \wBIn8[13] , \wBIn8[12] , \wBIn8[11] , \wBIn8[10] , 
        \wBIn8[9] , \wBIn8[8] , \wBIn8[7] , \wBIn8[6] , \wBIn8[5] , \wBIn8[4] , 
        \wBIn8[3] , \wBIn8[2] , \wBIn8[1] , \wBIn8[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_33 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink34[31] , \ScanLink34[30] , \ScanLink34[29] , 
        \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , \ScanLink34[25] , 
        \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , \ScanLink34[21] , 
        \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , \ScanLink34[17] , 
        \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , \ScanLink34[13] , 
        \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , \ScanLink34[9] , 
        \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , \ScanLink34[5] , 
        \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , \ScanLink34[1] , 
        \ScanLink34[0] }), .ScanOut({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA15[31] , \wRegInA15[30] , 
        \wRegInA15[29] , \wRegInA15[28] , \wRegInA15[27] , \wRegInA15[26] , 
        \wRegInA15[25] , \wRegInA15[24] , \wRegInA15[23] , \wRegInA15[22] , 
        \wRegInA15[21] , \wRegInA15[20] , \wRegInA15[19] , \wRegInA15[18] , 
        \wRegInA15[17] , \wRegInA15[16] , \wRegInA15[15] , \wRegInA15[14] , 
        \wRegInA15[13] , \wRegInA15[12] , \wRegInA15[11] , \wRegInA15[10] , 
        \wRegInA15[9] , \wRegInA15[8] , \wRegInA15[7] , \wRegInA15[6] , 
        \wRegInA15[5] , \wRegInA15[4] , \wRegInA15[3] , \wRegInA15[2] , 
        \wRegInA15[1] , \wRegInA15[0] }), .Out({\wAIn15[31] , \wAIn15[30] , 
        \wAIn15[29] , \wAIn15[28] , \wAIn15[27] , \wAIn15[26] , \wAIn15[25] , 
        \wAIn15[24] , \wAIn15[23] , \wAIn15[22] , \wAIn15[21] , \wAIn15[20] , 
        \wAIn15[19] , \wAIn15[18] , \wAIn15[17] , \wAIn15[16] , \wAIn15[15] , 
        \wAIn15[14] , \wAIn15[13] , \wAIn15[12] , \wAIn15[11] , \wAIn15[10] , 
        \wAIn15[9] , \wAIn15[8] , \wAIn15[7] , \wAIn15[6] , \wAIn15[5] , 
        \wAIn15[4] , \wAIn15[3] , \wAIn15[2] , \wAIn15[1] , \wAIn15[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_28 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink29[31] , \ScanLink29[30] , \ScanLink29[29] , 
        \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , \ScanLink29[25] , 
        \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , \ScanLink29[21] , 
        \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , \ScanLink29[17] , 
        \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , \ScanLink29[13] , 
        \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , \ScanLink29[9] , 
        \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , \ScanLink29[5] , 
        \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , \ScanLink29[1] , 
        \ScanLink29[0] }), .ScanOut({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB17[31] , \wRegInB17[30] , 
        \wRegInB17[29] , \wRegInB17[28] , \wRegInB17[27] , \wRegInB17[26] , 
        \wRegInB17[25] , \wRegInB17[24] , \wRegInB17[23] , \wRegInB17[22] , 
        \wRegInB17[21] , \wRegInB17[20] , \wRegInB17[19] , \wRegInB17[18] , 
        \wRegInB17[17] , \wRegInB17[16] , \wRegInB17[15] , \wRegInB17[14] , 
        \wRegInB17[13] , \wRegInB17[12] , \wRegInB17[11] , \wRegInB17[10] , 
        \wRegInB17[9] , \wRegInB17[8] , \wRegInB17[7] , \wRegInB17[6] , 
        \wRegInB17[5] , \wRegInB17[4] , \wRegInB17[3] , \wRegInB17[2] , 
        \wRegInB17[1] , \wRegInB17[0] }), .Out({\wBIn17[31] , \wBIn17[30] , 
        \wBIn17[29] , \wBIn17[28] , \wBIn17[27] , \wBIn17[26] , \wBIn17[25] , 
        \wBIn17[24] , \wBIn17[23] , \wBIn17[22] , \wBIn17[21] , \wBIn17[20] , 
        \wBIn17[19] , \wBIn17[18] , \wBIn17[17] , \wBIn17[16] , \wBIn17[15] , 
        \wBIn17[14] , \wBIn17[13] , \wBIn17[12] , \wBIn17[11] , \wBIn17[10] , 
        \wBIn17[9] , \wBIn17[8] , \wBIn17[7] , \wBIn17[6] , \wBIn17[5] , 
        \wBIn17[4] , \wBIn17[3] , \wBIn17[2] , \wBIn17[1] , \wBIn17[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_14 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[31] , \ScanLink15[30] , \ScanLink15[29] , 
        \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , \ScanLink15[25] , 
        \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , \ScanLink15[21] , 
        \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , \ScanLink15[17] , 
        \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , \ScanLink15[13] , 
        \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , \ScanLink15[9] , 
        \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB24[31] , \wRegInB24[30] , 
        \wRegInB24[29] , \wRegInB24[28] , \wRegInB24[27] , \wRegInB24[26] , 
        \wRegInB24[25] , \wRegInB24[24] , \wRegInB24[23] , \wRegInB24[22] , 
        \wRegInB24[21] , \wRegInB24[20] , \wRegInB24[19] , \wRegInB24[18] , 
        \wRegInB24[17] , \wRegInB24[16] , \wRegInB24[15] , \wRegInB24[14] , 
        \wRegInB24[13] , \wRegInB24[12] , \wRegInB24[11] , \wRegInB24[10] , 
        \wRegInB24[9] , \wRegInB24[8] , \wRegInB24[7] , \wRegInB24[6] , 
        \wRegInB24[5] , \wRegInB24[4] , \wRegInB24[3] , \wRegInB24[2] , 
        \wRegInB24[1] , \wRegInB24[0] }), .Out({\wBIn24[31] , \wBIn24[30] , 
        \wBIn24[29] , \wBIn24[28] , \wBIn24[27] , \wBIn24[26] , \wBIn24[25] , 
        \wBIn24[24] , \wBIn24[23] , \wBIn24[22] , \wBIn24[21] , \wBIn24[20] , 
        \wBIn24[19] , \wBIn24[18] , \wBIn24[17] , \wBIn24[16] , \wBIn24[15] , 
        \wBIn24[14] , \wBIn24[13] , \wBIn24[12] , \wBIn24[11] , \wBIn24[10] , 
        \wBIn24[9] , \wBIn24[8] , \wBIn24[7] , \wBIn24[6] , \wBIn24[5] , 
        \wBIn24[4] , \wBIn24[3] , \wBIn24[2] , \wBIn24[1] , \wBIn24[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn7[31] , 
        \wAIn7[30] , \wAIn7[29] , \wAIn7[28] , \wAIn7[27] , \wAIn7[26] , 
        \wAIn7[25] , \wAIn7[24] , \wAIn7[23] , \wAIn7[22] , \wAIn7[21] , 
        \wAIn7[20] , \wAIn7[19] , \wAIn7[18] , \wAIn7[17] , \wAIn7[16] , 
        \wAIn7[15] , \wAIn7[14] , \wAIn7[13] , \wAIn7[12] , \wAIn7[11] , 
        \wAIn7[10] , \wAIn7[9] , \wAIn7[8] , \wAIn7[7] , \wAIn7[6] , 
        \wAIn7[5] , \wAIn7[4] , \wAIn7[3] , \wAIn7[2] , \wAIn7[1] , \wAIn7[0] 
        }), .BIn({\wBIn7[31] , \wBIn7[30] , \wBIn7[29] , \wBIn7[28] , 
        \wBIn7[27] , \wBIn7[26] , \wBIn7[25] , \wBIn7[24] , \wBIn7[23] , 
        \wBIn7[22] , \wBIn7[21] , \wBIn7[20] , \wBIn7[19] , \wBIn7[18] , 
        \wBIn7[17] , \wBIn7[16] , \wBIn7[15] , \wBIn7[14] , \wBIn7[13] , 
        \wBIn7[12] , \wBIn7[11] , \wBIn7[10] , \wBIn7[9] , \wBIn7[8] , 
        \wBIn7[7] , \wBIn7[6] , \wBIn7[5] , \wBIn7[4] , \wBIn7[3] , \wBIn7[2] , 
        \wBIn7[1] , \wBIn7[0] }), .HiOut({\wBMid6[31] , \wBMid6[30] , 
        \wBMid6[29] , \wBMid6[28] , \wBMid6[27] , \wBMid6[26] , \wBMid6[25] , 
        \wBMid6[24] , \wBMid6[23] , \wBMid6[22] , \wBMid6[21] , \wBMid6[20] , 
        \wBMid6[19] , \wBMid6[18] , \wBMid6[17] , \wBMid6[16] , \wBMid6[15] , 
        \wBMid6[14] , \wBMid6[13] , \wBMid6[12] , \wBMid6[11] , \wBMid6[10] , 
        \wBMid6[9] , \wBMid6[8] , \wBMid6[7] , \wBMid6[6] , \wBMid6[5] , 
        \wBMid6[4] , \wBMid6[3] , \wBMid6[2] , \wBMid6[1] , \wBMid6[0] }), 
        .LoOut({\wAMid7[31] , \wAMid7[30] , \wAMid7[29] , \wAMid7[28] , 
        \wAMid7[27] , \wAMid7[26] , \wAMid7[25] , \wAMid7[24] , \wAMid7[23] , 
        \wAMid7[22] , \wAMid7[21] , \wAMid7[20] , \wAMid7[19] , \wAMid7[18] , 
        \wAMid7[17] , \wAMid7[16] , \wAMid7[15] , \wAMid7[14] , \wAMid7[13] , 
        \wAMid7[12] , \wAMid7[11] , \wAMid7[10] , \wAMid7[9] , \wAMid7[8] , 
        \wAMid7[7] , \wAMid7[6] , \wAMid7[5] , \wAMid7[4] , \wAMid7[3] , 
        \wAMid7[2] , \wAMid7[1] , \wAMid7[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn26[31] , \wAIn26[30] , \wAIn26[29] , \wAIn26[28] , \wAIn26[27] , 
        \wAIn26[26] , \wAIn26[25] , \wAIn26[24] , \wAIn26[23] , \wAIn26[22] , 
        \wAIn26[21] , \wAIn26[20] , \wAIn26[19] , \wAIn26[18] , \wAIn26[17] , 
        \wAIn26[16] , \wAIn26[15] , \wAIn26[14] , \wAIn26[13] , \wAIn26[12] , 
        \wAIn26[11] , \wAIn26[10] , \wAIn26[9] , \wAIn26[8] , \wAIn26[7] , 
        \wAIn26[6] , \wAIn26[5] , \wAIn26[4] , \wAIn26[3] , \wAIn26[2] , 
        \wAIn26[1] , \wAIn26[0] }), .BIn({\wBIn26[31] , \wBIn26[30] , 
        \wBIn26[29] , \wBIn26[28] , \wBIn26[27] , \wBIn26[26] , \wBIn26[25] , 
        \wBIn26[24] , \wBIn26[23] , \wBIn26[22] , \wBIn26[21] , \wBIn26[20] , 
        \wBIn26[19] , \wBIn26[18] , \wBIn26[17] , \wBIn26[16] , \wBIn26[15] , 
        \wBIn26[14] , \wBIn26[13] , \wBIn26[12] , \wBIn26[11] , \wBIn26[10] , 
        \wBIn26[9] , \wBIn26[8] , \wBIn26[7] , \wBIn26[6] , \wBIn26[5] , 
        \wBIn26[4] , \wBIn26[3] , \wBIn26[2] , \wBIn26[1] , \wBIn26[0] }), 
        .HiOut({\wBMid25[31] , \wBMid25[30] , \wBMid25[29] , \wBMid25[28] , 
        \wBMid25[27] , \wBMid25[26] , \wBMid25[25] , \wBMid25[24] , 
        \wBMid25[23] , \wBMid25[22] , \wBMid25[21] , \wBMid25[20] , 
        \wBMid25[19] , \wBMid25[18] , \wBMid25[17] , \wBMid25[16] , 
        \wBMid25[15] , \wBMid25[14] , \wBMid25[13] , \wBMid25[12] , 
        \wBMid25[11] , \wBMid25[10] , \wBMid25[9] , \wBMid25[8] , \wBMid25[7] , 
        \wBMid25[6] , \wBMid25[5] , \wBMid25[4] , \wBMid25[3] , \wBMid25[2] , 
        \wBMid25[1] , \wBMid25[0] }), .LoOut({\wAMid26[31] , \wAMid26[30] , 
        \wAMid26[29] , \wAMid26[28] , \wAMid26[27] , \wAMid26[26] , 
        \wAMid26[25] , \wAMid26[24] , \wAMid26[23] , \wAMid26[22] , 
        \wAMid26[21] , \wAMid26[20] , \wAMid26[19] , \wAMid26[18] , 
        \wAMid26[17] , \wAMid26[16] , \wAMid26[15] , \wAMid26[14] , 
        \wAMid26[13] , \wAMid26[12] , \wAMid26[11] , \wAMid26[10] , 
        \wAMid26[9] , \wAMid26[8] , \wAMid26[7] , \wAMid26[6] , \wAMid26[5] , 
        \wAMid26[4] , \wAMid26[3] , \wAMid26[2] , \wAMid26[1] , \wAMid26[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid0[31] , 
        \wAMid0[30] , \wAMid0[29] , \wAMid0[28] , \wAMid0[27] , \wAMid0[26] , 
        \wAMid0[25] , \wAMid0[24] , \wAMid0[23] , \wAMid0[22] , \wAMid0[21] , 
        \wAMid0[20] , \wAMid0[19] , \wAMid0[18] , \wAMid0[17] , \wAMid0[16] , 
        \wAMid0[15] , \wAMid0[14] , \wAMid0[13] , \wAMid0[12] , \wAMid0[11] , 
        \wAMid0[10] , \wAMid0[9] , \wAMid0[8] , \wAMid0[7] , \wAMid0[6] , 
        \wAMid0[5] , \wAMid0[4] , \wAMid0[3] , \wAMid0[2] , \wAMid0[1] , 
        \wAMid0[0] }), .BIn({\wBMid0[31] , \wBMid0[30] , \wBMid0[29] , 
        \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , \wBMid0[24] , 
        \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , \wBMid0[19] , 
        \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , \wBMid0[14] , 
        \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , \wBMid0[9] , 
        \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , \wBMid0[4] , 
        \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), .HiOut({
        \wRegInB0[31] , \wRegInB0[30] , \wRegInB0[29] , \wRegInB0[28] , 
        \wRegInB0[27] , \wRegInB0[26] , \wRegInB0[25] , \wRegInB0[24] , 
        \wRegInB0[23] , \wRegInB0[22] , \wRegInB0[21] , \wRegInB0[20] , 
        \wRegInB0[19] , \wRegInB0[18] , \wRegInB0[17] , \wRegInB0[16] , 
        \wRegInB0[15] , \wRegInB0[14] , \wRegInB0[13] , \wRegInB0[12] , 
        \wRegInB0[11] , \wRegInB0[10] , \wRegInB0[9] , \wRegInB0[8] , 
        \wRegInB0[7] , \wRegInB0[6] , \wRegInB0[5] , \wRegInB0[4] , 
        \wRegInB0[3] , \wRegInB0[2] , \wRegInB0[1] , \wRegInB0[0] }), .LoOut({
        \wRegInA1[31] , \wRegInA1[30] , \wRegInA1[29] , \wRegInA1[28] , 
        \wRegInA1[27] , \wRegInA1[26] , \wRegInA1[25] , \wRegInA1[24] , 
        \wRegInA1[23] , \wRegInA1[22] , \wRegInA1[21] , \wRegInA1[20] , 
        \wRegInA1[19] , \wRegInA1[18] , \wRegInA1[17] , \wRegInA1[16] , 
        \wRegInA1[15] , \wRegInA1[14] , \wRegInA1[13] , \wRegInA1[12] , 
        \wRegInA1[11] , \wRegInA1[10] , \wRegInA1[9] , \wRegInA1[8] , 
        \wRegInA1[7] , \wRegInA1[6] , \wRegInA1[5] , \wRegInA1[4] , 
        \wRegInA1[3] , \wRegInA1[2] , \wRegInA1[1] , \wRegInA1[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid16[31] , \wAMid16[30] , \wAMid16[29] , \wAMid16[28] , 
        \wAMid16[27] , \wAMid16[26] , \wAMid16[25] , \wAMid16[24] , 
        \wAMid16[23] , \wAMid16[22] , \wAMid16[21] , \wAMid16[20] , 
        \wAMid16[19] , \wAMid16[18] , \wAMid16[17] , \wAMid16[16] , 
        \wAMid16[15] , \wAMid16[14] , \wAMid16[13] , \wAMid16[12] , 
        \wAMid16[11] , \wAMid16[10] , \wAMid16[9] , \wAMid16[8] , \wAMid16[7] , 
        \wAMid16[6] , \wAMid16[5] , \wAMid16[4] , \wAMid16[3] , \wAMid16[2] , 
        \wAMid16[1] , \wAMid16[0] }), .BIn({\wBMid16[31] , \wBMid16[30] , 
        \wBMid16[29] , \wBMid16[28] , \wBMid16[27] , \wBMid16[26] , 
        \wBMid16[25] , \wBMid16[24] , \wBMid16[23] , \wBMid16[22] , 
        \wBMid16[21] , \wBMid16[20] , \wBMid16[19] , \wBMid16[18] , 
        \wBMid16[17] , \wBMid16[16] , \wBMid16[15] , \wBMid16[14] , 
        \wBMid16[13] , \wBMid16[12] , \wBMid16[11] , \wBMid16[10] , 
        \wBMid16[9] , \wBMid16[8] , \wBMid16[7] , \wBMid16[6] , \wBMid16[5] , 
        \wBMid16[4] , \wBMid16[3] , \wBMid16[2] , \wBMid16[1] , \wBMid16[0] }), 
        .HiOut({\wRegInB16[31] , \wRegInB16[30] , \wRegInB16[29] , 
        \wRegInB16[28] , \wRegInB16[27] , \wRegInB16[26] , \wRegInB16[25] , 
        \wRegInB16[24] , \wRegInB16[23] , \wRegInB16[22] , \wRegInB16[21] , 
        \wRegInB16[20] , \wRegInB16[19] , \wRegInB16[18] , \wRegInB16[17] , 
        \wRegInB16[16] , \wRegInB16[15] , \wRegInB16[14] , \wRegInB16[13] , 
        \wRegInB16[12] , \wRegInB16[11] , \wRegInB16[10] , \wRegInB16[9] , 
        \wRegInB16[8] , \wRegInB16[7] , \wRegInB16[6] , \wRegInB16[5] , 
        \wRegInB16[4] , \wRegInB16[3] , \wRegInB16[2] , \wRegInB16[1] , 
        \wRegInB16[0] }), .LoOut({\wRegInA17[31] , \wRegInA17[30] , 
        \wRegInA17[29] , \wRegInA17[28] , \wRegInA17[27] , \wRegInA17[26] , 
        \wRegInA17[25] , \wRegInA17[24] , \wRegInA17[23] , \wRegInA17[22] , 
        \wRegInA17[21] , \wRegInA17[20] , \wRegInA17[19] , \wRegInA17[18] , 
        \wRegInA17[17] , \wRegInA17[16] , \wRegInA17[15] , \wRegInA17[14] , 
        \wRegInA17[13] , \wRegInA17[12] , \wRegInA17[11] , \wRegInA17[10] , 
        \wRegInA17[9] , \wRegInA17[8] , \wRegInA17[7] , \wRegInA17[6] , 
        \wRegInA17[5] , \wRegInA17[4] , \wRegInA17[3] , \wRegInA17[2] , 
        \wRegInA17[1] , \wRegInA17[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_21 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink22[31] , \ScanLink22[30] , \ScanLink22[29] , 
        \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , \ScanLink22[25] , 
        \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , \ScanLink22[21] , 
        \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , \ScanLink22[17] , 
        \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , \ScanLink22[13] , 
        \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , \ScanLink22[9] , 
        \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , \ScanLink22[5] , 
        \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , \ScanLink22[1] , 
        \ScanLink22[0] }), .ScanOut({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA21[31] , \wRegInA21[30] , 
        \wRegInA21[29] , \wRegInA21[28] , \wRegInA21[27] , \wRegInA21[26] , 
        \wRegInA21[25] , \wRegInA21[24] , \wRegInA21[23] , \wRegInA21[22] , 
        \wRegInA21[21] , \wRegInA21[20] , \wRegInA21[19] , \wRegInA21[18] , 
        \wRegInA21[17] , \wRegInA21[16] , \wRegInA21[15] , \wRegInA21[14] , 
        \wRegInA21[13] , \wRegInA21[12] , \wRegInA21[11] , \wRegInA21[10] , 
        \wRegInA21[9] , \wRegInA21[8] , \wRegInA21[7] , \wRegInA21[6] , 
        \wRegInA21[5] , \wRegInA21[4] , \wRegInA21[3] , \wRegInA21[2] , 
        \wRegInA21[1] , \wRegInA21[0] }), .Out({\wAIn21[31] , \wAIn21[30] , 
        \wAIn21[29] , \wAIn21[28] , \wAIn21[27] , \wAIn21[26] , \wAIn21[25] , 
        \wAIn21[24] , \wAIn21[23] , \wAIn21[22] , \wAIn21[21] , \wAIn21[20] , 
        \wAIn21[19] , \wAIn21[18] , \wAIn21[17] , \wAIn21[16] , \wAIn21[15] , 
        \wAIn21[14] , \wAIn21[13] , \wAIn21[12] , \wAIn21[11] , \wAIn21[10] , 
        \wAIn21[9] , \wAIn21[8] , \wAIn21[7] , \wAIn21[6] , \wAIn21[5] , 
        \wAIn21[4] , \wAIn21[3] , \wAIn21[2] , \wAIn21[1] , \wAIn21[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_54 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink55[31] , \ScanLink55[30] , \ScanLink55[29] , 
        \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , \ScanLink55[25] , 
        \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , \ScanLink55[21] , 
        \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , \ScanLink55[17] , 
        \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , \ScanLink55[13] , 
        \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , \ScanLink55[9] , 
        \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , \ScanLink55[5] , 
        \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , \ScanLink55[1] , 
        \ScanLink55[0] }), .ScanOut({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB4[31] , \wRegInB4[30] , 
        \wRegInB4[29] , \wRegInB4[28] , \wRegInB4[27] , \wRegInB4[26] , 
        \wRegInB4[25] , \wRegInB4[24] , \wRegInB4[23] , \wRegInB4[22] , 
        \wRegInB4[21] , \wRegInB4[20] , \wRegInB4[19] , \wRegInB4[18] , 
        \wRegInB4[17] , \wRegInB4[16] , \wRegInB4[15] , \wRegInB4[14] , 
        \wRegInB4[13] , \wRegInB4[12] , \wRegInB4[11] , \wRegInB4[10] , 
        \wRegInB4[9] , \wRegInB4[8] , \wRegInB4[7] , \wRegInB4[6] , 
        \wRegInB4[5] , \wRegInB4[4] , \wRegInB4[3] , \wRegInB4[2] , 
        \wRegInB4[1] , \wRegInB4[0] }), .Out({\wBIn4[31] , \wBIn4[30] , 
        \wBIn4[29] , \wBIn4[28] , \wBIn4[27] , \wBIn4[26] , \wBIn4[25] , 
        \wBIn4[24] , \wBIn4[23] , \wBIn4[22] , \wBIn4[21] , \wBIn4[20] , 
        \wBIn4[19] , \wBIn4[18] , \wBIn4[17] , \wBIn4[16] , \wBIn4[15] , 
        \wBIn4[14] , \wBIn4[13] , \wBIn4[12] , \wBIn4[11] , \wBIn4[10] , 
        \wBIn4[9] , \wBIn4[8] , \wBIn4[7] , \wBIn4[6] , \wBIn4[5] , \wBIn4[4] , 
        \wBIn4[3] , \wBIn4[2] , \wBIn4[1] , \wBIn4[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn9[31] , 
        \wAIn9[30] , \wAIn9[29] , \wAIn9[28] , \wAIn9[27] , \wAIn9[26] , 
        \wAIn9[25] , \wAIn9[24] , \wAIn9[23] , \wAIn9[22] , \wAIn9[21] , 
        \wAIn9[20] , \wAIn9[19] , \wAIn9[18] , \wAIn9[17] , \wAIn9[16] , 
        \wAIn9[15] , \wAIn9[14] , \wAIn9[13] , \wAIn9[12] , \wAIn9[11] , 
        \wAIn9[10] , \wAIn9[9] , \wAIn9[8] , \wAIn9[7] , \wAIn9[6] , 
        \wAIn9[5] , \wAIn9[4] , \wAIn9[3] , \wAIn9[2] , \wAIn9[1] , \wAIn9[0] 
        }), .BIn({\wBIn9[31] , \wBIn9[30] , \wBIn9[29] , \wBIn9[28] , 
        \wBIn9[27] , \wBIn9[26] , \wBIn9[25] , \wBIn9[24] , \wBIn9[23] , 
        \wBIn9[22] , \wBIn9[21] , \wBIn9[20] , \wBIn9[19] , \wBIn9[18] , 
        \wBIn9[17] , \wBIn9[16] , \wBIn9[15] , \wBIn9[14] , \wBIn9[13] , 
        \wBIn9[12] , \wBIn9[11] , \wBIn9[10] , \wBIn9[9] , \wBIn9[8] , 
        \wBIn9[7] , \wBIn9[6] , \wBIn9[5] , \wBIn9[4] , \wBIn9[3] , \wBIn9[2] , 
        \wBIn9[1] , \wBIn9[0] }), .HiOut({\wBMid8[31] , \wBMid8[30] , 
        \wBMid8[29] , \wBMid8[28] , \wBMid8[27] , \wBMid8[26] , \wBMid8[25] , 
        \wBMid8[24] , \wBMid8[23] , \wBMid8[22] , \wBMid8[21] , \wBMid8[20] , 
        \wBMid8[19] , \wBMid8[18] , \wBMid8[17] , \wBMid8[16] , \wBMid8[15] , 
        \wBMid8[14] , \wBMid8[13] , \wBMid8[12] , \wBMid8[11] , \wBMid8[10] , 
        \wBMid8[9] , \wBMid8[8] , \wBMid8[7] , \wBMid8[6] , \wBMid8[5] , 
        \wBMid8[4] , \wBMid8[3] , \wBMid8[2] , \wBMid8[1] , \wBMid8[0] }), 
        .LoOut({\wAMid9[31] , \wAMid9[30] , \wAMid9[29] , \wAMid9[28] , 
        \wAMid9[27] , \wAMid9[26] , \wAMid9[25] , \wAMid9[24] , \wAMid9[23] , 
        \wAMid9[22] , \wAMid9[21] , \wAMid9[20] , \wAMid9[19] , \wAMid9[18] , 
        \wAMid9[17] , \wAMid9[16] , \wAMid9[15] , \wAMid9[14] , \wAMid9[13] , 
        \wAMid9[12] , \wAMid9[11] , \wAMid9[10] , \wAMid9[9] , \wAMid9[8] , 
        \wAMid9[7] , \wAMid9[6] , \wAMid9[5] , \wAMid9[4] , \wAMid9[3] , 
        \wAMid9[2] , \wAMid9[1] , \wAMid9[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn11[31] , \wAIn11[30] , \wAIn11[29] , \wAIn11[28] , \wAIn11[27] , 
        \wAIn11[26] , \wAIn11[25] , \wAIn11[24] , \wAIn11[23] , \wAIn11[22] , 
        \wAIn11[21] , \wAIn11[20] , \wAIn11[19] , \wAIn11[18] , \wAIn11[17] , 
        \wAIn11[16] , \wAIn11[15] , \wAIn11[14] , \wAIn11[13] , \wAIn11[12] , 
        \wAIn11[11] , \wAIn11[10] , \wAIn11[9] , \wAIn11[8] , \wAIn11[7] , 
        \wAIn11[6] , \wAIn11[5] , \wAIn11[4] , \wAIn11[3] , \wAIn11[2] , 
        \wAIn11[1] , \wAIn11[0] }), .BIn({\wBIn11[31] , \wBIn11[30] , 
        \wBIn11[29] , \wBIn11[28] , \wBIn11[27] , \wBIn11[26] , \wBIn11[25] , 
        \wBIn11[24] , \wBIn11[23] , \wBIn11[22] , \wBIn11[21] , \wBIn11[20] , 
        \wBIn11[19] , \wBIn11[18] , \wBIn11[17] , \wBIn11[16] , \wBIn11[15] , 
        \wBIn11[14] , \wBIn11[13] , \wBIn11[12] , \wBIn11[11] , \wBIn11[10] , 
        \wBIn11[9] , \wBIn11[8] , \wBIn11[7] , \wBIn11[6] , \wBIn11[5] , 
        \wBIn11[4] , \wBIn11[3] , \wBIn11[2] , \wBIn11[1] , \wBIn11[0] }), 
        .HiOut({\wBMid10[31] , \wBMid10[30] , \wBMid10[29] , \wBMid10[28] , 
        \wBMid10[27] , \wBMid10[26] , \wBMid10[25] , \wBMid10[24] , 
        \wBMid10[23] , \wBMid10[22] , \wBMid10[21] , \wBMid10[20] , 
        \wBMid10[19] , \wBMid10[18] , \wBMid10[17] , \wBMid10[16] , 
        \wBMid10[15] , \wBMid10[14] , \wBMid10[13] , \wBMid10[12] , 
        \wBMid10[11] , \wBMid10[10] , \wBMid10[9] , \wBMid10[8] , \wBMid10[7] , 
        \wBMid10[6] , \wBMid10[5] , \wBMid10[4] , \wBMid10[3] , \wBMid10[2] , 
        \wBMid10[1] , \wBMid10[0] }), .LoOut({\wAMid11[31] , \wAMid11[30] , 
        \wAMid11[29] , \wAMid11[28] , \wAMid11[27] , \wAMid11[26] , 
        \wAMid11[25] , \wAMid11[24] , \wAMid11[23] , \wAMid11[22] , 
        \wAMid11[21] , \wAMid11[20] , \wAMid11[19] , \wAMid11[18] , 
        \wAMid11[17] , \wAMid11[16] , \wAMid11[15] , \wAMid11[14] , 
        \wAMid11[13] , \wAMid11[12] , \wAMid11[11] , \wAMid11[10] , 
        \wAMid11[9] , \wAMid11[8] , \wAMid11[7] , \wAMid11[6] , \wAMid11[5] , 
        \wAMid11[4] , \wAMid11[3] , \wAMid11[2] , \wAMid11[1] , \wAMid11[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_31 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink32[31] , \ScanLink32[30] , \ScanLink32[29] , 
        \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , \ScanLink32[25] , 
        \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , \ScanLink32[21] , 
        \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , \ScanLink32[17] , 
        \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , \ScanLink32[13] , 
        \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , \ScanLink32[9] , 
        \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , \ScanLink32[5] , 
        \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , \ScanLink32[1] , 
        \ScanLink32[0] }), .ScanOut({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA16[31] , \wRegInA16[30] , 
        \wRegInA16[29] , \wRegInA16[28] , \wRegInA16[27] , \wRegInA16[26] , 
        \wRegInA16[25] , \wRegInA16[24] , \wRegInA16[23] , \wRegInA16[22] , 
        \wRegInA16[21] , \wRegInA16[20] , \wRegInA16[19] , \wRegInA16[18] , 
        \wRegInA16[17] , \wRegInA16[16] , \wRegInA16[15] , \wRegInA16[14] , 
        \wRegInA16[13] , \wRegInA16[12] , \wRegInA16[11] , \wRegInA16[10] , 
        \wRegInA16[9] , \wRegInA16[8] , \wRegInA16[7] , \wRegInA16[6] , 
        \wRegInA16[5] , \wRegInA16[4] , \wRegInA16[3] , \wRegInA16[2] , 
        \wRegInA16[1] , \wRegInA16[0] }), .Out({\wAIn16[31] , \wAIn16[30] , 
        \wAIn16[29] , \wAIn16[28] , \wAIn16[27] , \wAIn16[26] , \wAIn16[25] , 
        \wAIn16[24] , \wAIn16[23] , \wAIn16[22] , \wAIn16[21] , \wAIn16[20] , 
        \wAIn16[19] , \wAIn16[18] , \wAIn16[17] , \wAIn16[16] , \wAIn16[15] , 
        \wAIn16[14] , \wAIn16[13] , \wAIn16[12] , \wAIn16[11] , \wAIn16[10] , 
        \wAIn16[9] , \wAIn16[8] , \wAIn16[7] , \wAIn16[6] , \wAIn16[5] , 
        \wAIn16[4] , \wAIn16[3] , \wAIn16[2] , \wAIn16[1] , \wAIn16[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_16 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink17[31] , \ScanLink17[30] , \ScanLink17[29] , 
        \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , \ScanLink17[25] , 
        \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , \ScanLink17[21] , 
        \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , \ScanLink17[17] , 
        \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , \ScanLink17[13] , 
        \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , \ScanLink17[9] , 
        \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , \ScanLink17[5] , 
        \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , \ScanLink17[1] , 
        \ScanLink17[0] }), .ScanOut({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB23[31] , \wRegInB23[30] , 
        \wRegInB23[29] , \wRegInB23[28] , \wRegInB23[27] , \wRegInB23[26] , 
        \wRegInB23[25] , \wRegInB23[24] , \wRegInB23[23] , \wRegInB23[22] , 
        \wRegInB23[21] , \wRegInB23[20] , \wRegInB23[19] , \wRegInB23[18] , 
        \wRegInB23[17] , \wRegInB23[16] , \wRegInB23[15] , \wRegInB23[14] , 
        \wRegInB23[13] , \wRegInB23[12] , \wRegInB23[11] , \wRegInB23[10] , 
        \wRegInB23[9] , \wRegInB23[8] , \wRegInB23[7] , \wRegInB23[6] , 
        \wRegInB23[5] , \wRegInB23[4] , \wRegInB23[3] , \wRegInB23[2] , 
        \wRegInB23[1] , \wRegInB23[0] }), .Out({\wBIn23[31] , \wBIn23[30] , 
        \wBIn23[29] , \wBIn23[28] , \wBIn23[27] , \wBIn23[26] , \wBIn23[25] , 
        \wBIn23[24] , \wBIn23[23] , \wBIn23[22] , \wBIn23[21] , \wBIn23[20] , 
        \wBIn23[19] , \wBIn23[18] , \wBIn23[17] , \wBIn23[16] , \wBIn23[15] , 
        \wBIn23[14] , \wBIn23[13] , \wBIn23[12] , \wBIn23[11] , \wBIn23[10] , 
        \wBIn23[9] , \wBIn23[8] , \wBIn23[7] , \wBIn23[6] , \wBIn23[5] , 
        \wBIn23[4] , \wBIn23[3] , \wBIn23[2] , \wBIn23[1] , \wBIn23[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn18[31] , \wAIn18[30] , \wAIn18[29] , \wAIn18[28] , \wAIn18[27] , 
        \wAIn18[26] , \wAIn18[25] , \wAIn18[24] , \wAIn18[23] , \wAIn18[22] , 
        \wAIn18[21] , \wAIn18[20] , \wAIn18[19] , \wAIn18[18] , \wAIn18[17] , 
        \wAIn18[16] , \wAIn18[15] , \wAIn18[14] , \wAIn18[13] , \wAIn18[12] , 
        \wAIn18[11] , \wAIn18[10] , \wAIn18[9] , \wAIn18[8] , \wAIn18[7] , 
        \wAIn18[6] , \wAIn18[5] , \wAIn18[4] , \wAIn18[3] , \wAIn18[2] , 
        \wAIn18[1] , \wAIn18[0] }), .BIn({\wBIn18[31] , \wBIn18[30] , 
        \wBIn18[29] , \wBIn18[28] , \wBIn18[27] , \wBIn18[26] , \wBIn18[25] , 
        \wBIn18[24] , \wBIn18[23] , \wBIn18[22] , \wBIn18[21] , \wBIn18[20] , 
        \wBIn18[19] , \wBIn18[18] , \wBIn18[17] , \wBIn18[16] , \wBIn18[15] , 
        \wBIn18[14] , \wBIn18[13] , \wBIn18[12] , \wBIn18[11] , \wBIn18[10] , 
        \wBIn18[9] , \wBIn18[8] , \wBIn18[7] , \wBIn18[6] , \wBIn18[5] , 
        \wBIn18[4] , \wBIn18[3] , \wBIn18[2] , \wBIn18[1] , \wBIn18[0] }), 
        .HiOut({\wBMid17[31] , \wBMid17[30] , \wBMid17[29] , \wBMid17[28] , 
        \wBMid17[27] , \wBMid17[26] , \wBMid17[25] , \wBMid17[24] , 
        \wBMid17[23] , \wBMid17[22] , \wBMid17[21] , \wBMid17[20] , 
        \wBMid17[19] , \wBMid17[18] , \wBMid17[17] , \wBMid17[16] , 
        \wBMid17[15] , \wBMid17[14] , \wBMid17[13] , \wBMid17[12] , 
        \wBMid17[11] , \wBMid17[10] , \wBMid17[9] , \wBMid17[8] , \wBMid17[7] , 
        \wBMid17[6] , \wBMid17[5] , \wBMid17[4] , \wBMid17[3] , \wBMid17[2] , 
        \wBMid17[1] , \wBMid17[0] }), .LoOut({\wAMid18[31] , \wAMid18[30] , 
        \wAMid18[29] , \wAMid18[28] , \wAMid18[27] , \wAMid18[26] , 
        \wAMid18[25] , \wAMid18[24] , \wAMid18[23] , \wAMid18[22] , 
        \wAMid18[21] , \wAMid18[20] , \wAMid18[19] , \wAMid18[18] , 
        \wAMid18[17] , \wAMid18[16] , \wAMid18[15] , \wAMid18[14] , 
        \wAMid18[13] , \wAMid18[12] , \wAMid18[11] , \wAMid18[10] , 
        \wAMid18[9] , \wAMid18[8] , \wAMid18[7] , \wAMid18[6] , \wAMid18[5] , 
        \wAMid18[4] , \wAMid18[3] , \wAMid18[2] , \wAMid18[1] , \wAMid18[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn24[31] , \wAIn24[30] , \wAIn24[29] , \wAIn24[28] , \wAIn24[27] , 
        \wAIn24[26] , \wAIn24[25] , \wAIn24[24] , \wAIn24[23] , \wAIn24[22] , 
        \wAIn24[21] , \wAIn24[20] , \wAIn24[19] , \wAIn24[18] , \wAIn24[17] , 
        \wAIn24[16] , \wAIn24[15] , \wAIn24[14] , \wAIn24[13] , \wAIn24[12] , 
        \wAIn24[11] , \wAIn24[10] , \wAIn24[9] , \wAIn24[8] , \wAIn24[7] , 
        \wAIn24[6] , \wAIn24[5] , \wAIn24[4] , \wAIn24[3] , \wAIn24[2] , 
        \wAIn24[1] , \wAIn24[0] }), .BIn({\wBIn24[31] , \wBIn24[30] , 
        \wBIn24[29] , \wBIn24[28] , \wBIn24[27] , \wBIn24[26] , \wBIn24[25] , 
        \wBIn24[24] , \wBIn24[23] , \wBIn24[22] , \wBIn24[21] , \wBIn24[20] , 
        \wBIn24[19] , \wBIn24[18] , \wBIn24[17] , \wBIn24[16] , \wBIn24[15] , 
        \wBIn24[14] , \wBIn24[13] , \wBIn24[12] , \wBIn24[11] , \wBIn24[10] , 
        \wBIn24[9] , \wBIn24[8] , \wBIn24[7] , \wBIn24[6] , \wBIn24[5] , 
        \wBIn24[4] , \wBIn24[3] , \wBIn24[2] , \wBIn24[1] , \wBIn24[0] }), 
        .HiOut({\wBMid23[31] , \wBMid23[30] , \wBMid23[29] , \wBMid23[28] , 
        \wBMid23[27] , \wBMid23[26] , \wBMid23[25] , \wBMid23[24] , 
        \wBMid23[23] , \wBMid23[22] , \wBMid23[21] , \wBMid23[20] , 
        \wBMid23[19] , \wBMid23[18] , \wBMid23[17] , \wBMid23[16] , 
        \wBMid23[15] , \wBMid23[14] , \wBMid23[13] , \wBMid23[12] , 
        \wBMid23[11] , \wBMid23[10] , \wBMid23[9] , \wBMid23[8] , \wBMid23[7] , 
        \wBMid23[6] , \wBMid23[5] , \wBMid23[4] , \wBMid23[3] , \wBMid23[2] , 
        \wBMid23[1] , \wBMid23[0] }), .LoOut({\wAMid24[31] , \wAMid24[30] , 
        \wAMid24[29] , \wAMid24[28] , \wAMid24[27] , \wAMid24[26] , 
        \wAMid24[25] , \wAMid24[24] , \wAMid24[23] , \wAMid24[22] , 
        \wAMid24[21] , \wAMid24[20] , \wAMid24[19] , \wAMid24[18] , 
        \wAMid24[17] , \wAMid24[16] , \wAMid24[15] , \wAMid24[14] , 
        \wAMid24[13] , \wAMid24[12] , \wAMid24[11] , \wAMid24[10] , 
        \wAMid24[9] , \wAMid24[8] , \wAMid24[7] , \wAMid24[6] , \wAMid24[5] , 
        \wAMid24[4] , \wAMid24[3] , \wAMid24[2] , \wAMid24[1] , \wAMid24[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid21[31] , \wAMid21[30] , \wAMid21[29] , \wAMid21[28] , 
        \wAMid21[27] , \wAMid21[26] , \wAMid21[25] , \wAMid21[24] , 
        \wAMid21[23] , \wAMid21[22] , \wAMid21[21] , \wAMid21[20] , 
        \wAMid21[19] , \wAMid21[18] , \wAMid21[17] , \wAMid21[16] , 
        \wAMid21[15] , \wAMid21[14] , \wAMid21[13] , \wAMid21[12] , 
        \wAMid21[11] , \wAMid21[10] , \wAMid21[9] , \wAMid21[8] , \wAMid21[7] , 
        \wAMid21[6] , \wAMid21[5] , \wAMid21[4] , \wAMid21[3] , \wAMid21[2] , 
        \wAMid21[1] , \wAMid21[0] }), .BIn({\wBMid21[31] , \wBMid21[30] , 
        \wBMid21[29] , \wBMid21[28] , \wBMid21[27] , \wBMid21[26] , 
        \wBMid21[25] , \wBMid21[24] , \wBMid21[23] , \wBMid21[22] , 
        \wBMid21[21] , \wBMid21[20] , \wBMid21[19] , \wBMid21[18] , 
        \wBMid21[17] , \wBMid21[16] , \wBMid21[15] , \wBMid21[14] , 
        \wBMid21[13] , \wBMid21[12] , \wBMid21[11] , \wBMid21[10] , 
        \wBMid21[9] , \wBMid21[8] , \wBMid21[7] , \wBMid21[6] , \wBMid21[5] , 
        \wBMid21[4] , \wBMid21[3] , \wBMid21[2] , \wBMid21[1] , \wBMid21[0] }), 
        .HiOut({\wRegInB21[31] , \wRegInB21[30] , \wRegInB21[29] , 
        \wRegInB21[28] , \wRegInB21[27] , \wRegInB21[26] , \wRegInB21[25] , 
        \wRegInB21[24] , \wRegInB21[23] , \wRegInB21[22] , \wRegInB21[21] , 
        \wRegInB21[20] , \wRegInB21[19] , \wRegInB21[18] , \wRegInB21[17] , 
        \wRegInB21[16] , \wRegInB21[15] , \wRegInB21[14] , \wRegInB21[13] , 
        \wRegInB21[12] , \wRegInB21[11] , \wRegInB21[10] , \wRegInB21[9] , 
        \wRegInB21[8] , \wRegInB21[7] , \wRegInB21[6] , \wRegInB21[5] , 
        \wRegInB21[4] , \wRegInB21[3] , \wRegInB21[2] , \wRegInB21[1] , 
        \wRegInB21[0] }), .LoOut({\wRegInA22[31] , \wRegInA22[30] , 
        \wRegInA22[29] , \wRegInA22[28] , \wRegInA22[27] , \wRegInA22[26] , 
        \wRegInA22[25] , \wRegInA22[24] , \wRegInA22[23] , \wRegInA22[22] , 
        \wRegInA22[21] , \wRegInA22[20] , \wRegInA22[19] , \wRegInA22[18] , 
        \wRegInA22[17] , \wRegInA22[16] , \wRegInA22[15] , \wRegInA22[14] , 
        \wRegInA22[13] , \wRegInA22[12] , \wRegInA22[11] , \wRegInA22[10] , 
        \wRegInA22[9] , \wRegInA22[8] , \wRegInA22[7] , \wRegInA22[6] , 
        \wRegInA22[5] , \wRegInA22[4] , \wRegInA22[3] , \wRegInA22[2] , 
        \wRegInA22[1] , \wRegInA22[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_44 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink45[31] , \ScanLink45[30] , \ScanLink45[29] , 
        \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , \ScanLink45[25] , 
        \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , \ScanLink45[21] , 
        \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , \ScanLink45[17] , 
        \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , \ScanLink45[13] , 
        \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , \ScanLink45[9] , 
        \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , \ScanLink45[5] , 
        \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , \ScanLink45[1] , 
        \ScanLink45[0] }), .ScanOut({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB9[31] , \wRegInB9[30] , 
        \wRegInB9[29] , \wRegInB9[28] , \wRegInB9[27] , \wRegInB9[26] , 
        \wRegInB9[25] , \wRegInB9[24] , \wRegInB9[23] , \wRegInB9[22] , 
        \wRegInB9[21] , \wRegInB9[20] , \wRegInB9[19] , \wRegInB9[18] , 
        \wRegInB9[17] , \wRegInB9[16] , \wRegInB9[15] , \wRegInB9[14] , 
        \wRegInB9[13] , \wRegInB9[12] , \wRegInB9[11] , \wRegInB9[10] , 
        \wRegInB9[9] , \wRegInB9[8] , \wRegInB9[7] , \wRegInB9[6] , 
        \wRegInB9[5] , \wRegInB9[4] , \wRegInB9[3] , \wRegInB9[2] , 
        \wRegInB9[1] , \wRegInB9[0] }), .Out({\wBIn9[31] , \wBIn9[30] , 
        \wBIn9[29] , \wBIn9[28] , \wBIn9[27] , \wBIn9[26] , \wBIn9[25] , 
        \wBIn9[24] , \wBIn9[23] , \wBIn9[22] , \wBIn9[21] , \wBIn9[20] , 
        \wBIn9[19] , \wBIn9[18] , \wBIn9[17] , \wBIn9[16] , \wBIn9[15] , 
        \wBIn9[14] , \wBIn9[13] , \wBIn9[12] , \wBIn9[11] , \wBIn9[10] , 
        \wBIn9[9] , \wBIn9[8] , \wBIn9[7] , \wBIn9[6] , \wBIn9[5] , \wBIn9[4] , 
        \wBIn9[3] , \wBIn9[2] , \wBIn9[1] , \wBIn9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_63 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink64[31] , \ScanLink64[30] , \ScanLink64[29] , 
        \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , \ScanLink64[25] , 
        \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , \ScanLink64[21] , 
        \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , \ScanLink64[17] , 
        \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , \ScanLink64[13] , 
        \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , \ScanLink64[9] , 
        \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , \ScanLink64[5] , 
        \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , \ScanLink64[1] , 
        \ScanLink64[0] }), .ScanOut({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA0[31] , \wRegInA0[30] , 
        \wRegInA0[29] , \wRegInA0[28] , \wRegInA0[27] , \wRegInA0[26] , 
        \wRegInA0[25] , \wRegInA0[24] , \wRegInA0[23] , \wRegInA0[22] , 
        \wRegInA0[21] , \wRegInA0[20] , \wRegInA0[19] , \wRegInA0[18] , 
        \wRegInA0[17] , \wRegInA0[16] , \wRegInA0[15] , \wRegInA0[14] , 
        \wRegInA0[13] , \wRegInA0[12] , \wRegInA0[11] , \wRegInA0[10] , 
        \wRegInA0[9] , \wRegInA0[8] , \wRegInA0[7] , \wRegInA0[6] , 
        \wRegInA0[5] , \wRegInA0[4] , \wRegInA0[3] , \wRegInA0[2] , 
        \wRegInA0[1] , \wRegInA0[0] }), .Out({\wAIn0[31] , \wAIn0[30] , 
        \wAIn0[29] , \wAIn0[28] , \wAIn0[27] , \wAIn0[26] , \wAIn0[25] , 
        \wAIn0[24] , \wAIn0[23] , \wAIn0[22] , \wAIn0[21] , \wAIn0[20] , 
        \wAIn0[19] , \wAIn0[18] , \wAIn0[17] , \wAIn0[16] , \wAIn0[15] , 
        \wAIn0[14] , \wAIn0[13] , \wAIn0[12] , \wAIn0[11] , \wAIn0[10] , 
        \wAIn0[9] , \wAIn0[8] , \wAIn0[7] , \wAIn0[6] , \wAIn0[5] , \wAIn0[4] , 
        \wAIn0[3] , \wAIn0[2] , \wAIn0[1] , \wAIn0[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_7 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[31] , \ScanLink8[30] , \ScanLink8[29] , 
        \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , \ScanLink8[25] , 
        \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , \ScanLink8[21] , 
        \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , \ScanLink8[17] , 
        \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , \ScanLink8[13] , 
        \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , \ScanLink8[9] , 
        \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA28[31] , \wRegInA28[30] , 
        \wRegInA28[29] , \wRegInA28[28] , \wRegInA28[27] , \wRegInA28[26] , 
        \wRegInA28[25] , \wRegInA28[24] , \wRegInA28[23] , \wRegInA28[22] , 
        \wRegInA28[21] , \wRegInA28[20] , \wRegInA28[19] , \wRegInA28[18] , 
        \wRegInA28[17] , \wRegInA28[16] , \wRegInA28[15] , \wRegInA28[14] , 
        \wRegInA28[13] , \wRegInA28[12] , \wRegInA28[11] , \wRegInA28[10] , 
        \wRegInA28[9] , \wRegInA28[8] , \wRegInA28[7] , \wRegInA28[6] , 
        \wRegInA28[5] , \wRegInA28[4] , \wRegInA28[3] , \wRegInA28[2] , 
        \wRegInA28[1] , \wRegInA28[0] }), .Out({\wAIn28[31] , \wAIn28[30] , 
        \wAIn28[29] , \wAIn28[28] , \wAIn28[27] , \wAIn28[26] , \wAIn28[25] , 
        \wAIn28[24] , \wAIn28[23] , \wAIn28[22] , \wAIn28[21] , \wAIn28[20] , 
        \wAIn28[19] , \wAIn28[18] , \wAIn28[17] , \wAIn28[16] , \wAIn28[15] , 
        \wAIn28[14] , \wAIn28[13] , \wAIn28[12] , \wAIn28[11] , \wAIn28[10] , 
        \wAIn28[9] , \wAIn28[8] , \wAIn28[7] , \wAIn28[6] , \wAIn28[5] , 
        \wAIn28[4] , \wAIn28[3] , \wAIn28[2] , \wAIn28[1] , \wAIn28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_56 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink57[31] , \ScanLink57[30] , \ScanLink57[29] , 
        \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , \ScanLink57[25] , 
        \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , \ScanLink57[21] , 
        \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , \ScanLink57[17] , 
        \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , \ScanLink57[13] , 
        \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , \ScanLink57[9] , 
        \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , \ScanLink57[5] , 
        \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , \ScanLink57[1] , 
        \ScanLink57[0] }), .ScanOut({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB3[31] , \wRegInB3[30] , 
        \wRegInB3[29] , \wRegInB3[28] , \wRegInB3[27] , \wRegInB3[26] , 
        \wRegInB3[25] , \wRegInB3[24] , \wRegInB3[23] , \wRegInB3[22] , 
        \wRegInB3[21] , \wRegInB3[20] , \wRegInB3[19] , \wRegInB3[18] , 
        \wRegInB3[17] , \wRegInB3[16] , \wRegInB3[15] , \wRegInB3[14] , 
        \wRegInB3[13] , \wRegInB3[12] , \wRegInB3[11] , \wRegInB3[10] , 
        \wRegInB3[9] , \wRegInB3[8] , \wRegInB3[7] , \wRegInB3[6] , 
        \wRegInB3[5] , \wRegInB3[4] , \wRegInB3[3] , \wRegInB3[2] , 
        \wRegInB3[1] , \wRegInB3[0] }), .Out({\wBIn3[31] , \wBIn3[30] , 
        \wBIn3[29] , \wBIn3[28] , \wBIn3[27] , \wBIn3[26] , \wBIn3[25] , 
        \wBIn3[24] , \wBIn3[23] , \wBIn3[22] , \wBIn3[21] , \wBIn3[20] , 
        \wBIn3[19] , \wBIn3[18] , \wBIn3[17] , \wBIn3[16] , \wBIn3[15] , 
        \wBIn3[14] , \wBIn3[13] , \wBIn3[12] , \wBIn3[11] , \wBIn3[10] , 
        \wBIn3[9] , \wBIn3[8] , \wBIn3[7] , \wBIn3[6] , \wBIn3[5] , \wBIn3[4] , 
        \wBIn3[3] , \wBIn3[2] , \wBIn3[1] , \wBIn3[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid14[31] , \wAMid14[30] , \wAMid14[29] , \wAMid14[28] , 
        \wAMid14[27] , \wAMid14[26] , \wAMid14[25] , \wAMid14[24] , 
        \wAMid14[23] , \wAMid14[22] , \wAMid14[21] , \wAMid14[20] , 
        \wAMid14[19] , \wAMid14[18] , \wAMid14[17] , \wAMid14[16] , 
        \wAMid14[15] , \wAMid14[14] , \wAMid14[13] , \wAMid14[12] , 
        \wAMid14[11] , \wAMid14[10] , \wAMid14[9] , \wAMid14[8] , \wAMid14[7] , 
        \wAMid14[6] , \wAMid14[5] , \wAMid14[4] , \wAMid14[3] , \wAMid14[2] , 
        \wAMid14[1] , \wAMid14[0] }), .BIn({\wBMid14[31] , \wBMid14[30] , 
        \wBMid14[29] , \wBMid14[28] , \wBMid14[27] , \wBMid14[26] , 
        \wBMid14[25] , \wBMid14[24] , \wBMid14[23] , \wBMid14[22] , 
        \wBMid14[21] , \wBMid14[20] , \wBMid14[19] , \wBMid14[18] , 
        \wBMid14[17] , \wBMid14[16] , \wBMid14[15] , \wBMid14[14] , 
        \wBMid14[13] , \wBMid14[12] , \wBMid14[11] , \wBMid14[10] , 
        \wBMid14[9] , \wBMid14[8] , \wBMid14[7] , \wBMid14[6] , \wBMid14[5] , 
        \wBMid14[4] , \wBMid14[3] , \wBMid14[2] , \wBMid14[1] , \wBMid14[0] }), 
        .HiOut({\wRegInB14[31] , \wRegInB14[30] , \wRegInB14[29] , 
        \wRegInB14[28] , \wRegInB14[27] , \wRegInB14[26] , \wRegInB14[25] , 
        \wRegInB14[24] , \wRegInB14[23] , \wRegInB14[22] , \wRegInB14[21] , 
        \wRegInB14[20] , \wRegInB14[19] , \wRegInB14[18] , \wRegInB14[17] , 
        \wRegInB14[16] , \wRegInB14[15] , \wRegInB14[14] , \wRegInB14[13] , 
        \wRegInB14[12] , \wRegInB14[11] , \wRegInB14[10] , \wRegInB14[9] , 
        \wRegInB14[8] , \wRegInB14[7] , \wRegInB14[6] , \wRegInB14[5] , 
        \wRegInB14[4] , \wRegInB14[3] , \wRegInB14[2] , \wRegInB14[1] , 
        \wRegInB14[0] }), .LoOut({\wRegInA15[31] , \wRegInA15[30] , 
        \wRegInA15[29] , \wRegInA15[28] , \wRegInA15[27] , \wRegInA15[26] , 
        \wRegInA15[25] , \wRegInA15[24] , \wRegInA15[23] , \wRegInA15[22] , 
        \wRegInA15[21] , \wRegInA15[20] , \wRegInA15[19] , \wRegInA15[18] , 
        \wRegInA15[17] , \wRegInA15[16] , \wRegInA15[15] , \wRegInA15[14] , 
        \wRegInA15[13] , \wRegInA15[12] , \wRegInA15[11] , \wRegInA15[10] , 
        \wRegInA15[9] , \wRegInA15[8] , \wRegInA15[7] , \wRegInA15[6] , 
        \wRegInA15[5] , \wRegInA15[4] , \wRegInA15[3] , \wRegInA15[2] , 
        \wRegInA15[1] , \wRegInA15[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid28[31] , \wAMid28[30] , \wAMid28[29] , \wAMid28[28] , 
        \wAMid28[27] , \wAMid28[26] , \wAMid28[25] , \wAMid28[24] , 
        \wAMid28[23] , \wAMid28[22] , \wAMid28[21] , \wAMid28[20] , 
        \wAMid28[19] , \wAMid28[18] , \wAMid28[17] , \wAMid28[16] , 
        \wAMid28[15] , \wAMid28[14] , \wAMid28[13] , \wAMid28[12] , 
        \wAMid28[11] , \wAMid28[10] , \wAMid28[9] , \wAMid28[8] , \wAMid28[7] , 
        \wAMid28[6] , \wAMid28[5] , \wAMid28[4] , \wAMid28[3] , \wAMid28[2] , 
        \wAMid28[1] , \wAMid28[0] }), .BIn({\wBMid28[31] , \wBMid28[30] , 
        \wBMid28[29] , \wBMid28[28] , \wBMid28[27] , \wBMid28[26] , 
        \wBMid28[25] , \wBMid28[24] , \wBMid28[23] , \wBMid28[22] , 
        \wBMid28[21] , \wBMid28[20] , \wBMid28[19] , \wBMid28[18] , 
        \wBMid28[17] , \wBMid28[16] , \wBMid28[15] , \wBMid28[14] , 
        \wBMid28[13] , \wBMid28[12] , \wBMid28[11] , \wBMid28[10] , 
        \wBMid28[9] , \wBMid28[8] , \wBMid28[7] , \wBMid28[6] , \wBMid28[5] , 
        \wBMid28[4] , \wBMid28[3] , \wBMid28[2] , \wBMid28[1] , \wBMid28[0] }), 
        .HiOut({\wRegInB28[31] , \wRegInB28[30] , \wRegInB28[29] , 
        \wRegInB28[28] , \wRegInB28[27] , \wRegInB28[26] , \wRegInB28[25] , 
        \wRegInB28[24] , \wRegInB28[23] , \wRegInB28[22] , \wRegInB28[21] , 
        \wRegInB28[20] , \wRegInB28[19] , \wRegInB28[18] , \wRegInB28[17] , 
        \wRegInB28[16] , \wRegInB28[15] , \wRegInB28[14] , \wRegInB28[13] , 
        \wRegInB28[12] , \wRegInB28[11] , \wRegInB28[10] , \wRegInB28[9] , 
        \wRegInB28[8] , \wRegInB28[7] , \wRegInB28[6] , \wRegInB28[5] , 
        \wRegInB28[4] , \wRegInB28[3] , \wRegInB28[2] , \wRegInB28[1] , 
        \wRegInB28[0] }), .LoOut({\wRegInA29[31] , \wRegInA29[30] , 
        \wRegInA29[29] , \wRegInA29[28] , \wRegInA29[27] , \wRegInA29[26] , 
        \wRegInA29[25] , \wRegInA29[24] , \wRegInA29[23] , \wRegInA29[22] , 
        \wRegInA29[21] , \wRegInA29[20] , \wRegInA29[19] , \wRegInA29[18] , 
        \wRegInA29[17] , \wRegInA29[16] , \wRegInA29[15] , \wRegInA29[14] , 
        \wRegInA29[13] , \wRegInA29[12] , \wRegInA29[11] , \wRegInA29[10] , 
        \wRegInA29[9] , \wRegInA29[8] , \wRegInA29[7] , \wRegInA29[6] , 
        \wRegInA29[5] , \wRegInA29[4] , \wRegInA29[3] , \wRegInA29[2] , 
        \wRegInA29[1] , \wRegInA29[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_38 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink39[31] , \ScanLink39[30] , \ScanLink39[29] , 
        \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , \ScanLink39[25] , 
        \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , \ScanLink39[21] , 
        \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , \ScanLink39[17] , 
        \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , \ScanLink39[13] , 
        \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , \ScanLink39[9] , 
        \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , \ScanLink39[5] , 
        \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , \ScanLink39[1] , 
        \ScanLink39[0] }), .ScanOut({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB12[31] , \wRegInB12[30] , 
        \wRegInB12[29] , \wRegInB12[28] , \wRegInB12[27] , \wRegInB12[26] , 
        \wRegInB12[25] , \wRegInB12[24] , \wRegInB12[23] , \wRegInB12[22] , 
        \wRegInB12[21] , \wRegInB12[20] , \wRegInB12[19] , \wRegInB12[18] , 
        \wRegInB12[17] , \wRegInB12[16] , \wRegInB12[15] , \wRegInB12[14] , 
        \wRegInB12[13] , \wRegInB12[12] , \wRegInB12[11] , \wRegInB12[10] , 
        \wRegInB12[9] , \wRegInB12[8] , \wRegInB12[7] , \wRegInB12[6] , 
        \wRegInB12[5] , \wRegInB12[4] , \wRegInB12[3] , \wRegInB12[2] , 
        \wRegInB12[1] , \wRegInB12[0] }), .Out({\wBIn12[31] , \wBIn12[30] , 
        \wBIn12[29] , \wBIn12[28] , \wBIn12[27] , \wBIn12[26] , \wBIn12[25] , 
        \wBIn12[24] , \wBIn12[23] , \wBIn12[22] , \wBIn12[21] , \wBIn12[20] , 
        \wBIn12[19] , \wBIn12[18] , \wBIn12[17] , \wBIn12[16] , \wBIn12[15] , 
        \wBIn12[14] , \wBIn12[13] , \wBIn12[12] , \wBIn12[11] , \wBIn12[10] , 
        \wBIn12[9] , \wBIn12[8] , \wBIn12[7] , \wBIn12[6] , \wBIn12[5] , 
        \wBIn12[4] , \wBIn12[3] , \wBIn12[2] , \wBIn12[1] , \wBIn12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_23 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink24[31] , \ScanLink24[30] , \ScanLink24[29] , 
        \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , \ScanLink24[25] , 
        \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , \ScanLink24[21] , 
        \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , \ScanLink24[17] , 
        \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , \ScanLink24[13] , 
        \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , \ScanLink24[9] , 
        \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , \ScanLink24[5] , 
        \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , \ScanLink24[1] , 
        \ScanLink24[0] }), .ScanOut({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA20[31] , \wRegInA20[30] , 
        \wRegInA20[29] , \wRegInA20[28] , \wRegInA20[27] , \wRegInA20[26] , 
        \wRegInA20[25] , \wRegInA20[24] , \wRegInA20[23] , \wRegInA20[22] , 
        \wRegInA20[21] , \wRegInA20[20] , \wRegInA20[19] , \wRegInA20[18] , 
        \wRegInA20[17] , \wRegInA20[16] , \wRegInA20[15] , \wRegInA20[14] , 
        \wRegInA20[13] , \wRegInA20[12] , \wRegInA20[11] , \wRegInA20[10] , 
        \wRegInA20[9] , \wRegInA20[8] , \wRegInA20[7] , \wRegInA20[6] , 
        \wRegInA20[5] , \wRegInA20[4] , \wRegInA20[3] , \wRegInA20[2] , 
        \wRegInA20[1] , \wRegInA20[0] }), .Out({\wAIn20[31] , \wAIn20[30] , 
        \wAIn20[29] , \wAIn20[28] , \wAIn20[27] , \wAIn20[26] , \wAIn20[25] , 
        \wAIn20[24] , \wAIn20[23] , \wAIn20[22] , \wAIn20[21] , \wAIn20[20] , 
        \wAIn20[19] , \wAIn20[18] , \wAIn20[17] , \wAIn20[16] , \wAIn20[15] , 
        \wAIn20[14] , \wAIn20[13] , \wAIn20[12] , \wAIn20[11] , \wAIn20[10] , 
        \wAIn20[9] , \wAIn20[8] , \wAIn20[7] , \wAIn20[6] , \wAIn20[5] , 
        \wAIn20[4] , \wAIn20[3] , \wAIn20[2] , \wAIn20[1] , \wAIn20[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid2[31] , 
        \wAMid2[30] , \wAMid2[29] , \wAMid2[28] , \wAMid2[27] , \wAMid2[26] , 
        \wAMid2[25] , \wAMid2[24] , \wAMid2[23] , \wAMid2[22] , \wAMid2[21] , 
        \wAMid2[20] , \wAMid2[19] , \wAMid2[18] , \wAMid2[17] , \wAMid2[16] , 
        \wAMid2[15] , \wAMid2[14] , \wAMid2[13] , \wAMid2[12] , \wAMid2[11] , 
        \wAMid2[10] , \wAMid2[9] , \wAMid2[8] , \wAMid2[7] , \wAMid2[6] , 
        \wAMid2[5] , \wAMid2[4] , \wAMid2[3] , \wAMid2[2] , \wAMid2[1] , 
        \wAMid2[0] }), .BIn({\wBMid2[31] , \wBMid2[30] , \wBMid2[29] , 
        \wBMid2[28] , \wBMid2[27] , \wBMid2[26] , \wBMid2[25] , \wBMid2[24] , 
        \wBMid2[23] , \wBMid2[22] , \wBMid2[21] , \wBMid2[20] , \wBMid2[19] , 
        \wBMid2[18] , \wBMid2[17] , \wBMid2[16] , \wBMid2[15] , \wBMid2[14] , 
        \wBMid2[13] , \wBMid2[12] , \wBMid2[11] , \wBMid2[10] , \wBMid2[9] , 
        \wBMid2[8] , \wBMid2[7] , \wBMid2[6] , \wBMid2[5] , \wBMid2[4] , 
        \wBMid2[3] , \wBMid2[2] , \wBMid2[1] , \wBMid2[0] }), .HiOut({
        \wRegInB2[31] , \wRegInB2[30] , \wRegInB2[29] , \wRegInB2[28] , 
        \wRegInB2[27] , \wRegInB2[26] , \wRegInB2[25] , \wRegInB2[24] , 
        \wRegInB2[23] , \wRegInB2[22] , \wRegInB2[21] , \wRegInB2[20] , 
        \wRegInB2[19] , \wRegInB2[18] , \wRegInB2[17] , \wRegInB2[16] , 
        \wRegInB2[15] , \wRegInB2[14] , \wRegInB2[13] , \wRegInB2[12] , 
        \wRegInB2[11] , \wRegInB2[10] , \wRegInB2[9] , \wRegInB2[8] , 
        \wRegInB2[7] , \wRegInB2[6] , \wRegInB2[5] , \wRegInB2[4] , 
        \wRegInB2[3] , \wRegInB2[2] , \wRegInB2[1] , \wRegInB2[0] }), .LoOut({
        \wRegInA3[31] , \wRegInA3[30] , \wRegInA3[29] , \wRegInA3[28] , 
        \wRegInA3[27] , \wRegInA3[26] , \wRegInA3[25] , \wRegInA3[24] , 
        \wRegInA3[23] , \wRegInA3[22] , \wRegInA3[21] , \wRegInA3[20] , 
        \wRegInA3[19] , \wRegInA3[18] , \wRegInA3[17] , \wRegInA3[16] , 
        \wRegInA3[15] , \wRegInA3[14] , \wRegInA3[13] , \wRegInA3[12] , 
        \wRegInA3[11] , \wRegInA3[10] , \wRegInA3[9] , \wRegInA3[8] , 
        \wRegInA3[7] , \wRegInA3[6] , \wRegInA3[5] , \wRegInA3[4] , 
        \wRegInA3[3] , \wRegInA3[2] , \wRegInA3[1] , \wRegInA3[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid5[31] , 
        \wAMid5[30] , \wAMid5[29] , \wAMid5[28] , \wAMid5[27] , \wAMid5[26] , 
        \wAMid5[25] , \wAMid5[24] , \wAMid5[23] , \wAMid5[22] , \wAMid5[21] , 
        \wAMid5[20] , \wAMid5[19] , \wAMid5[18] , \wAMid5[17] , \wAMid5[16] , 
        \wAMid5[15] , \wAMid5[14] , \wAMid5[13] , \wAMid5[12] , \wAMid5[11] , 
        \wAMid5[10] , \wAMid5[9] , \wAMid5[8] , \wAMid5[7] , \wAMid5[6] , 
        \wAMid5[5] , \wAMid5[4] , \wAMid5[3] , \wAMid5[2] , \wAMid5[1] , 
        \wAMid5[0] }), .BIn({\wBMid5[31] , \wBMid5[30] , \wBMid5[29] , 
        \wBMid5[28] , \wBMid5[27] , \wBMid5[26] , \wBMid5[25] , \wBMid5[24] , 
        \wBMid5[23] , \wBMid5[22] , \wBMid5[21] , \wBMid5[20] , \wBMid5[19] , 
        \wBMid5[18] , \wBMid5[17] , \wBMid5[16] , \wBMid5[15] , \wBMid5[14] , 
        \wBMid5[13] , \wBMid5[12] , \wBMid5[11] , \wBMid5[10] , \wBMid5[9] , 
        \wBMid5[8] , \wBMid5[7] , \wBMid5[6] , \wBMid5[5] , \wBMid5[4] , 
        \wBMid5[3] , \wBMid5[2] , \wBMid5[1] , \wBMid5[0] }), .HiOut({
        \wRegInB5[31] , \wRegInB5[30] , \wRegInB5[29] , \wRegInB5[28] , 
        \wRegInB5[27] , \wRegInB5[26] , \wRegInB5[25] , \wRegInB5[24] , 
        \wRegInB5[23] , \wRegInB5[22] , \wRegInB5[21] , \wRegInB5[20] , 
        \wRegInB5[19] , \wRegInB5[18] , \wRegInB5[17] , \wRegInB5[16] , 
        \wRegInB5[15] , \wRegInB5[14] , \wRegInB5[13] , \wRegInB5[12] , 
        \wRegInB5[11] , \wRegInB5[10] , \wRegInB5[9] , \wRegInB5[8] , 
        \wRegInB5[7] , \wRegInB5[6] , \wRegInB5[5] , \wRegInB5[4] , 
        \wRegInB5[3] , \wRegInB5[2] , \wRegInB5[1] , \wRegInB5[0] }), .LoOut({
        \wRegInA6[31] , \wRegInA6[30] , \wRegInA6[29] , \wRegInA6[28] , 
        \wRegInA6[27] , \wRegInA6[26] , \wRegInA6[25] , \wRegInA6[24] , 
        \wRegInA6[23] , \wRegInA6[22] , \wRegInA6[21] , \wRegInA6[20] , 
        \wRegInA6[19] , \wRegInA6[18] , \wRegInA6[17] , \wRegInA6[16] , 
        \wRegInA6[15] , \wRegInA6[14] , \wRegInA6[13] , \wRegInA6[12] , 
        \wRegInA6[11] , \wRegInA6[10] , \wRegInA6[9] , \wRegInA6[8] , 
        \wRegInA6[7] , \wRegInA6[6] , \wRegInA6[5] , \wRegInA6[4] , 
        \wRegInA6[3] , \wRegInA6[2] , \wRegInA6[1] , \wRegInA6[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_9 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[31] , \ScanLink10[30] , \ScanLink10[29] , 
        \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , \ScanLink10[25] , 
        \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , \ScanLink10[21] , 
        \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , \ScanLink10[17] , 
        \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , \ScanLink10[13] , 
        \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , \ScanLink10[9] , 
        \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA27[31] , \wRegInA27[30] , 
        \wRegInA27[29] , \wRegInA27[28] , \wRegInA27[27] , \wRegInA27[26] , 
        \wRegInA27[25] , \wRegInA27[24] , \wRegInA27[23] , \wRegInA27[22] , 
        \wRegInA27[21] , \wRegInA27[20] , \wRegInA27[19] , \wRegInA27[18] , 
        \wRegInA27[17] , \wRegInA27[16] , \wRegInA27[15] , \wRegInA27[14] , 
        \wRegInA27[13] , \wRegInA27[12] , \wRegInA27[11] , \wRegInA27[10] , 
        \wRegInA27[9] , \wRegInA27[8] , \wRegInA27[7] , \wRegInA27[6] , 
        \wRegInA27[5] , \wRegInA27[4] , \wRegInA27[3] , \wRegInA27[2] , 
        \wRegInA27[1] , \wRegInA27[0] }), .Out({\wAIn27[31] , \wAIn27[30] , 
        \wAIn27[29] , \wAIn27[28] , \wAIn27[27] , \wAIn27[26] , \wAIn27[25] , 
        \wAIn27[24] , \wAIn27[23] , \wAIn27[22] , \wAIn27[21] , \wAIn27[20] , 
        \wAIn27[19] , \wAIn27[18] , \wAIn27[17] , \wAIn27[16] , \wAIn27[15] , 
        \wAIn27[14] , \wAIn27[13] , \wAIn27[12] , \wAIn27[11] , \wAIn27[10] , 
        \wAIn27[9] , \wAIn27[8] , \wAIn27[7] , \wAIn27[6] , \wAIn27[5] , 
        \wAIn27[4] , \wAIn27[3] , \wAIn27[2] , \wAIn27[1] , \wAIn27[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_24 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink25[31] , \ScanLink25[30] , \ScanLink25[29] , 
        \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , \ScanLink25[25] , 
        \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , \ScanLink25[21] , 
        \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , \ScanLink25[17] , 
        \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , \ScanLink25[13] , 
        \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , \ScanLink25[9] , 
        \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , \ScanLink25[5] , 
        \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , \ScanLink25[1] , 
        \ScanLink25[0] }), .ScanOut({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB19[31] , \wRegInB19[30] , 
        \wRegInB19[29] , \wRegInB19[28] , \wRegInB19[27] , \wRegInB19[26] , 
        \wRegInB19[25] , \wRegInB19[24] , \wRegInB19[23] , \wRegInB19[22] , 
        \wRegInB19[21] , \wRegInB19[20] , \wRegInB19[19] , \wRegInB19[18] , 
        \wRegInB19[17] , \wRegInB19[16] , \wRegInB19[15] , \wRegInB19[14] , 
        \wRegInB19[13] , \wRegInB19[12] , \wRegInB19[11] , \wRegInB19[10] , 
        \wRegInB19[9] , \wRegInB19[8] , \wRegInB19[7] , \wRegInB19[6] , 
        \wRegInB19[5] , \wRegInB19[4] , \wRegInB19[3] , \wRegInB19[2] , 
        \wRegInB19[1] , \wRegInB19[0] }), .Out({\wBIn19[31] , \wBIn19[30] , 
        \wBIn19[29] , \wBIn19[28] , \wBIn19[27] , \wBIn19[26] , \wBIn19[25] , 
        \wBIn19[24] , \wBIn19[23] , \wBIn19[22] , \wBIn19[21] , \wBIn19[20] , 
        \wBIn19[19] , \wBIn19[18] , \wBIn19[17] , \wBIn19[16] , \wBIn19[15] , 
        \wBIn19[14] , \wBIn19[13] , \wBIn19[12] , \wBIn19[11] , \wBIn19[10] , 
        \wBIn19[9] , \wBIn19[8] , \wBIn19[7] , \wBIn19[6] , \wBIn19[5] , 
        \wBIn19[4] , \wBIn19[3] , \wBIn19[2] , \wBIn19[1] , \wBIn19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_18 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink19[31] , \ScanLink19[30] , \ScanLink19[29] , 
        \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , \ScanLink19[25] , 
        \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , \ScanLink19[21] , 
        \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , \ScanLink19[17] , 
        \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , \ScanLink19[13] , 
        \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , \ScanLink19[9] , 
        \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , \ScanLink19[5] , 
        \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , \ScanLink19[1] , 
        \ScanLink19[0] }), .ScanOut({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB22[31] , \wRegInB22[30] , 
        \wRegInB22[29] , \wRegInB22[28] , \wRegInB22[27] , \wRegInB22[26] , 
        \wRegInB22[25] , \wRegInB22[24] , \wRegInB22[23] , \wRegInB22[22] , 
        \wRegInB22[21] , \wRegInB22[20] , \wRegInB22[19] , \wRegInB22[18] , 
        \wRegInB22[17] , \wRegInB22[16] , \wRegInB22[15] , \wRegInB22[14] , 
        \wRegInB22[13] , \wRegInB22[12] , \wRegInB22[11] , \wRegInB22[10] , 
        \wRegInB22[9] , \wRegInB22[8] , \wRegInB22[7] , \wRegInB22[6] , 
        \wRegInB22[5] , \wRegInB22[4] , \wRegInB22[3] , \wRegInB22[2] , 
        \wRegInB22[1] , \wRegInB22[0] }), .Out({\wBIn22[31] , \wBIn22[30] , 
        \wBIn22[29] , \wBIn22[28] , \wBIn22[27] , \wBIn22[26] , \wBIn22[25] , 
        \wBIn22[24] , \wBIn22[23] , \wBIn22[22] , \wBIn22[21] , \wBIn22[20] , 
        \wBIn22[19] , \wBIn22[18] , \wBIn22[17] , \wBIn22[16] , \wBIn22[15] , 
        \wBIn22[14] , \wBIn22[13] , \wBIn22[12] , \wBIn22[11] , \wBIn22[10] , 
        \wBIn22[9] , \wBIn22[8] , \wBIn22[7] , \wBIn22[6] , \wBIn22[5] , 
        \wBIn22[4] , \wBIn22[3] , \wBIn22[2] , \wBIn22[1] , \wBIn22[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn16[31] , \wAIn16[30] , \wAIn16[29] , \wAIn16[28] , \wAIn16[27] , 
        \wAIn16[26] , \wAIn16[25] , \wAIn16[24] , \wAIn16[23] , \wAIn16[22] , 
        \wAIn16[21] , \wAIn16[20] , \wAIn16[19] , \wAIn16[18] , \wAIn16[17] , 
        \wAIn16[16] , \wAIn16[15] , \wAIn16[14] , \wAIn16[13] , \wAIn16[12] , 
        \wAIn16[11] , \wAIn16[10] , \wAIn16[9] , \wAIn16[8] , \wAIn16[7] , 
        \wAIn16[6] , \wAIn16[5] , \wAIn16[4] , \wAIn16[3] , \wAIn16[2] , 
        \wAIn16[1] , \wAIn16[0] }), .BIn({\wBIn16[31] , \wBIn16[30] , 
        \wBIn16[29] , \wBIn16[28] , \wBIn16[27] , \wBIn16[26] , \wBIn16[25] , 
        \wBIn16[24] , \wBIn16[23] , \wBIn16[22] , \wBIn16[21] , \wBIn16[20] , 
        \wBIn16[19] , \wBIn16[18] , \wBIn16[17] , \wBIn16[16] , \wBIn16[15] , 
        \wBIn16[14] , \wBIn16[13] , \wBIn16[12] , \wBIn16[11] , \wBIn16[10] , 
        \wBIn16[9] , \wBIn16[8] , \wBIn16[7] , \wBIn16[6] , \wBIn16[5] , 
        \wBIn16[4] , \wBIn16[3] , \wBIn16[2] , \wBIn16[1] , \wBIn16[0] }), 
        .HiOut({\wBMid15[31] , \wBMid15[30] , \wBMid15[29] , \wBMid15[28] , 
        \wBMid15[27] , \wBMid15[26] , \wBMid15[25] , \wBMid15[24] , 
        \wBMid15[23] , \wBMid15[22] , \wBMid15[21] , \wBMid15[20] , 
        \wBMid15[19] , \wBMid15[18] , \wBMid15[17] , \wBMid15[16] , 
        \wBMid15[15] , \wBMid15[14] , \wBMid15[13] , \wBMid15[12] , 
        \wBMid15[11] , \wBMid15[10] , \wBMid15[9] , \wBMid15[8] , \wBMid15[7] , 
        \wBMid15[6] , \wBMid15[5] , \wBMid15[4] , \wBMid15[3] , \wBMid15[2] , 
        \wBMid15[1] , \wBMid15[0] }), .LoOut({\wAMid16[31] , \wAMid16[30] , 
        \wAMid16[29] , \wAMid16[28] , \wAMid16[27] , \wAMid16[26] , 
        \wAMid16[25] , \wAMid16[24] , \wAMid16[23] , \wAMid16[22] , 
        \wAMid16[21] , \wAMid16[20] , \wAMid16[19] , \wAMid16[18] , 
        \wAMid16[17] , \wAMid16[16] , \wAMid16[15] , \wAMid16[14] , 
        \wAMid16[13] , \wAMid16[12] , \wAMid16[11] , \wAMid16[10] , 
        \wAMid16[9] , \wAMid16[8] , \wAMid16[7] , \wAMid16[6] , \wAMid16[5] , 
        \wAMid16[4] , \wAMid16[3] , \wAMid16[2] , \wAMid16[1] , \wAMid16[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn23[31] , \wAIn23[30] , \wAIn23[29] , \wAIn23[28] , \wAIn23[27] , 
        \wAIn23[26] , \wAIn23[25] , \wAIn23[24] , \wAIn23[23] , \wAIn23[22] , 
        \wAIn23[21] , \wAIn23[20] , \wAIn23[19] , \wAIn23[18] , \wAIn23[17] , 
        \wAIn23[16] , \wAIn23[15] , \wAIn23[14] , \wAIn23[13] , \wAIn23[12] , 
        \wAIn23[11] , \wAIn23[10] , \wAIn23[9] , \wAIn23[8] , \wAIn23[7] , 
        \wAIn23[6] , \wAIn23[5] , \wAIn23[4] , \wAIn23[3] , \wAIn23[2] , 
        \wAIn23[1] , \wAIn23[0] }), .BIn({\wBIn23[31] , \wBIn23[30] , 
        \wBIn23[29] , \wBIn23[28] , \wBIn23[27] , \wBIn23[26] , \wBIn23[25] , 
        \wBIn23[24] , \wBIn23[23] , \wBIn23[22] , \wBIn23[21] , \wBIn23[20] , 
        \wBIn23[19] , \wBIn23[18] , \wBIn23[17] , \wBIn23[16] , \wBIn23[15] , 
        \wBIn23[14] , \wBIn23[13] , \wBIn23[12] , \wBIn23[11] , \wBIn23[10] , 
        \wBIn23[9] , \wBIn23[8] , \wBIn23[7] , \wBIn23[6] , \wBIn23[5] , 
        \wBIn23[4] , \wBIn23[3] , \wBIn23[2] , \wBIn23[1] , \wBIn23[0] }), 
        .HiOut({\wBMid22[31] , \wBMid22[30] , \wBMid22[29] , \wBMid22[28] , 
        \wBMid22[27] , \wBMid22[26] , \wBMid22[25] , \wBMid22[24] , 
        \wBMid22[23] , \wBMid22[22] , \wBMid22[21] , \wBMid22[20] , 
        \wBMid22[19] , \wBMid22[18] , \wBMid22[17] , \wBMid22[16] , 
        \wBMid22[15] , \wBMid22[14] , \wBMid22[13] , \wBMid22[12] , 
        \wBMid22[11] , \wBMid22[10] , \wBMid22[9] , \wBMid22[8] , \wBMid22[7] , 
        \wBMid22[6] , \wBMid22[5] , \wBMid22[4] , \wBMid22[3] , \wBMid22[2] , 
        \wBMid22[1] , \wBMid22[0] }), .LoOut({\wAMid23[31] , \wAMid23[30] , 
        \wAMid23[29] , \wAMid23[28] , \wAMid23[27] , \wAMid23[26] , 
        \wAMid23[25] , \wAMid23[24] , \wAMid23[23] , \wAMid23[22] , 
        \wAMid23[21] , \wAMid23[20] , \wAMid23[19] , \wAMid23[18] , 
        \wAMid23[17] , \wAMid23[16] , \wAMid23[15] , \wAMid23[14] , 
        \wAMid23[13] , \wAMid23[12] , \wAMid23[11] , \wAMid23[10] , 
        \wAMid23[9] , \wAMid23[8] , \wAMid23[7] , \wAMid23[6] , \wAMid23[5] , 
        \wAMid23[4] , \wAMid23[3] , \wAMid23[2] , \wAMid23[1] , \wAMid23[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid13[31] , \wAMid13[30] , \wAMid13[29] , \wAMid13[28] , 
        \wAMid13[27] , \wAMid13[26] , \wAMid13[25] , \wAMid13[24] , 
        \wAMid13[23] , \wAMid13[22] , \wAMid13[21] , \wAMid13[20] , 
        \wAMid13[19] , \wAMid13[18] , \wAMid13[17] , \wAMid13[16] , 
        \wAMid13[15] , \wAMid13[14] , \wAMid13[13] , \wAMid13[12] , 
        \wAMid13[11] , \wAMid13[10] , \wAMid13[9] , \wAMid13[8] , \wAMid13[7] , 
        \wAMid13[6] , \wAMid13[5] , \wAMid13[4] , \wAMid13[3] , \wAMid13[2] , 
        \wAMid13[1] , \wAMid13[0] }), .BIn({\wBMid13[31] , \wBMid13[30] , 
        \wBMid13[29] , \wBMid13[28] , \wBMid13[27] , \wBMid13[26] , 
        \wBMid13[25] , \wBMid13[24] , \wBMid13[23] , \wBMid13[22] , 
        \wBMid13[21] , \wBMid13[20] , \wBMid13[19] , \wBMid13[18] , 
        \wBMid13[17] , \wBMid13[16] , \wBMid13[15] , \wBMid13[14] , 
        \wBMid13[13] , \wBMid13[12] , \wBMid13[11] , \wBMid13[10] , 
        \wBMid13[9] , \wBMid13[8] , \wBMid13[7] , \wBMid13[6] , \wBMid13[5] , 
        \wBMid13[4] , \wBMid13[3] , \wBMid13[2] , \wBMid13[1] , \wBMid13[0] }), 
        .HiOut({\wRegInB13[31] , \wRegInB13[30] , \wRegInB13[29] , 
        \wRegInB13[28] , \wRegInB13[27] , \wRegInB13[26] , \wRegInB13[25] , 
        \wRegInB13[24] , \wRegInB13[23] , \wRegInB13[22] , \wRegInB13[21] , 
        \wRegInB13[20] , \wRegInB13[19] , \wRegInB13[18] , \wRegInB13[17] , 
        \wRegInB13[16] , \wRegInB13[15] , \wRegInB13[14] , \wRegInB13[13] , 
        \wRegInB13[12] , \wRegInB13[11] , \wRegInB13[10] , \wRegInB13[9] , 
        \wRegInB13[8] , \wRegInB13[7] , \wRegInB13[6] , \wRegInB13[5] , 
        \wRegInB13[4] , \wRegInB13[3] , \wRegInB13[2] , \wRegInB13[1] , 
        \wRegInB13[0] }), .LoOut({\wRegInA14[31] , \wRegInA14[30] , 
        \wRegInA14[29] , \wRegInA14[28] , \wRegInA14[27] , \wRegInA14[26] , 
        \wRegInA14[25] , \wRegInA14[24] , \wRegInA14[23] , \wRegInA14[22] , 
        \wRegInA14[21] , \wRegInA14[20] , \wRegInA14[19] , \wRegInA14[18] , 
        \wRegInA14[17] , \wRegInA14[16] , \wRegInA14[15] , \wRegInA14[14] , 
        \wRegInA14[13] , \wRegInA14[12] , \wRegInA14[11] , \wRegInA14[10] , 
        \wRegInA14[9] , \wRegInA14[8] , \wRegInA14[7] , \wRegInA14[6] , 
        \wRegInA14[5] , \wRegInA14[4] , \wRegInA14[3] , \wRegInA14[2] , 
        \wRegInA14[1] , \wRegInA14[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn31[31] , \wAIn31[30] , \wAIn31[29] , \wAIn31[28] , \wAIn31[27] , 
        \wAIn31[26] , \wAIn31[25] , \wAIn31[24] , \wAIn31[23] , \wAIn31[22] , 
        \wAIn31[21] , \wAIn31[20] , \wAIn31[19] , \wAIn31[18] , \wAIn31[17] , 
        \wAIn31[16] , \wAIn31[15] , \wAIn31[14] , \wAIn31[13] , \wAIn31[12] , 
        \wAIn31[11] , \wAIn31[10] , \wAIn31[9] , \wAIn31[8] , \wAIn31[7] , 
        \wAIn31[6] , \wAIn31[5] , \wAIn31[4] , \wAIn31[3] , \wAIn31[2] , 
        \wAIn31[1] , \wAIn31[0] }), .BIn({\wBIn31[31] , \wBIn31[30] , 
        \wBIn31[29] , \wBIn31[28] , \wBIn31[27] , \wBIn31[26] , \wBIn31[25] , 
        \wBIn31[24] , \wBIn31[23] , \wBIn31[22] , \wBIn31[21] , \wBIn31[20] , 
        \wBIn31[19] , \wBIn31[18] , \wBIn31[17] , \wBIn31[16] , \wBIn31[15] , 
        \wBIn31[14] , \wBIn31[13] , \wBIn31[12] , \wBIn31[11] , \wBIn31[10] , 
        \wBIn31[9] , \wBIn31[8] , \wBIn31[7] , \wBIn31[6] , \wBIn31[5] , 
        \wBIn31[4] , \wBIn31[3] , \wBIn31[2] , \wBIn31[1] , \wBIn31[0] }), 
        .HiOut({\wBMid30[31] , \wBMid30[30] , \wBMid30[29] , \wBMid30[28] , 
        \wBMid30[27] , \wBMid30[26] , \wBMid30[25] , \wBMid30[24] , 
        \wBMid30[23] , \wBMid30[22] , \wBMid30[21] , \wBMid30[20] , 
        \wBMid30[19] , \wBMid30[18] , \wBMid30[17] , \wBMid30[16] , 
        \wBMid30[15] , \wBMid30[14] , \wBMid30[13] , \wBMid30[12] , 
        \wBMid30[11] , \wBMid30[10] , \wBMid30[9] , \wBMid30[8] , \wBMid30[7] , 
        \wBMid30[6] , \wBMid30[5] , \wBMid30[4] , \wBMid30[3] , \wBMid30[2] , 
        \wBMid30[1] , \wBMid30[0] }), .LoOut({\wRegInB31[31] , \wRegInB31[30] , 
        \wRegInB31[29] , \wRegInB31[28] , \wRegInB31[27] , \wRegInB31[26] , 
        \wRegInB31[25] , \wRegInB31[24] , \wRegInB31[23] , \wRegInB31[22] , 
        \wRegInB31[21] , \wRegInB31[20] , \wRegInB31[19] , \wRegInB31[18] , 
        \wRegInB31[17] , \wRegInB31[16] , \wRegInB31[15] , \wRegInB31[14] , 
        \wRegInB31[13] , \wRegInB31[12] , \wRegInB31[11] , \wRegInB31[10] , 
        \wRegInB31[9] , \wRegInB31[8] , \wRegInB31[7] , \wRegInB31[6] , 
        \wRegInB31[5] , \wRegInB31[4] , \wRegInB31[3] , \wRegInB31[2] , 
        \wRegInB31[1] , \wRegInB31[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_51 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink52[31] , \ScanLink52[30] , \ScanLink52[29] , 
        \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , \ScanLink52[25] , 
        \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , \ScanLink52[21] , 
        \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , \ScanLink52[17] , 
        \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , \ScanLink52[13] , 
        \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , \ScanLink52[9] , 
        \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , \ScanLink52[5] , 
        \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , \ScanLink52[1] , 
        \ScanLink52[0] }), .ScanOut({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA6[31] , \wRegInA6[30] , 
        \wRegInA6[29] , \wRegInA6[28] , \wRegInA6[27] , \wRegInA6[26] , 
        \wRegInA6[25] , \wRegInA6[24] , \wRegInA6[23] , \wRegInA6[22] , 
        \wRegInA6[21] , \wRegInA6[20] , \wRegInA6[19] , \wRegInA6[18] , 
        \wRegInA6[17] , \wRegInA6[16] , \wRegInA6[15] , \wRegInA6[14] , 
        \wRegInA6[13] , \wRegInA6[12] , \wRegInA6[11] , \wRegInA6[10] , 
        \wRegInA6[9] , \wRegInA6[8] , \wRegInA6[7] , \wRegInA6[6] , 
        \wRegInA6[5] , \wRegInA6[4] , \wRegInA6[3] , \wRegInA6[2] , 
        \wRegInA6[1] , \wRegInA6[0] }), .Out({\wAIn6[31] , \wAIn6[30] , 
        \wAIn6[29] , \wAIn6[28] , \wAIn6[27] , \wAIn6[26] , \wAIn6[25] , 
        \wAIn6[24] , \wAIn6[23] , \wAIn6[22] , \wAIn6[21] , \wAIn6[20] , 
        \wAIn6[19] , \wAIn6[18] , \wAIn6[17] , \wAIn6[16] , \wAIn6[15] , 
        \wAIn6[14] , \wAIn6[13] , \wAIn6[12] , \wAIn6[11] , \wAIn6[10] , 
        \wAIn6[9] , \wAIn6[8] , \wAIn6[7] , \wAIn6[6] , \wAIn6[5] , \wAIn6[4] , 
        \wAIn6[3] , \wAIn6[2] , \wAIn6[1] , \wAIn6[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid26[31] , \wAMid26[30] , \wAMid26[29] , \wAMid26[28] , 
        \wAMid26[27] , \wAMid26[26] , \wAMid26[25] , \wAMid26[24] , 
        \wAMid26[23] , \wAMid26[22] , \wAMid26[21] , \wAMid26[20] , 
        \wAMid26[19] , \wAMid26[18] , \wAMid26[17] , \wAMid26[16] , 
        \wAMid26[15] , \wAMid26[14] , \wAMid26[13] , \wAMid26[12] , 
        \wAMid26[11] , \wAMid26[10] , \wAMid26[9] , \wAMid26[8] , \wAMid26[7] , 
        \wAMid26[6] , \wAMid26[5] , \wAMid26[4] , \wAMid26[3] , \wAMid26[2] , 
        \wAMid26[1] , \wAMid26[0] }), .BIn({\wBMid26[31] , \wBMid26[30] , 
        \wBMid26[29] , \wBMid26[28] , \wBMid26[27] , \wBMid26[26] , 
        \wBMid26[25] , \wBMid26[24] , \wBMid26[23] , \wBMid26[22] , 
        \wBMid26[21] , \wBMid26[20] , \wBMid26[19] , \wBMid26[18] , 
        \wBMid26[17] , \wBMid26[16] , \wBMid26[15] , \wBMid26[14] , 
        \wBMid26[13] , \wBMid26[12] , \wBMid26[11] , \wBMid26[10] , 
        \wBMid26[9] , \wBMid26[8] , \wBMid26[7] , \wBMid26[6] , \wBMid26[5] , 
        \wBMid26[4] , \wBMid26[3] , \wBMid26[2] , \wBMid26[1] , \wBMid26[0] }), 
        .HiOut({\wRegInB26[31] , \wRegInB26[30] , \wRegInB26[29] , 
        \wRegInB26[28] , \wRegInB26[27] , \wRegInB26[26] , \wRegInB26[25] , 
        \wRegInB26[24] , \wRegInB26[23] , \wRegInB26[22] , \wRegInB26[21] , 
        \wRegInB26[20] , \wRegInB26[19] , \wRegInB26[18] , \wRegInB26[17] , 
        \wRegInB26[16] , \wRegInB26[15] , \wRegInB26[14] , \wRegInB26[13] , 
        \wRegInB26[12] , \wRegInB26[11] , \wRegInB26[10] , \wRegInB26[9] , 
        \wRegInB26[8] , \wRegInB26[7] , \wRegInB26[6] , \wRegInB26[5] , 
        \wRegInB26[4] , \wRegInB26[3] , \wRegInB26[2] , \wRegInB26[1] , 
        \wRegInB26[0] }), .LoOut({\wRegInA27[31] , \wRegInA27[30] , 
        \wRegInA27[29] , \wRegInA27[28] , \wRegInA27[27] , \wRegInA27[26] , 
        \wRegInA27[25] , \wRegInA27[24] , \wRegInA27[23] , \wRegInA27[22] , 
        \wRegInA27[21] , \wRegInA27[20] , \wRegInA27[19] , \wRegInA27[18] , 
        \wRegInA27[17] , \wRegInA27[16] , \wRegInA27[15] , \wRegInA27[14] , 
        \wRegInA27[13] , \wRegInA27[12] , \wRegInA27[11] , \wRegInA27[10] , 
        \wRegInA27[9] , \wRegInA27[8] , \wRegInA27[7] , \wRegInA27[6] , 
        \wRegInA27[5] , \wRegInA27[4] , \wRegInA27[3] , \wRegInA27[2] , 
        \wRegInA27[1] , \wRegInA27[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_43 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink44[31] , \ScanLink44[30] , \ScanLink44[29] , 
        \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , \ScanLink44[25] , 
        \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , \ScanLink44[21] , 
        \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , \ScanLink44[17] , 
        \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , \ScanLink44[13] , 
        \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , \ScanLink44[9] , 
        \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , \ScanLink44[5] , 
        \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , \ScanLink44[1] , 
        \ScanLink44[0] }), .ScanOut({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA10[31] , \wRegInA10[30] , 
        \wRegInA10[29] , \wRegInA10[28] , \wRegInA10[27] , \wRegInA10[26] , 
        \wRegInA10[25] , \wRegInA10[24] , \wRegInA10[23] , \wRegInA10[22] , 
        \wRegInA10[21] , \wRegInA10[20] , \wRegInA10[19] , \wRegInA10[18] , 
        \wRegInA10[17] , \wRegInA10[16] , \wRegInA10[15] , \wRegInA10[14] , 
        \wRegInA10[13] , \wRegInA10[12] , \wRegInA10[11] , \wRegInA10[10] , 
        \wRegInA10[9] , \wRegInA10[8] , \wRegInA10[7] , \wRegInA10[6] , 
        \wRegInA10[5] , \wRegInA10[4] , \wRegInA10[3] , \wRegInA10[2] , 
        \wRegInA10[1] , \wRegInA10[0] }), .Out({\wAIn10[31] , \wAIn10[30] , 
        \wAIn10[29] , \wAIn10[28] , \wAIn10[27] , \wAIn10[26] , \wAIn10[25] , 
        \wAIn10[24] , \wAIn10[23] , \wAIn10[22] , \wAIn10[21] , \wAIn10[20] , 
        \wAIn10[19] , \wAIn10[18] , \wAIn10[17] , \wAIn10[16] , \wAIn10[15] , 
        \wAIn10[14] , \wAIn10[13] , \wAIn10[12] , \wAIn10[11] , \wAIn10[10] , 
        \wAIn10[9] , \wAIn10[8] , \wAIn10[7] , \wAIn10[6] , \wAIn10[5] , 
        \wAIn10[4] , \wAIn10[3] , \wAIn10[2] , \wAIn10[1] , \wAIn10[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_0 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[31] , \ScanLink1[30] , \ScanLink1[29] , 
        \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , \ScanLink1[25] , 
        \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , \ScanLink1[21] , 
        \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , \ScanLink1[17] , 
        \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , \ScanLink1[13] , 
        \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , \ScanLink1[9] , 
        \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB31[31] , \wRegInB31[30] , 
        \wRegInB31[29] , \wRegInB31[28] , \wRegInB31[27] , \wRegInB31[26] , 
        \wRegInB31[25] , \wRegInB31[24] , \wRegInB31[23] , \wRegInB31[22] , 
        \wRegInB31[21] , \wRegInB31[20] , \wRegInB31[19] , \wRegInB31[18] , 
        \wRegInB31[17] , \wRegInB31[16] , \wRegInB31[15] , \wRegInB31[14] , 
        \wRegInB31[13] , \wRegInB31[12] , \wRegInB31[11] , \wRegInB31[10] , 
        \wRegInB31[9] , \wRegInB31[8] , \wRegInB31[7] , \wRegInB31[6] , 
        \wRegInB31[5] , \wRegInB31[4] , \wRegInB31[3] , \wRegInB31[2] , 
        \wRegInB31[1] , \wRegInB31[0] }), .Out({\wBIn31[31] , \wBIn31[30] , 
        \wBIn31[29] , \wBIn31[28] , \wBIn31[27] , \wBIn31[26] , \wBIn31[25] , 
        \wBIn31[24] , \wBIn31[23] , \wBIn31[22] , \wBIn31[21] , \wBIn31[20] , 
        \wBIn31[19] , \wBIn31[18] , \wBIn31[17] , \wBIn31[16] , \wBIn31[15] , 
        \wBIn31[14] , \wBIn31[13] , \wBIn31[12] , \wBIn31[11] , \wBIn31[10] , 
        \wBIn31[9] , \wBIn31[8] , \wBIn31[7] , \wBIn31[6] , \wBIn31[5] , 
        \wBIn31[4] , \wBIn31[3] , \wBIn31[2] , \wBIn31[1] , \wBIn31[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_36 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink37[31] , \ScanLink37[30] , \ScanLink37[29] , 
        \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , \ScanLink37[25] , 
        \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , \ScanLink37[21] , 
        \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , \ScanLink37[17] , 
        \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , \ScanLink37[13] , 
        \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , \ScanLink37[9] , 
        \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , \ScanLink37[5] , 
        \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , \ScanLink37[1] , 
        \ScanLink37[0] }), .ScanOut({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB13[31] , \wRegInB13[30] , 
        \wRegInB13[29] , \wRegInB13[28] , \wRegInB13[27] , \wRegInB13[26] , 
        \wRegInB13[25] , \wRegInB13[24] , \wRegInB13[23] , \wRegInB13[22] , 
        \wRegInB13[21] , \wRegInB13[20] , \wRegInB13[19] , \wRegInB13[18] , 
        \wRegInB13[17] , \wRegInB13[16] , \wRegInB13[15] , \wRegInB13[14] , 
        \wRegInB13[13] , \wRegInB13[12] , \wRegInB13[11] , \wRegInB13[10] , 
        \wRegInB13[9] , \wRegInB13[8] , \wRegInB13[7] , \wRegInB13[6] , 
        \wRegInB13[5] , \wRegInB13[4] , \wRegInB13[3] , \wRegInB13[2] , 
        \wRegInB13[1] , \wRegInB13[0] }), .Out({\wBIn13[31] , \wBIn13[30] , 
        \wBIn13[29] , \wBIn13[28] , \wBIn13[27] , \wBIn13[26] , \wBIn13[25] , 
        \wBIn13[24] , \wBIn13[23] , \wBIn13[22] , \wBIn13[21] , \wBIn13[20] , 
        \wBIn13[19] , \wBIn13[18] , \wBIn13[17] , \wBIn13[16] , \wBIn13[15] , 
        \wBIn13[14] , \wBIn13[13] , \wBIn13[12] , \wBIn13[11] , \wBIn13[10] , 
        \wBIn13[9] , \wBIn13[8] , \wBIn13[7] , \wBIn13[6] , \wBIn13[5] , 
        \wBIn13[4] , \wBIn13[3] , \wBIn13[2] , \wBIn13[1] , \wBIn13[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_11 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[31] , \ScanLink12[30] , \ScanLink12[29] , 
        \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , \ScanLink12[25] , 
        \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , \ScanLink12[21] , 
        \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , \ScanLink12[17] , 
        \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , \ScanLink12[13] , 
        \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , \ScanLink12[9] , 
        \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA26[31] , \wRegInA26[30] , 
        \wRegInA26[29] , \wRegInA26[28] , \wRegInA26[27] , \wRegInA26[26] , 
        \wRegInA26[25] , \wRegInA26[24] , \wRegInA26[23] , \wRegInA26[22] , 
        \wRegInA26[21] , \wRegInA26[20] , \wRegInA26[19] , \wRegInA26[18] , 
        \wRegInA26[17] , \wRegInA26[16] , \wRegInA26[15] , \wRegInA26[14] , 
        \wRegInA26[13] , \wRegInA26[12] , \wRegInA26[11] , \wRegInA26[10] , 
        \wRegInA26[9] , \wRegInA26[8] , \wRegInA26[7] , \wRegInA26[6] , 
        \wRegInA26[5] , \wRegInA26[4] , \wRegInA26[3] , \wRegInA26[2] , 
        \wRegInA26[1] , \wRegInA26[0] }), .Out({\wAIn26[31] , \wAIn26[30] , 
        \wAIn26[29] , \wAIn26[28] , \wAIn26[27] , \wAIn26[26] , \wAIn26[25] , 
        \wAIn26[24] , \wAIn26[23] , \wAIn26[22] , \wAIn26[21] , \wAIn26[20] , 
        \wAIn26[19] , \wAIn26[18] , \wAIn26[17] , \wAIn26[16] , \wAIn26[15] , 
        \wAIn26[14] , \wAIn26[13] , \wAIn26[12] , \wAIn26[11] , \wAIn26[10] , 
        \wAIn26[9] , \wAIn26[8] , \wAIn26[7] , \wAIn26[6] , \wAIn26[5] , 
        \wAIn26[4] , \wAIn26[3] , \wAIn26[2] , \wAIn26[1] , \wAIn26[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn1[31] , 
        \wAIn1[30] , \wAIn1[29] , \wAIn1[28] , \wAIn1[27] , \wAIn1[26] , 
        \wAIn1[25] , \wAIn1[24] , \wAIn1[23] , \wAIn1[22] , \wAIn1[21] , 
        \wAIn1[20] , \wAIn1[19] , \wAIn1[18] , \wAIn1[17] , \wAIn1[16] , 
        \wAIn1[15] , \wAIn1[14] , \wAIn1[13] , \wAIn1[12] , \wAIn1[11] , 
        \wAIn1[10] , \wAIn1[9] , \wAIn1[8] , \wAIn1[7] , \wAIn1[6] , 
        \wAIn1[5] , \wAIn1[4] , \wAIn1[3] , \wAIn1[2] , \wAIn1[1] , \wAIn1[0] 
        }), .BIn({\wBIn1[31] , \wBIn1[30] , \wBIn1[29] , \wBIn1[28] , 
        \wBIn1[27] , \wBIn1[26] , \wBIn1[25] , \wBIn1[24] , \wBIn1[23] , 
        \wBIn1[22] , \wBIn1[21] , \wBIn1[20] , \wBIn1[19] , \wBIn1[18] , 
        \wBIn1[17] , \wBIn1[16] , \wBIn1[15] , \wBIn1[14] , \wBIn1[13] , 
        \wBIn1[12] , \wBIn1[11] , \wBIn1[10] , \wBIn1[9] , \wBIn1[8] , 
        \wBIn1[7] , \wBIn1[6] , \wBIn1[5] , \wBIn1[4] , \wBIn1[3] , \wBIn1[2] , 
        \wBIn1[1] , \wBIn1[0] }), .HiOut({\wBMid0[31] , \wBMid0[30] , 
        \wBMid0[29] , \wBMid0[28] , \wBMid0[27] , \wBMid0[26] , \wBMid0[25] , 
        \wBMid0[24] , \wBMid0[23] , \wBMid0[22] , \wBMid0[21] , \wBMid0[20] , 
        \wBMid0[19] , \wBMid0[18] , \wBMid0[17] , \wBMid0[16] , \wBMid0[15] , 
        \wBMid0[14] , \wBMid0[13] , \wBMid0[12] , \wBMid0[11] , \wBMid0[10] , 
        \wBMid0[9] , \wBMid0[8] , \wBMid0[7] , \wBMid0[6] , \wBMid0[5] , 
        \wBMid0[4] , \wBMid0[3] , \wBMid0[2] , \wBMid0[1] , \wBMid0[0] }), 
        .LoOut({\wAMid1[31] , \wAMid1[30] , \wAMid1[29] , \wAMid1[28] , 
        \wAMid1[27] , \wAMid1[26] , \wAMid1[25] , \wAMid1[24] , \wAMid1[23] , 
        \wAMid1[22] , \wAMid1[21] , \wAMid1[20] , \wAMid1[19] , \wAMid1[18] , 
        \wAMid1[17] , \wAMid1[16] , \wAMid1[15] , \wAMid1[14] , \wAMid1[13] , 
        \wAMid1[12] , \wAMid1[11] , \wAMid1[10] , \wAMid1[9] , \wAMid1[8] , 
        \wAMid1[7] , \wAMid1[6] , \wAMid1[5] , \wAMid1[4] , \wAMid1[3] , 
        \wAMid1[2] , \wAMid1[1] , \wAMid1[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn8[31] , 
        \wAIn8[30] , \wAIn8[29] , \wAIn8[28] , \wAIn8[27] , \wAIn8[26] , 
        \wAIn8[25] , \wAIn8[24] , \wAIn8[23] , \wAIn8[22] , \wAIn8[21] , 
        \wAIn8[20] , \wAIn8[19] , \wAIn8[18] , \wAIn8[17] , \wAIn8[16] , 
        \wAIn8[15] , \wAIn8[14] , \wAIn8[13] , \wAIn8[12] , \wAIn8[11] , 
        \wAIn8[10] , \wAIn8[9] , \wAIn8[8] , \wAIn8[7] , \wAIn8[6] , 
        \wAIn8[5] , \wAIn8[4] , \wAIn8[3] , \wAIn8[2] , \wAIn8[1] , \wAIn8[0] 
        }), .BIn({\wBIn8[31] , \wBIn8[30] , \wBIn8[29] , \wBIn8[28] , 
        \wBIn8[27] , \wBIn8[26] , \wBIn8[25] , \wBIn8[24] , \wBIn8[23] , 
        \wBIn8[22] , \wBIn8[21] , \wBIn8[20] , \wBIn8[19] , \wBIn8[18] , 
        \wBIn8[17] , \wBIn8[16] , \wBIn8[15] , \wBIn8[14] , \wBIn8[13] , 
        \wBIn8[12] , \wBIn8[11] , \wBIn8[10] , \wBIn8[9] , \wBIn8[8] , 
        \wBIn8[7] , \wBIn8[6] , \wBIn8[5] , \wBIn8[4] , \wBIn8[3] , \wBIn8[2] , 
        \wBIn8[1] , \wBIn8[0] }), .HiOut({\wBMid7[31] , \wBMid7[30] , 
        \wBMid7[29] , \wBMid7[28] , \wBMid7[27] , \wBMid7[26] , \wBMid7[25] , 
        \wBMid7[24] , \wBMid7[23] , \wBMid7[22] , \wBMid7[21] , \wBMid7[20] , 
        \wBMid7[19] , \wBMid7[18] , \wBMid7[17] , \wBMid7[16] , \wBMid7[15] , 
        \wBMid7[14] , \wBMid7[13] , \wBMid7[12] , \wBMid7[11] , \wBMid7[10] , 
        \wBMid7[9] , \wBMid7[8] , \wBMid7[7] , \wBMid7[6] , \wBMid7[5] , 
        \wBMid7[4] , \wBMid7[3] , \wBMid7[2] , \wBMid7[1] , \wBMid7[0] }), 
        .LoOut({\wAMid8[31] , \wAMid8[30] , \wAMid8[29] , \wAMid8[28] , 
        \wAMid8[27] , \wAMid8[26] , \wAMid8[25] , \wAMid8[24] , \wAMid8[23] , 
        \wAMid8[22] , \wAMid8[21] , \wAMid8[20] , \wAMid8[19] , \wAMid8[18] , 
        \wAMid8[17] , \wAMid8[16] , \wAMid8[15] , \wAMid8[14] , \wAMid8[13] , 
        \wAMid8[12] , \wAMid8[11] , \wAMid8[10] , \wAMid8[9] , \wAMid8[8] , 
        \wAMid8[7] , \wAMid8[6] , \wAMid8[5] , \wAMid8[4] , \wAMid8[3] , 
        \wAMid8[2] , \wAMid8[1] , \wAMid8[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_58 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink59[31] , \ScanLink59[30] , \ScanLink59[29] , 
        \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , \ScanLink59[25] , 
        \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , \ScanLink59[21] , 
        \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , \ScanLink59[17] , 
        \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , \ScanLink59[13] , 
        \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , \ScanLink59[9] , 
        \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , \ScanLink59[5] , 
        \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , \ScanLink59[1] , 
        \ScanLink59[0] }), .ScanOut({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB2[31] , \wRegInB2[30] , 
        \wRegInB2[29] , \wRegInB2[28] , \wRegInB2[27] , \wRegInB2[26] , 
        \wRegInB2[25] , \wRegInB2[24] , \wRegInB2[23] , \wRegInB2[22] , 
        \wRegInB2[21] , \wRegInB2[20] , \wRegInB2[19] , \wRegInB2[18] , 
        \wRegInB2[17] , \wRegInB2[16] , \wRegInB2[15] , \wRegInB2[14] , 
        \wRegInB2[13] , \wRegInB2[12] , \wRegInB2[11] , \wRegInB2[10] , 
        \wRegInB2[9] , \wRegInB2[8] , \wRegInB2[7] , \wRegInB2[6] , 
        \wRegInB2[5] , \wRegInB2[4] , \wRegInB2[3] , \wRegInB2[2] , 
        \wRegInB2[1] , \wRegInB2[0] }), .Out({\wBIn2[31] , \wBIn2[30] , 
        \wBIn2[29] , \wBIn2[28] , \wBIn2[27] , \wBIn2[26] , \wBIn2[25] , 
        \wBIn2[24] , \wBIn2[23] , \wBIn2[22] , \wBIn2[21] , \wBIn2[20] , 
        \wBIn2[19] , \wBIn2[18] , \wBIn2[17] , \wBIn2[16] , \wBIn2[15] , 
        \wBIn2[14] , \wBIn2[13] , \wBIn2[12] , \wBIn2[11] , \wBIn2[10] , 
        \wBIn2[9] , \wBIn2[8] , \wBIn2[7] , \wBIn2[6] , \wBIn2[5] , \wBIn2[4] , 
        \wBIn2[3] , \wBIn2[2] , \wBIn2[1] , \wBIn2[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn22[31] , \wAIn22[30] , \wAIn22[29] , \wAIn22[28] , \wAIn22[27] , 
        \wAIn22[26] , \wAIn22[25] , \wAIn22[24] , \wAIn22[23] , \wAIn22[22] , 
        \wAIn22[21] , \wAIn22[20] , \wAIn22[19] , \wAIn22[18] , \wAIn22[17] , 
        \wAIn22[16] , \wAIn22[15] , \wAIn22[14] , \wAIn22[13] , \wAIn22[12] , 
        \wAIn22[11] , \wAIn22[10] , \wAIn22[9] , \wAIn22[8] , \wAIn22[7] , 
        \wAIn22[6] , \wAIn22[5] , \wAIn22[4] , \wAIn22[3] , \wAIn22[2] , 
        \wAIn22[1] , \wAIn22[0] }), .BIn({\wBIn22[31] , \wBIn22[30] , 
        \wBIn22[29] , \wBIn22[28] , \wBIn22[27] , \wBIn22[26] , \wBIn22[25] , 
        \wBIn22[24] , \wBIn22[23] , \wBIn22[22] , \wBIn22[21] , \wBIn22[20] , 
        \wBIn22[19] , \wBIn22[18] , \wBIn22[17] , \wBIn22[16] , \wBIn22[15] , 
        \wBIn22[14] , \wBIn22[13] , \wBIn22[12] , \wBIn22[11] , \wBIn22[10] , 
        \wBIn22[9] , \wBIn22[8] , \wBIn22[7] , \wBIn22[6] , \wBIn22[5] , 
        \wBIn22[4] , \wBIn22[3] , \wBIn22[2] , \wBIn22[1] , \wBIn22[0] }), 
        .HiOut({\wBMid21[31] , \wBMid21[30] , \wBMid21[29] , \wBMid21[28] , 
        \wBMid21[27] , \wBMid21[26] , \wBMid21[25] , \wBMid21[24] , 
        \wBMid21[23] , \wBMid21[22] , \wBMid21[21] , \wBMid21[20] , 
        \wBMid21[19] , \wBMid21[18] , \wBMid21[17] , \wBMid21[16] , 
        \wBMid21[15] , \wBMid21[14] , \wBMid21[13] , \wBMid21[12] , 
        \wBMid21[11] , \wBMid21[10] , \wBMid21[9] , \wBMid21[8] , \wBMid21[7] , 
        \wBMid21[6] , \wBMid21[5] , \wBMid21[4] , \wBMid21[3] , \wBMid21[2] , 
        \wBMid21[1] , \wBMid21[0] }), .LoOut({\wAMid22[31] , \wAMid22[30] , 
        \wAMid22[29] , \wAMid22[28] , \wAMid22[27] , \wAMid22[26] , 
        \wAMid22[25] , \wAMid22[24] , \wAMid22[23] , \wAMid22[22] , 
        \wAMid22[21] , \wAMid22[20] , \wAMid22[19] , \wAMid22[18] , 
        \wAMid22[17] , \wAMid22[16] , \wAMid22[15] , \wAMid22[14] , 
        \wAMid22[13] , \wAMid22[12] , \wAMid22[11] , \wAMid22[10] , 
        \wAMid22[9] , \wAMid22[8] , \wAMid22[7] , \wAMid22[6] , \wAMid22[5] , 
        \wAMid22[4] , \wAMid22[3] , \wAMid22[2] , \wAMid22[1] , \wAMid22[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid4[31] , 
        \wAMid4[30] , \wAMid4[29] , \wAMid4[28] , \wAMid4[27] , \wAMid4[26] , 
        \wAMid4[25] , \wAMid4[24] , \wAMid4[23] , \wAMid4[22] , \wAMid4[21] , 
        \wAMid4[20] , \wAMid4[19] , \wAMid4[18] , \wAMid4[17] , \wAMid4[16] , 
        \wAMid4[15] , \wAMid4[14] , \wAMid4[13] , \wAMid4[12] , \wAMid4[11] , 
        \wAMid4[10] , \wAMid4[9] , \wAMid4[8] , \wAMid4[7] , \wAMid4[6] , 
        \wAMid4[5] , \wAMid4[4] , \wAMid4[3] , \wAMid4[2] , \wAMid4[1] , 
        \wAMid4[0] }), .BIn({\wBMid4[31] , \wBMid4[30] , \wBMid4[29] , 
        \wBMid4[28] , \wBMid4[27] , \wBMid4[26] , \wBMid4[25] , \wBMid4[24] , 
        \wBMid4[23] , \wBMid4[22] , \wBMid4[21] , \wBMid4[20] , \wBMid4[19] , 
        \wBMid4[18] , \wBMid4[17] , \wBMid4[16] , \wBMid4[15] , \wBMid4[14] , 
        \wBMid4[13] , \wBMid4[12] , \wBMid4[11] , \wBMid4[10] , \wBMid4[9] , 
        \wBMid4[8] , \wBMid4[7] , \wBMid4[6] , \wBMid4[5] , \wBMid4[4] , 
        \wBMid4[3] , \wBMid4[2] , \wBMid4[1] , \wBMid4[0] }), .HiOut({
        \wRegInB4[31] , \wRegInB4[30] , \wRegInB4[29] , \wRegInB4[28] , 
        \wRegInB4[27] , \wRegInB4[26] , \wRegInB4[25] , \wRegInB4[24] , 
        \wRegInB4[23] , \wRegInB4[22] , \wRegInB4[21] , \wRegInB4[20] , 
        \wRegInB4[19] , \wRegInB4[18] , \wRegInB4[17] , \wRegInB4[16] , 
        \wRegInB4[15] , \wRegInB4[14] , \wRegInB4[13] , \wRegInB4[12] , 
        \wRegInB4[11] , \wRegInB4[10] , \wRegInB4[9] , \wRegInB4[8] , 
        \wRegInB4[7] , \wRegInB4[6] , \wRegInB4[5] , \wRegInB4[4] , 
        \wRegInB4[3] , \wRegInB4[2] , \wRegInB4[1] , \wRegInB4[0] }), .LoOut({
        \wRegInA5[31] , \wRegInA5[30] , \wRegInA5[29] , \wRegInA5[28] , 
        \wRegInA5[27] , \wRegInA5[26] , \wRegInA5[25] , \wRegInA5[24] , 
        \wRegInA5[23] , \wRegInA5[22] , \wRegInA5[21] , \wRegInA5[20] , 
        \wRegInA5[19] , \wRegInA5[18] , \wRegInA5[17] , \wRegInA5[16] , 
        \wRegInA5[15] , \wRegInA5[14] , \wRegInA5[13] , \wRegInA5[12] , 
        \wRegInA5[11] , \wRegInA5[10] , \wRegInA5[9] , \wRegInA5[8] , 
        \wRegInA5[7] , \wRegInA5[6] , \wRegInA5[5] , \wRegInA5[4] , 
        \wRegInA5[3] , \wRegInA5[2] , \wRegInA5[1] , \wRegInA5[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid12[31] , \wAMid12[30] , \wAMid12[29] , \wAMid12[28] , 
        \wAMid12[27] , \wAMid12[26] , \wAMid12[25] , \wAMid12[24] , 
        \wAMid12[23] , \wAMid12[22] , \wAMid12[21] , \wAMid12[20] , 
        \wAMid12[19] , \wAMid12[18] , \wAMid12[17] , \wAMid12[16] , 
        \wAMid12[15] , \wAMid12[14] , \wAMid12[13] , \wAMid12[12] , 
        \wAMid12[11] , \wAMid12[10] , \wAMid12[9] , \wAMid12[8] , \wAMid12[7] , 
        \wAMid12[6] , \wAMid12[5] , \wAMid12[4] , \wAMid12[3] , \wAMid12[2] , 
        \wAMid12[1] , \wAMid12[0] }), .BIn({\wBMid12[31] , \wBMid12[30] , 
        \wBMid12[29] , \wBMid12[28] , \wBMid12[27] , \wBMid12[26] , 
        \wBMid12[25] , \wBMid12[24] , \wBMid12[23] , \wBMid12[22] , 
        \wBMid12[21] , \wBMid12[20] , \wBMid12[19] , \wBMid12[18] , 
        \wBMid12[17] , \wBMid12[16] , \wBMid12[15] , \wBMid12[14] , 
        \wBMid12[13] , \wBMid12[12] , \wBMid12[11] , \wBMid12[10] , 
        \wBMid12[9] , \wBMid12[8] , \wBMid12[7] , \wBMid12[6] , \wBMid12[5] , 
        \wBMid12[4] , \wBMid12[3] , \wBMid12[2] , \wBMid12[1] , \wBMid12[0] }), 
        .HiOut({\wRegInB12[31] , \wRegInB12[30] , \wRegInB12[29] , 
        \wRegInB12[28] , \wRegInB12[27] , \wRegInB12[26] , \wRegInB12[25] , 
        \wRegInB12[24] , \wRegInB12[23] , \wRegInB12[22] , \wRegInB12[21] , 
        \wRegInB12[20] , \wRegInB12[19] , \wRegInB12[18] , \wRegInB12[17] , 
        \wRegInB12[16] , \wRegInB12[15] , \wRegInB12[14] , \wRegInB12[13] , 
        \wRegInB12[12] , \wRegInB12[11] , \wRegInB12[10] , \wRegInB12[9] , 
        \wRegInB12[8] , \wRegInB12[7] , \wRegInB12[6] , \wRegInB12[5] , 
        \wRegInB12[4] , \wRegInB12[3] , \wRegInB12[2] , \wRegInB12[1] , 
        \wRegInB12[0] }), .LoOut({\wRegInA13[31] , \wRegInA13[30] , 
        \wRegInA13[29] , \wRegInA13[28] , \wRegInA13[27] , \wRegInA13[26] , 
        \wRegInA13[25] , \wRegInA13[24] , \wRegInA13[23] , \wRegInA13[22] , 
        \wRegInA13[21] , \wRegInA13[20] , \wRegInA13[19] , \wRegInA13[18] , 
        \wRegInA13[17] , \wRegInA13[16] , \wRegInA13[15] , \wRegInA13[14] , 
        \wRegInA13[13] , \wRegInA13[12] , \wRegInA13[11] , \wRegInA13[10] , 
        \wRegInA13[9] , \wRegInA13[8] , \wRegInA13[7] , \wRegInA13[6] , 
        \wRegInA13[5] , \wRegInA13[4] , \wRegInA13[3] , \wRegInA13[2] , 
        \wRegInA13[1] , \wRegInA13[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_50 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink51[31] , \ScanLink51[30] , \ScanLink51[29] , 
        \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , \ScanLink51[25] , 
        \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , \ScanLink51[21] , 
        \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , \ScanLink51[17] , 
        \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , \ScanLink51[13] , 
        \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , \ScanLink51[9] , 
        \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , \ScanLink51[5] , 
        \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , \ScanLink51[1] , 
        \ScanLink51[0] }), .ScanOut({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB6[31] , \wRegInB6[30] , 
        \wRegInB6[29] , \wRegInB6[28] , \wRegInB6[27] , \wRegInB6[26] , 
        \wRegInB6[25] , \wRegInB6[24] , \wRegInB6[23] , \wRegInB6[22] , 
        \wRegInB6[21] , \wRegInB6[20] , \wRegInB6[19] , \wRegInB6[18] , 
        \wRegInB6[17] , \wRegInB6[16] , \wRegInB6[15] , \wRegInB6[14] , 
        \wRegInB6[13] , \wRegInB6[12] , \wRegInB6[11] , \wRegInB6[10] , 
        \wRegInB6[9] , \wRegInB6[8] , \wRegInB6[7] , \wRegInB6[6] , 
        \wRegInB6[5] , \wRegInB6[4] , \wRegInB6[3] , \wRegInB6[2] , 
        \wRegInB6[1] , \wRegInB6[0] }), .Out({\wBIn6[31] , \wBIn6[30] , 
        \wBIn6[29] , \wBIn6[28] , \wBIn6[27] , \wBIn6[26] , \wBIn6[25] , 
        \wBIn6[24] , \wBIn6[23] , \wBIn6[22] , \wBIn6[21] , \wBIn6[20] , 
        \wBIn6[19] , \wBIn6[18] , \wBIn6[17] , \wBIn6[16] , \wBIn6[15] , 
        \wBIn6[14] , \wBIn6[13] , \wBIn6[12] , \wBIn6[11] , \wBIn6[10] , 
        \wBIn6[9] , \wBIn6[8] , \wBIn6[7] , \wBIn6[6] , \wBIn6[5] , \wBIn6[4] , 
        \wBIn6[3] , \wBIn6[2] , \wBIn6[1] , \wBIn6[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_25 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink26[31] , \ScanLink26[30] , \ScanLink26[29] , 
        \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , \ScanLink26[25] , 
        \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , \ScanLink26[21] , 
        \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , \ScanLink26[17] , 
        \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , \ScanLink26[13] , 
        \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , \ScanLink26[9] , 
        \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , \ScanLink26[5] , 
        \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , \ScanLink26[1] , 
        \ScanLink26[0] }), .ScanOut({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA19[31] , \wRegInA19[30] , 
        \wRegInA19[29] , \wRegInA19[28] , \wRegInA19[27] , \wRegInA19[26] , 
        \wRegInA19[25] , \wRegInA19[24] , \wRegInA19[23] , \wRegInA19[22] , 
        \wRegInA19[21] , \wRegInA19[20] , \wRegInA19[19] , \wRegInA19[18] , 
        \wRegInA19[17] , \wRegInA19[16] , \wRegInA19[15] , \wRegInA19[14] , 
        \wRegInA19[13] , \wRegInA19[12] , \wRegInA19[11] , \wRegInA19[10] , 
        \wRegInA19[9] , \wRegInA19[8] , \wRegInA19[7] , \wRegInA19[6] , 
        \wRegInA19[5] , \wRegInA19[4] , \wRegInA19[3] , \wRegInA19[2] , 
        \wRegInA19[1] , \wRegInA19[0] }), .Out({\wAIn19[31] , \wAIn19[30] , 
        \wAIn19[29] , \wAIn19[28] , \wAIn19[27] , \wAIn19[26] , \wAIn19[25] , 
        \wAIn19[24] , \wAIn19[23] , \wAIn19[22] , \wAIn19[21] , \wAIn19[20] , 
        \wAIn19[19] , \wAIn19[18] , \wAIn19[17] , \wAIn19[16] , \wAIn19[15] , 
        \wAIn19[14] , \wAIn19[13] , \wAIn19[12] , \wAIn19[11] , \wAIn19[10] , 
        \wAIn19[9] , \wAIn19[8] , \wAIn19[7] , \wAIn19[6] , \wAIn19[5] , 
        \wAIn19[4] , \wAIn19[3] , \wAIn19[2] , \wAIn19[1] , \wAIn19[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_19 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink20[31] , \ScanLink20[30] , \ScanLink20[29] , 
        \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , \ScanLink20[25] , 
        \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , \ScanLink20[21] , 
        \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , \ScanLink20[17] , 
        \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , \ScanLink20[13] , 
        \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , \ScanLink20[9] , 
        \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , \ScanLink20[5] , 
        \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , \ScanLink20[1] , 
        \ScanLink20[0] }), .ScanOut({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA22[31] , \wRegInA22[30] , 
        \wRegInA22[29] , \wRegInA22[28] , \wRegInA22[27] , \wRegInA22[26] , 
        \wRegInA22[25] , \wRegInA22[24] , \wRegInA22[23] , \wRegInA22[22] , 
        \wRegInA22[21] , \wRegInA22[20] , \wRegInA22[19] , \wRegInA22[18] , 
        \wRegInA22[17] , \wRegInA22[16] , \wRegInA22[15] , \wRegInA22[14] , 
        \wRegInA22[13] , \wRegInA22[12] , \wRegInA22[11] , \wRegInA22[10] , 
        \wRegInA22[9] , \wRegInA22[8] , \wRegInA22[7] , \wRegInA22[6] , 
        \wRegInA22[5] , \wRegInA22[4] , \wRegInA22[3] , \wRegInA22[2] , 
        \wRegInA22[1] , \wRegInA22[0] }), .Out({\wAIn22[31] , \wAIn22[30] , 
        \wAIn22[29] , \wAIn22[28] , \wAIn22[27] , \wAIn22[26] , \wAIn22[25] , 
        \wAIn22[24] , \wAIn22[23] , \wAIn22[22] , \wAIn22[21] , \wAIn22[20] , 
        \wAIn22[19] , \wAIn22[18] , \wAIn22[17] , \wAIn22[16] , \wAIn22[15] , 
        \wAIn22[14] , \wAIn22[13] , \wAIn22[12] , \wAIn22[11] , \wAIn22[10] , 
        \wAIn22[9] , \wAIn22[8] , \wAIn22[7] , \wAIn22[6] , \wAIn22[5] , 
        \wAIn22[4] , \wAIn22[3] , \wAIn22[2] , \wAIn22[1] , \wAIn22[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_8 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[31] , \ScanLink9[30] , \ScanLink9[29] , 
        \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , \ScanLink9[25] , 
        \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , \ScanLink9[21] , 
        \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , \ScanLink9[17] , 
        \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , \ScanLink9[13] , 
        \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , \ScanLink9[9] , 
        \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB27[31] , \wRegInB27[30] , 
        \wRegInB27[29] , \wRegInB27[28] , \wRegInB27[27] , \wRegInB27[26] , 
        \wRegInB27[25] , \wRegInB27[24] , \wRegInB27[23] , \wRegInB27[22] , 
        \wRegInB27[21] , \wRegInB27[20] , \wRegInB27[19] , \wRegInB27[18] , 
        \wRegInB27[17] , \wRegInB27[16] , \wRegInB27[15] , \wRegInB27[14] , 
        \wRegInB27[13] , \wRegInB27[12] , \wRegInB27[11] , \wRegInB27[10] , 
        \wRegInB27[9] , \wRegInB27[8] , \wRegInB27[7] , \wRegInB27[6] , 
        \wRegInB27[5] , \wRegInB27[4] , \wRegInB27[3] , \wRegInB27[2] , 
        \wRegInB27[1] , \wRegInB27[0] }), .Out({\wBIn27[31] , \wBIn27[30] , 
        \wBIn27[29] , \wBIn27[28] , \wBIn27[27] , \wBIn27[26] , \wBIn27[25] , 
        \wBIn27[24] , \wBIn27[23] , \wBIn27[22] , \wBIn27[21] , \wBIn27[20] , 
        \wBIn27[19] , \wBIn27[18] , \wBIn27[17] , \wBIn27[16] , \wBIn27[15] , 
        \wBIn27[14] , \wBIn27[13] , \wBIn27[12] , \wBIn27[11] , \wBIn27[10] , 
        \wBIn27[9] , \wBIn27[8] , \wBIn27[7] , \wBIn27[6] , \wBIn27[5] , 
        \wBIn27[4] , \wBIn27[3] , \wBIn27[2] , \wBIn27[1] , \wBIn27[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAIn6[31] , 
        \wAIn6[30] , \wAIn6[29] , \wAIn6[28] , \wAIn6[27] , \wAIn6[26] , 
        \wAIn6[25] , \wAIn6[24] , \wAIn6[23] , \wAIn6[22] , \wAIn6[21] , 
        \wAIn6[20] , \wAIn6[19] , \wAIn6[18] , \wAIn6[17] , \wAIn6[16] , 
        \wAIn6[15] , \wAIn6[14] , \wAIn6[13] , \wAIn6[12] , \wAIn6[11] , 
        \wAIn6[10] , \wAIn6[9] , \wAIn6[8] , \wAIn6[7] , \wAIn6[6] , 
        \wAIn6[5] , \wAIn6[4] , \wAIn6[3] , \wAIn6[2] , \wAIn6[1] , \wAIn6[0] 
        }), .BIn({\wBIn6[31] , \wBIn6[30] , \wBIn6[29] , \wBIn6[28] , 
        \wBIn6[27] , \wBIn6[26] , \wBIn6[25] , \wBIn6[24] , \wBIn6[23] , 
        \wBIn6[22] , \wBIn6[21] , \wBIn6[20] , \wBIn6[19] , \wBIn6[18] , 
        \wBIn6[17] , \wBIn6[16] , \wBIn6[15] , \wBIn6[14] , \wBIn6[13] , 
        \wBIn6[12] , \wBIn6[11] , \wBIn6[10] , \wBIn6[9] , \wBIn6[8] , 
        \wBIn6[7] , \wBIn6[6] , \wBIn6[5] , \wBIn6[4] , \wBIn6[3] , \wBIn6[2] , 
        \wBIn6[1] , \wBIn6[0] }), .HiOut({\wBMid5[31] , \wBMid5[30] , 
        \wBMid5[29] , \wBMid5[28] , \wBMid5[27] , \wBMid5[26] , \wBMid5[25] , 
        \wBMid5[24] , \wBMid5[23] , \wBMid5[22] , \wBMid5[21] , \wBMid5[20] , 
        \wBMid5[19] , \wBMid5[18] , \wBMid5[17] , \wBMid5[16] , \wBMid5[15] , 
        \wBMid5[14] , \wBMid5[13] , \wBMid5[12] , \wBMid5[11] , \wBMid5[10] , 
        \wBMid5[9] , \wBMid5[8] , \wBMid5[7] , \wBMid5[6] , \wBMid5[5] , 
        \wBMid5[4] , \wBMid5[3] , \wBMid5[2] , \wBMid5[1] , \wBMid5[0] }), 
        .LoOut({\wAMid6[31] , \wAMid6[30] , \wAMid6[29] , \wAMid6[28] , 
        \wAMid6[27] , \wAMid6[26] , \wAMid6[25] , \wAMid6[24] , \wAMid6[23] , 
        \wAMid6[22] , \wAMid6[21] , \wAMid6[20] , \wAMid6[19] , \wAMid6[18] , 
        \wAMid6[17] , \wAMid6[16] , \wAMid6[15] , \wAMid6[14] , \wAMid6[13] , 
        \wAMid6[12] , \wAMid6[11] , \wAMid6[10] , \wAMid6[9] , \wAMid6[8] , 
        \wAMid6[7] , \wAMid6[6] , \wAMid6[5] , \wAMid6[4] , \wAMid6[3] , 
        \wAMid6[2] , \wAMid6[1] , \wAMid6[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn10[31] , \wAIn10[30] , \wAIn10[29] , \wAIn10[28] , \wAIn10[27] , 
        \wAIn10[26] , \wAIn10[25] , \wAIn10[24] , \wAIn10[23] , \wAIn10[22] , 
        \wAIn10[21] , \wAIn10[20] , \wAIn10[19] , \wAIn10[18] , \wAIn10[17] , 
        \wAIn10[16] , \wAIn10[15] , \wAIn10[14] , \wAIn10[13] , \wAIn10[12] , 
        \wAIn10[11] , \wAIn10[10] , \wAIn10[9] , \wAIn10[8] , \wAIn10[7] , 
        \wAIn10[6] , \wAIn10[5] , \wAIn10[4] , \wAIn10[3] , \wAIn10[2] , 
        \wAIn10[1] , \wAIn10[0] }), .BIn({\wBIn10[31] , \wBIn10[30] , 
        \wBIn10[29] , \wBIn10[28] , \wBIn10[27] , \wBIn10[26] , \wBIn10[25] , 
        \wBIn10[24] , \wBIn10[23] , \wBIn10[22] , \wBIn10[21] , \wBIn10[20] , 
        \wBIn10[19] , \wBIn10[18] , \wBIn10[17] , \wBIn10[16] , \wBIn10[15] , 
        \wBIn10[14] , \wBIn10[13] , \wBIn10[12] , \wBIn10[11] , \wBIn10[10] , 
        \wBIn10[9] , \wBIn10[8] , \wBIn10[7] , \wBIn10[6] , \wBIn10[5] , 
        \wBIn10[4] , \wBIn10[3] , \wBIn10[2] , \wBIn10[1] , \wBIn10[0] }), 
        .HiOut({\wBMid9[31] , \wBMid9[30] , \wBMid9[29] , \wBMid9[28] , 
        \wBMid9[27] , \wBMid9[26] , \wBMid9[25] , \wBMid9[24] , \wBMid9[23] , 
        \wBMid9[22] , \wBMid9[21] , \wBMid9[20] , \wBMid9[19] , \wBMid9[18] , 
        \wBMid9[17] , \wBMid9[16] , \wBMid9[15] , \wBMid9[14] , \wBMid9[13] , 
        \wBMid9[12] , \wBMid9[11] , \wBMid9[10] , \wBMid9[9] , \wBMid9[8] , 
        \wBMid9[7] , \wBMid9[6] , \wBMid9[5] , \wBMid9[4] , \wBMid9[3] , 
        \wBMid9[2] , \wBMid9[1] , \wBMid9[0] }), .LoOut({\wAMid10[31] , 
        \wAMid10[30] , \wAMid10[29] , \wAMid10[28] , \wAMid10[27] , 
        \wAMid10[26] , \wAMid10[25] , \wAMid10[24] , \wAMid10[23] , 
        \wAMid10[22] , \wAMid10[21] , \wAMid10[20] , \wAMid10[19] , 
        \wAMid10[18] , \wAMid10[17] , \wAMid10[16] , \wAMid10[15] , 
        \wAMid10[14] , \wAMid10[13] , \wAMid10[12] , \wAMid10[11] , 
        \wAMid10[10] , \wAMid10[9] , \wAMid10[8] , \wAMid10[7] , \wAMid10[6] , 
        \wAMid10[5] , \wAMid10[4] , \wAMid10[3] , \wAMid10[2] , \wAMid10[1] , 
        \wAMid10[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn17[31] , \wAIn17[30] , \wAIn17[29] , \wAIn17[28] , \wAIn17[27] , 
        \wAIn17[26] , \wAIn17[25] , \wAIn17[24] , \wAIn17[23] , \wAIn17[22] , 
        \wAIn17[21] , \wAIn17[20] , \wAIn17[19] , \wAIn17[18] , \wAIn17[17] , 
        \wAIn17[16] , \wAIn17[15] , \wAIn17[14] , \wAIn17[13] , \wAIn17[12] , 
        \wAIn17[11] , \wAIn17[10] , \wAIn17[9] , \wAIn17[8] , \wAIn17[7] , 
        \wAIn17[6] , \wAIn17[5] , \wAIn17[4] , \wAIn17[3] , \wAIn17[2] , 
        \wAIn17[1] , \wAIn17[0] }), .BIn({\wBIn17[31] , \wBIn17[30] , 
        \wBIn17[29] , \wBIn17[28] , \wBIn17[27] , \wBIn17[26] , \wBIn17[25] , 
        \wBIn17[24] , \wBIn17[23] , \wBIn17[22] , \wBIn17[21] , \wBIn17[20] , 
        \wBIn17[19] , \wBIn17[18] , \wBIn17[17] , \wBIn17[16] , \wBIn17[15] , 
        \wBIn17[14] , \wBIn17[13] , \wBIn17[12] , \wBIn17[11] , \wBIn17[10] , 
        \wBIn17[9] , \wBIn17[8] , \wBIn17[7] , \wBIn17[6] , \wBIn17[5] , 
        \wBIn17[4] , \wBIn17[3] , \wBIn17[2] , \wBIn17[1] , \wBIn17[0] }), 
        .HiOut({\wBMid16[31] , \wBMid16[30] , \wBMid16[29] , \wBMid16[28] , 
        \wBMid16[27] , \wBMid16[26] , \wBMid16[25] , \wBMid16[24] , 
        \wBMid16[23] , \wBMid16[22] , \wBMid16[21] , \wBMid16[20] , 
        \wBMid16[19] , \wBMid16[18] , \wBMid16[17] , \wBMid16[16] , 
        \wBMid16[15] , \wBMid16[14] , \wBMid16[13] , \wBMid16[12] , 
        \wBMid16[11] , \wBMid16[10] , \wBMid16[9] , \wBMid16[8] , \wBMid16[7] , 
        \wBMid16[6] , \wBMid16[5] , \wBMid16[4] , \wBMid16[3] , \wBMid16[2] , 
        \wBMid16[1] , \wBMid16[0] }), .LoOut({\wAMid17[31] , \wAMid17[30] , 
        \wAMid17[29] , \wAMid17[28] , \wAMid17[27] , \wAMid17[26] , 
        \wAMid17[25] , \wAMid17[24] , \wAMid17[23] , \wAMid17[22] , 
        \wAMid17[21] , \wAMid17[20] , \wAMid17[19] , \wAMid17[18] , 
        \wAMid17[17] , \wAMid17[16] , \wAMid17[15] , \wAMid17[14] , 
        \wAMid17[13] , \wAMid17[12] , \wAMid17[11] , \wAMid17[10] , 
        \wAMid17[9] , \wAMid17[8] , \wAMid17[7] , \wAMid17[6] , \wAMid17[5] , 
        \wAMid17[4] , \wAMid17[3] , \wAMid17[2] , \wAMid17[1] , \wAMid17[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn30[31] , \wAIn30[30] , \wAIn30[29] , \wAIn30[28] , \wAIn30[27] , 
        \wAIn30[26] , \wAIn30[25] , \wAIn30[24] , \wAIn30[23] , \wAIn30[22] , 
        \wAIn30[21] , \wAIn30[20] , \wAIn30[19] , \wAIn30[18] , \wAIn30[17] , 
        \wAIn30[16] , \wAIn30[15] , \wAIn30[14] , \wAIn30[13] , \wAIn30[12] , 
        \wAIn30[11] , \wAIn30[10] , \wAIn30[9] , \wAIn30[8] , \wAIn30[7] , 
        \wAIn30[6] , \wAIn30[5] , \wAIn30[4] , \wAIn30[3] , \wAIn30[2] , 
        \wAIn30[1] , \wAIn30[0] }), .BIn({\wBIn30[31] , \wBIn30[30] , 
        \wBIn30[29] , \wBIn30[28] , \wBIn30[27] , \wBIn30[26] , \wBIn30[25] , 
        \wBIn30[24] , \wBIn30[23] , \wBIn30[22] , \wBIn30[21] , \wBIn30[20] , 
        \wBIn30[19] , \wBIn30[18] , \wBIn30[17] , \wBIn30[16] , \wBIn30[15] , 
        \wBIn30[14] , \wBIn30[13] , \wBIn30[12] , \wBIn30[11] , \wBIn30[10] , 
        \wBIn30[9] , \wBIn30[8] , \wBIn30[7] , \wBIn30[6] , \wBIn30[5] , 
        \wBIn30[4] , \wBIn30[3] , \wBIn30[2] , \wBIn30[1] , \wBIn30[0] }), 
        .HiOut({\wBMid29[31] , \wBMid29[30] , \wBMid29[29] , \wBMid29[28] , 
        \wBMid29[27] , \wBMid29[26] , \wBMid29[25] , \wBMid29[24] , 
        \wBMid29[23] , \wBMid29[22] , \wBMid29[21] , \wBMid29[20] , 
        \wBMid29[19] , \wBMid29[18] , \wBMid29[17] , \wBMid29[16] , 
        \wBMid29[15] , \wBMid29[14] , \wBMid29[13] , \wBMid29[12] , 
        \wBMid29[11] , \wBMid29[10] , \wBMid29[9] , \wBMid29[8] , \wBMid29[7] , 
        \wBMid29[6] , \wBMid29[5] , \wBMid29[4] , \wBMid29[3] , \wBMid29[2] , 
        \wBMid29[1] , \wBMid29[0] }), .LoOut({\wAMid30[31] , \wAMid30[30] , 
        \wAMid30[29] , \wAMid30[28] , \wAMid30[27] , \wAMid30[26] , 
        \wAMid30[25] , \wAMid30[24] , \wAMid30[23] , \wAMid30[22] , 
        \wAMid30[21] , \wAMid30[20] , \wAMid30[19] , \wAMid30[18] , 
        \wAMid30[17] , \wAMid30[16] , \wAMid30[15] , \wAMid30[14] , 
        \wAMid30[13] , \wAMid30[12] , \wAMid30[11] , \wAMid30[10] , 
        \wAMid30[9] , \wAMid30[8] , \wAMid30[7] , \wAMid30[6] , \wAMid30[5] , 
        \wAMid30[4] , \wAMid30[3] , \wAMid30[2] , \wAMid30[1] , \wAMid30[0] })
         );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_59 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink60[31] , \ScanLink60[30] , \ScanLink60[29] , 
        \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , \ScanLink60[25] , 
        \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , \ScanLink60[21] , 
        \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , \ScanLink60[17] , 
        \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , \ScanLink60[13] , 
        \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , \ScanLink60[9] , 
        \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , \ScanLink60[5] , 
        \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , \ScanLink60[1] , 
        \ScanLink60[0] }), .ScanOut({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA2[31] , \wRegInA2[30] , 
        \wRegInA2[29] , \wRegInA2[28] , \wRegInA2[27] , \wRegInA2[26] , 
        \wRegInA2[25] , \wRegInA2[24] , \wRegInA2[23] , \wRegInA2[22] , 
        \wRegInA2[21] , \wRegInA2[20] , \wRegInA2[19] , \wRegInA2[18] , 
        \wRegInA2[17] , \wRegInA2[16] , \wRegInA2[15] , \wRegInA2[14] , 
        \wRegInA2[13] , \wRegInA2[12] , \wRegInA2[11] , \wRegInA2[10] , 
        \wRegInA2[9] , \wRegInA2[8] , \wRegInA2[7] , \wRegInA2[6] , 
        \wRegInA2[5] , \wRegInA2[4] , \wRegInA2[3] , \wRegInA2[2] , 
        \wRegInA2[1] , \wRegInA2[0] }), .Out({\wAIn2[31] , \wAIn2[30] , 
        \wAIn2[29] , \wAIn2[28] , \wAIn2[27] , \wAIn2[26] , \wAIn2[25] , 
        \wAIn2[24] , \wAIn2[23] , \wAIn2[22] , \wAIn2[21] , \wAIn2[20] , 
        \wAIn2[19] , \wAIn2[18] , \wAIn2[17] , \wAIn2[16] , \wAIn2[15] , 
        \wAIn2[14] , \wAIn2[13] , \wAIn2[12] , \wAIn2[11] , \wAIn2[10] , 
        \wAIn2[9] , \wAIn2[8] , \wAIn2[7] , \wAIn2[6] , \wAIn2[5] , \wAIn2[4] , 
        \wAIn2[3] , \wAIn2[2] , \wAIn2[1] , \wAIn2[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_37 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink38[31] , \ScanLink38[30] , \ScanLink38[29] , 
        \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , \ScanLink38[25] , 
        \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , \ScanLink38[21] , 
        \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , \ScanLink38[17] , 
        \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , \ScanLink38[13] , 
        \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , \ScanLink38[9] , 
        \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , \ScanLink38[5] , 
        \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , \ScanLink38[1] , 
        \ScanLink38[0] }), .ScanOut({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA13[31] , \wRegInA13[30] , 
        \wRegInA13[29] , \wRegInA13[28] , \wRegInA13[27] , \wRegInA13[26] , 
        \wRegInA13[25] , \wRegInA13[24] , \wRegInA13[23] , \wRegInA13[22] , 
        \wRegInA13[21] , \wRegInA13[20] , \wRegInA13[19] , \wRegInA13[18] , 
        \wRegInA13[17] , \wRegInA13[16] , \wRegInA13[15] , \wRegInA13[14] , 
        \wRegInA13[13] , \wRegInA13[12] , \wRegInA13[11] , \wRegInA13[10] , 
        \wRegInA13[9] , \wRegInA13[8] , \wRegInA13[7] , \wRegInA13[6] , 
        \wRegInA13[5] , \wRegInA13[4] , \wRegInA13[3] , \wRegInA13[2] , 
        \wRegInA13[1] , \wRegInA13[0] }), .Out({\wAIn13[31] , \wAIn13[30] , 
        \wAIn13[29] , \wAIn13[28] , \wAIn13[27] , \wAIn13[26] , \wAIn13[25] , 
        \wAIn13[24] , \wAIn13[23] , \wAIn13[22] , \wAIn13[21] , \wAIn13[20] , 
        \wAIn13[19] , \wAIn13[18] , \wAIn13[17] , \wAIn13[16] , \wAIn13[15] , 
        \wAIn13[14] , \wAIn13[13] , \wAIn13[12] , \wAIn13[11] , \wAIn13[10] , 
        \wAIn13[9] , \wAIn13[8] , \wAIn13[7] , \wAIn13[6] , \wAIn13[5] , 
        \wAIn13[4] , \wAIn13[3] , \wAIn13[2] , \wAIn13[1] , \wAIn13[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_10 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[31] , \ScanLink11[30] , \ScanLink11[29] , 
        \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , \ScanLink11[25] , 
        \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , \ScanLink11[21] , 
        \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , \ScanLink11[17] , 
        \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , \ScanLink11[13] , 
        \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , \ScanLink11[9] , 
        \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB26[31] , \wRegInB26[30] , 
        \wRegInB26[29] , \wRegInB26[28] , \wRegInB26[27] , \wRegInB26[26] , 
        \wRegInB26[25] , \wRegInB26[24] , \wRegInB26[23] , \wRegInB26[22] , 
        \wRegInB26[21] , \wRegInB26[20] , \wRegInB26[19] , \wRegInB26[18] , 
        \wRegInB26[17] , \wRegInB26[16] , \wRegInB26[15] , \wRegInB26[14] , 
        \wRegInB26[13] , \wRegInB26[12] , \wRegInB26[11] , \wRegInB26[10] , 
        \wRegInB26[9] , \wRegInB26[8] , \wRegInB26[7] , \wRegInB26[6] , 
        \wRegInB26[5] , \wRegInB26[4] , \wRegInB26[3] , \wRegInB26[2] , 
        \wRegInB26[1] , \wRegInB26[0] }), .Out({\wBIn26[31] , \wBIn26[30] , 
        \wBIn26[29] , \wBIn26[28] , \wBIn26[27] , \wBIn26[26] , \wBIn26[25] , 
        \wBIn26[24] , \wBIn26[23] , \wBIn26[22] , \wBIn26[21] , \wBIn26[20] , 
        \wBIn26[19] , \wBIn26[18] , \wBIn26[17] , \wBIn26[16] , \wBIn26[15] , 
        \wBIn26[14] , \wBIn26[13] , \wBIn26[12] , \wBIn26[11] , \wBIn26[10] , 
        \wBIn26[9] , \wBIn26[8] , \wBIn26[7] , \wBIn26[6] , \wBIn26[5] , 
        \wBIn26[4] , \wBIn26[3] , \wBIn26[2] , \wBIn26[1] , \wBIn26[0] }) );
    BubbleSort_Control_CWIDTH6_IDWIDTH1_WIDTH32_SCAN1 U_BSC ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink64[31] , 
        \ScanLink64[30] , \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , 
        \ScanLink64[26] , \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , 
        \ScanLink64[22] , \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , 
        \ScanLink64[18] , \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , 
        \ScanLink64[14] , \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , 
        \ScanLink64[10] , \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , 
        \ScanLink64[6] , \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , 
        \ScanLink64[2] , \ScanLink64[1] , \ScanLink64[0] }), .ScanEnable(
        \ScanEnable[0] ), .ScanId(1'b0), .Id(1'b1), .Enable(\wEnable[0] ) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_1 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[31] , \ScanLink2[30] , \ScanLink2[29] , 
        \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , \ScanLink2[25] , 
        \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , \ScanLink2[21] , 
        \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , \ScanLink2[17] , 
        \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , \ScanLink2[13] , 
        \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , \ScanLink2[9] , 
        \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA31[31] , \wRegInA31[30] , 
        \wRegInA31[29] , \wRegInA31[28] , \wRegInA31[27] , \wRegInA31[26] , 
        \wRegInA31[25] , \wRegInA31[24] , \wRegInA31[23] , \wRegInA31[22] , 
        \wRegInA31[21] , \wRegInA31[20] , \wRegInA31[19] , \wRegInA31[18] , 
        \wRegInA31[17] , \wRegInA31[16] , \wRegInA31[15] , \wRegInA31[14] , 
        \wRegInA31[13] , \wRegInA31[12] , \wRegInA31[11] , \wRegInA31[10] , 
        \wRegInA31[9] , \wRegInA31[8] , \wRegInA31[7] , \wRegInA31[6] , 
        \wRegInA31[5] , \wRegInA31[4] , \wRegInA31[3] , \wRegInA31[2] , 
        \wRegInA31[1] , \wRegInA31[0] }), .Out({\wAIn31[31] , \wAIn31[30] , 
        \wAIn31[29] , \wAIn31[28] , \wAIn31[27] , \wAIn31[26] , \wAIn31[25] , 
        \wAIn31[24] , \wAIn31[23] , \wAIn31[22] , \wAIn31[21] , \wAIn31[20] , 
        \wAIn31[19] , \wAIn31[18] , \wAIn31[17] , \wAIn31[16] , \wAIn31[15] , 
        \wAIn31[14] , \wAIn31[13] , \wAIn31[12] , \wAIn31[11] , \wAIn31[10] , 
        \wAIn31[9] , \wAIn31[8] , \wAIn31[7] , \wAIn31[6] , \wAIn31[5] , 
        \wAIn31[4] , \wAIn31[3] , \wAIn31[2] , \wAIn31[1] , \wAIn31[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid20[31] , \wAMid20[30] , \wAMid20[29] , \wAMid20[28] , 
        \wAMid20[27] , \wAMid20[26] , \wAMid20[25] , \wAMid20[24] , 
        \wAMid20[23] , \wAMid20[22] , \wAMid20[21] , \wAMid20[20] , 
        \wAMid20[19] , \wAMid20[18] , \wAMid20[17] , \wAMid20[16] , 
        \wAMid20[15] , \wAMid20[14] , \wAMid20[13] , \wAMid20[12] , 
        \wAMid20[11] , \wAMid20[10] , \wAMid20[9] , \wAMid20[8] , \wAMid20[7] , 
        \wAMid20[6] , \wAMid20[5] , \wAMid20[4] , \wAMid20[3] , \wAMid20[2] , 
        \wAMid20[1] , \wAMid20[0] }), .BIn({\wBMid20[31] , \wBMid20[30] , 
        \wBMid20[29] , \wBMid20[28] , \wBMid20[27] , \wBMid20[26] , 
        \wBMid20[25] , \wBMid20[24] , \wBMid20[23] , \wBMid20[22] , 
        \wBMid20[21] , \wBMid20[20] , \wBMid20[19] , \wBMid20[18] , 
        \wBMid20[17] , \wBMid20[16] , \wBMid20[15] , \wBMid20[14] , 
        \wBMid20[13] , \wBMid20[12] , \wBMid20[11] , \wBMid20[10] , 
        \wBMid20[9] , \wBMid20[8] , \wBMid20[7] , \wBMid20[6] , \wBMid20[5] , 
        \wBMid20[4] , \wBMid20[3] , \wBMid20[2] , \wBMid20[1] , \wBMid20[0] }), 
        .HiOut({\wRegInB20[31] , \wRegInB20[30] , \wRegInB20[29] , 
        \wRegInB20[28] , \wRegInB20[27] , \wRegInB20[26] , \wRegInB20[25] , 
        \wRegInB20[24] , \wRegInB20[23] , \wRegInB20[22] , \wRegInB20[21] , 
        \wRegInB20[20] , \wRegInB20[19] , \wRegInB20[18] , \wRegInB20[17] , 
        \wRegInB20[16] , \wRegInB20[15] , \wRegInB20[14] , \wRegInB20[13] , 
        \wRegInB20[12] , \wRegInB20[11] , \wRegInB20[10] , \wRegInB20[9] , 
        \wRegInB20[8] , \wRegInB20[7] , \wRegInB20[6] , \wRegInB20[5] , 
        \wRegInB20[4] , \wRegInB20[3] , \wRegInB20[2] , \wRegInB20[1] , 
        \wRegInB20[0] }), .LoOut({\wRegInA21[31] , \wRegInA21[30] , 
        \wRegInA21[29] , \wRegInA21[28] , \wRegInA21[27] , \wRegInA21[26] , 
        \wRegInA21[25] , \wRegInA21[24] , \wRegInA21[23] , \wRegInA21[22] , 
        \wRegInA21[21] , \wRegInA21[20] , \wRegInA21[19] , \wRegInA21[18] , 
        \wRegInA21[17] , \wRegInA21[16] , \wRegInA21[15] , \wRegInA21[14] , 
        \wRegInA21[13] , \wRegInA21[12] , \wRegInA21[11] , \wRegInA21[10] , 
        \wRegInA21[9] , \wRegInA21[8] , \wRegInA21[7] , \wRegInA21[6] , 
        \wRegInA21[5] , \wRegInA21[4] , \wRegInA21[3] , \wRegInA21[2] , 
        \wRegInA21[1] , \wRegInA21[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid27[31] , \wAMid27[30] , \wAMid27[29] , \wAMid27[28] , 
        \wAMid27[27] , \wAMid27[26] , \wAMid27[25] , \wAMid27[24] , 
        \wAMid27[23] , \wAMid27[22] , \wAMid27[21] , \wAMid27[20] , 
        \wAMid27[19] , \wAMid27[18] , \wAMid27[17] , \wAMid27[16] , 
        \wAMid27[15] , \wAMid27[14] , \wAMid27[13] , \wAMid27[12] , 
        \wAMid27[11] , \wAMid27[10] , \wAMid27[9] , \wAMid27[8] , \wAMid27[7] , 
        \wAMid27[6] , \wAMid27[5] , \wAMid27[4] , \wAMid27[3] , \wAMid27[2] , 
        \wAMid27[1] , \wAMid27[0] }), .BIn({\wBMid27[31] , \wBMid27[30] , 
        \wBMid27[29] , \wBMid27[28] , \wBMid27[27] , \wBMid27[26] , 
        \wBMid27[25] , \wBMid27[24] , \wBMid27[23] , \wBMid27[22] , 
        \wBMid27[21] , \wBMid27[20] , \wBMid27[19] , \wBMid27[18] , 
        \wBMid27[17] , \wBMid27[16] , \wBMid27[15] , \wBMid27[14] , 
        \wBMid27[13] , \wBMid27[12] , \wBMid27[11] , \wBMid27[10] , 
        \wBMid27[9] , \wBMid27[8] , \wBMid27[7] , \wBMid27[6] , \wBMid27[5] , 
        \wBMid27[4] , \wBMid27[3] , \wBMid27[2] , \wBMid27[1] , \wBMid27[0] }), 
        .HiOut({\wRegInB27[31] , \wRegInB27[30] , \wRegInB27[29] , 
        \wRegInB27[28] , \wRegInB27[27] , \wRegInB27[26] , \wRegInB27[25] , 
        \wRegInB27[24] , \wRegInB27[23] , \wRegInB27[22] , \wRegInB27[21] , 
        \wRegInB27[20] , \wRegInB27[19] , \wRegInB27[18] , \wRegInB27[17] , 
        \wRegInB27[16] , \wRegInB27[15] , \wRegInB27[14] , \wRegInB27[13] , 
        \wRegInB27[12] , \wRegInB27[11] , \wRegInB27[10] , \wRegInB27[9] , 
        \wRegInB27[8] , \wRegInB27[7] , \wRegInB27[6] , \wRegInB27[5] , 
        \wRegInB27[4] , \wRegInB27[3] , \wRegInB27[2] , \wRegInB27[1] , 
        \wRegInB27[0] }), .LoOut({\wRegInA28[31] , \wRegInA28[30] , 
        \wRegInA28[29] , \wRegInA28[28] , \wRegInA28[27] , \wRegInA28[26] , 
        \wRegInA28[25] , \wRegInA28[24] , \wRegInA28[23] , \wRegInA28[22] , 
        \wRegInA28[21] , \wRegInA28[20] , \wRegInA28[19] , \wRegInA28[18] , 
        \wRegInA28[17] , \wRegInA28[16] , \wRegInA28[15] , \wRegInA28[14] , 
        \wRegInA28[13] , \wRegInA28[12] , \wRegInA28[11] , \wRegInA28[10] , 
        \wRegInA28[9] , \wRegInA28[8] , \wRegInA28[7] , \wRegInA28[6] , 
        \wRegInA28[5] , \wRegInA28[4] , \wRegInA28[3] , \wRegInA28[2] , 
        \wRegInA28[1] , \wRegInA28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_42 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink43[31] , \ScanLink43[30] , \ScanLink43[29] , 
        \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , \ScanLink43[25] , 
        \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , \ScanLink43[21] , 
        \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , \ScanLink43[17] , 
        \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , \ScanLink43[13] , 
        \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , \ScanLink43[9] , 
        \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , \ScanLink43[5] , 
        \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , \ScanLink43[1] , 
        \ScanLink43[0] }), .ScanOut({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB10[31] , \wRegInB10[30] , 
        \wRegInB10[29] , \wRegInB10[28] , \wRegInB10[27] , \wRegInB10[26] , 
        \wRegInB10[25] , \wRegInB10[24] , \wRegInB10[23] , \wRegInB10[22] , 
        \wRegInB10[21] , \wRegInB10[20] , \wRegInB10[19] , \wRegInB10[18] , 
        \wRegInB10[17] , \wRegInB10[16] , \wRegInB10[15] , \wRegInB10[14] , 
        \wRegInB10[13] , \wRegInB10[12] , \wRegInB10[11] , \wRegInB10[10] , 
        \wRegInB10[9] , \wRegInB10[8] , \wRegInB10[7] , \wRegInB10[6] , 
        \wRegInB10[5] , \wRegInB10[4] , \wRegInB10[3] , \wRegInB10[2] , 
        \wRegInB10[1] , \wRegInB10[0] }), .Out({\wBIn10[31] , \wBIn10[30] , 
        \wBIn10[29] , \wBIn10[28] , \wBIn10[27] , \wBIn10[26] , \wBIn10[25] , 
        \wBIn10[24] , \wBIn10[23] , \wBIn10[22] , \wBIn10[21] , \wBIn10[20] , 
        \wBIn10[19] , \wBIn10[18] , \wBIn10[17] , \wBIn10[16] , \wBIn10[15] , 
        \wBIn10[14] , \wBIn10[13] , \wBIn10[12] , \wBIn10[11] , \wBIn10[10] , 
        \wBIn10[9] , \wBIn10[8] , \wBIn10[7] , \wBIn10[6] , \wBIn10[5] , 
        \wBIn10[4] , \wBIn10[3] , \wBIn10[2] , \wBIn10[1] , \wBIn10[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_45 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink46[31] , \ScanLink46[30] , \ScanLink46[29] , 
        \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , \ScanLink46[25] , 
        \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , \ScanLink46[21] , 
        \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , \ScanLink46[17] , 
        \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , \ScanLink46[13] , 
        \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , \ScanLink46[9] , 
        \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , \ScanLink46[5] , 
        \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , \ScanLink46[1] , 
        \ScanLink46[0] }), .ScanOut({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA9[31] , \wRegInA9[30] , 
        \wRegInA9[29] , \wRegInA9[28] , \wRegInA9[27] , \wRegInA9[26] , 
        \wRegInA9[25] , \wRegInA9[24] , \wRegInA9[23] , \wRegInA9[22] , 
        \wRegInA9[21] , \wRegInA9[20] , \wRegInA9[19] , \wRegInA9[18] , 
        \wRegInA9[17] , \wRegInA9[16] , \wRegInA9[15] , \wRegInA9[14] , 
        \wRegInA9[13] , \wRegInA9[12] , \wRegInA9[11] , \wRegInA9[10] , 
        \wRegInA9[9] , \wRegInA9[8] , \wRegInA9[7] , \wRegInA9[6] , 
        \wRegInA9[5] , \wRegInA9[4] , \wRegInA9[3] , \wRegInA9[2] , 
        \wRegInA9[1] , \wRegInA9[0] }), .Out({\wAIn9[31] , \wAIn9[30] , 
        \wAIn9[29] , \wAIn9[28] , \wAIn9[27] , \wAIn9[26] , \wAIn9[25] , 
        \wAIn9[24] , \wAIn9[23] , \wAIn9[22] , \wAIn9[21] , \wAIn9[20] , 
        \wAIn9[19] , \wAIn9[18] , \wAIn9[17] , \wAIn9[16] , \wAIn9[15] , 
        \wAIn9[14] , \wAIn9[13] , \wAIn9[12] , \wAIn9[11] , \wAIn9[10] , 
        \wAIn9[9] , \wAIn9[8] , \wAIn9[7] , \wAIn9[6] , \wAIn9[5] , \wAIn9[4] , 
        \wAIn9[3] , \wAIn9[2] , \wAIn9[1] , \wAIn9[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_62 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink63[31] , \ScanLink63[30] , \ScanLink63[29] , 
        \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , \ScanLink63[25] , 
        \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , \ScanLink63[21] , 
        \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , \ScanLink63[17] , 
        \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , \ScanLink63[13] , 
        \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , \ScanLink63[9] , 
        \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , \ScanLink63[5] , 
        \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , \ScanLink63[1] , 
        \ScanLink63[0] }), .ScanOut({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB0[31] , \wRegInB0[30] , 
        \wRegInB0[29] , \wRegInB0[28] , \wRegInB0[27] , \wRegInB0[26] , 
        \wRegInB0[25] , \wRegInB0[24] , \wRegInB0[23] , \wRegInB0[22] , 
        \wRegInB0[21] , \wRegInB0[20] , \wRegInB0[19] , \wRegInB0[18] , 
        \wRegInB0[17] , \wRegInB0[16] , \wRegInB0[15] , \wRegInB0[14] , 
        \wRegInB0[13] , \wRegInB0[12] , \wRegInB0[11] , \wRegInB0[10] , 
        \wRegInB0[9] , \wRegInB0[8] , \wRegInB0[7] , \wRegInB0[6] , 
        \wRegInB0[5] , \wRegInB0[4] , \wRegInB0[3] , \wRegInB0[2] , 
        \wRegInB0[1] , \wRegInB0[0] }), .Out({\wBIn0[31] , \wBIn0[30] , 
        \wBIn0[29] , \wBIn0[28] , \wBIn0[27] , \wBIn0[26] , \wBIn0[25] , 
        \wBIn0[24] , \wBIn0[23] , \wBIn0[22] , \wBIn0[21] , \wBIn0[20] , 
        \wBIn0[19] , \wBIn0[18] , \wBIn0[17] , \wBIn0[16] , \wBIn0[15] , 
        \wBIn0[14] , \wBIn0[13] , \wBIn0[12] , \wBIn0[11] , \wBIn0[10] , 
        \wBIn0[9] , \wBIn0[8] , \wBIn0[7] , \wBIn0[6] , \wBIn0[5] , \wBIn0[4] , 
        \wBIn0[3] , \wBIn0[2] , \wBIn0[1] , \wBIn0[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_6 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[31] , \ScanLink7[30] , \ScanLink7[29] , 
        \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , \ScanLink7[25] , 
        \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , \ScanLink7[21] , 
        \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , \ScanLink7[17] , 
        \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , \ScanLink7[13] , 
        \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , \ScanLink7[9] , 
        \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB28[31] , \wRegInB28[30] , 
        \wRegInB28[29] , \wRegInB28[28] , \wRegInB28[27] , \wRegInB28[26] , 
        \wRegInB28[25] , \wRegInB28[24] , \wRegInB28[23] , \wRegInB28[22] , 
        \wRegInB28[21] , \wRegInB28[20] , \wRegInB28[19] , \wRegInB28[18] , 
        \wRegInB28[17] , \wRegInB28[16] , \wRegInB28[15] , \wRegInB28[14] , 
        \wRegInB28[13] , \wRegInB28[12] , \wRegInB28[11] , \wRegInB28[10] , 
        \wRegInB28[9] , \wRegInB28[8] , \wRegInB28[7] , \wRegInB28[6] , 
        \wRegInB28[5] , \wRegInB28[4] , \wRegInB28[3] , \wRegInB28[2] , 
        \wRegInB28[1] , \wRegInB28[0] }), .Out({\wBIn28[31] , \wBIn28[30] , 
        \wBIn28[29] , \wBIn28[28] , \wBIn28[27] , \wBIn28[26] , \wBIn28[25] , 
        \wBIn28[24] , \wBIn28[23] , \wBIn28[22] , \wBIn28[21] , \wBIn28[20] , 
        \wBIn28[19] , \wBIn28[18] , \wBIn28[17] , \wBIn28[16] , \wBIn28[15] , 
        \wBIn28[14] , \wBIn28[13] , \wBIn28[12] , \wBIn28[11] , \wBIn28[10] , 
        \wBIn28[9] , \wBIn28[8] , \wBIn28[7] , \wBIn28[6] , \wBIn28[5] , 
        \wBIn28[4] , \wBIn28[3] , \wBIn28[2] , \wBIn28[1] , \wBIn28[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_30 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink31[31] , \ScanLink31[30] , \ScanLink31[29] , 
        \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , \ScanLink31[25] , 
        \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , \ScanLink31[21] , 
        \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , \ScanLink31[17] , 
        \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , \ScanLink31[13] , 
        \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , \ScanLink31[9] , 
        \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , \ScanLink31[5] , 
        \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , \ScanLink31[1] , 
        \ScanLink31[0] }), .ScanOut({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB16[31] , \wRegInB16[30] , 
        \wRegInB16[29] , \wRegInB16[28] , \wRegInB16[27] , \wRegInB16[26] , 
        \wRegInB16[25] , \wRegInB16[24] , \wRegInB16[23] , \wRegInB16[22] , 
        \wRegInB16[21] , \wRegInB16[20] , \wRegInB16[19] , \wRegInB16[18] , 
        \wRegInB16[17] , \wRegInB16[16] , \wRegInB16[15] , \wRegInB16[14] , 
        \wRegInB16[13] , \wRegInB16[12] , \wRegInB16[11] , \wRegInB16[10] , 
        \wRegInB16[9] , \wRegInB16[8] , \wRegInB16[7] , \wRegInB16[6] , 
        \wRegInB16[5] , \wRegInB16[4] , \wRegInB16[3] , \wRegInB16[2] , 
        \wRegInB16[1] , \wRegInB16[0] }), .Out({\wBIn16[31] , \wBIn16[30] , 
        \wBIn16[29] , \wBIn16[28] , \wBIn16[27] , \wBIn16[26] , \wBIn16[25] , 
        \wBIn16[24] , \wBIn16[23] , \wBIn16[22] , \wBIn16[21] , \wBIn16[20] , 
        \wBIn16[19] , \wBIn16[18] , \wBIn16[17] , \wBIn16[16] , \wBIn16[15] , 
        \wBIn16[14] , \wBIn16[13] , \wBIn16[12] , \wBIn16[11] , \wBIn16[10] , 
        \wBIn16[9] , \wBIn16[8] , \wBIn16[7] , \wBIn16[6] , \wBIn16[5] , 
        \wBIn16[4] , \wBIn16[3] , \wBIn16[2] , \wBIn16[1] , \wBIn16[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_17 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink18[31] , \ScanLink18[30] , \ScanLink18[29] , 
        \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , \ScanLink18[25] , 
        \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , \ScanLink18[21] , 
        \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , \ScanLink18[17] , 
        \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , \ScanLink18[13] , 
        \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , \ScanLink18[9] , 
        \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , \ScanLink18[5] , 
        \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , \ScanLink18[1] , 
        \ScanLink18[0] }), .ScanOut({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA23[31] , \wRegInA23[30] , 
        \wRegInA23[29] , \wRegInA23[28] , \wRegInA23[27] , \wRegInA23[26] , 
        \wRegInA23[25] , \wRegInA23[24] , \wRegInA23[23] , \wRegInA23[22] , 
        \wRegInA23[21] , \wRegInA23[20] , \wRegInA23[19] , \wRegInA23[18] , 
        \wRegInA23[17] , \wRegInA23[16] , \wRegInA23[15] , \wRegInA23[14] , 
        \wRegInA23[13] , \wRegInA23[12] , \wRegInA23[11] , \wRegInA23[10] , 
        \wRegInA23[9] , \wRegInA23[8] , \wRegInA23[7] , \wRegInA23[6] , 
        \wRegInA23[5] , \wRegInA23[4] , \wRegInA23[3] , \wRegInA23[2] , 
        \wRegInA23[1] , \wRegInA23[0] }), .Out({\wAIn23[31] , \wAIn23[30] , 
        \wAIn23[29] , \wAIn23[28] , \wAIn23[27] , \wAIn23[26] , \wAIn23[25] , 
        \wAIn23[24] , \wAIn23[23] , \wAIn23[22] , \wAIn23[21] , \wAIn23[20] , 
        \wAIn23[19] , \wAIn23[18] , \wAIn23[17] , \wAIn23[16] , \wAIn23[15] , 
        \wAIn23[14] , \wAIn23[13] , \wAIn23[12] , \wAIn23[11] , \wAIn23[10] , 
        \wAIn23[9] , \wAIn23[8] , \wAIn23[7] , \wAIn23[6] , \wAIn23[5] , 
        \wAIn23[4] , \wAIn23[3] , \wAIn23[2] , \wAIn23[1] , \wAIn23[0] }) );
    BubbleSort_Node_WIDTH32 BSN1_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn19[31] , \wAIn19[30] , \wAIn19[29] , \wAIn19[28] , \wAIn19[27] , 
        \wAIn19[26] , \wAIn19[25] , \wAIn19[24] , \wAIn19[23] , \wAIn19[22] , 
        \wAIn19[21] , \wAIn19[20] , \wAIn19[19] , \wAIn19[18] , \wAIn19[17] , 
        \wAIn19[16] , \wAIn19[15] , \wAIn19[14] , \wAIn19[13] , \wAIn19[12] , 
        \wAIn19[11] , \wAIn19[10] , \wAIn19[9] , \wAIn19[8] , \wAIn19[7] , 
        \wAIn19[6] , \wAIn19[5] , \wAIn19[4] , \wAIn19[3] , \wAIn19[2] , 
        \wAIn19[1] , \wAIn19[0] }), .BIn({\wBIn19[31] , \wBIn19[30] , 
        \wBIn19[29] , \wBIn19[28] , \wBIn19[27] , \wBIn19[26] , \wBIn19[25] , 
        \wBIn19[24] , \wBIn19[23] , \wBIn19[22] , \wBIn19[21] , \wBIn19[20] , 
        \wBIn19[19] , \wBIn19[18] , \wBIn19[17] , \wBIn19[16] , \wBIn19[15] , 
        \wBIn19[14] , \wBIn19[13] , \wBIn19[12] , \wBIn19[11] , \wBIn19[10] , 
        \wBIn19[9] , \wBIn19[8] , \wBIn19[7] , \wBIn19[6] , \wBIn19[5] , 
        \wBIn19[4] , \wBIn19[3] , \wBIn19[2] , \wBIn19[1] , \wBIn19[0] }), 
        .HiOut({\wBMid18[31] , \wBMid18[30] , \wBMid18[29] , \wBMid18[28] , 
        \wBMid18[27] , \wBMid18[26] , \wBMid18[25] , \wBMid18[24] , 
        \wBMid18[23] , \wBMid18[22] , \wBMid18[21] , \wBMid18[20] , 
        \wBMid18[19] , \wBMid18[18] , \wBMid18[17] , \wBMid18[16] , 
        \wBMid18[15] , \wBMid18[14] , \wBMid18[13] , \wBMid18[12] , 
        \wBMid18[11] , \wBMid18[10] , \wBMid18[9] , \wBMid18[8] , \wBMid18[7] , 
        \wBMid18[6] , \wBMid18[5] , \wBMid18[4] , \wBMid18[3] , \wBMid18[2] , 
        \wBMid18[1] , \wBMid18[0] }), .LoOut({\wAMid19[31] , \wAMid19[30] , 
        \wAMid19[29] , \wAMid19[28] , \wAMid19[27] , \wAMid19[26] , 
        \wAMid19[25] , \wAMid19[24] , \wAMid19[23] , \wAMid19[22] , 
        \wAMid19[21] , \wAMid19[20] , \wAMid19[19] , \wAMid19[18] , 
        \wAMid19[17] , \wAMid19[16] , \wAMid19[15] , \wAMid19[14] , 
        \wAMid19[13] , \wAMid19[12] , \wAMid19[11] , \wAMid19[10] , 
        \wAMid19[9] , \wAMid19[8] , \wAMid19[7] , \wAMid19[6] , \wAMid19[5] , 
        \wAMid19[4] , \wAMid19[3] , \wAMid19[2] , \wAMid19[1] , \wAMid19[0] })
         );
    BubbleSort_Node_WIDTH32 BSN1_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAIn25[31] , \wAIn25[30] , \wAIn25[29] , \wAIn25[28] , \wAIn25[27] , 
        \wAIn25[26] , \wAIn25[25] , \wAIn25[24] , \wAIn25[23] , \wAIn25[22] , 
        \wAIn25[21] , \wAIn25[20] , \wAIn25[19] , \wAIn25[18] , \wAIn25[17] , 
        \wAIn25[16] , \wAIn25[15] , \wAIn25[14] , \wAIn25[13] , \wAIn25[12] , 
        \wAIn25[11] , \wAIn25[10] , \wAIn25[9] , \wAIn25[8] , \wAIn25[7] , 
        \wAIn25[6] , \wAIn25[5] , \wAIn25[4] , \wAIn25[3] , \wAIn25[2] , 
        \wAIn25[1] , \wAIn25[0] }), .BIn({\wBIn25[31] , \wBIn25[30] , 
        \wBIn25[29] , \wBIn25[28] , \wBIn25[27] , \wBIn25[26] , \wBIn25[25] , 
        \wBIn25[24] , \wBIn25[23] , \wBIn25[22] , \wBIn25[21] , \wBIn25[20] , 
        \wBIn25[19] , \wBIn25[18] , \wBIn25[17] , \wBIn25[16] , \wBIn25[15] , 
        \wBIn25[14] , \wBIn25[13] , \wBIn25[12] , \wBIn25[11] , \wBIn25[10] , 
        \wBIn25[9] , \wBIn25[8] , \wBIn25[7] , \wBIn25[6] , \wBIn25[5] , 
        \wBIn25[4] , \wBIn25[3] , \wBIn25[2] , \wBIn25[1] , \wBIn25[0] }), 
        .HiOut({\wBMid24[31] , \wBMid24[30] , \wBMid24[29] , \wBMid24[28] , 
        \wBMid24[27] , \wBMid24[26] , \wBMid24[25] , \wBMid24[24] , 
        \wBMid24[23] , \wBMid24[22] , \wBMid24[21] , \wBMid24[20] , 
        \wBMid24[19] , \wBMid24[18] , \wBMid24[17] , \wBMid24[16] , 
        \wBMid24[15] , \wBMid24[14] , \wBMid24[13] , \wBMid24[12] , 
        \wBMid24[11] , \wBMid24[10] , \wBMid24[9] , \wBMid24[8] , \wBMid24[7] , 
        \wBMid24[6] , \wBMid24[5] , \wBMid24[4] , \wBMid24[3] , \wBMid24[2] , 
        \wBMid24[1] , \wBMid24[0] }), .LoOut({\wAMid25[31] , \wAMid25[30] , 
        \wAMid25[29] , \wAMid25[28] , \wAMid25[27] , \wAMid25[26] , 
        \wAMid25[25] , \wAMid25[24] , \wAMid25[23] , \wAMid25[22] , 
        \wAMid25[21] , \wAMid25[20] , \wAMid25[19] , \wAMid25[18] , 
        \wAMid25[17] , \wAMid25[16] , \wAMid25[15] , \wAMid25[14] , 
        \wAMid25[13] , \wAMid25[12] , \wAMid25[11] , \wAMid25[10] , 
        \wAMid25[9] , \wAMid25[8] , \wAMid25[7] , \wAMid25[6] , \wAMid25[5] , 
        \wAMid25[4] , \wAMid25[3] , \wAMid25[2] , \wAMid25[1] , \wAMid25[0] })
         );
    BubbleSort_Node_WIDTH32 BSN2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR
        ), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({\wAMid3[31] , 
        \wAMid3[30] , \wAMid3[29] , \wAMid3[28] , \wAMid3[27] , \wAMid3[26] , 
        \wAMid3[25] , \wAMid3[24] , \wAMid3[23] , \wAMid3[22] , \wAMid3[21] , 
        \wAMid3[20] , \wAMid3[19] , \wAMid3[18] , \wAMid3[17] , \wAMid3[16] , 
        \wAMid3[15] , \wAMid3[14] , \wAMid3[13] , \wAMid3[12] , \wAMid3[11] , 
        \wAMid3[10] , \wAMid3[9] , \wAMid3[8] , \wAMid3[7] , \wAMid3[6] , 
        \wAMid3[5] , \wAMid3[4] , \wAMid3[3] , \wAMid3[2] , \wAMid3[1] , 
        \wAMid3[0] }), .BIn({\wBMid3[31] , \wBMid3[30] , \wBMid3[29] , 
        \wBMid3[28] , \wBMid3[27] , \wBMid3[26] , \wBMid3[25] , \wBMid3[24] , 
        \wBMid3[23] , \wBMid3[22] , \wBMid3[21] , \wBMid3[20] , \wBMid3[19] , 
        \wBMid3[18] , \wBMid3[17] , \wBMid3[16] , \wBMid3[15] , \wBMid3[14] , 
        \wBMid3[13] , \wBMid3[12] , \wBMid3[11] , \wBMid3[10] , \wBMid3[9] , 
        \wBMid3[8] , \wBMid3[7] , \wBMid3[6] , \wBMid3[5] , \wBMid3[4] , 
        \wBMid3[3] , \wBMid3[2] , \wBMid3[1] , \wBMid3[0] }), .HiOut({
        \wRegInB3[31] , \wRegInB3[30] , \wRegInB3[29] , \wRegInB3[28] , 
        \wRegInB3[27] , \wRegInB3[26] , \wRegInB3[25] , \wRegInB3[24] , 
        \wRegInB3[23] , \wRegInB3[22] , \wRegInB3[21] , \wRegInB3[20] , 
        \wRegInB3[19] , \wRegInB3[18] , \wRegInB3[17] , \wRegInB3[16] , 
        \wRegInB3[15] , \wRegInB3[14] , \wRegInB3[13] , \wRegInB3[12] , 
        \wRegInB3[11] , \wRegInB3[10] , \wRegInB3[9] , \wRegInB3[8] , 
        \wRegInB3[7] , \wRegInB3[6] , \wRegInB3[5] , \wRegInB3[4] , 
        \wRegInB3[3] , \wRegInB3[2] , \wRegInB3[1] , \wRegInB3[0] }), .LoOut({
        \wRegInA4[31] , \wRegInA4[30] , \wRegInA4[29] , \wRegInA4[28] , 
        \wRegInA4[27] , \wRegInA4[26] , \wRegInA4[25] , \wRegInA4[24] , 
        \wRegInA4[23] , \wRegInA4[22] , \wRegInA4[21] , \wRegInA4[20] , 
        \wRegInA4[19] , \wRegInA4[18] , \wRegInA4[17] , \wRegInA4[16] , 
        \wRegInA4[15] , \wRegInA4[14] , \wRegInA4[13] , \wRegInA4[12] , 
        \wRegInA4[11] , \wRegInA4[10] , \wRegInA4[9] , \wRegInA4[8] , 
        \wRegInA4[7] , \wRegInA4[6] , \wRegInA4[5] , \wRegInA4[4] , 
        \wRegInA4[3] , \wRegInA4[2] , \wRegInA4[1] , \wRegInA4[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid29[31] , \wAMid29[30] , \wAMid29[29] , \wAMid29[28] , 
        \wAMid29[27] , \wAMid29[26] , \wAMid29[25] , \wAMid29[24] , 
        \wAMid29[23] , \wAMid29[22] , \wAMid29[21] , \wAMid29[20] , 
        \wAMid29[19] , \wAMid29[18] , \wAMid29[17] , \wAMid29[16] , 
        \wAMid29[15] , \wAMid29[14] , \wAMid29[13] , \wAMid29[12] , 
        \wAMid29[11] , \wAMid29[10] , \wAMid29[9] , \wAMid29[8] , \wAMid29[7] , 
        \wAMid29[6] , \wAMid29[5] , \wAMid29[4] , \wAMid29[3] , \wAMid29[2] , 
        \wAMid29[1] , \wAMid29[0] }), .BIn({\wBMid29[31] , \wBMid29[30] , 
        \wBMid29[29] , \wBMid29[28] , \wBMid29[27] , \wBMid29[26] , 
        \wBMid29[25] , \wBMid29[24] , \wBMid29[23] , \wBMid29[22] , 
        \wBMid29[21] , \wBMid29[20] , \wBMid29[19] , \wBMid29[18] , 
        \wBMid29[17] , \wBMid29[16] , \wBMid29[15] , \wBMid29[14] , 
        \wBMid29[13] , \wBMid29[12] , \wBMid29[11] , \wBMid29[10] , 
        \wBMid29[9] , \wBMid29[8] , \wBMid29[7] , \wBMid29[6] , \wBMid29[5] , 
        \wBMid29[4] , \wBMid29[3] , \wBMid29[2] , \wBMid29[1] , \wBMid29[0] }), 
        .HiOut({\wRegInB29[31] , \wRegInB29[30] , \wRegInB29[29] , 
        \wRegInB29[28] , \wRegInB29[27] , \wRegInB29[26] , \wRegInB29[25] , 
        \wRegInB29[24] , \wRegInB29[23] , \wRegInB29[22] , \wRegInB29[21] , 
        \wRegInB29[20] , \wRegInB29[19] , \wRegInB29[18] , \wRegInB29[17] , 
        \wRegInB29[16] , \wRegInB29[15] , \wRegInB29[14] , \wRegInB29[13] , 
        \wRegInB29[12] , \wRegInB29[11] , \wRegInB29[10] , \wRegInB29[9] , 
        \wRegInB29[8] , \wRegInB29[7] , \wRegInB29[6] , \wRegInB29[5] , 
        \wRegInB29[4] , \wRegInB29[3] , \wRegInB29[2] , \wRegInB29[1] , 
        \wRegInB29[0] }), .LoOut({\wRegInA30[31] , \wRegInA30[30] , 
        \wRegInA30[29] , \wRegInA30[28] , \wRegInA30[27] , \wRegInA30[26] , 
        \wRegInA30[25] , \wRegInA30[24] , \wRegInA30[23] , \wRegInA30[22] , 
        \wRegInA30[21] , \wRegInA30[20] , \wRegInA30[19] , \wRegInA30[18] , 
        \wRegInA30[17] , \wRegInA30[16] , \wRegInA30[15] , \wRegInA30[14] , 
        \wRegInA30[13] , \wRegInA30[12] , \wRegInA30[11] , \wRegInA30[10] , 
        \wRegInA30[9] , \wRegInA30[8] , \wRegInA30[7] , \wRegInA30[6] , 
        \wRegInA30[5] , \wRegInA30[4] , \wRegInA30[3] , \wRegInA30[2] , 
        \wRegInA30[1] , \wRegInA30[0] }) );
    BubbleSort_Node_WIDTH32 BSN2_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(
        WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn({
        \wAMid15[31] , \wAMid15[30] , \wAMid15[29] , \wAMid15[28] , 
        \wAMid15[27] , \wAMid15[26] , \wAMid15[25] , \wAMid15[24] , 
        \wAMid15[23] , \wAMid15[22] , \wAMid15[21] , \wAMid15[20] , 
        \wAMid15[19] , \wAMid15[18] , \wAMid15[17] , \wAMid15[16] , 
        \wAMid15[15] , \wAMid15[14] , \wAMid15[13] , \wAMid15[12] , 
        \wAMid15[11] , \wAMid15[10] , \wAMid15[9] , \wAMid15[8] , \wAMid15[7] , 
        \wAMid15[6] , \wAMid15[5] , \wAMid15[4] , \wAMid15[3] , \wAMid15[2] , 
        \wAMid15[1] , \wAMid15[0] }), .BIn({\wBMid15[31] , \wBMid15[30] , 
        \wBMid15[29] , \wBMid15[28] , \wBMid15[27] , \wBMid15[26] , 
        \wBMid15[25] , \wBMid15[24] , \wBMid15[23] , \wBMid15[22] , 
        \wBMid15[21] , \wBMid15[20] , \wBMid15[19] , \wBMid15[18] , 
        \wBMid15[17] , \wBMid15[16] , \wBMid15[15] , \wBMid15[14] , 
        \wBMid15[13] , \wBMid15[12] , \wBMid15[11] , \wBMid15[10] , 
        \wBMid15[9] , \wBMid15[8] , \wBMid15[7] , \wBMid15[6] , \wBMid15[5] , 
        \wBMid15[4] , \wBMid15[3] , \wBMid15[2] , \wBMid15[1] , \wBMid15[0] }), 
        .HiOut({\wRegInB15[31] , \wRegInB15[30] , \wRegInB15[29] , 
        \wRegInB15[28] , \wRegInB15[27] , \wRegInB15[26] , \wRegInB15[25] , 
        \wRegInB15[24] , \wRegInB15[23] , \wRegInB15[22] , \wRegInB15[21] , 
        \wRegInB15[20] , \wRegInB15[19] , \wRegInB15[18] , \wRegInB15[17] , 
        \wRegInB15[16] , \wRegInB15[15] , \wRegInB15[14] , \wRegInB15[13] , 
        \wRegInB15[12] , \wRegInB15[11] , \wRegInB15[10] , \wRegInB15[9] , 
        \wRegInB15[8] , \wRegInB15[7] , \wRegInB15[6] , \wRegInB15[5] , 
        \wRegInB15[4] , \wRegInB15[3] , \wRegInB15[2] , \wRegInB15[1] , 
        \wRegInB15[0] }), .LoOut({\wRegInA16[31] , \wRegInA16[30] , 
        \wRegInA16[29] , \wRegInA16[28] , \wRegInA16[27] , \wRegInA16[26] , 
        \wRegInA16[25] , \wRegInA16[24] , \wRegInA16[23] , \wRegInA16[22] , 
        \wRegInA16[21] , \wRegInA16[20] , \wRegInA16[19] , \wRegInA16[18] , 
        \wRegInA16[17] , \wRegInA16[16] , \wRegInA16[15] , \wRegInA16[14] , 
        \wRegInA16[13] , \wRegInA16[12] , \wRegInA16[11] , \wRegInA16[10] , 
        \wRegInA16[9] , \wRegInA16[8] , \wRegInA16[7] , \wRegInA16[6] , 
        \wRegInA16[5] , \wRegInA16[4] , \wRegInA16[3] , \wRegInA16[2] , 
        \wRegInA16[1] , \wRegInA16[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_57 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink58[31] , \ScanLink58[30] , \ScanLink58[29] , 
        \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , \ScanLink58[25] , 
        \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , \ScanLink58[21] , 
        \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , \ScanLink58[17] , 
        \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , \ScanLink58[13] , 
        \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , \ScanLink58[9] , 
        \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , \ScanLink58[5] , 
        \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , \ScanLink58[1] , 
        \ScanLink58[0] }), .ScanOut({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA3[31] , \wRegInA3[30] , 
        \wRegInA3[29] , \wRegInA3[28] , \wRegInA3[27] , \wRegInA3[26] , 
        \wRegInA3[25] , \wRegInA3[24] , \wRegInA3[23] , \wRegInA3[22] , 
        \wRegInA3[21] , \wRegInA3[20] , \wRegInA3[19] , \wRegInA3[18] , 
        \wRegInA3[17] , \wRegInA3[16] , \wRegInA3[15] , \wRegInA3[14] , 
        \wRegInA3[13] , \wRegInA3[12] , \wRegInA3[11] , \wRegInA3[10] , 
        \wRegInA3[9] , \wRegInA3[8] , \wRegInA3[7] , \wRegInA3[6] , 
        \wRegInA3[5] , \wRegInA3[4] , \wRegInA3[3] , \wRegInA3[2] , 
        \wRegInA3[1] , \wRegInA3[0] }), .Out({\wAIn3[31] , \wAIn3[30] , 
        \wAIn3[29] , \wAIn3[28] , \wAIn3[27] , \wAIn3[26] , \wAIn3[25] , 
        \wAIn3[24] , \wAIn3[23] , \wAIn3[22] , \wAIn3[21] , \wAIn3[20] , 
        \wAIn3[19] , \wAIn3[18] , \wAIn3[17] , \wAIn3[16] , \wAIn3[15] , 
        \wAIn3[14] , \wAIn3[13] , \wAIn3[12] , \wAIn3[11] , \wAIn3[10] , 
        \wAIn3[9] , \wAIn3[8] , \wAIn3[7] , \wAIn3[6] , \wAIn3[5] , \wAIn3[4] , 
        \wAIn3[3] , \wAIn3[2] , \wAIn3[1] , \wAIn3[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_39 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink40[31] , \ScanLink40[30] , \ScanLink40[29] , 
        \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , \ScanLink40[25] , 
        \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , \ScanLink40[21] , 
        \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , \ScanLink40[17] , 
        \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , \ScanLink40[13] , 
        \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , \ScanLink40[9] , 
        \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , \ScanLink40[5] , 
        \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , \ScanLink40[1] , 
        \ScanLink40[0] }), .ScanOut({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInA12[31] , \wRegInA12[30] , 
        \wRegInA12[29] , \wRegInA12[28] , \wRegInA12[27] , \wRegInA12[26] , 
        \wRegInA12[25] , \wRegInA12[24] , \wRegInA12[23] , \wRegInA12[22] , 
        \wRegInA12[21] , \wRegInA12[20] , \wRegInA12[19] , \wRegInA12[18] , 
        \wRegInA12[17] , \wRegInA12[16] , \wRegInA12[15] , \wRegInA12[14] , 
        \wRegInA12[13] , \wRegInA12[12] , \wRegInA12[11] , \wRegInA12[10] , 
        \wRegInA12[9] , \wRegInA12[8] , \wRegInA12[7] , \wRegInA12[6] , 
        \wRegInA12[5] , \wRegInA12[4] , \wRegInA12[3] , \wRegInA12[2] , 
        \wRegInA12[1] , \wRegInA12[0] }), .Out({\wAIn12[31] , \wAIn12[30] , 
        \wAIn12[29] , \wAIn12[28] , \wAIn12[27] , \wAIn12[26] , \wAIn12[25] , 
        \wAIn12[24] , \wAIn12[23] , \wAIn12[22] , \wAIn12[21] , \wAIn12[20] , 
        \wAIn12[19] , \wAIn12[18] , \wAIn12[17] , \wAIn12[16] , \wAIn12[15] , 
        \wAIn12[14] , \wAIn12[13] , \wAIn12[12] , \wAIn12[11] , \wAIn12[10] , 
        \wAIn12[9] , \wAIn12[8] , \wAIn12[7] , \wAIn12[6] , \wAIn12[5] , 
        \wAIn12[4] , \wAIn12[3] , \wAIn12[2] , \wAIn12[1] , \wAIn12[0] }) );
    BubbleSort_Reg_WIDTH32_IDWIDTH1_SCAN1 U_BSR_22 ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink23[31] , \ScanLink23[30] , \ScanLink23[29] , 
        \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , \ScanLink23[25] , 
        \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , \ScanLink23[21] , 
        \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , \ScanLink23[17] , 
        \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , \ScanLink23[13] , 
        \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , \ScanLink23[9] , 
        \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , \ScanLink23[5] , 
        \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , \ScanLink23[1] , 
        \ScanLink23[0] }), .ScanOut({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(\ScanEnable[0] ), .Id(
        1'b0), .Enable(\wEnable[0] ), .In({\wRegInB20[31] , \wRegInB20[30] , 
        \wRegInB20[29] , \wRegInB20[28] , \wRegInB20[27] , \wRegInB20[26] , 
        \wRegInB20[25] , \wRegInB20[24] , \wRegInB20[23] , \wRegInB20[22] , 
        \wRegInB20[21] , \wRegInB20[20] , \wRegInB20[19] , \wRegInB20[18] , 
        \wRegInB20[17] , \wRegInB20[16] , \wRegInB20[15] , \wRegInB20[14] , 
        \wRegInB20[13] , \wRegInB20[12] , \wRegInB20[11] , \wRegInB20[10] , 
        \wRegInB20[9] , \wRegInB20[8] , \wRegInB20[7] , \wRegInB20[6] , 
        \wRegInB20[5] , \wRegInB20[4] , \wRegInB20[3] , \wRegInB20[2] , 
        \wRegInB20[1] , \wRegInB20[0] }), .Out({\wBIn20[31] , \wBIn20[30] , 
        \wBIn20[29] , \wBIn20[28] , \wBIn20[27] , \wBIn20[26] , \wBIn20[25] , 
        \wBIn20[24] , \wBIn20[23] , \wBIn20[22] , \wBIn20[21] , \wBIn20[20] , 
        \wBIn20[19] , \wBIn20[18] , \wBIn20[17] , \wBIn20[16] , \wBIn20[15] , 
        \wBIn20[14] , \wBIn20[13] , \wBIn20[12] , \wBIn20[11] , \wBIn20[10] , 
        \wBIn20[9] , \wBIn20[8] , \wBIn20[7] , \wBIn20[6] , \wBIn20[5] , 
        \wBIn20[4] , \wBIn20[3] , \wBIn20[2] , \wBIn20[1] , \wBIn20[0] }) );
endmodule

