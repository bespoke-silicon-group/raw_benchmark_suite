
module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_31 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15;
    VMW_NOR2 U3 ( .A(A[5]), .B(n15), .Z(LT_LE) );
    VMW_AND5 U4 ( .A(A[1]), .B(A[2]), .C(A[4]), .D(A[0]), .E(A[3]), .Z(n15) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_30 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n16;
    VMW_NOR4 U3 ( .A(n16), .B(A[0]), .C(A[2]), .D(A[1]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[5]), .B(A[4]), .C(A[3]), .Z(n16) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_29 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n17;
    VMW_NOR4 U3 ( .A(A[5]), .B(A[4]), .C(A[3]), .D(n17), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n17) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_28 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n18, n19;
    VMW_NOR2 U3 ( .A(n18), .B(A[5]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n19), .Z(n18) );
    VMW_OAI211 U4 ( .A(A[2]), .B(A[1]), .C(A[4]), .D(A[3]), .Z(n19) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_27 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n20, n21;
    VMW_NOR4 U3 ( .A(A[5]), .B(A[4]), .C(A[3]), .D(n20), .Z(LT_LE) );
    VMW_INV U5 ( .A(n21), .Z(n20) );
    VMW_OAI21 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .Z(n21) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_26 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n22;
    VMW_AOI211 U3 ( .A(A[3]), .B(n22), .C(A[4]), .D(A[5]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[2]), .B(A[1]), .Z(n22) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_25 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n23;
    VMW_NOR3 U3 ( .A(n23), .B(A[5]), .C(A[4]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[1]), .B(A[2]), .C(A[3]), .Z(n23) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_24 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n24, n25;
    VMW_AOI21 U3 ( .A(A[4]), .B(n24), .C(A[5]), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[2]), .B(n25), .C(A[3]), .Z(n24) );
    VMW_OR2 U4 ( .A(A[1]), .B(A[0]), .Z(n25) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_23 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n27, n26;
    VMW_NOR2 U3 ( .A(A[5]), .B(n26), .Z(LT_LE) );
    VMW_OR3 U5 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n27) );
    VMW_AND3 U4 ( .A(A[4]), .B(n27), .C(A[3]), .Z(n26) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_22 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n29, n28;
    VMW_NOR2 U3 ( .A(A[5]), .B(n28), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[1]), .B(A[0]), .Z(n29) );
    VMW_AND4 U4 ( .A(A[3]), .B(A[4]), .C(A[2]), .D(n29), .Z(n28) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_21 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR3 U3 ( .A(A[3]), .B(A[5]), .C(A[4]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_20 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n31, n30;
    VMW_AOI21 U3 ( .A(A[4]), .B(n30), .C(A[5]), .Z(LT_LE) );
    VMW_INV U5 ( .A(n31), .Z(n30) );
    VMW_AOI211 U4 ( .A(A[0]), .B(A[1]), .C(A[3]), .D(A[2]), .Z(n31) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_19 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI211 U3 ( .A(A[2]), .B(A[3]), .C(A[5]), .D(A[4]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_18 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n32;
    VMW_AOI211 U3 ( .A(A[0]), .B(A[1]), .C(n32), .D(A[2]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[5]), .B(A[4]), .C(A[3]), .Z(n32) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_17 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n33;
    VMW_NOR3 U3 ( .A(n33), .B(A[5]), .C(A[4]), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n33) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_16 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n35, n34;
    VMW_AOI21 U3 ( .A(A[4]), .B(n34), .C(A[5]), .Z(LT_LE) );
    VMW_OR2 U5 ( .A(A[3]), .B(n35), .Z(n34) );
    VMW_AND3 U4 ( .A(A[1]), .B(A[2]), .C(A[0]), .Z(n35) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_15 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n36;
    VMW_AOI21 U3 ( .A(A[4]), .B(n36), .C(A[5]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[3]), .B(A[2]), .C(A[1]), .Z(n36) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_14 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n37, n38;
    VMW_NOR3 U3 ( .A(A[4]), .B(A[5]), .C(n37), .Z(LT_LE) );
    VMW_INV U5 ( .A(n38), .Z(n37) );
    VMW_OAI211 U4 ( .A(A[1]), .B(A[0]), .C(A[2]), .D(A[3]), .Z(n38) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_13 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR5 U3 ( .A(A[2]), .B(A[1]), .C(A[3]), .D(A[5]), .E(A[4]), .Z(LT_LE)
         );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_12 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n39;
    VMW_NOR2 U3 ( .A(A[5]), .B(n39), .Z(LT_LE) );
    VMW_AND3 U4 ( .A(A[3]), .B(A[4]), .C(A[2]), .Z(n39) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_11 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_AOI21 U3 ( .A(A[3]), .B(A[4]), .C(A[5]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_10 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n40;
    VMW_AOI211 U3 ( .A(A[3]), .B(n40), .C(A[5]), .D(A[4]), .Z(LT_LE) );
    VMW_OR3 U4 ( .A(A[2]), .B(A[1]), .C(A[0]), .Z(n40) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_9 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n41;
    VMW_AOI21 U3 ( .A(A[4]), .B(n41), .C(A[5]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[1]), .B(A[2]), .C(A[3]), .Z(n41) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_8 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR4 U3 ( .A(A[5]), .B(A[4]), .C(A[3]), .D(A[2]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_7 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n42;
    VMW_AOI21 U3 ( .A(A[4]), .B(n42), .C(A[5]), .Z(LT_LE) );
    VMW_OR4 U4 ( .A(A[1]), .B(A[0]), .C(A[3]), .D(A[2]), .Z(n42) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_6 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n43;
    VMW_NOR2 U3 ( .A(A[5]), .B(n43), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[1]), .B(A[3]), .C(A[4]), .D(A[2]), .Z(n43) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_5 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    VMW_NOR2 U3 ( .A(A[5]), .B(A[4]), .Z(LT_LE) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_4 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n44;
    VMW_AOI211 U3 ( .A(A[3]), .B(n44), .C(A[4]), .D(A[5]), .Z(LT_LE) );
    VMW_AO21 U4 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n44) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_3 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n45;
    VMW_AOI21 U3 ( .A(A[4]), .B(n45), .C(A[5]), .Z(LT_LE) );
    VMW_OR2 U4 ( .A(A[3]), .B(A[2]), .Z(n45) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_2 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n47, n46;
    VMW_NOR2 U3 ( .A(A[5]), .B(n46), .Z(LT_LE) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(A[2]), .Z(n47) );
    VMW_AND3 U4 ( .A(A[4]), .B(n47), .C(A[3]), .Z(n46) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [5:0] A;
input  [5:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n48;
    VMW_NOR3 U3 ( .A(n48), .B(A[5]), .C(A[4]), .Z(LT_LE) );
    VMW_AND4 U4 ( .A(A[0]), .B(A[3]), .C(A[1]), .D(A[2]), .Z(n48) );
endmodule


module NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, CallIn, ReturnIn, ColIn, PDiagIn, 
    NDiagIn, CallOut, ReturnOut, ColOut, PDiagOut, NDiagOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [5:0] Id;
input  [31:0] ColIn;
output [31:0] ColOut;
input  [5:0] ScanIn;
output [5:0] ScanOut;
input  [31:0] NDiagIn;
output [31:0] PDiagOut;
output [31:0] NDiagOut;
input  [31:0] PDiagIn;
input  Clk, Reset, RD, WR, ScanEnable, CallIn, ReturnIn;
output CallOut, ReturnOut;
    wire \NDiagOut[0] , n2791, n2943, n2964, n2981, n2858, n2811, n2753, n2774, 
        n658, n2836, n2936, n2881, n2911, n2726, n2748, n2843, n2864, n2701, 
        n2958, n2734, n2798, n866, n2876, n2713, n2851, n2818, n546, n2924, 
        Logic11, n2888, n2893, n2903, n2918, n834, n2956, n2971, n2976, n2698, 
        n2708, n2741, n2803, n2766, n2824, n898, n514, n2783, n2951, n2728, 
        n946, n466, n2784, n738, n2823, n2938, n2761, n2746, n2804, n2838, 
        n914, n2894, n2904, n2923, n2714, n2856, n498, n2871, n2696, n2706, 
        n2733, n2844, n2978, n2863, n2721, n2886, n2916, n2931, n2768, n2754, 
        n2773, n2831, n2816, n2715, n2963, n2796, n2944, n2878, n786, n722, 
        n2732, n2857, n2870, n2839, n2895, n2905, n2922, n2939, n770, n2747, 
        n2760, n2822, n2805, n2729, n2957, n2970, n482, n2962, n2785, n2945, 
        n2755, n2772, n2797, n2830, n2879, n2817, n2769, n2887, n2917, n2930, 
        n2959, n2979, n2697, \n1108[3] , n2707, n2720, n2845, n2862, 
        \n1108[1] , n2700, n2727, n2842, n2865, n2880, n2937, n2910, n642, 
        n2749, n2980, n2810, n2752, n2775, n2837, n2965, n2790, n2942, n2699, 
        n2859, n610, n2709, n2977, ReturnOut1063, n2950, n2782, \n1108[5] , 
        n2889, n2919, n2740, n2802, n2767, n2825, n2819, n882, n2925, n2892, 
        n2902, n2712, n2735, n2799, n2850, n2877, n2719, n2967, n2982, 
        \n1108[4] , n2792, n2940, n2777, n2899, n802, n2909, n2812, n2835, 
        \n1108[0] , n2750, n2809, n2882, n2912, n2702, n2789, n2935, n2840, 
        n850, n2710, n2725, n2852, n2867, n2737, n2875, n690, n2949, n2890, 
        n2900, n2927, n2759, n2742, n2765, n562, n2800, n2827, n2955, n2975, 
        n2952, n2780, n2849, n530, n2972, n2787, n2745, n2869, n2762, n2807, 
        n2820, n2779, n2897, n2920, n2907, CallOut1070, n2969, n2717, n2730, 
        n2872, n930, n2855, n2985, n2695, \n1108[2] , n2722, n2860, n2705, 
        n2829, n2847, n2885, n2915, n2932, n2757, n2929, n2770, n2815, n2832, 
        n2739, n2960, n2795, n2947, n2873, n2968, n2731, n2716, n2854, n2744, 
        n706, n2778, n2896, n2906, n2921, n2806, n2821, n2763, n2954, n754, 
        n2786, n2973, n2961, n2738, n2868, n2794, n2946, n2984, n2928, n2756, 
        n2814, n2833, n2771, n2828, n2861, n2884, n2933, n2914, n2694, n2704, 
        n2723, n2788, n2846, n594, n2703, n2841, n2724, n2808, n2866, n2883, 
        n2913, n818, n2934, n2776, n2898, n2908, n2834, n2966, n2983, n2718, 
        n2813, n2751, n2974, n2793, n2941, n2781, n2953, n2764, n2848, n626, 
        n2801, n2826, n578, n2743, n2891, n2901, n2758, n674, n2926, n2853, 
        n2711, n2736, n2874, n2948;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 , 
	UNCONNECTED_5 , UNCONNECTED_6 , UNCONNECTED_7 , UNCONNECTED_8 , 
	UNCONNECTED_9 , UNCONNECTED_10 , UNCONNECTED_11 , UNCONNECTED_12 , 
	UNCONNECTED_13 , UNCONNECTED_14 , UNCONNECTED_15 , UNCONNECTED_16 , 
	UNCONNECTED_17 , UNCONNECTED_18 , UNCONNECTED_19 , UNCONNECTED_20 , 
	UNCONNECTED_21 , UNCONNECTED_22 , UNCONNECTED_23 , UNCONNECTED_24 , 
	UNCONNECTED_25 , UNCONNECTED_26 ;
    assign PDiagOut[31] = \NDiagOut[0] ;
    assign NDiagOut[0] = \NDiagOut[0] ;
    VMW_PULLDOWN U719 ( .Z(n2970) );
    VMW_PULLDOWN U725 ( .Z(n2976) );
    VMW_OR3 U840 ( .A(n2769), .B(n2772), .C(n2773), .Z(n2953) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_2 gt_104_4 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , Logic11, 
        Logic11}), .LEQ(n2956), .TC(n2956), .LT_LE(n530) );
    VMW_NAND2 U750 ( .A(n2711), .B(n2712), .Z(PDiagOut[23]) );
    VMW_OR2 U777 ( .A(ColIn[28]), .B(n2704), .Z(ColOut[28]) );
    VMW_OR2 U789 ( .A(ColIn[16]), .B(n2724), .Z(ColOut[16]) );
    VMW_OR4 U867 ( .A(n2833), .B(NDiagIn[14]), .C(ColIn[14]), .D(PDiagIn[14]), 
        .Z(n2832) );
    VMW_INV U1047 ( .A(PDiagIn[12]), .Z(n2729) );
    VMW_NAND2 U809 ( .A(n2706), .B(n2755), .Z(NDiagOut[28]) );
    VMW_NAND3 U882 ( .A(n2866), .B(n2783), .C(n2801), .Z(n2865) );
    VMW_MUX2I U912 ( .A(ScanOut[5]), .B(ScanIn[5]), .S(ScanEnable), .Z(n2695)
         );
    VMW_INV U1060 ( .A(NDiagIn[27]), .Z(n2755) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_24 gt_104_10 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        Logic11}), .LEQ(n2978), .TC(n2978), .LT_LE(n626) );
    VMW_OR2 U935 ( .A(n2912), .B(n2886), .Z(n2706) );
    VMW_NOR2 U999 ( .A(CallIn), .B(n882), .Z(n2926) );
    VMW_NAND2 U1029 ( .A(n2819), .B(n2942), .Z(n2944) );
    VMW_INV U1085 ( .A(n2768), .Z(n2767) );
    VMW_NAND2 U812 ( .A(n2712), .B(n2758), .Z(NDiagOut[25]) );
    VMW_OR2 U835 ( .A(NDiagIn[1]), .B(n2742), .Z(NDiagOut[2]) );
    VMW_AND4 U982 ( .A(n2918), .B(n2758), .C(n2746), .D(n2711), .Z(n2810) );
    VMW_OR2 U792 ( .A(ColIn[13]), .B(n2728), .Z(ColOut[13]) );
    VMW_NOR2 U899 ( .A(n2881), .B(n2884), .Z(n2888) );
    VMW_NAND4 U909 ( .A(n2898), .B(n2765), .C(n2753), .D(n2739), .Z(n2897) );
    VMW_OR4 U1015 ( .A(NDiagIn[31]), .B(n2780), .C(ColIn[31]), .D(PDiagIn[31]), 
        .Z(n2902) );
    VMW_AO21 U1032 ( .A(n2946), .B(n2862), .C(n2947), .Z(n2812) );
    VMW_NAND4 U967 ( .A(n2913), .B(n2763), .C(n2751), .D(n2725), .Z(n2817) );
    VMW_OR2 U940 ( .A(n2830), .B(n2887), .Z(n2716) );
    VMW_PULLDOWN U705 ( .Z(n2956) );
    VMW_PULLDOWN U710 ( .Z(n2961) );
    VMW_NAND2 U742 ( .A(n2694), .B(n2700), .Z(\n1108[0] ) );
    VMW_OR2 U765 ( .A(n2733), .B(PDiagIn[9]), .Z(PDiagOut[8]) );
    VMW_NAND2 U780 ( .A(n2710), .B(n2745), .Z(ColOut[25]) );
    VMW_AOI211 U849 ( .A(n2796), .B(n2797), .C(n2798), .D(n2799), .Z(n2795) );
    VMW_NAND4 U975 ( .A(n2915), .B(n2762), .C(n2750), .D(n2719), .Z(n2845) );
    VMW_INV U1069 ( .A(NDiagIn[12]), .Z(n2764) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_19 gt_104_19 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , UNCONNECTED_1, 
        UNCONNECTED_2}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2973), .TC(n2973), .LT_LE(n770)
         );
    VMW_NOR2 U952 ( .A(n2829), .B(n2830), .Z(n2732) );
    VMW_OR4 U1007 ( .A(n2930), .B(NDiagIn[7]), .C(ColIn[7]), .D(PDiagIn[7]), 
        .Z(n2863) );
    VMW_OAI211 U1020 ( .A(n2809), .B(n2849), .C(n2817), .D(n2834), .Z(n2903)
         );
    VMW_OR2 U800 ( .A(ColIn[5]), .B(n2737), .Z(ColOut[5]) );
    VMW_OR2 U827 ( .A(NDiagIn[9]), .B(n2733), .Z(NDiagOut[10]) );
    VMW_NOR2 U990 ( .A(CallIn), .B(n754), .Z(n2901) );
    VMW_NAND2 U759 ( .A(n2725), .B(n2726), .Z(PDiagOut[14]) );
    VMW_AOI211 U852 ( .A(n2807), .B(n2808), .C(n2809), .D(n2810), .Z(n2806) );
    VMW_OR2 U890 ( .A(ScanOut[1]), .B(ScanOut[0]), .Z(n2878) );
    VMW_INV U1097 ( .A(n2933), .Z(n2861) );
    VMW_NOR2 U900 ( .A(n2767), .B(n2890), .Z(n2889) );
    VMW_AO21 U927 ( .A(n2816), .B(n2906), .C(n2859), .Z(n2803) );
    VMW_NOR2 U949 ( .A(n2825), .B(n2877), .Z(n2728) );
    VMW_INV U1055 ( .A(ColIn[21]), .Z(n2749) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_25 gt_104_25 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_3}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11, \NDiagOut[0] }), .LEQ(n2979), .TC(n2979), .LT_LE(
        n866) );
    VMW_INV U1072 ( .A(ReturnIn), .Z(n2876) );
    VMW_PULLDOWN U717 ( .Z(n2968) );
    VMW_PULLDOWN U730 ( .Z(n2981) );
    VMW_NAND2 U737 ( .A(n2694), .B(n2695), .Z(\n1108[5] ) );
    VMW_NAND3 U872 ( .A(n2847), .B(n2817), .C(n2848), .Z(n2846) );
    VMW_NAND2 U875 ( .A(n2851), .B(n2852), .Z(n2797) );
    VMW_NOR4 U969 ( .A(n2914), .B(NDiagIn[16]), .C(ColIn[16]), .D(PDiagIn[16]), 
        .Z(n2841) );
    VMW_INV U1075 ( .A(n2834), .Z(n2874) );
    VMW_INV U1052 ( .A(ColIn[24]), .Z(n2746) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_10 gt_104_22 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11}), .LEQ(n2964), .TC(n2964), .LT_LE(n818) );
    VMW_PULLDOWN U722 ( .Z(n2973) );
    VMW_NAND2 U739 ( .A(n2694), .B(n2697), .Z(\n1108[3] ) );
    VMW_OR2 U745 ( .A(n2703), .B(PDiagIn[29]), .Z(PDiagOut[28]) );
    VMW_NAND2 U779 ( .A(n2708), .B(n2744), .Z(ColOut[26]) );
    VMW_AND5 U855 ( .A(n2816), .B(n2817), .C(n2818), .D(n2767), .E(n2819), .Z(
        n2778) );
    VMW_OR2 U897 ( .A(n2827), .B(n2881), .Z(n2886) );
    VMW_OR4 U907 ( .A(n2895), .B(NDiagIn[18]), .C(ColIn[18]), .D(PDiagIn[18]), 
        .Z(n2894) );
    VMW_AO22 U920 ( .A(n2890), .B(ScanOut[4]), .C(n2889), .D(ScanIn[4]), .Z(
        n2779) );
    VMW_INV U1090 ( .A(n2897), .Z(n2860) );
    VMW_NOR4 U1000 ( .A(n2926), .B(NDiagIn[5]), .C(ColIn[5]), .D(PDiagIn[5]), 
        .Z(n2856) );
    VMW_AO21 U1027 ( .A(n2847), .B(n2940), .C(n2839), .Z(n2941) );
    VMW_NAND2 U762 ( .A(n2729), .B(n2730), .Z(PDiagOut[11]) );
    VMW_OR2 U807 ( .A(NDiagIn[29]), .B(n2703), .Z(NDiagOut[30]) );
    VMW_NOR2 U997 ( .A(CallIn), .B(n802), .Z(n2925) );
    VMW_OR2 U820 ( .A(NDiagIn[16]), .B(n2724), .Z(NDiagOut[17]) );
    VMW_OR2 U787 ( .A(ColIn[18]), .B(n2722), .Z(ColOut[18]) );
    VMW_NAND2 U869 ( .A(n2837), .B(n2838), .Z(n2836) );
    VMW_NOR2 U955 ( .A(n2912), .B(n2880), .Z(n2735) );
    VMW_INV U1049 ( .A(ColIn[27]), .Z(n2743) );
    VMW_OR2 U795 ( .A(ColIn[10]), .B(n2732), .Z(ColOut[10]) );
    VMW_OR2 U947 ( .A(n2912), .B(n2825), .Z(n2726) );
    VMW_NOR2 U972 ( .A(CallIn), .B(n674), .Z(n2895) );
    VMW_NOR2 U960 ( .A(n2830), .B(n2885), .Z(n2741) );
    VMW_OR2 U757 ( .A(n2723), .B(PDiagIn[17]), .Z(PDiagOut[16]) );
    VMW_OR2 U770 ( .A(n2738), .B(PDiagIn[4]), .Z(PDiagOut[3]) );
    VMW_NAND2 U815 ( .A(n2718), .B(n2761), .Z(NDiagOut[22]) );
    VMW_INV U1099 ( .A(n2870), .Z(n2939) );
    VMW_OR2 U832 ( .A(NDiagIn[4]), .B(n2738), .Z(NDiagOut[5]) );
    VMW_OR2 U985 ( .A(CallIn), .B(n530), .Z(n2920) );
    VMW_OR2 U829 ( .A(NDiagIn[7]), .B(n2735), .Z(NDiagOut[8]) );
    VMW_AND2 U885 ( .A(n2872), .B(n2822), .Z(n2818) );
    VMW_AO22 U929 ( .A(n2890), .B(ScanOut[1]), .C(n2889), .D(ScanIn[1]), .Z(
        n2773) );
    VMW_NOR2 U1012 ( .A(CallIn), .B(n834), .Z(n2934) );
    VMW_AND2 U932 ( .A(n2883), .B(n2909), .Z(n2702) );
    VMW_INV U1035 ( .A(ScanOut[4]), .Z(n2882) );
    VMW_OR4 U1009 ( .A(n2931), .B(NDiagIn[6]), .C(ColIn[6]), .D(PDiagIn[6]), 
        .Z(n2813) );
    VMW_MUX2I U915 ( .A(ScanOut[2]), .B(ScanIn[2]), .S(ScanEnable), .Z(n2698)
         );
    VMW_NAND2 U860 ( .A(ScanOut[3]), .B(ScanOut[2]), .Z(n2823) );
    VMW_INV U1082 ( .A(n2865), .Z(n2867) );
    VMW_OR2 U744 ( .A(n2702), .B(PDiagIn[30]), .Z(PDiagOut[29]) );
    VMW_OR2 U786 ( .A(ColIn[19]), .B(n2721), .Z(ColOut[19]) );
    VMW_AND2 U847 ( .A(n2789), .B(n2790), .Z(n2788) );
    VMW_AND2 U868 ( .A(n2832), .B(n2835), .Z(n2834) );
    VMW_INV U1040 ( .A(PDiagIn[25]), .Z(n2709) );
    VMW_INV U1067 ( .A(NDiagIn[20]), .Z(n2762) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_12 gt_104_3 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , UNCONNECTED_4, 
        UNCONNECTED_5}), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2966), .TC(n2966), .LT_LE(n514)
         );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_17 gt_104_17 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_6}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        Logic11, \NDiagOut[0] }), .LEQ(n2971), .TC(n2971), .LT_LE(n738) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_30 gt_104_30 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11}), .LEQ(n2984), .TC(n2984), .LT_LE(n946) );
    VMW_NOR2 U954 ( .A(n2829), .B(n2878), .Z(n2734) );
    VMW_INV U1048 ( .A(PDiagIn[3]), .Z(n2739) );
    VMW_OR3 U973 ( .A(n2840), .B(n2841), .C(n2894), .Z(n2905) );
    VMW_NOR2 U1001 ( .A(CallIn), .B(n898), .Z(n2927) );
    VMW_OAI21 U1026 ( .A(n2806), .B(n2907), .C(n2845), .Z(n2940) );
    VMW_OR2 U763 ( .A(n2731), .B(PDiagIn[11]), .Z(PDiagOut[10]) );
    VMW_OR2 U806 ( .A(NDiagIn[30]), .B(n2702), .Z(NDiagOut[31]) );
    VMW_NAND2 U821 ( .A(n2726), .B(n2763), .Z(NDiagOut[16]) );
    VMW_OR4 U996 ( .A(PDiagIn[0]), .B(n2694), .C(ColIn[0]), .D(NDiagIn[0]), 
        .Z(n2822) );
    VMW_PULLDOWN U704 ( .Z(n2955) );
    VMW_PULLDOWN U716 ( .Z(n2967) );
    VMW_PULLDOWN U731 ( .Z(n2982) );
    VMW_NAND2 U778 ( .A(n2706), .B(n2743), .Z(ColOut[27]) );
    VMW_NAND2 U873 ( .A(n2789), .B(n2790), .Z(n2809) );
    VMW_OR2 U896 ( .A(n2824), .B(n2884), .Z(n2885) );
    VMW_AO22 U921 ( .A(n2867), .B(n2891), .C(n2792), .D(n2903), .Z(n2786) );
    VMW_INV U1091 ( .A(n2840), .Z(n2943) );
    VMW_OAI21 U906 ( .A(n2788), .B(n2849), .C(n2817), .Z(n2799) );
    VMW_NOR2 U968 ( .A(CallIn), .B(n706), .Z(n2914) );
    VMW_INV U1053 ( .A(ColIn[23]), .Z(n2747) );
    VMW_INV U1074 ( .A(n2830), .Z(n2909) );
    VMW_FD CallOut_reg ( .D(CallOut1070), .CP(Clk), .Q(CallOut) );
    VMW_FD \MyColumn_reg[5]  ( .D(n2949), .CP(Clk), .Q(ScanOut[5]) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_21 gt_104_23 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , UNCONNECTED_7, UNCONNECTED_8, 
        UNCONNECTED_9}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2975), .TC(n2975), 
        .LT_LE(n834) );
    VMW_PULLDOWN U723 ( .Z(n2974) );
    VMW_AOI211 U854 ( .A(n2767), .B(n2766), .C(n2815), .D(n2769), .Z(n2814) );
    VMW_OR2 U861 ( .A(ScanOut[5]), .B(ScanOut[4]), .Z(n2824) );
    VMW_PULLDOWN U711 ( .Z(n2962) );
    VMW_PULLDOWN U718 ( .Z(n2969) );
    VMW_NAND2 U738 ( .A(n2694), .B(n2696), .Z(\n1108[4] ) );
    VMW_OR2 U756 ( .A(n2722), .B(PDiagIn[18]), .Z(PDiagOut[17]) );
    VMW_OR2 U828 ( .A(NDiagIn[8]), .B(n2734), .Z(NDiagOut[9]) );
    VMW_NOR3 U846 ( .A(n2786), .B(n2787), .C(n2781), .Z(n2785) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_22 gt_104_2 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, \NDiagOut[0] , 
        Logic11}), .LEQ(n2976), .TC(n2976), .LT_LE(n498) );
    VMW_OR4 U884 ( .A(n2853), .B(n2797), .C(n2870), .D(n2871), .Z(n2869) );
    VMW_MUX2I U914 ( .A(ScanOut[3]), .B(ScanIn[3]), .S(ScanEnable), .Z(n2697)
         );
    VMW_AND2 U933 ( .A(n2883), .B(n2910), .Z(n2703) );
    VMW_INV U1041 ( .A(PDiagIn[24]), .Z(n2711) );
    VMW_INV U1066 ( .A(NDiagIn[21]), .Z(n2761) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_1 gt_104_16 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, Logic11, 
        Logic11}), .LEQ(n2955), .TC(n2955), .LT_LE(n722) );
    VMW_NOR2 U1008 ( .A(CallIn), .B(n866), .Z(n2931) );
    VMW_INV U1083 ( .A(n2818), .Z(n2820) );
    VMW_NAND2 U771 ( .A(n2739), .B(n2740), .Z(PDiagOut[2]) );
    VMW_NAND2 U814 ( .A(n2716), .B(n2760), .Z(NDiagOut[23]) );
    VMW_AND4 U984 ( .A(n2919), .B(n2757), .C(n2745), .D(n2709), .Z(n2854) );
    VMW_NAND2 U833 ( .A(n2740), .B(n2765), .Z(NDiagOut[4]) );
    VMW_INV U1098 ( .A(n2863), .Z(n2947) );
    VMW_OR2 U794 ( .A(ColIn[11]), .B(n2731), .Z(ColOut[11]) );
    VMW_AO21 U928 ( .A(n2891), .B(n2867), .C(n2860), .Z(n2802) );
    VMW_OR4 U1013 ( .A(n2934), .B(NDiagIn[8]), .C(ColIn[8]), .D(PDiagIn[8]), 
        .Z(n2862) );
    VMW_FD \MyColumn_reg[1]  ( .D(n2953), .CP(Clk), .Q(ScanOut[1]) );
    VMW_OAI211 U1034 ( .A(n2859), .B(n2897), .C(n2948), .D(n2872), .Z(n2821)
         );
    VMW_AND2 U946 ( .A(n2888), .B(n2911), .Z(n2724) );
    VMW_NOR2 U961 ( .A(n2877), .B(n2885), .Z(n2742) );
    VMW_NAND2 U793 ( .A(n2730), .B(n2752), .Z(ColOut[12]) );
    VMW_OR2 U966 ( .A(CallIn), .B(n722), .Z(n2913) );
    VMW_OR2 U941 ( .A(n2877), .B(n2887), .Z(n2718) );
    VMW_PULLDOWN U724 ( .Z(n2975) );
    VMW_NAND2 U751 ( .A(n2713), .B(n2714), .Z(PDiagOut[22]) );
    VMW_OR2 U776 ( .A(ColIn[29]), .B(n2703), .Z(ColOut[29]) );
    VMW_NAND2 U813 ( .A(n2714), .B(n2759), .Z(NDiagOut[24]) );
    VMW_OR2 U834 ( .A(NDiagIn[2]), .B(n2741), .Z(NDiagOut[3]) );
    VMW_OR2 U983 ( .A(CallIn), .B(n562), .Z(n2919) );
    VMW_OR2 U808 ( .A(NDiagIn[28]), .B(n2704), .Z(NDiagOut[29]) );
    VMW_AND2 U883 ( .A(n2867), .B(n2868), .Z(n2816) );
    VMW_OR2 U898 ( .A(n2879), .B(n2881), .Z(n2887) );
    VMW_OAI211 U1033 ( .A(n2811), .B(n2856), .C(n2928), .D(n2858), .Z(n2948)
         );
    VMW_FD \MyColumn_reg[3]  ( .D(n2951), .CP(Clk), .Q(ScanOut[3]) );
    VMW_OR4 U908 ( .A(n2896), .B(NDiagIn[19]), .C(ColIn[19]), .D(PDiagIn[19]), 
        .Z(n2847) );
    VMW_NOR2 U1014 ( .A(CallIn), .B(n482), .Z(n2805) );
    VMW_MUX2I U913 ( .A(ScanOut[4]), .B(ScanIn[4]), .S(ScanEnable), .Z(n2696)
         );
    VMW_AND2 U934 ( .A(n2883), .B(n2911), .Z(n2704) );
    VMW_OAI211 U1028 ( .A(n2841), .B(n2943), .C(n2941), .D(n2817), .Z(n2942)
         );
    VMW_OR3 U841 ( .A(n2769), .B(n2774), .C(n2775), .Z(n2952) );
    VMW_OR4 U998 ( .A(n2925), .B(NDiagIn[10]), .C(ColIn[10]), .D(PDiagIn[10]), 
        .Z(n2868) );
    VMW_INV U1084 ( .A(n2873), .Z(n2819) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_28 gt_104_5 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_10}), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        Logic11, \NDiagOut[0] }), .LEQ(n2982), .TC(n2982), .LT_LE(n546) );
    VMW_OR2 U788 ( .A(ColIn[17]), .B(n2723), .Z(ColOut[17]) );
    VMW_OR2 U866 ( .A(n2831), .B(ScanOut[0]), .Z(n2830) );
    VMW_INV U1046 ( .A(PDiagIn[15]), .Z(n2725) );
    VMW_AND2 U853 ( .A(n2812), .B(n2813), .Z(n2811) );
    VMW_NOR2 U948 ( .A(n2825), .B(n2830), .Z(n2727) );
    VMW_INV U1054 ( .A(ColIn[22]), .Z(n2748) );
    VMW_INV U1061 ( .A(NDiagIn[26]), .Z(n2756) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_3 gt_104_11 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , UNCONNECTED_11, 
        UNCONNECTED_12}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2957), .TC(n2957), .LT_LE(n642)
         );
    VMW_INV U1073 ( .A(n2826), .Z(n2912) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_29 gt_104_24 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, 
        Logic11}), .LEQ(n2983), .TC(n2983), .LT_LE(n850) );
    VMW_PULLDOWN U736 ( .Z(\NDiagOut[0] ) );
    VMW_OR2 U743 ( .A(n2701), .B(PDiagIn[31]), .Z(PDiagOut[30]) );
    VMW_OR2 U758 ( .A(n2724), .B(PDiagIn[16]), .Z(PDiagOut[15]) );
    VMW_NAND2 U874 ( .A(n2843), .B(n2850), .Z(n2849) );
    VMW_OR2 U764 ( .A(n2732), .B(PDiagIn[10]), .Z(PDiagOut[9]) );
    VMW_NAND2 U891 ( .A(n2828), .B(ScanOut[2]), .Z(n2879) );
    VMW_NOR3 U901 ( .A(CallIn), .B(ScanEnable), .C(n2767), .Z(n2890) );
    VMW_INV U1096 ( .A(n2928), .Z(n2857) );
    VMW_OAI211 U926 ( .A(n2839), .B(n2847), .C(n2905), .D(n2869), .Z(n2798) );
    VMW_NOR2 U1006 ( .A(CallIn), .B(n850), .Z(n2930) );
    VMW_OR3 U1021 ( .A(n2874), .B(n2799), .C(n2904), .Z(n2793) );
    VMW_OR2 U801 ( .A(ColIn[4]), .B(n2738), .Z(ColOut[4]) );
    VMW_OR2 U826 ( .A(NDiagIn[10]), .B(n2732), .Z(NDiagOut[11]) );
    VMW_NOR2 U991 ( .A(CallIn), .B(n786), .Z(n2923) );
    VMW_PULLDOWN U706 ( .Z(n2957) );
    VMW_PULLDOWN U708 ( .Z(n2959) );
    VMW_PULLDOWN U726 ( .Z(n2977) );
    VMW_NAND2 U781 ( .A(n2712), .B(n2746), .Z(ColOut[24]) );
    VMW_AOI211 U848 ( .A(n2792), .B(n2793), .C(n2794), .D(n2787), .Z(n2791) );
    VMW_OR2 U974 ( .A(CallIn), .B(n642), .Z(n2915) );
    VMW_INV U1068 ( .A(NDiagIn[15]), .Z(n2763) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_14 gt_104_18 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        Logic11}), .LEQ(n2968), .TC(n2968), .LT_LE(n754) );
    VMW_NOR2 U953 ( .A(n2829), .B(n2877), .Z(n2733) );
    VMW_NOR2 U958 ( .A(n2878), .B(n2880), .Z(n2738) );
    VMW_INV U1063 ( .A(NDiagIn[24]), .Z(n2758) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_15 gt_104_13 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_13}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n2969), .TC(n2969), 
        .LT_LE(n674) );
    VMW_INV U1044 ( .A(PDiagIn[21]), .Z(n2717) );
    VMW_NAND2 U748 ( .A(n2707), .B(n2708), .Z(PDiagOut[25]) );
    VMW_OR3 U843 ( .A(n2769), .B(n2778), .C(n2779), .Z(n2950) );
    VMW_OR2 U864 ( .A(ScanOut[2]), .B(n2828), .Z(n2827) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_11 gt_104_7 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , UNCONNECTED_14, UNCONNECTED_15, 
        UNCONNECTED_16}), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2965), .TC(n2965), .LT_LE(n578)
         );
    VMW_NAND2 U753 ( .A(n2717), .B(n2718), .Z(PDiagOut[20]) );
    VMW_NAND2 U811 ( .A(n2710), .B(n2757), .Z(NDiagOut[26]) );
    VMW_NAND2 U881 ( .A(n2864), .B(n2858), .Z(n2784) );
    VMW_OR2 U936 ( .A(n2830), .B(n2886), .Z(n2708) );
    VMW_INV U1086 ( .A(n2814), .Z(n2949) );
    VMW_NOR4 U911 ( .A(n2901), .B(NDiagIn[13]), .C(ColIn[13]), .D(PDiagIn[13]), 
        .Z(n2900) );
    VMW_NOR2 U1016 ( .A(CallIn), .B(n498), .Z(n2935) );
    VMW_AO21 U1031 ( .A(n2945), .B(n2868), .C(n2933), .Z(n2946) );
    VMW_OR2 U981 ( .A(CallIn), .B(n578), .Z(n2918) );
    VMW_OR2 U774 ( .A(n2701), .B(ColIn[31]), .Z(ColOut[31]) );
    VMW_NAND2 U783 ( .A(n2716), .B(n2748), .Z(ColOut[22]) );
    VMW_OR2 U791 ( .A(ColIn[14]), .B(n2727), .Z(ColOut[14]) );
    VMW_OR2 U836 ( .A(NDiagIn[0]), .B(n2754), .Z(NDiagOut[1]) );
    VMW_NOR3 U858 ( .A(n2768), .B(n2800), .C(n2820), .Z(n2772) );
    VMW_AND2 U943 ( .A(n2888), .B(n2826), .Z(n2721) );
    VMW_NOR2 U964 ( .A(n2885), .B(n2878), .Z(n2754) );
    VMW_INV U1078 ( .A(n2853), .Z(n2796) );
    VMW_NOR2 U951 ( .A(n2912), .B(n2829), .Z(n2731) );
    VMW_OR2 U976 ( .A(CallIn), .B(n626), .Z(n2916) );
    VMW_PULLDOWN U713 ( .Z(n2964) );
    VMW_PULLDOWN U734 ( .Z(n2985) );
    VMW_NAND2 U741 ( .A(n2694), .B(n2699), .Z(\n1108[1] ) );
    VMW_OR2 U803 ( .A(ColIn[2]), .B(n2741), .Z(ColOut[2]) );
    VMW_OR2 U993 ( .A(CallIn), .B(n770), .Z(n2892) );
    VMW_OR2 U766 ( .A(n2734), .B(PDiagIn[8]), .Z(PDiagOut[7]) );
    VMW_OR2 U818 ( .A(NDiagIn[18]), .B(n2722), .Z(NDiagOut[19]) );
    VMW_NAND2 U824 ( .A(n2730), .B(n2764), .Z(NDiagOut[13]) );
    VMW_AO21 U888 ( .A(n2876), .B(n2694), .C(Reset), .Z(n2768) );
    VMW_NAND3 U918 ( .A(n2902), .B(n2804), .C(n2816), .Z(n2875) );
    VMW_NOR4 U1004 ( .A(n2929), .B(NDiagIn[2]), .C(ColIn[2]), .D(PDiagIn[2]), 
        .Z(n2859) );
    VMW_OR2 U893 ( .A(n2882), .B(ScanOut[5]), .Z(n2881) );
    VMW_NAND4 U903 ( .A(n2892), .B(n2764), .C(n2752), .D(n2729), .Z(n2838) );
    VMW_AO22 U924 ( .A(n2801), .B(n2782), .C(n2858), .D(n2855), .Z(n2794) );
    VMW_OAI21 U1023 ( .A(n2795), .B(n2873), .C(n2937), .Z(n2906) );
    VMW_FD \MyColumn_reg[2]  ( .D(n2952), .CP(Clk), .Q(ScanOut[2]) );
    VMW_INV U1038 ( .A(PDiagIn[27]), .Z(n2705) );
    VMW_AND4 U988 ( .A(n2921), .B(n2756), .C(n2744), .D(n2707), .Z(n2922) );
    VMW_INV U1094 ( .A(n2854), .Z(n2807) );
    VMW_OR4 U851 ( .A(n2805), .B(NDiagIn[30]), .C(ColIn[30]), .D(PDiagIn[30]), 
        .Z(n2804) );
    VMW_OR4 U876 ( .A(n2849), .B(n2809), .C(n2854), .D(n2810), .Z(n2853) );
    VMW_PULLDOWN U714 ( .Z(n2965) );
    VMW_OR2 U798 ( .A(ColIn[7]), .B(n2735), .Z(ColOut[7]) );
    VMW_INV U1056 ( .A(ColIn[20]), .Z(n2750) );
    VMW_INV U1071 ( .A(CallIn), .Z(n2694) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_27 gt_104_26 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11}), .LEQ(n2981), .TC(n2981), .LT_LE(n882) );
    VMW_PULLDOWN U728 ( .Z(n2979) );
    VMW_PULLDOWN U733 ( .Z(n2984) );
    VMW_NOR3 U856 ( .A(n2768), .B(n2785), .C(n2820), .Z(n2776) );
    VMW_AND2 U871 ( .A(n2844), .B(n2845), .Z(n2843) );
    VMW_OR2 U746 ( .A(n2704), .B(PDiagIn[28]), .Z(PDiagOut[27]) );
    VMW_OR2 U761 ( .A(n2728), .B(PDiagIn[13]), .Z(PDiagOut[12]) );
    VMW_OR2 U823 ( .A(NDiagIn[13]), .B(n2728), .Z(NDiagOut[14]) );
    VMW_NOR2 U838 ( .A(n2768), .B(n2766), .Z(CallOut1070) );
    VMW_NOR2 U894 ( .A(n2823), .B(n2881), .Z(n2883) );
    VMW_NOR2 U1018 ( .A(CallIn), .B(n514), .Z(n2936) );
    VMW_INV U1051 ( .A(ColIn[25]), .Z(n2745) );
    VMW_INV U1076 ( .A(n2839), .Z(n2848) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_26 gt_104_21 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_17}), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n2980), .TC(n2980), 
        .LT_LE(n802) );
    VMW_NOR2 U904 ( .A(n2891), .B(n2865), .Z(n2792) );
    VMW_OAI22 U923 ( .A(n2797), .B(n2853), .C(n2843), .D(n2846), .Z(n2904) );
    VMW_INV U1093 ( .A(n2894), .Z(n2842) );
    VMW_NAND2 U784 ( .A(n2718), .B(n2749), .Z(ColOut[21]) );
    VMW_OR2 U804 ( .A(ColIn[1]), .B(n2742), .Z(ColOut[1]) );
    VMW_INV U1088 ( .A(n2878), .Z(n2911) );
    VMW_OR2 U938 ( .A(n2878), .B(n2886), .Z(n2712) );
    VMW_NOR2 U994 ( .A(CallIn), .B(n946), .Z(n2924) );
    VMW_NOR2 U956 ( .A(n2830), .B(n2880), .Z(n2736) );
    VMW_NOR2 U971 ( .A(CallIn), .B(n690), .Z(n2899) );
    VMW_NOR2 U1003 ( .A(CallIn), .B(n930), .Z(n2929) );
    VMW_OAI21 U1024 ( .A(n2804), .B(n2871), .C(n2939), .Z(n2938) );
    VMW_FD \MyColumn_reg[0]  ( .D(n2954), .CP(Clk), .Q(ScanOut[0]) );
    VMW_NAND2 U754 ( .A(n2719), .B(n2720), .Z(PDiagOut[19]) );
    VMW_OR2 U773 ( .A(n2742), .B(PDiagIn[1]), .Z(PDiagOut[0]) );
    VMW_OR2 U796 ( .A(ColIn[9]), .B(n2733), .Z(ColOut[9]) );
    VMW_NOR2 U878 ( .A(n2859), .B(n2860), .Z(n2858) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_9 gt_104_9 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_18}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        Logic11, \NDiagOut[0] }), .LEQ(n2963), .TC(n2963), .LT_LE(n610) );
    VMW_AND2 U944 ( .A(n2888), .B(n2909), .Z(n2722) );
    VMW_AND2 U963 ( .A(n2883), .B(n2826), .Z(n2701) );
    VMW_INV U1058 ( .A(ColIn[12]), .Z(n2752) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_18 gt_104_28 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, Logic11}), .LEQ(n2972), .TC(n2972), .LT_LE(n914) );
    VMW_OR2 U831 ( .A(NDiagIn[5]), .B(n2737), .Z(NDiagOut[6]) );
    VMW_NOR4 U1011 ( .A(n2932), .B(NDiagIn[9]), .C(ColIn[9]), .D(PDiagIn[9]), 
        .Z(n2933) );
    VMW_INV U1036 ( .A(ScanOut[3]), .Z(n2828) );
    VMW_OR2 U768 ( .A(n2736), .B(PDiagIn[6]), .Z(PDiagOut[5]) );
    VMW_NAND2 U816 ( .A(n2720), .B(n2762), .Z(NDiagOut[21]) );
    VMW_NAND4 U986 ( .A(n2920), .B(n2755), .C(n2743), .D(n2705), .Z(n2851) );
    VMW_INV U1081 ( .A(n2855), .Z(n2864) );
    VMW_OR2 U886 ( .A(n2874), .B(n2836), .Z(n2873) );
    VMW_MUX2I U916 ( .A(ScanOut[1]), .B(ScanIn[1]), .S(ScanEnable), .Z(n2699)
         );
    VMW_AO22 U931 ( .A(n2890), .B(ScanOut[0]), .C(n2889), .D(ScanIn[0]), .Z(
        n2771) );
    VMW_OR2 U978 ( .A(CallIn), .B(n610), .Z(n2917) );
    VMW_INV U1043 ( .A(PDiagIn[22]), .Z(n2715) );
    VMW_FD \MyColumn_reg[4]  ( .D(n2950), .CP(Clk), .Q(ScanOut[4]) );
    VMW_INV U1064 ( .A(NDiagIn[23]), .Z(n2759) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_7 gt_104_14 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11}), .LEQ(n2961), .TC(n2961), .LT_LE(n690) );
    VMW_PULLDOWN U707 ( .Z(n2958) );
    VMW_PULLDOWN U715 ( .Z(n2966) );
    VMW_PULLDOWN U721 ( .Z(n2972) );
    VMW_NOR2 U844 ( .A(CallIn), .B(n466), .Z(n2780) );
    VMW_AND2 U863 ( .A(ScanOut[1]), .B(ScanOut[0]), .Z(n2826) );
    VMW_PULLDOWN U729 ( .Z(n2980) );
    VMW_NAND2 U785 ( .A(n2720), .B(n2750), .Z(ColOut[20]) );
    VMW_NOR2 U957 ( .A(n2877), .B(n2880), .Z(n2737) );
    VMW_NOR2 U970 ( .A(CallIn), .B(n658), .Z(n2896) );
    VMW_NAND2 U747 ( .A(n2705), .B(n2706), .Z(PDiagOut[26]) );
    VMW_OR2 U760 ( .A(n2727), .B(PDiagIn[14]), .Z(PDiagOut[13]) );
    VMW_OR2 U822 ( .A(NDiagIn[14]), .B(n2727), .Z(NDiagOut[15]) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_16 gt_104_8 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, Logic11, 
        Logic11}), .LEQ(n2970), .TC(n2970), .LT_LE(n594) );
    VMW_OR2 U805 ( .A(ColIn[0]), .B(n2754), .Z(ColOut[0]) );
    VMW_OR4 U995 ( .A(n2924), .B(NDiagIn[1]), .C(ColIn[1]), .D(PDiagIn[1]), 
        .Z(n2872) );
    VMW_OR3 U839 ( .A(n2769), .B(n2770), .C(n2771), .Z(n2954) );
    VMW_OR2 U895 ( .A(ScanOut[3]), .B(ScanOut[2]), .Z(n2884) );
    VMW_NAND4 U905 ( .A(n2893), .B(n2759), .C(n2747), .D(n2713), .Z(n2790) );
    VMW_OR2 U939 ( .A(n2912), .B(n2887), .Z(n2714) );
    VMW_AO21 U1025 ( .A(n2851), .B(n2938), .C(n2922), .Z(n2808) );
    VMW_INV U1089 ( .A(n2908), .Z(n2789) );
    VMW_OR4 U1002 ( .A(n2927), .B(NDiagIn[4]), .C(ColIn[4]), .D(PDiagIn[4]), 
        .Z(n2928) );
    VMW_AO22 U922 ( .A(n2890), .B(ScanOut[3]), .C(n2889), .D(ScanIn[3]), .Z(
        n2777) );
    VMW_NOR4 U1019 ( .A(n2936), .B(NDiagIn[28]), .C(ColIn[28]), .D(PDiagIn[28]
        ), .Z(n2870) );
    VMW_INV U1092 ( .A(n2900), .Z(n2835) );
    VMW_PULLDOWN U732 ( .Z(n2983) );
    VMW_NOR3 U857 ( .A(n2768), .B(n2791), .C(n2820), .Z(n2774) );
    VMW_OR3 U870 ( .A(n2840), .B(n2841), .C(n2842), .Z(n2839) );
    VMW_AND4 U979 ( .A(n2917), .B(n2760), .C(n2748), .D(n2715), .Z(n2908) );
    VMW_INV U1042 ( .A(PDiagIn[23]), .Z(n2713) );
    VMW_INV U1050 ( .A(ColIn[26]), .Z(n2744) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_4 gt_104_20 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , \NDiagOut[0] , Logic11, \NDiagOut[0] , Logic11, 
        Logic11}), .LEQ(n2958), .TC(n2958), .LT_LE(n786) );
    VMW_INV U1077 ( .A(n2846), .Z(n2850) );
    VMW_INV U1065 ( .A(NDiagIn[22]), .Z(n2760) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_5 gt_104_15 ( .A({
        \n1108[5] , \n1108[4] , UNCONNECTED_19, UNCONNECTED_20, UNCONNECTED_21, 
        UNCONNECTED_22}), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , 
        \NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2959), .TC(n2959), 
        .LT_LE(n706) );
    VMW_PULLDOWN U709 ( .Z(n2960) );
    VMW_PULLDOWN U712 ( .Z(n2963) );
    VMW_PULLDOWN U720 ( .Z(n2971) );
    VMW_NOR3 U845 ( .A(n2782), .B(n2783), .C(n2784), .Z(n2781) );
    VMW_OR2 U862 ( .A(n2823), .B(n2824), .Z(n2825) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_6 gt_104_1 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_23}), .B({\NDiagOut[0] , Logic11, Logic11, Logic11, 
        Logic11, \NDiagOut[0] }), .LEQ(n2960), .TC(n2960), .LT_LE(n482) );
    VMW_PULLDOWN U727 ( .Z(n2978) );
    VMW_NAND2 U749 ( .A(n2709), .B(n2710), .Z(PDiagOut[24]) );
    VMW_NAND2 U752 ( .A(n2715), .B(n2716), .Z(PDiagOut[21]) );
    VMW_OR2 U755 ( .A(n2721), .B(PDiagIn[19]), .Z(PDiagOut[18]) );
    VMW_OR2 U769 ( .A(n2737), .B(PDiagIn[5]), .Z(PDiagOut[4]) );
    VMW_INV U1080 ( .A(n2784), .Z(n2801) );
    VMW_OR2 U772 ( .A(n2741), .B(PDiagIn[2]), .Z(PDiagOut[1]) );
    VMW_OR2 U830 ( .A(NDiagIn[6]), .B(n2736), .Z(NDiagOut[7]) );
    VMW_NOR4 U887 ( .A(n2820), .B(n2869), .C(n2873), .D(n2875), .Z(n2766) );
    VMW_MUX2I U917 ( .A(ScanOut[0]), .B(ScanIn[0]), .S(ScanEnable), .Z(n2700)
         );
    VMW_OAI21 U930 ( .A(n2908), .B(n2790), .C(n2844), .Z(n2907) );
    VMW_NOR2 U1010 ( .A(CallIn), .B(n818), .Z(n2932) );
    VMW_INV U1037 ( .A(ScanOut[1]), .Z(n2831) );
    VMW_NAND2 U790 ( .A(n2726), .B(n2751), .Z(ColOut[15]) );
    VMW_OR2 U797 ( .A(ColIn[8]), .B(n2734), .Z(ColOut[8]) );
    VMW_OR2 U817 ( .A(NDiagIn[19]), .B(n2721), .Z(NDiagOut[20]) );
    VMW_AND2 U879 ( .A(n2861), .B(n2862), .Z(n2783) );
    VMW_OR2 U987 ( .A(CallIn), .B(n546), .Z(n2921) );
    VMW_AND2 U945 ( .A(n2888), .B(n2910), .Z(n2723) );
    VMW_AND2 U962 ( .A(n2889), .B(CallIn), .Z(n2769) );
    VMW_INV U1059 ( .A(ColIn[3]), .Z(n2753) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_13 gt_104_29 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , 
        UNCONNECTED_24}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        \NDiagOut[0] , Logic11, \NDiagOut[0] }), .LEQ(n2967), .TC(n2967), 
        .LT_LE(n930) );
    VMW_AND3 U859 ( .A(n2821), .B(n2822), .C(n2767), .Z(n2770) );
    VMW_NAND2 U810 ( .A(n2708), .B(n2756), .Z(NDiagOut[27]) );
    VMW_OR2 U942 ( .A(n2878), .B(n2887), .Z(n2720) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_31 gt_104 ( .A({\n1108[5] , 
        \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] }), .B({
        \NDiagOut[0] , Logic11, Logic11, Logic11, Logic11, Logic11}), .LEQ(
        n2985), .TC(n2985), .LT_LE(n466) );
    VMW_NOR3 U965 ( .A(n2891), .B(n2865), .C(n2838), .Z(n2787) );
    VMW_OR2 U980 ( .A(CallIn), .B(n594), .Z(n2893) );
    VMW_NOR4 U1017 ( .A(n2935), .B(NDiagIn[29]), .C(ColIn[29]), .D(PDiagIn[29]
        ), .Z(n2871) );
    VMW_INV U1079 ( .A(n2782), .Z(n2866) );
    VMW_OAI211 U1030 ( .A(n2836), .B(n2835), .C(n2944), .D(n2837), .Z(n2945)
         );
    VMW_OR2 U775 ( .A(ColIn[30]), .B(n2702), .Z(ColOut[30]) );
    VMW_AND2 U837 ( .A(n2766), .B(n2767), .Z(ReturnOut1063) );
    VMW_FD ReturnOut_reg ( .D(ReturnOut1063), .CP(Clk), .Q(ReturnOut) );
    VMW_NAND2 U880 ( .A(n2813), .B(n2863), .Z(n2782) );
    VMW_NOR4 U910 ( .A(n2899), .B(NDiagIn[17]), .C(ColIn[17]), .D(PDiagIn[17]), 
        .Z(n2840) );
    VMW_OR2 U937 ( .A(n2877), .B(n2886), .Z(n2710) );
    VMW_INV U1087 ( .A(n2877), .Z(n2910) );
    VMW_OR2 U959 ( .A(n2885), .B(n2912), .Z(n2740) );
    VMW_INV U1045 ( .A(PDiagIn[20]), .Z(n2719) );
    VMW_INV U1062 ( .A(NDiagIn[25]), .Z(n2757) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_20 gt_104_12 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, \NDiagOut[0] , \NDiagOut[0] , Logic11, 
        Logic11}), .LEQ(n2974), .TC(n2974), .LT_LE(n658) );
    VMW_PULLUP U735 ( .Z(Logic11) );
    VMW_OR3 U842 ( .A(n2769), .B(n2776), .C(n2777), .Z(n2951) );
    VMW_OR2 U865 ( .A(n2827), .B(n2824), .Z(n2829) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_23 gt_104_6 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , \n1108[1] , \n1108[0] 
        }), .B({\NDiagOut[0] , Logic11, Logic11, \NDiagOut[0] , \NDiagOut[0] , 
        Logic11}), .LEQ(n2977), .TC(n2977), .LT_LE(n562) );
    VMW_AOI211 U850 ( .A(n2801), .B(n2782), .C(n2802), .D(n2803), .Z(n2800) );
    VMW_OR2 U877 ( .A(n2856), .B(n2857), .Z(n2855) );
    VMW_NAND2 U740 ( .A(n2694), .B(n2698), .Z(\n1108[2] ) );
    VMW_OR2 U799 ( .A(ColIn[6]), .B(n2736), .Z(ColOut[6]) );
    VMW_INV U1057 ( .A(ColIn[15]), .Z(n2751) );
    VMW_INV U1070 ( .A(NDiagIn[3]), .Z(n2765) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1_DW01_cmp2_6_8 gt_104_27 ( .A({
        \n1108[5] , \n1108[4] , \n1108[3] , \n1108[2] , UNCONNECTED_25, 
        UNCONNECTED_26}), .B({\NDiagOut[0] , \NDiagOut[0] , \NDiagOut[0] , 
        Logic11, \NDiagOut[0] , \NDiagOut[0] }), .LEQ(n2962), .TC(n2962), 
        .LT_LE(n898) );
    VMW_NAND2 U802 ( .A(n2740), .B(n2753), .Z(ColOut[3]) );
    VMW_OR2 U819 ( .A(NDiagIn[17]), .B(n2723), .Z(NDiagOut[18]) );
    VMW_OR2 U892 ( .A(n2879), .B(n2824), .Z(n2880) );
    VMW_AO22 U925 ( .A(n2890), .B(ScanOut[2]), .C(n2889), .D(ScanIn[2]), .Z(
        n2775) );
    VMW_INV U1039 ( .A(PDiagIn[26]), .Z(n2707) );
    VMW_NAND2 U902 ( .A(n2868), .B(n2837), .Z(n2891) );
    VMW_NOR2 U989 ( .A(CallIn), .B(n738), .Z(n2833) );
    VMW_INV U1095 ( .A(n2922), .Z(n2852) );
    VMW_OR4 U992 ( .A(n2923), .B(NDiagIn[11]), .C(ColIn[11]), .D(PDiagIn[11]), 
        .Z(n2837) );
    VMW_OR2 U767 ( .A(n2735), .B(PDiagIn[7]), .Z(PDiagOut[6]) );
    VMW_NAND2 U782 ( .A(n2714), .B(n2747), .Z(ColOut[23]) );
    VMW_OR2 U825 ( .A(NDiagIn[11]), .B(n2731), .Z(NDiagOut[12]) );
    VMW_NAND2 U889 ( .A(ScanOut[0]), .B(n2831), .Z(n2877) );
    VMW_AO22 U919 ( .A(n2890), .B(ScanOut[5]), .C(n2889), .D(ScanIn[5]), .Z(
        n2815) );
    VMW_OR2 U1005 ( .A(CallIn), .B(n914), .Z(n2898) );
    VMW_OR3 U1022 ( .A(n2832), .B(n2900), .C(n2836), .Z(n2937) );
    VMW_OR2 U950 ( .A(n2878), .B(n2825), .Z(n2730) );
    VMW_NAND4 U977 ( .A(n2916), .B(n2761), .C(n2749), .D(n2717), .Z(n2844) );
endmodule


module NQueens_Control_IDWIDTH6_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, CallIn, ReturnIn, 
    CallOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [5:0] Id;
input  [5:0] ScanIn;
output [5:0] ScanOut;
input  [5:0] ScanId;
input  Clk, Reset, RD, WR, CallIn, ReturnIn;
output ScanEnable, CallOut;
    wire n421, n433, n387, n406, n414, n395, n446, n428, n441, n389, n408, 
        n434, n392, n413, n426, n401, n448, n412, n393, \status[4] , n435, 
        n440, \ScanReg[2] , n388, n409, n449, n452, \status[0] , n427, n400, 
        n420, \ScanReg[4] , n386, n407, \status[2] , n429, n447, \ScanReg[0] , 
        n432, n415, n394, \status[6] , n439, \ScanReg[1] , n422, n405, 
        \status[7] , \ScanReg[5] , n430, n417, n396, \status[3] , n445, 
        \status[1] , n442, n425, n437, n391, n410, n402, \status[5] , n450, 
        n419, n398, \ScanReg[3] , n436, n390, n411, n443, n451, n399, n418, 
        n424, n403, n423, n385, n404, Logic01, n438, n444, n416, n397, n431;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    assign ScanOut[5] = Logic01;
    assign ScanOut[4] = Logic01;
    assign ScanOut[3] = Logic01;
    assign ScanOut[2] = Logic01;
    assign ScanOut[1] = Logic01;
    assign ScanOut[0] = Logic01;
    VMW_PULLDOWN U96 ( .Z(n437) );
    VMW_OAI21 U113 ( .A(n395), .B(n393), .C(n396), .Z(n452) );
    VMW_XNOR2 U134 ( .A(Addr[5]), .B(Id[5]), .Z(n409) );
    VMW_AND2 U108 ( .A(n387), .B(\status[7] ), .Z(n438) );
    VMW_INV U141 ( .A(\status[2] ), .Z(n403) );
    VMW_BUFIZ U166 ( .A(n431), .E(n417), .Z(\arr[29] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_PULLDOWN U83 ( .Z(n421) );
    VMW_PULLDOWN U84 ( .Z(n422) );
    VMW_BUFIZ U148 ( .A(n412), .E(n417), .Z(\arr[19] ) );
    VMW_BUFIZ U153 ( .A(n418), .E(n417), .Z(\arr[4] ) );
    VMW_BUFIZ U174 ( .A(n439), .E(n417), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U101 ( .Z(Logic01) );
    VMW_AND2 U106 ( .A(\status[6] ), .B(n386), .Z(n446) );
    VMW_AO22 U121 ( .A(\status[4] ), .B(n387), .C(\ScanReg[4] ), .D(n385), .Z(
        n418) );
    VMW_AND3 U126 ( .A(n408), .B(n409), .C(n410), .Z(n400) );
    VMW_BUFIZ U168 ( .A(n433), .E(n417), .Z(\arr[24] ) );
    VMW_PULLDOWN U91 ( .Z(n431) );
    VMW_PULLDOWN U98 ( .Z(n441) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_NAND2 U128 ( .A(n387), .B(WR), .Z(n391) );
    VMW_BUFIZ U154 ( .A(n419), .E(n417), .Z(\arr[27] ) );
    VMW_BUFIZ U173 ( .A(n438), .E(n417), .Z(\arr[7] ) );
    VMW_INV U146 ( .A(n405), .Z(n411) );
    VMW_BUFIZ U161 ( .A(n426), .E(n417), .Z(\arr[21] ) );
    VMW_PULLDOWN U99 ( .Z(n442) );
    VMW_AND4 U114 ( .A(n397), .B(n398), .C(n399), .D(n400), .Z(n387) );
    VMW_AO21 U133 ( .A(n389), .B(n391), .C(Reset), .Z(n396) );
    VMW_FD \status_reg[7]  ( .D(n445), .CP(Clk), .Q(\status[7] ) );
    VMW_BUFIZ U155 ( .A(n420), .E(n417), .Z(\arr[14] ) );
    VMW_BUFIZ U172 ( .A(n437), .E(n417), .Z(\arr[15] ) );
    VMW_PULLDOWN U82 ( .Z(n420) );
    VMW_BUFIZ U169 ( .A(n434), .E(n417), .Z(\arr[17] ) );
    VMW_PULLDOWN U85 ( .Z(n423) );
    VMW_PULLDOWN U90 ( .Z(n430) );
    VMW_AND2 U107 ( .A(\status[7] ), .B(n386), .Z(n445) );
    VMW_AO22 U120 ( .A(\status[5] ), .B(n387), .C(\ScanReg[5] ), .D(n385), .Z(
        n439) );
    VMW_NOR5 U115 ( .A(\status[6] ), .B(\status[7] ), .C(\status[5] ), .D(
        \status[3] ), .E(\status[4] ), .Z(n401) );
    VMW_NAND3 U132 ( .A(n390), .B(n391), .C(n411), .Z(n394) );
    VMW_FD \status_reg[3]  ( .D(n449), .CP(Clk), .Q(\status[3] ) );
    VMW_PULLDOWN U97 ( .Z(n440) );
    VMW_AND2 U109 ( .A(n387), .B(\status[6] ), .Z(n424) );
    VMW_AND2 U129 ( .A(n402), .B(CallIn), .Z(n406) );
    VMW_INV U147 ( .A(n406), .Z(n389) );
    VMW_BUFIZ U160 ( .A(n425), .E(n417), .Z(\arr[31] ) );
    VMW_INV U140 ( .A(n387), .Z(n385) );
    VMW_BUFIZ U167 ( .A(n432), .E(n417), .Z(\arr[20] ) );
    VMW_PULLDOWN U100 ( .Z(n444) );
    VMW_OAI21 U112 ( .A(n392), .B(n393), .C(n394), .Z(n451) );
    VMW_XNOR2 U135 ( .A(Addr[3]), .B(Id[3]), .Z(n408) );
    VMW_FD \status_reg[1]  ( .D(n451), .CP(Clk), .Q(\status[1] ) );
    VMW_AND2 U127 ( .A(n403), .B(n404), .Z(CallOut) );
    VMW_BUFIZ U149 ( .A(n413), .E(n417), .Z(\arr[0] ) );
    VMW_BUFIZ U152 ( .A(n416), .E(n417), .Z(\arr[9] ) );
    VMW_BUFIZ U175 ( .A(n440), .E(n417), .Z(\arr[22] ) );
    VMW_FD \status_reg[5]  ( .D(n447), .CP(Clk), .Q(\status[5] ) );
    VMW_PULLDOWN U77 ( .Z(n412) );
    VMW_PULLDOWN U79 ( .Z(n415) );
    VMW_PULLDOWN U95 ( .Z(n436) );
    VMW_OR2 U110 ( .A(n387), .B(RD), .Z(n417) );
    VMW_XNOR2 U137 ( .A(Addr[0]), .B(Id[0]), .Z(n398) );
    VMW_BUFIZ U159 ( .A(n424), .E(n417), .Z(\arr[6] ) );
    VMW_AND4 U119 ( .A(n405), .B(n407), .C(n390), .D(n391), .Z(n386) );
    VMW_INV U142 ( .A(\status[1] ), .Z(n392) );
    VMW_FD \status_reg[4]  ( .D(n448), .CP(Clk), .Q(\status[4] ) );
    VMW_BUFIZ U165 ( .A(n430), .E(n417), .Z(\arr[30] ) );
    VMW_PULLDOWN U80 ( .Z(n416) );
    VMW_PULLDOWN U87 ( .Z(n426) );
    VMW_BUFIZ U150 ( .A(n414), .E(n417), .Z(\arr[23] ) );
    VMW_BUFIZ U177 ( .A(n442), .E(n417), .Z(\arr[11] ) );
    VMW_AND2 U102 ( .A(RD), .B(n385), .Z(ScanEnable) );
    VMW_AO22 U125 ( .A(\status[0] ), .B(n387), .C(\ScanReg[0] ), .D(n385), .Z(
        n413) );
    VMW_AND2 U105 ( .A(\status[5] ), .B(n386), .Z(n447) );
    VMW_FD \status_reg[0]  ( .D(n452), .CP(Clk), .Q(\status[0] ) );
    VMW_AO22 U122 ( .A(\status[3] ), .B(n387), .C(\ScanReg[3] ), .D(n385), .Z(
        n435) );
    VMW_FD \status_reg[2]  ( .D(n450), .CP(Clk), .Q(\status[2] ) );
    VMW_PULLDOWN U89 ( .Z(n429) );
    VMW_XNOR2 U139 ( .A(Addr[1]), .B(Id[1]), .Z(n399) );
    VMW_BUFIZ U157 ( .A(n422), .E(n417), .Z(\arr[16] ) );
    VMW_BUFIZ U170 ( .A(n435), .E(n417), .Z(\arr[3] ) );
    VMW_PULLDOWN U92 ( .Z(n432) );
    VMW_INV U145 ( .A(n386), .Z(n393) );
    VMW_BUFIZ U162 ( .A(n427), .E(n417), .Z(\arr[28] ) );
    VMW_FD \status_reg[6]  ( .D(n446), .CP(Clk), .Q(\status[6] ) );
    VMW_BUFIZ U179 ( .A(n444), .E(n417), .Z(\arr[8] ) );
    VMW_AND3 U117 ( .A(n401), .B(n392), .C(\status[0] ), .Z(n404) );
    VMW_PULLDOWN U78 ( .Z(n414) );
    VMW_PULLDOWN U81 ( .Z(n419) );
    VMW_NAND2 U130 ( .A(ReturnIn), .B(n402), .Z(n407) );
    VMW_XNOR2 U138 ( .A(Addr[2]), .B(Id[2]), .Z(n397) );
    VMW_BUFIZ U156 ( .A(n421), .E(n417), .Z(\arr[25] ) );
    VMW_BUFIZ U171 ( .A(n436), .E(n417), .Z(\arr[26] ) );
    VMW_PULLDOWN U86 ( .Z(n425) );
    VMW_PULLDOWN U88 ( .Z(n427) );
    VMW_PULLDOWN U93 ( .Z(n433) );
    VMW_AND2 U104 ( .A(\status[4] ), .B(n386), .Z(n448) );
    VMW_AND4 U116 ( .A(\status[1] ), .B(n401), .C(n395), .D(n403), .Z(n402) );
    VMW_AO22 U123 ( .A(\status[2] ), .B(n387), .C(\ScanReg[2] ), .D(n385), .Z(
        n428) );
    VMW_OAI21 U131 ( .A(n404), .B(n386), .C(n403), .Z(n388) );
    VMW_BUFIZ U178 ( .A(n443), .E(n417), .Z(\arr[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_PULLDOWN U94 ( .Z(n434) );
    VMW_INV U143 ( .A(\status[0] ), .Z(n395) );
    VMW_INV U144 ( .A(Reset), .Z(n390) );
    VMW_BUFIZ U163 ( .A(n428), .E(n417), .Z(\arr[2] ) );
    VMW_BUFIZ U158 ( .A(n423), .E(n417), .Z(\arr[12] ) );
    VMW_BUFIZ U164 ( .A(n429), .E(n417), .Z(\arr[13] ) );
    VMW_AND2 U103 ( .A(\status[3] ), .B(n386), .Z(n449) );
    VMW_AND4 U111 ( .A(n388), .B(n389), .C(n390), .D(n391), .Z(n450) );
    VMW_XNOR2 U136 ( .A(Addr[4]), .B(Id[4]), .Z(n410) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AO22 U124 ( .A(\status[1] ), .B(n387), .C(\ScanReg[1] ), .D(n385), .Z(
        n443) );
    VMW_NOR2 U118 ( .A(n406), .B(CallOut), .Z(n405) );
    VMW_BUFIZ U151 ( .A(n415), .E(n417), .Z(\arr[10] ) );
    VMW_BUFIZ U176 ( .A(n441), .E(n417), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \wColumn_13[27] , \wNDiag_29[0] , \wColumn_30[16] , \wColumn_6[31] , 
        \wPDiag_12[18] , \wColumn_25[22] , \wPDiag_31[30] , \wPDiag_31[29] , 
        \wColumn_30[0] , \wColumn_6[28] , \wPDiag_8[4] , \wPDiag_18[9] , 
        \wColumn_25[11] , \wPDiag_1[21] , \wPDiag_5[23] , \wNDiag_10[22] , 
        \wColumn_13[14] , \wColumn_30[25] , \wNDiag_26[27] , \wPDiag_5[10] , 
        \wColumn_18[18] , \wScan_19[0] , \wPDiag_19[27] , \wColumn_28[2] , 
        \wNDiag_31[2] , \wNDiag_10[11] , \wPDiag_19[14] , \wNDiag_26[14] , 
        \wPDiag_1[12] , \wColumn_3[4] , \wColumn_9[26] , \wNDiag_14[20] , 
        \wNDiag_22[25] , \wColumn_9[15] , \wColumn_12[8] , \wNDiag_15[4] , 
        \wNDiag_22[16] , \wNDiag_14[13] , \wNDiag_1[30] , \wColumn_2[19] , 
        \wNDiag_4[21] , \wNDiag_16[7] , \wPDiag_22[3] , \wScan_3[5] , 
        \wColumn_3[20] , \wNDiag_4[12] , \wColumn_6[9] , \wColumn_17[25] , 
        \wColumn_21[20] , \wPDiag_21[0] , \wColumn_14[6] , \wPDiag_16[30] , 
        \wPDiag_16[29] , \wNDiag_9[4] , \wColumn_17[16] , \wColumn_17[5] , 
        \wColumn_21[13] , \wNDiag_10[9] , \wReturn_13[0] , \wNDiag_15[19] , 
        \wScan_25[4] , \wNDiag_29[29] , \wNDiag_29[30] , \wNDiag_18[1] , 
        \wScan_30[3] , \wPDiag_29[8] , \wColumn_3[13] , \wNDiag_4[1] , 
        \wNDiag_28[23] , \wNDiag_5[18] , \wNDiag_7[2] , \wColumn_20[19] , 
        \wScan_28[1] , \wPDiag_17[23] , \wColumn_19[3] , \wPDiag_21[26] , 
        \wPDiag_6[2] , \wPDiag_17[10] , \wNDiag_28[10] , \wPDiag_21[15] , 
        \wPDiag_13[21] , \wPDiag_25[24] , \wPDiag_30[10] , \wPDiag_5[1] , 
        \wColumn_7[22] , \wNDiag_1[29] , \wColumn_7[11] , \wPDiag_13[12] , 
        \wPDiag_25[17] , \wNDiag_27[6] , \wNDiag_24[5] , \wPDiag_30[23] , 
        \wPDiag_10[1] , \wColumn_23[9] , \wColumn_24[31] , \wColumn_24[28] , 
        \wPDiag_13[2] , \wScan_14[5] , \wColumn_19[21] , \wNDiag_21[8] , 
        \wColumn_26[4] , \wNDiag_1[20] , \wNDiag_1[5] , \wNDiag_2[6] , 
        \wColumn_3[30] , \wColumn_3[29] , \wPDiag_4[30] , \wPDiag_4[29] , 
        \wNDiag_5[22] , \wCall_11[0] , \wColumn_19[12] , \wNDiag_11[31] , 
        \wColumn_25[7] , \wNDiag_11[28] , \wColumn_16[26] , \wPDiag_17[19] , 
        \wColumn_20[23] , \wNDiag_28[19] , \wPDiag_31[3] , \wNDiag_4[8] , 
        \wColumn_8[6] , \wColumn_16[15] , \wColumn_20[10] , \wNDiag_5[11] , 
        \wColumn_8[25] , \wNDiag_15[23] , \wNDiag_23[26] , \wNDiag_15[10] , 
        \wCall_28[0] , \wPDiag_29[1] , \wColumn_8[16] , \wNDiag_18[8] , 
        \wNDiag_23[15] , \wPDiag_3[6] , \wPDiag_4[20] , \wPDiag_18[24] , 
        \wNDiag_21[1] , \wPDiag_4[13] , \wScan_5[2] , \wPDiag_10[8] , 
        \wNDiag_11[21] , \wNDiag_22[2] , \wPDiag_18[17] , \wNDiag_27[24] , 
        \wScan_6[1] , \wNDiag_11[12] , \wNDiag_27[17] , \wColumn_19[31] , 
        \wColumn_19[28] , \wColumn_20[3] , \wNDiag_1[13] , \wColumn_7[18] , 
        \wScan_12[2] , \wScan_11[1] , \wColumn_12[24] , \wColumn_23[0] , 
        \wColumn_24[21] , \wPDiag_13[31] , \wPDiag_13[28] , \wColumn_31[15] , 
        \wPDiag_16[6] , \wPDiag_30[19] , \wColumn_2[23] , \wPDiag_5[19] , 
        \wPDiag_5[8] , \wColumn_12[17] , \wPDiag_15[5] , \wColumn_24[12] , 
        \wColumn_31[26] , \wColumn_6[21] , \wNDiag_10[18] , \wColumn_18[22] , 
        \wColumn_18[11] , \wPDiag_18[0] , \wColumn_6[12] , \wPDiag_12[22] , 
        \wPDiag_24[27] , \wColumn_25[18] , \wPDiag_31[13] , \wNDiag_29[9] , 
        \wColumn_6[0] , \wPDiag_12[11] , \wPDiag_31[20] , \wNDiag_13[3] , 
        \wPDiag_24[14] , \wColumn_30[9] , \wPDiag_16[20] , \wNDiag_10[0] , 
        \wPDiag_20[25] , \wNDiag_29[20] , \wNDiag_4[31] , \wNDiag_4[28] , 
        \wColumn_5[3] , \wCall_6[0] , \wPDiag_1[31] , \wColumn_2[10] , 
        \wPDiag_16[13] , \wPDiag_20[16] , \wNDiag_29[13] , \wColumn_11[2] , 
        \wColumn_12[1] , \wScan_20[0] , \wColumn_21[30] , \wColumn_21[29] , 
        \wPDiag_21[9] , \wScan_23[3] , \wPDiag_24[4] , \wPDiag_1[28] , 
        \wPDiag_10[5] , \wPDiag_13[6] , \wNDiag_14[30] , \wNDiag_14[29] , 
        \wPDiag_27[7] , \wColumn_19[25] , \wScan_17[2] , \wColumn_19[16] , 
        \wColumn_25[3] , \wNDiag_27[30] , \wNDiag_27[29] , \wScan_0[2] , 
        \wScan_14[1] , \wPDiag_18[30] , \wColumn_26[0] , \wPDiag_18[29] , 
        \wPDiag_5[5] , \wColumn_7[26] , \wPDiag_15[8] , \wPDiag_1[25] , 
        \wNDiag_1[8] , \wScan_3[1] , \wColumn_3[24] , \wNDiag_4[5] , 
        \wPDiag_6[6] , \wPDiag_25[20] , \wPDiag_30[14] , \wColumn_7[15] , 
        \wColumn_12[30] , \wPDiag_13[25] , \wColumn_31[18] , \wColumn_12[29] , 
        \wNDiag_7[6] , \wPDiag_13[16] , \wNDiag_24[1] , \wPDiag_30[27] , 
        \wPDiag_17[27] , \wPDiag_25[13] , \wNDiag_27[2] , \wColumn_19[7] , 
        \wPDiag_21[22] , \wScan_28[5] , \wColumn_16[18] , \wNDiag_28[27] , 
        \wColumn_3[17] , \wPDiag_17[14] , \wPDiag_21[11] , \wNDiag_28[14] , 
        \wNDiag_18[5] , \wNDiag_4[25] , \wColumn_8[31] , \wNDiag_23[18] , 
        \wColumn_8[28] , \wColumn_17[21] , \wColumn_21[24] , \wPDiag_21[4] , 
        \wPDiag_22[7] , \wNDiag_4[16] , \wNDiag_9[0] , \wScan_25[0] , 
        \wColumn_17[12] , \wColumn_21[17] , \wColumn_17[1] , \wColumn_9[22] , 
        \wColumn_14[2] , \wPDiag_20[31] , \wPDiag_20[28] , \wScan_26[3] , 
        \wNDiag_14[24] , \wNDiag_22[21] , \wPDiag_1[16] , \wColumn_3[0] , 
        \wNDiag_16[3] , \wPDiag_24[9] , \wCall_3[0] , \wColumn_9[11] , 
        \wNDiag_14[17] , \wNDiag_15[0] , \wNDiag_22[12] , \wPDiag_5[27] , 
        \wScan_19[4] , \wPDiag_19[23] , \wColumn_28[6] , \wNDiag_31[6] , 
        \wPDiag_5[14] , \wNDiag_10[26] , \wNDiag_10[15] , \wPDiag_19[10] , 
        \wNDiag_26[23] , \wNDiag_26[10] , \wPDiag_24[19] , \wColumn_30[4] , 
        \wColumn_13[23] , \wColumn_25[26] , \wNDiag_29[4] , \wColumn_13[10] , 
        \wColumn_30[12] , \wColumn_25[15] , \wColumn_30[21] , \wColumn_2[27] , 
        \wColumn_3[9] , \wPDiag_8[0] , \wColumn_5[7] , \wColumn_9[18] , 
        \wColumn_11[6] , \wColumn_12[5] , \wNDiag_15[9] , \wScan_20[4] , 
        \wNDiag_22[31] , \wPDiag_27[3] , \wNDiag_22[28] , \wPDiag_24[0] , 
        \wNDiag_9[9] , \wColumn_2[14] , \wColumn_6[4] , \wNDiag_10[4] , 
        \wColumn_17[8] , \wNDiag_29[24] , \wNDiag_13[7] , \wPDiag_20[21] , 
        \wPDiag_16[24] , \wColumn_17[31] , \wColumn_17[28] , \wPDiag_12[26] , 
        \wPDiag_16[17] , \wNDiag_29[17] , \wPDiag_20[12] , \wPDiag_24[23] , 
        \wPDiag_31[17] , \wNDiag_1[24] , \wColumn_6[25] , \wPDiag_8[9] , 
        \wColumn_13[19] , \wColumn_30[31] , \wColumn_30[28] , \wColumn_6[16] , 
        \wPDiag_12[15] , \wPDiag_18[4] , \wPDiag_24[10] , \wPDiag_31[24] , 
        \wScan_8[3] , \wScan_11[5] , \wColumn_12[20] , \wColumn_18[26] , 
        \wPDiag_19[19] , \wNDiag_26[19] , \wColumn_18[15] , \wColumn_31[11] , 
        \wColumn_23[4] , \wColumn_24[25] , \wNDiag_24[8] , \wNDiag_1[17] , 
        \wColumn_12[13] , \wCall_14[0] , \wColumn_20[7] , \wColumn_24[16] , 
        \wColumn_31[22] , \wPDiag_15[1] , \wPDiag_4[24] , \wNDiag_11[25] , 
        \wPDiag_16[2] , \wPDiag_25[30] , \wPDiag_25[29] , \wNDiag_27[20] , 
        \wNDiag_22[6] , \wNDiag_1[26] , \wNDiag_1[1] , \wPDiag_3[2] , 
        \wPDiag_18[20] , \wNDiag_21[5] , \wColumn_26[9] , \wPDiag_4[17] , 
        \wScan_6[5] , \wNDiag_11[16] , \wColumn_8[21] , \wNDiag_15[27] , 
        \wPDiag_18[13] , \wNDiag_27[13] , \wPDiag_29[5] , \wNDiag_23[22] , 
        \wNDiag_2[2] , \wNDiag_23[11] , \wNDiag_5[26] , \wColumn_8[12] , 
        \wNDiag_15[14] , \wNDiag_5[15] , \wReturn_16[0] , \wColumn_16[22] , 
        \wColumn_20[27] , \wPDiag_21[18] , \wPDiag_31[7] , \wColumn_8[2] , 
        \wColumn_16[11] , \wColumn_20[14] , \wNDiag_1[15] , \wScan_12[4] , 
        \wColumn_20[5] , \wColumn_12[22] , \wColumn_23[6] , \wPDiag_25[18] , 
        \wNDiag_27[9] , \wColumn_24[27] , \wColumn_31[13] , \wPDiag_16[0] , 
        \wNDiag_1[3] , \wNDiag_2[0] , \wPDiag_3[0] , \wPDiag_4[26] , 
        \wColumn_12[11] , \wPDiag_15[3] , \wColumn_31[20] , \wPDiag_18[22] , 
        \wColumn_24[14] , \wNDiag_21[7] , \wNDiag_22[4] , \wPDiag_4[15] , 
        \wScan_5[4] , \wNDiag_11[27] , \wPDiag_18[11] , \wColumn_25[8] , 
        \wNDiag_27[22] , \wNDiag_11[14] , \wNDiag_27[11] , \wColumn_8[23] , 
        \wNDiag_23[20] , \wColumn_8[10] , \wNDiag_15[25] , \wNDiag_15[16] , 
        \wPDiag_29[7] , \wNDiag_23[13] , \wColumn_2[25] , \wNDiag_5[24] , 
        \wColumn_16[20] , \wColumn_20[25] , \wPDiag_31[5] , \wNDiag_5[17] , 
        \wColumn_8[0] , \wColumn_20[16] , \wColumn_16[13] , \wColumn_6[6] , 
        \wCall_8[0] , \wColumn_9[30] , \wColumn_9[29] , \wColumn_11[4] , 
        \wColumn_12[7] , \wPDiag_21[30] , \wPDiag_21[29] , \wCall_26[0] , 
        \wNDiag_16[8] , \wNDiag_22[19] , \wScan_23[5] , \wPDiag_24[2] , 
        \wNDiag_13[5] , \wPDiag_27[1] , \wPDiag_16[26] , \wPDiag_20[23] , 
        \wColumn_14[9] , \wColumn_17[19] , \wColumn_2[16] , \wColumn_5[5] , 
        \wNDiag_10[6] , \wNDiag_29[26] , \wPDiag_16[15] , \wPDiag_20[10] , 
        \wColumn_6[27] , \wPDiag_18[6] , \wNDiag_29[15] , \wPDiag_12[24] , 
        \wPDiag_24[21] , \wPDiag_31[15] , \wReturn_0[0] , \wPDiag_1[27] , 
        \wNDiag_4[27] , \wColumn_6[14] , \wColumn_13[31] , \wColumn_13[28] , 
        \wColumn_30[19] , \wScan_8[1] , \wPDiag_12[17] , \wColumn_18[24] , 
        \wPDiag_24[12] , \wPDiag_31[26] , \wReturn_24[0] , \wColumn_18[17] , 
        \wNDiag_26[31] , \wNDiag_26[28] , \wPDiag_19[31] , \wPDiag_19[28] , 
        \wPDiag_22[5] , \wNDiag_4[14] , \wColumn_14[0] , \wColumn_17[23] , 
        \wPDiag_20[19] , \wColumn_21[26] , \wPDiag_21[6] , \wScan_26[1] , 
        \wNDiag_9[2] , \wColumn_17[10] , \wColumn_17[3] , \wColumn_21[15] , 
        \wScan_25[2] , \wPDiag_1[14] , \wColumn_9[20] , \wNDiag_14[26] , 
        \wPDiag_27[8] , \wColumn_9[13] , \wNDiag_15[2] , \wNDiag_22[23] , 
        \wNDiag_14[15] , \wNDiag_22[10] , \wColumn_3[2] , \wPDiag_5[25] , 
        \wNDiag_10[24] , \wNDiag_16[1] , \wNDiag_26[21] , \wPDiag_5[16] , 
        \wPDiag_19[21] , \wColumn_28[4] , \wNDiag_31[4] , \wNDiag_10[17] , 
        \wNDiag_26[12] , \wColumn_13[21] , \wPDiag_19[12] , \wColumn_25[24] , 
        \wNDiag_29[6] , \wColumn_30[10] , \wColumn_30[6] , \wPDiag_3[9] , 
        \wPDiag_8[2] , \wColumn_25[17] , \wPDiag_10[7] , \wColumn_13[12] , 
        \wPDiag_18[18] , \wPDiag_24[31] , \wPDiag_24[28] , \wColumn_30[23] , 
        \wPDiag_13[4] , \wColumn_19[27] , \wNDiag_27[18] , \wColumn_26[2] , 
        \wScan_0[0] , \wScan_3[3] , \wPDiag_6[4] , \wPDiag_13[27] , 
        \wScan_14[3] , \wScan_17[0] , \wColumn_19[14] , \wColumn_25[1] , 
        \wPDiag_30[16] , \wPDiag_25[22] , \wPDiag_16[9] , \wColumn_2[21] , 
        \wNDiag_2[9] , \wColumn_3[26] , \wPDiag_5[7] , \wColumn_12[18] , 
        \wColumn_31[30] , \wColumn_31[29] , \wColumn_7[24] , \wColumn_7[17] , 
        \wPDiag_13[14] , \wPDiag_25[11] , \wNDiag_27[0] , \wPDiag_30[25] , 
        \wNDiag_24[3] , \wNDiag_28[25] , \wColumn_3[15] , \wNDiag_4[7] , 
        \wColumn_8[9] , \wNDiag_7[4] , \wColumn_16[30] , \wPDiag_17[25] , 
        \wColumn_19[5] , \wPDiag_21[20] , \wColumn_16[29] , \wNDiag_28[16] , 
        \wColumn_8[19] , \wPDiag_17[16] , \wPDiag_21[13] , \wReturn_5[0] , 
        \wPDiag_5[31] , \wScan_8[5] , \wNDiag_18[7] , \wNDiag_23[30] , 
        \wNDiag_23[29] , \wScan_30[5] , \wColumn_18[20] , \wNDiag_31[9] , 
        \wPDiag_5[28] , \wNDiag_10[30] , \wNDiag_10[29] , \wColumn_18[13] , 
        \wColumn_28[9] , \wPDiag_12[20] , \wPDiag_31[11] , \wPDiag_24[25] , 
        \wColumn_5[1] , \wColumn_6[23] , \wColumn_6[10] , \wPDiag_12[13] , 
        \wPDiag_18[2] , \wPDiag_24[16] , \wPDiag_31[22] , \wColumn_25[30] , 
        \wColumn_25[29] , \wNDiag_10[2] , \wNDiag_29[22] , \wColumn_2[12] , 
        \wNDiag_4[19] , \wColumn_21[18] , \wColumn_6[2] , \wPDiag_20[27] , 
        \wNDiag_13[1] , \wPDiag_16[22] , \wNDiag_29[11] , \wPDiag_16[11] , 
        \wReturn_18[0] , \wScan_0[4] , \wPDiag_1[19] , \wPDiag_20[14] , 
        \wPDiag_22[8] , \wNDiag_1[22] , \wNDiag_1[7] , \wColumn_3[18] , 
        \wNDiag_5[20] , \wColumn_11[0] , \wScan_23[1] , \wColumn_12[3] , 
        \wNDiag_14[18] , \wScan_20[2] , \wPDiag_24[6] , \wPDiag_27[5] , 
        \wNDiag_5[13] , \wNDiag_7[9] , \wColumn_16[24] , \wColumn_20[21] , 
        \wPDiag_31[1] , \wPDiag_17[31] , \wPDiag_17[28] , \wColumn_19[8] , 
        \wCall_30[0] , \wColumn_8[27] , \wColumn_8[4] , \wColumn_16[17] , 
        \wNDiag_15[21] , \wColumn_20[12] , \wNDiag_28[31] , \wNDiag_28[28] , 
        \wPDiag_29[3] , \wNDiag_23[24] , \wNDiag_2[4] , \wColumn_8[14] , 
        \wPDiag_3[4] , \wPDiag_4[22] , \wNDiag_11[23] , \wNDiag_15[12] , 
        \wNDiag_23[17] , \wNDiag_27[26] , \wPDiag_18[26] , \wColumn_19[19] , 
        \wNDiag_22[0] , \wNDiag_21[3] , \wPDiag_4[11] , \wScan_5[0] , 
        \wScan_6[3] , \wNDiag_11[10] , \wPDiag_13[9] , \wNDiag_27[15] , 
        \wScan_11[3] , \wColumn_12[26] , \wPDiag_18[15] , \wColumn_23[2] , 
        \wColumn_24[23] , \wColumn_31[17] , \wScan_12[0] , \wPDiag_13[19] , 
        \wColumn_20[1] , \wPDiag_30[31] , \wPDiag_30[28] , \wNDiag_1[11] , 
        \wColumn_7[30] , \wColumn_7[29] , \wColumn_12[15] , \wPDiag_15[7] , 
        \wColumn_24[10] , \wColumn_31[24] , \wColumn_3[22] , \wNDiag_4[3] , 
        \wPDiag_6[9] , \wPDiag_16[4] , \wNDiag_7[0] , \wNDiag_15[31] , 
        \wNDiag_18[3] , \wScan_30[1] , \wNDiag_15[28] , \wPDiag_17[21] , 
        \wColumn_19[1] , \wPDiag_21[24] , \wScan_28[3] , \wColumn_3[11] , 
        \wNDiag_5[30] , \wNDiag_28[21] , \wNDiag_5[29] , \wPDiag_17[12] , 
        \wPDiag_21[17] , \wPDiag_5[3] , \wColumn_7[20] , \wColumn_20[31] , 
        \wColumn_20[28] , \wNDiag_28[12] , \wPDiag_31[8] , \wNDiag_1[18] , 
        \wColumn_24[19] , \wPDiag_4[18] , \wPDiag_6[0] , \wPDiag_13[23] , 
        \wPDiag_25[26] , \wColumn_7[13] , \wPDiag_30[12] , \wPDiag_13[10] , 
        \wNDiag_24[7] , \wColumn_20[8] , \wPDiag_25[15] , \wPDiag_30[21] , 
        \wNDiag_27[4] , \wPDiag_10[3] , \wNDiag_11[19] , \wPDiag_13[0] , 
        \wColumn_19[23] , \wScan_17[4] , \wColumn_19[10] , \wColumn_25[5] , 
        \wNDiag_22[9] , \wColumn_6[19] , \wColumn_26[6] , \wColumn_30[2] , 
        \wColumn_25[20] , \wPDiag_8[6] , \wPDiag_12[30] , \wColumn_13[25] , 
        \wColumn_30[14] , \wNDiag_29[2] , \wPDiag_31[18] , \wPDiag_12[29] , 
        \wColumn_13[16] , \wColumn_30[27] , \wColumn_1[8] , \wPDiag_1[23] , 
        \wPDiag_5[21] , \wScan_19[2] , \wReturn_21[0] , \wColumn_25[13] , 
        \wPDiag_19[25] , \wColumn_28[0] , \wNDiag_31[0] , \wPDiag_5[12] , 
        \wNDiag_10[20] , \wNDiag_10[13] , \wPDiag_19[16] , \wNDiag_26[25] , 
        \wNDiag_26[16] , \wColumn_9[24] , \wColumn_18[30] , \wColumn_18[29] , 
        \wNDiag_22[27] , \wNDiag_14[22] , \wPDiag_1[10] , \wNDiag_16[5] , 
        \wColumn_2[31] , \wColumn_3[6] , \wNDiag_4[23] , \wColumn_9[17] , 
        \wColumn_11[9] , \wNDiag_14[11] , \wNDiag_22[14] , \wNDiag_15[6] , 
        \wPDiag_16[18] , \wColumn_17[27] , \wColumn_21[22] , \wPDiag_21[2] , 
        \wNDiag_29[18] , \wPDiag_22[1] , \wColumn_2[28] , \wNDiag_2[27] , 
        \wNDiag_2[14] , \wNDiag_4[10] , \wColumn_5[8] , \wNDiag_9[6] , 
        \wColumn_17[14] , \wColumn_17[7] , \wColumn_21[11] , \wCall_23[0] , 
        \wNDiag_13[8] , \wColumn_14[4] , \wScan_26[5] , \wColumn_11[10] , 
        \wPDiag_25[2] , \wPDiag_26[1] , \wColumn_27[15] , \wColumn_10[4] , 
        \wNDiag_17[8] , \wScan_22[5] , \wNDiag_19[19] , \wPDiag_26[19] , 
        \wPDiag_3[25] , \wPDiag_3[16] , \wColumn_4[5] , \wPDiag_7[14] , 
        \wColumn_11[23] , \wNDiag_12[15] , \wColumn_13[7] , \wCall_27[0] , 
        \wColumn_27[26] , \wNDiag_24[10] , \wNDiag_31[24] , \wNDiag_9[18] , 
        \wNDiag_11[6] , \wColumn_7[6] , \wPDiag_7[27] , \wNDiag_12[5] , 
        \wNDiag_12[26] , \wNDiag_24[23] , \wColumn_15[9] , \wNDiag_31[17] , 
        \wColumn_28[31] , \wColumn_28[28] , \wNDiag_16[24] , \wNDiag_16[17] , 
        \wNDiag_20[12] , \wPDiag_29[17] , \wNDiag_20[21] , \wNDiag_6[16] , 
        \wPDiag_8[30] , \wColumn_15[12] , \wPDiag_19[6] , \wPDiag_29[24] , 
        \wPDiag_8[29] , \wColumn_23[17] , \wScan_9[1] , \wColumn_15[21] , 
        \wPDiag_22[31] , \wPDiag_22[28] , \wColumn_23[24] , \wReturn_25[0] , 
        \wColumn_1[17] , \wPDiag_2[0] , \wNDiag_6[25] , \wScan_13[4] , 
        \wPDiag_14[3] , \wPDiag_17[0] , \wColumn_29[11] , \wColumn_21[5] , 
        \wColumn_22[6] , \wNDiag_21[18] , \wColumn_29[22] , \wPDiag_15[14] , 
        \wNDiag_26[9] , \wPDiag_23[11] , \wPDiag_1[3] , \wScan_4[4] , 
        \wPDiag_9[10] , \wPDiag_15[27] , \wPDiag_23[22] , \wNDiag_23[4] , 
        \wColumn_24[8] , \wColumn_1[24] , \wPDiag_9[23] , \wColumn_14[18] , 
        \wColumn_10[30] , \wColumn_10[29] , \wNDiag_20[7] , \wNDiag_3[0] , 
        \wColumn_5[15] , \wNDiag_18[13] , \wPDiag_11[16] , \wPDiag_27[13] , 
        \wColumn_5[26] , \wNDiag_18[20] , \wPDiag_28[7] , \wScan_1[0] , 
        \wPDiag_2[15] , \wPDiag_2[9] , \wNDiag_7[26] , \wNDiag_7[15] , 
        \wNDiag_8[21] , \wNDiag_8[12] , \wCall_9[0] , \wPDiag_11[25] , 
        \wNDiag_25[30] , \wPDiag_27[20] , \wNDiag_25[29] , \wColumn_9[0] , 
        \wPDiag_30[5] , \wScan_16[0] , \wPDiag_12[4] , \wColumn_14[11] , 
        \wColumn_22[14] , \wColumn_24[1] , \wColumn_27[2] , \wScan_15[3] , 
        \wPDiag_23[18] , \wPDiag_9[19] , \wColumn_14[22] , \wColumn_22[27] , 
        \wPDiag_11[7] , \wNDiag_17[14] , \wNDiag_25[3] , \wPDiag_28[14] , 
        \wNDiag_21[11] , \wNDiag_26[0] , \wScan_2[3] , \wPDiag_2[26] , 
        \wPDiag_4[7] , \wPDiag_28[27] , \wPDiag_7[4] , \wColumn_29[18] , 
        \wNDiag_5[7] , \wPDiag_6[24] , \wPDiag_6[17] , \wPDiag_17[9] , 
        \wNDiag_21[22] , \wNDiag_17[27] , \wNDiag_6[4] , \wNDiag_8[31] , 
        \wNDiag_13[16] , \wNDiag_25[13] , \wNDiag_30[27] , \wNDiag_8[28] , 
        \wNDiag_13[25] , \wNDiag_30[14] , \wColumn_18[5] , \wNDiag_25[20] , 
        \wColumn_9[9] , \wColumn_10[13] , \wNDiag_18[30] , \wNDiag_18[29] , 
        \wColumn_26[16] , \wNDiag_3[17] , \wColumn_10[20] , \wColumn_26[25] , 
        \wPDiag_27[30] , \wPDiag_27[29] , \wNDiag_19[7] , \wScan_31[5] , 
        \wReturn_1[0] , \wColumn_1[1] , \wColumn_2[2] , \wNDiag_3[24] , 
        \wNDiag_3[9] , \wNDiag_8[2] , \wColumn_16[3] , \wNDiag_9[22] , 
        \wNDiag_9[11] , \wColumn_15[0] , \wScan_24[2] , \wScan_27[1] , 
        \wPDiag_20[6] , \wPDiag_23[5] , \wNDiag_24[19] , \wColumn_4[16] , 
        \wPDiag_10[15] , \wNDiag_17[1] , \wPDiag_26[10] , \wColumn_4[25] , 
        \wPDiag_10[26] , \wNDiag_14[2] , \wNDiag_19[10] , \wPDiag_26[23] , 
        \wColumn_11[19] , \wPDiag_26[8] , \wNDiag_19[23] , \wColumn_15[31] , 
        \wNDiag_3[30] , \wNDiag_3[29] , \wPDiag_6[30] , \wPDiag_8[20] , 
        \wPDiag_8[13] , \wColumn_15[28] , \wPDiag_14[17] , \wPDiag_22[12] , 
        \wNDiag_30[4] , \wNDiag_8[16] , \wColumn_9[4] , \wPDiag_9[2] , 
        \wPDiag_14[24] , \wNDiag_20[31] , \wNDiag_20[28] , \wPDiag_22[21] , 
        \wColumn_29[4] , \wColumn_28[12] , \wColumn_28[21] , \wNDiag_28[6] , 
        \wColumn_31[6] , \wColumn_18[8] , \wPDiag_6[29] , \wNDiag_6[9] , 
        \wNDiag_13[28] , \wNDiag_8[25] , \wNDiag_13[31] , \wNDiag_30[19] , 
        \wCall_31[0] , \wPDiag_30[1] , \wNDiag_3[4] , \wColumn_5[11] , 
        \wPDiag_11[12] , \wPDiag_27[17] , \wNDiag_18[17] , \wColumn_26[31] , 
        \wPDiag_11[21] , \wColumn_26[28] , \wPDiag_27[24] , \wColumn_1[20] , 
        \wColumn_1[13] , \wPDiag_1[7] , \wScan_4[0] , \wColumn_5[22] , 
        \wNDiag_18[24] , \wPDiag_28[3] , \wPDiag_9[14] , \wPDiag_2[4] , 
        \wScan_7[3] , \wPDiag_15[10] , \wPDiag_23[15] , \wPDiag_12[9] , 
        \wNDiag_20[3] , \wPDiag_2[18] , \wPDiag_7[9] , \wNDiag_7[18] , 
        \wPDiag_9[27] , \wColumn_22[19] , \wPDiag_15[23] , \wPDiag_17[4] , 
        \wPDiag_23[26] , \wNDiag_23[0] , \wScan_13[0] , \wPDiag_14[7] , 
        \wColumn_29[15] , \wNDiag_6[21] , \wNDiag_6[12] , \wScan_10[3] , 
        \wNDiag_17[19] , \wColumn_29[26] , \wColumn_21[1] , \wColumn_22[2] , 
        \wPDiag_28[19] , \wPDiag_14[30] , \wPDiag_14[29] , \wColumn_29[9] , 
        \wColumn_15[16] , \wColumn_23[13] , \wNDiag_30[9] , \wColumn_1[5] , 
        \wNDiag_2[23] , \wNDiag_2[10] , \wPDiag_3[21] , \wPDiag_3[12] , 
        \wScan_9[5] , \wColumn_15[25] , \wNDiag_16[13] , \wColumn_23[20] , 
        \wPDiag_29[13] , \wNDiag_20[16] , \wReturn_4[0] , \wPDiag_19[2] , 
        \wPDiag_29[20] , \wColumn_4[31] , \wColumn_4[28] , \wColumn_4[1] , 
        \wColumn_7[2] , \wPDiag_7[10] , \wNDiag_16[20] , \wNDiag_20[25] , 
        \wNDiag_12[22] , \wNDiag_12[11] , \wPDiag_23[8] , \wNDiag_24[14] , 
        \wNDiag_31[20] , \wReturn_19[0] , \wNDiag_31[13] , \wNDiag_24[27] , 
        \wPDiag_7[23] , \wNDiag_12[1] , \wNDiag_11[2] , \wColumn_11[14] , 
        \wPDiag_25[6] , \wPDiag_26[5] , \wColumn_27[11] , \wColumn_10[0] , 
        \wPDiag_10[18] , \wColumn_11[27] , \wColumn_13[3] , \wColumn_27[22] , 
        \wScan_21[2] , \wScan_22[1] , \wPDiag_3[31] , \wPDiag_3[28] , 
        \wPDiag_9[6] , \wPDiag_29[30] , \wPDiag_29[29] , \wReturn_20[0] , 
        \wColumn_28[16] , \wColumn_4[12] , \wNDiag_6[31] , \wNDiag_16[30] , 
        \wNDiag_16[29] , \wColumn_28[25] , \wNDiag_28[2] , \wColumn_31[2] , 
        \wNDiag_6[28] , \wPDiag_8[24] , \wPDiag_8[17] , \wPDiag_14[13] , 
        \wPDiag_22[16] , \wPDiag_14[20] , \wPDiag_22[25] , \wColumn_23[30] , 
        \wColumn_23[29] , \wColumn_29[0] , \wNDiag_14[6] , \wScan_18[2] , 
        \wNDiag_30[0] , \wNDiag_19[14] , \wColumn_2[6] , \wPDiag_10[11] , 
        \wNDiag_17[5] , \wPDiag_26[14] , \wNDiag_2[19] , \wColumn_4[21] , 
        \wColumn_10[9] , \wNDiag_19[27] , \wColumn_27[18] , \wNDiag_3[20] , 
        \wNDiag_3[13] , \wColumn_4[8] , \wNDiag_9[15] , \wPDiag_10[22] , 
        \wNDiag_12[8] , \wColumn_15[4] , \wPDiag_26[27] , \wScan_27[5] , 
        \wPDiag_7[19] , \wNDiag_8[6] , \wColumn_16[7] , \wCall_22[0] , 
        \wNDiag_9[26] , \wNDiag_12[18] , \wNDiag_31[29] , \wPDiag_20[2] , 
        \wPDiag_23[1] , \wNDiag_31[30] , \wPDiag_11[31] , \wPDiag_11[28] , 
        \wColumn_10[17] , \wColumn_26[12] , \wScan_32[2] , \wPDiag_2[11] , 
        \wColumn_5[18] , \wScan_31[1] , \wNDiag_5[3] , \wPDiag_6[13] , 
        \wColumn_10[24] , \wNDiag_13[12] , \wNDiag_19[3] , \wColumn_26[21] , 
        \wPDiag_30[8] , \wNDiag_25[17] , \wNDiag_30[23] , \wScan_29[3] , 
        \wPDiag_6[20] , \wNDiag_6[0] , \wNDiag_13[21] , \wColumn_18[1] , 
        \wNDiag_25[24] , \wNDiag_30[10] , \wColumn_21[8] , \wNDiag_26[4] , 
        \wNDiag_21[15] , \wScan_1[4] , \wPDiag_2[22] , \wPDiag_7[0] , 
        \wNDiag_17[23] , \wNDiag_17[10] , \wNDiag_25[7] , \wPDiag_28[10] , 
        \wNDiag_21[26] , \wPDiag_4[3] , \wPDiag_28[23] , \wColumn_1[30] , 
        \wColumn_1[29] , \wNDiag_3[11] , \wColumn_5[30] , \wNDiag_7[22] , 
        \wNDiag_7[11] , \wColumn_14[15] , \wColumn_27[6] , \wColumn_22[10] , 
        \wColumn_24[5] , \wPDiag_11[3] , \wScan_16[4] , \wNDiag_23[9] , 
        \wColumn_14[26] , \wColumn_22[23] , \wPDiag_15[19] , \wPDiag_12[0] , 
        \wPDiag_28[8] , \wColumn_5[29] , \wColumn_10[15] , \wReturn_12[0] , 
        \wColumn_26[10] , \wColumn_10[26] , \wNDiag_19[1] , \wColumn_26[23] , 
        \wScan_31[3] , \wColumn_1[18] , \wScan_2[5] , \wPDiag_2[20] , 
        \wPDiag_2[13] , \wNDiag_3[22] , \wPDiag_11[19] , \wScan_32[0] , 
        \wNDiag_5[1] , \wPDiag_6[22] , \wPDiag_6[11] , \wNDiag_6[2] , 
        \wNDiag_13[10] , \wNDiag_25[15] , \wNDiag_30[21] , \wNDiag_13[23] , 
        \wColumn_18[3] , \wNDiag_25[26] , \wNDiag_30[12] , \wNDiag_17[12] , 
        \wColumn_22[9] , \wNDiag_25[5] , \wScan_29[1] , \wPDiag_28[12] , 
        \wNDiag_21[17] , \wNDiag_26[6] , \wPDiag_4[1] , \wPDiag_28[21] , 
        \wPDiag_7[2] , \wNDiag_21[24] , \wNDiag_7[20] , \wNDiag_7[13] , 
        \wPDiag_15[31] , \wNDiag_17[21] , \wPDiag_15[28] , \wCall_10[0] , 
        \wColumn_14[17] , \wColumn_22[12] , \wColumn_24[7] , \wScan_15[5] , 
        \wNDiag_20[8] , \wColumn_27[4] , \wPDiag_12[2] , \wPDiag_3[19] , 
        \wPDiag_9[4] , \wPDiag_11[1] , \wColumn_14[24] , \wPDiag_19[9] , 
        \wColumn_22[21] , \wColumn_28[14] , \wColumn_28[27] , \wPDiag_8[15] , 
        \wNDiag_16[18] , \wNDiag_28[0] , \wPDiag_29[18] , \wColumn_31[0] , 
        \wColumn_1[7] , \wColumn_2[4] , \wNDiag_2[31] , \wNDiag_6[19] , 
        \wPDiag_8[26] , \wPDiag_14[11] , \wPDiag_22[14] , \wNDiag_30[2] , 
        \wScan_18[0] , \wColumn_23[18] , \wPDiag_14[22] , \wPDiag_22[27] , 
        \wColumn_29[2] , \wNDiag_2[28] , \wPDiag_10[13] , \wNDiag_17[7] , 
        \wPDiag_26[16] , \wColumn_4[23] , \wColumn_4[10] , \wPDiag_10[20] , 
        \wColumn_13[8] , \wNDiag_14[4] , \wNDiag_19[16] , \wColumn_27[29] , 
        \wPDiag_26[25] , \wColumn_27[30] , \wNDiag_19[25] , \wNDiag_6[10] , 
        \wColumn_7[9] , \wNDiag_8[4] , \wColumn_16[5] , \wNDiag_9[17] , 
        \wNDiag_11[9] , \wScan_24[4] , \wPDiag_7[31] , \wPDiag_7[28] , 
        \wNDiag_9[24] , \wNDiag_12[30] , \wNDiag_12[29] , \wColumn_15[6] , 
        \wNDiag_31[18] , \wColumn_15[14] , \wPDiag_20[0] , \wPDiag_23[3] , 
        \wColumn_23[11] , \wColumn_15[27] , \wColumn_23[22] , \wPDiag_3[10] , 
        \wNDiag_6[23] , \wPDiag_14[18] , \wNDiag_16[22] , \wNDiag_16[11] , 
        \wNDiag_20[14] , \wColumn_31[9] , \wNDiag_28[9] , \wPDiag_29[11] , 
        \wScanEnable[0] , \wNDiag_2[21] , \wNDiag_2[12] , \wPDiag_3[23] , 
        \wNDiag_20[27] , \wColumn_4[3] , \wPDiag_7[12] , \wNDiag_12[13] , 
        \wPDiag_19[0] , \wPDiag_20[9] , \wPDiag_29[22] , \wNDiag_31[22] , 
        \wNDiag_24[16] , \wNDiag_11[0] , \wCall_7[0] , \wColumn_7[0] , 
        \wPDiag_7[21] , \wNDiag_12[3] , \wPDiag_10[30] , \wPDiag_10[29] , 
        \wNDiag_12[20] , \wNDiag_24[25] , \wNDiag_31[11] , \wColumn_10[2] , 
        \wColumn_11[16] , \wPDiag_26[7] , \wColumn_27[13] , \wPDiag_25[4] , 
        \wColumn_4[19] , \wScan_21[0] , \wScan_22[3] , \wNDiag_5[8] , 
        \wNDiag_8[14] , \wColumn_11[25] , \wColumn_13[1] , \wColumn_27[20] , 
        \wColumn_9[6] , \wPDiag_6[18] , \wNDiag_8[27] , \wNDiag_13[19] , 
        \wNDiag_30[31] , \wPDiag_30[3] , \wNDiag_30[28] , \wNDiag_19[8] , 
        \wNDiag_3[6] , \wColumn_5[13] , \wNDiag_18[15] , \wPDiag_11[10] , 
        \wPDiag_27[15] , \wCall_29[0] , \wColumn_5[20] , \wNDiag_18[26] , 
        \wPDiag_28[1] , \wScan_1[2] , \wColumn_1[22] , \wColumn_1[11] , 
        \wPDiag_2[6] , \wNDiag_3[18] , \wColumn_26[19] , \wScan_7[1] , 
        \wNDiag_7[30] , \wNDiag_7[29] , \wPDiag_11[23] , \wPDiag_27[26] , 
        \wPDiag_15[12] , \wPDiag_23[17] , \wPDiag_1[5] , \wScan_4[2] , 
        \wPDiag_9[16] , \wPDiag_11[8] , \wColumn_22[31] , \wColumn_22[28] , 
        \wPDiag_9[25] , \wPDiag_15[21] , \wPDiag_23[24] , \wNDiag_23[2] , 
        \wNDiag_20[1] , \wColumn_1[3] , \wCall_2[0] , \wPDiag_2[30] , 
        \wPDiag_4[8] , \wPDiag_14[5] , \wPDiag_28[31] , \wPDiag_28[28] , 
        \wPDiag_2[29] , \wNDiag_8[0] , \wNDiag_9[13] , \wScan_10[1] , 
        \wPDiag_17[6] , \wNDiag_17[31] , \wNDiag_17[28] , \wColumn_29[17] , 
        \wScan_13[2] , \wColumn_21[3] , \wColumn_22[0] , \wColumn_29[24] , 
        \wColumn_15[2] , \wNDiag_24[31] , \wNDiag_24[28] , \wScan_27[3] , 
        \wScan_24[0] , \wNDiag_9[20] , \wColumn_16[1] , \wPDiag_20[4] , 
        \wPDiag_23[7] , \wColumn_11[31] , \wColumn_11[28] , \wNDiag_14[0] , 
        \wNDiag_19[12] , \wPDiag_1[8] , \wColumn_2[0] , \wColumn_4[14] , 
        \wNDiag_17[3] , \wPDiag_26[12] , \wColumn_4[27] , \wPDiag_10[17] , 
        \wNDiag_7[17] , \wPDiag_8[22] , \wPDiag_8[11] , \wPDiag_10[24] , 
        \wNDiag_19[21] , \wPDiag_25[9] , \wPDiag_14[15] , \wPDiag_26[21] , 
        \wPDiag_22[10] , \wPDiag_14[26] , \wPDiag_22[23] , \wColumn_29[6] , 
        \wColumn_15[19] , \wScan_18[4] , \wPDiag_9[31] , \wPDiag_9[28] , 
        \wPDiag_9[0] , \wNDiag_30[6] , \wColumn_14[13] , \wScan_15[1] , 
        \wNDiag_20[19] , \wColumn_28[10] , \wNDiag_28[4] , \wColumn_28[23] , 
        \wColumn_31[4] , \wColumn_22[16] , \wColumn_27[0] , \wColumn_24[3] , 
        \wPDiag_11[5] , \wScan_16[2] , \wPDiag_23[30] , \wPDiag_23[29] , 
        \wColumn_22[25] , \wColumn_14[20] , \wScan_2[1] , \wPDiag_2[17] , 
        \wNDiag_7[24] , \wPDiag_12[6] , \wNDiag_17[25] , \wNDiag_17[16] , 
        \wNDiag_21[13] , \wNDiag_26[2] , \wColumn_29[30] , \wColumn_29[29] , 
        \wNDiag_25[1] , \wPDiag_28[16] , \wPDiag_2[24] , \wNDiag_21[20] , 
        \wPDiag_4[5] , \wPDiag_7[6] , \wPDiag_14[8] , \wPDiag_28[25] , 
        \wNDiag_3[26] , \wNDiag_3[15] , \wNDiag_5[5] , \wPDiag_6[15] , 
        \wNDiag_13[14] , \wNDiag_30[25] , \wNDiag_25[11] , \wScan_29[5] , 
        \wPDiag_6[26] , \wNDiag_8[19] , \wNDiag_6[6] , \wColumn_18[7] , 
        \wNDiag_25[22] , \wNDiag_30[16] , \wNDiag_13[27] , \wColumn_10[11] , 
        \wColumn_26[14] , \wPDiag_27[18] , \wScan_32[4] , \wColumn_10[22] , 
        \wNDiag_18[18] , \wNDiag_19[5] , \wColumn_26[27] , \wColumn_1[26] , 
        \wColumn_1[15] , \wPDiag_1[1] , \wPDiag_9[12] , \wScan_10[5] , 
        \wPDiag_14[1] , \wPDiag_17[2] , \wNDiag_21[30] , \wNDiag_21[29] , 
        \wColumn_29[13] , \wCall_15[0] , \wColumn_29[20] , \wColumn_21[7] , 
        \wColumn_22[4] , \wNDiag_25[8] , \wColumn_14[30] , \wColumn_14[29] , 
        \wPDiag_2[2] , \wPDiag_23[13] , \wScan_7[5] , \wPDiag_15[16] , 
        \wNDiag_3[2] , \wPDiag_9[21] , \wNDiag_20[5] , \wPDiag_15[25] , 
        \wColumn_27[9] , \wPDiag_23[20] , \wNDiag_23[6] , \wPDiag_11[14] , 
        \wColumn_5[17] , \wPDiag_27[11] , \wNDiag_18[11] , \wColumn_10[18] , 
        \wPDiag_11[27] , \wPDiag_27[22] , \wColumn_2[9] , \wNDiag_2[16] , 
        \wColumn_5[24] , \wNDiag_18[22] , \wPDiag_28[5] , \wNDiag_8[23] , 
        \wNDiag_8[10] , \wColumn_9[2] , \wColumn_11[12] , \wReturn_17[0] , 
        \wNDiag_25[18] , \wPDiag_30[7] , \wNDiag_19[31] , \wNDiag_19[28] , 
        \wPDiag_25[0] , \wPDiag_26[3] , \wColumn_27[17] , \wColumn_11[21] , 
        \wColumn_13[5] , \wPDiag_26[31] , \wPDiag_26[28] , \wColumn_27[24] , 
        \wNDiag_14[9] , \wScan_21[4] , \wNDiag_2[25] , \wPDiag_3[27] , 
        \wPDiag_3[14] , \wColumn_4[7] , \wColumn_7[4] , \wPDiag_7[16] , 
        \wColumn_10[6] , \wNDiag_9[30] , \wNDiag_9[29] , \wNDiag_12[17] , 
        \wNDiag_24[12] , \wNDiag_31[26] , \wNDiag_12[24] , \wNDiag_24[21] , 
        \wNDiag_31[15] , \wPDiag_7[25] , \wNDiag_12[7] , \wNDiag_8[9] , 
        \wNDiag_11[4] , \wColumn_16[8] , \wNDiag_16[15] , \wPDiag_29[15] , 
        \wNDiag_20[10] , \wPDiag_9[9] , \wPDiag_19[4] , \wPDiag_29[26] , 
        \wColumn_28[19] , \wNDiag_6[27] , \wNDiag_6[14] , \wNDiag_16[26] , 
        \wNDiag_20[23] , \wColumn_15[10] , \wColumn_23[15] , \wScan_9[3] , 
        \wPDiag_22[19] , \wScan_1[3] , \wColumn_1[2] , \wColumn_2[1] , 
        \wPDiag_8[18] , \wColumn_15[23] , \wPDiag_10[16] , \wColumn_23[26] , 
        \wColumn_11[30] , \wColumn_11[29] , \wNDiag_17[2] , \wPDiag_26[13] , 
        \wReturn_2[0] , \wColumn_4[26] , \wColumn_4[15] , \wPDiag_10[25] , 
        \wNDiag_14[1] , \wNDiag_19[13] , \wPDiag_26[20] , \wNDiag_19[20] , 
        \wPDiag_8[10] , \wNDiag_8[1] , \wPDiag_25[8] , \wPDiag_9[1] , 
        \wNDiag_9[21] , \wNDiag_9[12] , \wScan_24[1] , \wColumn_15[3] , 
        \wColumn_16[0] , \wPDiag_20[5] , \wNDiag_24[30] , \wNDiag_24[29] , 
        \wScan_27[2] , \wPDiag_23[6] , \wColumn_28[11] , \wNDiag_20[18] , 
        \wColumn_28[22] , \wColumn_31[5] , \wNDiag_28[5] , \wPDiag_2[16] , 
        \wPDiag_8[23] , \wPDiag_14[14] , \wPDiag_22[11] , \wPDiag_14[27] , 
        \wColumn_15[18] , \wScan_18[5] , \wNDiag_30[7] , \wPDiag_22[22] , 
        \wNDiag_25[0] , \wPDiag_28[17] , \wColumn_29[7] , \wNDiag_26[3] , 
        \wColumn_29[31] , \wPDiag_4[4] , \wNDiag_17[17] , \wColumn_29[28] , 
        \wNDiag_21[12] , \wPDiag_1[9] , \wScan_2[0] , \wPDiag_14[9] , 
        \wNDiag_21[21] , \wPDiag_28[24] , \wPDiag_2[25] , \wPDiag_7[7] , 
        \wNDiag_17[24] , \wNDiag_7[25] , \wNDiag_7[16] , \wPDiag_9[30] , 
        \wScan_15[0] , \wScan_16[3] , \wColumn_24[2] , \wPDiag_23[31] , 
        \wPDiag_23[28] , \wPDiag_9[29] , \wColumn_22[17] , \wColumn_14[12] , 
        \wColumn_27[1] , \wPDiag_11[4] , \wPDiag_12[7] , \wColumn_14[21] , 
        \wColumn_22[24] , \wNDiag_3[14] , \wColumn_10[10] , \wColumn_26[15] , 
        \wNDiag_18[19] , \wNDiag_3[27] , \wColumn_10[23] , \wNDiag_19[4] , 
        \wColumn_26[26] , \wColumn_1[27] , \wColumn_1[14] , \wPDiag_2[3] , 
        \wNDiag_5[4] , \wPDiag_6[27] , \wPDiag_6[14] , \wNDiag_13[15] , 
        \wNDiag_25[10] , \wPDiag_27[19] , \wScan_32[5] , \wNDiag_30[24] , 
        \wColumn_18[6] , \wNDiag_6[7] , \wNDiag_13[26] , \wNDiag_25[23] , 
        \wNDiag_30[17] , \wNDiag_8[18] , \wScan_29[4] , \wPDiag_15[17] , 
        \wScan_7[4] , \wPDiag_23[12] , \wPDiag_9[13] , \wColumn_14[31] , 
        \wColumn_14[28] , \wPDiag_1[0] , \wPDiag_15[24] , \wPDiag_23[21] , 
        \wNDiag_23[7] , \wNDiag_20[4] , \wColumn_5[16] , \wNDiag_8[22] , 
        \wNDiag_8[11] , \wColumn_9[3] , \wPDiag_9[20] , \wColumn_27[8] , 
        \wScan_10[4] , \wPDiag_14[0] , \wPDiag_17[3] , \wNDiag_21[31] , 
        \wNDiag_21[28] , \wColumn_22[5] , \wColumn_29[12] , \wNDiag_25[9] , 
        \wColumn_21[6] , \wColumn_29[21] , \wNDiag_25[19] , \wNDiag_18[10] , 
        \wPDiag_30[6] , \wNDiag_3[3] , \wPDiag_27[10] , \wPDiag_11[15] , 
        \wColumn_2[8] , \wNDiag_2[17] , \wColumn_4[6] , \wColumn_5[25] , 
        \wColumn_10[19] , \wPDiag_7[17] , \wNDiag_9[31] , \wPDiag_11[26] , 
        \wNDiag_18[23] , \wPDiag_28[4] , \wPDiag_27[23] , \wNDiag_9[28] , 
        \wNDiag_11[5] , \wNDiag_12[16] , \wNDiag_31[27] , \wNDiag_24[13] , 
        \wColumn_7[5] , \wPDiag_7[24] , \wNDiag_8[8] , \wNDiag_12[25] , 
        \wColumn_16[9] , \wNDiag_24[20] , \wNDiag_31[14] , \wNDiag_12[6] , 
        \wColumn_11[13] , \wNDiag_19[30] , \wPDiag_26[30] , \wPDiag_26[29] , 
        \wPDiag_26[2] , \wNDiag_19[29] , \wColumn_27[16] , \wPDiag_25[1] , 
        \wNDiag_2[24] , \wColumn_10[7] , \wCall_24[0] , \wNDiag_6[15] , 
        \wColumn_11[20] , \wColumn_13[4] , \wColumn_27[25] , \wNDiag_14[8] , 
        \wColumn_15[11] , \wScan_21[5] , \wColumn_23[14] , \wPDiag_3[26] , 
        \wPDiag_3[15] , \wNDiag_6[26] , \wPDiag_8[19] , \wScan_9[2] , 
        \wColumn_15[22] , \wColumn_23[27] , \wNDiag_16[14] , \wNDiag_20[11] , 
        \wPDiag_22[18] , \wReturn_26[0] , \wColumn_28[18] , \wPDiag_29[14] , 
        \wNDiag_3[10] , \wNDiag_5[0] , \wPDiag_6[10] , \wPDiag_9[8] , 
        \wNDiag_16[27] , \wNDiag_20[22] , \wPDiag_29[27] , \wPDiag_19[5] , 
        \wNDiag_13[11] , \wNDiag_30[20] , \wNDiag_25[14] , \wScan_29[0] , 
        \wPDiag_6[23] , \wNDiag_6[3] , \wNDiag_25[27] , \wNDiag_30[13] , 
        \wNDiag_13[22] , \wColumn_18[2] , \wColumn_5[31] , \wColumn_5[28] , 
        \wColumn_10[14] , \wColumn_26[11] , \wPDiag_28[9] , \wPDiag_11[18] , 
        \wScan_32[1] , \wColumn_1[19] , \wNDiag_3[23] , \wNDiag_7[12] , 
        \wColumn_10[27] , \wNDiag_19[0] , \wColumn_14[16] , \wColumn_26[22] , 
        \wScan_31[2] , \wScan_15[4] , \wNDiag_20[9] , \wColumn_22[13] , 
        \wColumn_27[5] , \wPDiag_15[30] , \wPDiag_15[29] , \wColumn_24[6] , 
        \wScan_2[4] , \wPDiag_2[21] , \wPDiag_2[12] , \wNDiag_7[21] , 
        \wPDiag_11[0] , \wColumn_22[20] , \wPDiag_12[3] , \wColumn_14[25] , 
        \wNDiag_17[13] , \wNDiag_21[16] , \wColumn_22[8] , \wNDiag_25[4] , 
        \wNDiag_26[7] , \wPDiag_28[13] , \wPDiag_7[3] , \wNDiag_17[20] , 
        \wPDiag_4[0] , \wNDiag_21[25] , \wPDiag_28[20] , \wPDiag_8[14] , 
        \wPDiag_14[10] , \wPDiag_22[15] , \wColumn_1[6] , \wPDiag_3[18] , 
        \wNDiag_6[18] , \wPDiag_8[27] , \wPDiag_14[23] , \wPDiag_22[26] , 
        \wColumn_29[3] , \wScan_18[1] , \wNDiag_30[3] , \wPDiag_9[5] , 
        \wPDiag_19[8] , \wColumn_23[19] , \wReturn_23[0] , \wColumn_28[26] , 
        \wColumn_28[15] , \wNDiag_28[1] , \wPDiag_29[19] , \wColumn_7[8] , 
        \wPDiag_7[30] , \wNDiag_16[19] , \wColumn_31[1] , \wPDiag_7[29] , 
        \wNDiag_8[5] , \wNDiag_9[16] , \wNDiag_12[31] , \wNDiag_12[28] , 
        \wCall_21[0] , \wColumn_15[7] , \wColumn_16[4] , \wNDiag_31[19] , 
        \wNDiag_11[8] , \wScan_24[5] , \wNDiag_9[25] , \wPDiag_23[2] , 
        \wNDiag_14[5] , \wNDiag_19[17] , \wPDiag_20[1] , \wColumn_2[5] , 
        \wNDiag_2[30] , \wNDiag_2[29] , \wColumn_4[11] , \wColumn_13[9] , 
        \wColumn_27[31] , \wColumn_27[28] , \wNDiag_17[6] , \wPDiag_26[17] , 
        \wPDiag_3[22] , \wPDiag_3[11] , \wColumn_4[22] , \wPDiag_10[12] , 
        \wPDiag_10[21] , \wNDiag_19[24] , \wCall_18[0] , \wPDiag_26[24] , 
        \wNDiag_28[8] , \wPDiag_29[10] , \wReturn_7[0] , \wNDiag_16[10] , 
        \wPDiag_19[1] , \wNDiag_20[15] , \wColumn_31[8] , \wNDiag_20[26] , 
        \wPDiag_29[23] , \wNDiag_16[23] , \wNDiag_6[22] , \wNDiag_6[11] , 
        \wPDiag_14[19] , \wColumn_15[15] , \wColumn_23[10] , \wColumn_15[26] , 
        \wColumn_23[23] , \wNDiag_2[20] , \wNDiag_2[13] , \wPDiag_10[31] , 
        \wColumn_11[17] , \wPDiag_25[5] , \wColumn_27[12] , \wPDiag_10[28] , 
        \wPDiag_26[6] , \wColumn_4[18] , \wColumn_11[24] , \wColumn_13[0] , 
        \wScan_21[1] , \wColumn_27[21] , \wNDiag_3[7] , \wColumn_4[2] , 
        \wColumn_7[1] , \wPDiag_7[13] , \wColumn_10[3] , \wNDiag_12[12] , 
        \wScan_22[2] , \wNDiag_24[17] , \wNDiag_31[23] , \wPDiag_20[8] , 
        \wPDiag_7[20] , \wNDiag_12[2] , \wNDiag_12[21] , \wNDiag_24[24] , 
        \wNDiag_31[10] , \wPDiag_11[11] , \wNDiag_11[1] , \wPDiag_27[14] , 
        \wNDiag_3[19] , \wColumn_5[12] , \wNDiag_19[9] , \wNDiag_18[14] , 
        \wColumn_5[21] , \wPDiag_11[22] , \wPDiag_27[27] , \wNDiag_18[27] , 
        \wPDiag_28[0] , \wColumn_26[18] , \wColumn_1[23] , \wColumn_1[10] , 
        \wPDiag_1[4] , \wPDiag_2[31] , \wPDiag_2[28] , \wNDiag_5[9] , 
        \wNDiag_8[15] , \wColumn_9[7] , \wPDiag_6[19] , \wNDiag_8[26] , 
        \wPDiag_30[2] , \wCall_32[0] , \wNDiag_13[18] , \wNDiag_30[30] , 
        \wNDiag_30[29] , \wColumn_29[16] , \wPDiag_4[9] , \wPDiag_14[4] , 
        \wPDiag_17[7] , \wNDiag_17[30] , \wNDiag_17[29] , \wPDiag_28[30] , 
        \wPDiag_28[29] , \wReturn_30[0] , \wScan_10[0] , \wScan_13[3] , 
        \wColumn_21[2] , \wColumn_29[25] , \wColumn_22[1] , \wPDiag_2[7] , 
        \wScan_4[3] , \wScan_7[0] , \wPDiag_9[17] , \wColumn_22[29] , 
        \wPDiag_11[9] , \wColumn_22[30] , \wNDiag_7[31] , \wNDiag_7[28] , 
        \wPDiag_23[16] , \wPDiag_9[24] , \wPDiag_15[13] , \wColumn_5[10] , 
        \wPDiag_15[20] , \wNDiag_20[0] , \wNDiag_23[3] , \wNDiag_18[16] , 
        \wPDiag_23[25] , \wColumn_26[30] , \wColumn_26[29] , \wNDiag_3[31] , 
        \wNDiag_3[28] , \wNDiag_3[5] , \wPDiag_11[13] , \wPDiag_27[16] , 
        \wColumn_1[21] , \wColumn_1[12] , \wPDiag_2[19] , \wColumn_5[23] , 
        \wPDiag_6[31] , \wPDiag_6[28] , \wPDiag_11[20] , \wNDiag_18[25] , 
        \wPDiag_28[2] , \wPDiag_27[25] , \wNDiag_6[8] , \wNDiag_13[30] , 
        \wColumn_18[9] , \wNDiag_30[18] , \wNDiag_13[29] , \wPDiag_7[8] , 
        \wNDiag_8[24] , \wNDiag_8[17] , \wColumn_9[5] , \wPDiag_14[6] , 
        \wPDiag_30[0] , \wPDiag_17[5] , \wColumn_29[14] , \wScan_10[2] , 
        \wColumn_22[3] , \wPDiag_28[18] , \wPDiag_2[5] , \wScan_13[1] , 
        \wColumn_29[27] , \wPDiag_15[11] , \wNDiag_17[18] , \wColumn_21[0] , 
        \wPDiag_23[14] , \wScan_4[1] , \wScan_7[2] , \wPDiag_12[8] , 
        \wPDiag_9[15] , \wPDiag_1[6] , \wNDiag_7[19] , \wReturn_28[0] , 
        \wPDiag_15[22] , \wPDiag_23[27] , \wNDiag_23[1] , \wPDiag_3[20] , 
        \wPDiag_3[13] , \wPDiag_9[26] , \wNDiag_20[2] , \wColumn_22[18] , 
        \wNDiag_16[12] , \wNDiag_20[17] , \wPDiag_29[12] , \wNDiag_6[13] , 
        \wPDiag_14[31] , \wColumn_15[17] , \wNDiag_16[21] , \wPDiag_19[3] , 
        \wNDiag_20[24] , \wPDiag_29[21] , \wColumn_23[12] , \wColumn_29[8] , 
        \wNDiag_30[8] , \wPDiag_14[28] , \wScan_9[4] , \wColumn_1[4] , 
        \wColumn_2[7] , \wNDiag_2[22] , \wNDiag_2[11] , \wNDiag_6[20] , 
        \wColumn_15[24] , \wColumn_23[21] , \wColumn_4[30] , \wPDiag_26[4] , 
        \wColumn_4[29] , \wPDiag_10[19] , \wColumn_11[15] , \wPDiag_25[7] , 
        \wColumn_27[10] , \wScan_22[0] , \wPDiag_3[30] , \wCall_4[0] , 
        \wColumn_4[0] , \wPDiag_7[11] , \wColumn_10[1] , \wColumn_11[26] , 
        \wColumn_13[2] , \wScan_21[3] , \wColumn_27[23] , \wNDiag_11[3] , 
        \wNDiag_12[10] , \wPDiag_23[9] , \wNDiag_31[21] , \wNDiag_24[15] , 
        \wColumn_7[3] , \wPDiag_7[22] , \wNDiag_12[23] , \wNDiag_24[26] , 
        \wNDiag_12[0] , \wNDiag_31[12] , \wNDiag_6[30] , \wNDiag_6[29] , 
        \wPDiag_8[16] , \wColumn_23[31] , \wColumn_23[28] , \wPDiag_8[25] , 
        \wPDiag_14[12] , \wPDiag_22[17] , \wScan_18[3] , \wPDiag_14[21] , 
        \wNDiag_30[1] , \wPDiag_22[24] , \wColumn_29[1] , \wPDiag_3[29] , 
        \wColumn_28[17] , \wColumn_4[9] , \wPDiag_9[7] , \wNDiag_16[31] , 
        \wNDiag_16[28] , \wColumn_28[24] , \wPDiag_29[31] , \wPDiag_29[28] , 
        \wColumn_31[3] , \wNDiag_28[3] , \wPDiag_7[18] , \wNDiag_8[7] , 
        \wNDiag_9[27] , \wNDiag_9[14] , \wNDiag_12[9] , \wColumn_15[5] , 
        \wColumn_16[6] , \wScan_27[4] , \wPDiag_20[3] , \wNDiag_12[19] , 
        \wPDiag_23[0] , \wNDiag_31[31] , \wNDiag_31[28] , \wColumn_4[13] , 
        \wColumn_10[8] , \wPDiag_10[10] , \wNDiag_17[4] , \wPDiag_26[15] , 
        \wNDiag_2[18] , \wNDiag_14[7] , \wNDiag_19[15] , \wColumn_4[20] , 
        \wPDiag_10[23] , \wPDiag_26[26] , \wNDiag_19[26] , \wPDiag_6[12] , 
        \wNDiag_13[13] , \wNDiag_25[16] , \wColumn_27[19] , \wNDiag_30[22] , 
        \wPDiag_30[9] , \wNDiag_3[21] , \wNDiag_3[12] , \wNDiag_5[2] , 
        \wPDiag_6[21] , \wColumn_18[0] , \wNDiag_6[1] , \wNDiag_13[20] , 
        \wNDiag_30[11] , \wNDiag_25[25] , \wColumn_10[16] , \wScan_29[2] , 
        \wReturn_11[0] , \wColumn_26[13] , \wPDiag_11[30] , \wPDiag_11[29] , 
        \wColumn_5[19] , \wColumn_10[25] , \wColumn_26[20] , \wScan_31[0] , 
        \wNDiag_19[2] , \wScan_1[5] , \wColumn_1[31] , \wColumn_1[28] , 
        \wNDiag_7[10] , \wScan_32[3] , \wScan_16[5] , \wColumn_24[4] , 
        \wNDiag_23[8] , \wPDiag_2[10] , \wNDiag_7[23] , \wPDiag_12[1] , 
        \wCall_13[0] , \wColumn_22[11] , \wColumn_27[7] , \wColumn_14[14] , 
        \wPDiag_15[18] , \wPDiag_11[2] , \wColumn_14[27] , \wColumn_22[22] , 
        \wNDiag_25[6] , \wPDiag_28[11] , \wNDiag_26[5] , \wPDiag_4[2] , 
        \wNDiag_17[11] , \wColumn_21[9] , \wNDiag_21[14] , \wColumn_1[9] , 
        \wPDiag_2[23] , \wNDiag_17[22] , \wNDiag_21[27] , \wPDiag_28[22] , 
        \wNDiag_2[15] , \wColumn_4[4] , \wColumn_7[7] , \wPDiag_7[15] , 
        \wPDiag_7[1] , \wNDiag_12[14] , \wNDiag_24[11] , \wNDiag_31[25] , 
        \wPDiag_7[26] , \wNDiag_12[27] , \wNDiag_12[4] , \wColumn_15[8] , 
        \wNDiag_31[16] , \wNDiag_24[22] , \wNDiag_9[19] , \wNDiag_11[7] , 
        \wColumn_11[11] , \wPDiag_25[3] , \wPDiag_26[0] , \wColumn_27[14] , 
        \wNDiag_2[26] , \wColumn_10[5] , \wColumn_11[22] , \wColumn_13[6] , 
        \wNDiag_19[18] , \wColumn_27[27] , \wNDiag_6[24] , \wNDiag_6[17] , 
        \wNDiag_17[9] , \wScan_22[4] , \wPDiag_26[18] , \wPDiag_8[31] , 
        \wPDiag_8[28] , \wPDiag_22[30] , \wPDiag_22[29] , \wColumn_23[16] , 
        \wColumn_15[13] , \wColumn_15[20] , \wColumn_23[25] , \wColumn_1[25] , 
        \wColumn_1[16] , \wPDiag_1[2] , \wPDiag_3[24] , \wPDiag_3[17] , 
        \wScan_9[0] , \wColumn_28[29] , \wPDiag_29[16] , \wNDiag_16[25] , 
        \wNDiag_16[16] , \wColumn_28[30] , \wPDiag_19[7] , \wNDiag_20[13] , 
        \wNDiag_20[20] , \wPDiag_29[25] , \wPDiag_2[1] , \wScan_4[5] , 
        \wPDiag_9[11] , \wPDiag_9[22] , \wPDiag_15[15] , \wPDiag_23[10] , 
        \wColumn_14[19] , \wNDiag_20[6] , \wNDiag_3[1] , \wNDiag_8[20] , 
        \wNDiag_8[13] , \wReturn_9[0] , \wPDiag_14[2] , \wPDiag_15[26] , 
        \wNDiag_23[5] , \wPDiag_17[1] , \wPDiag_23[23] , \wColumn_24[9] , 
        \wColumn_29[10] , \wScan_13[5] , \wColumn_21[4] , \wNDiag_21[19] , 
        \wCall_16[0] , \wColumn_22[7] , \wNDiag_26[8] , \wColumn_29[23] , 
        \wColumn_9[1] , \wReturn_14[0] , \wNDiag_25[31] , \wNDiag_25[28] , 
        \wPDiag_30[4] , \wPDiag_11[17] , \wPDiag_27[12] , \wColumn_5[27] , 
        \wColumn_5[14] , \wColumn_10[31] , \wColumn_10[28] , \wPDiag_11[24] , 
        \wNDiag_18[12] , \wPDiag_27[21] , \wNDiag_18[21] , \wPDiag_28[6] , 
        \wScan_1[1] , \wScan_2[2] , \wPDiag_2[27] , \wPDiag_2[14] , 
        \wNDiag_17[15] , \wNDiag_21[10] , \wPDiag_7[5] , \wNDiag_25[2] , 
        \wNDiag_26[1] , \wPDiag_28[15] , \wPDiag_17[8] , \wNDiag_17[26] , 
        \wColumn_29[19] , \wNDiag_21[23] , \wPDiag_28[26] , \wPDiag_2[8] , 
        \wPDiag_4[6] , \wNDiag_7[27] , \wNDiag_7[14] , \wColumn_14[10] , 
        \wColumn_27[3] , \wScan_15[2] , \wColumn_22[15] , \wScan_16[1] , 
        \wColumn_24[0] , \wPDiag_9[18] , \wPDiag_11[6] , \wColumn_22[26] , 
        \wColumn_14[23] , \wPDiag_12[5] , \wNDiag_3[16] , \wPDiag_23[19] , 
        \wNDiag_18[31] , \wNDiag_18[28] , \wPDiag_27[31] , \wPDiag_27[28] , 
        \wColumn_10[12] , \wColumn_26[17] , \wCall_1[0] , \wColumn_1[0] , 
        \wNDiag_3[25] , \wNDiag_3[8] , \wColumn_4[17] , \wNDiag_5[6] , 
        \wPDiag_6[16] , \wNDiag_8[30] , \wNDiag_8[29] , \wColumn_10[21] , 
        \wNDiag_19[6] , \wColumn_26[24] , \wScan_31[4] , \wColumn_9[8] , 
        \wNDiag_13[17] , \wNDiag_25[12] , \wNDiag_30[26] , \wPDiag_6[25] , 
        \wNDiag_6[5] , \wNDiag_13[24] , \wNDiag_25[21] , \wNDiag_30[15] , 
        \wNDiag_14[3] , \wColumn_18[4] , \wNDiag_19[11] , \wPDiag_10[14] , 
        \wNDiag_17[0] , \wPDiag_26[11] , \wPDiag_1[18] , \wColumn_2[3] , 
        \wColumn_4[24] , \wColumn_11[18] , \wPDiag_5[30] , \wPDiag_5[29] , 
        \wColumn_6[22] , \wPDiag_8[21] , \wPDiag_8[12] , \wNDiag_8[3] , 
        \wNDiag_9[10] , \wPDiag_10[27] , \wNDiag_19[22] , \wColumn_15[1] , 
        \wPDiag_26[22] , \wPDiag_26[9] , \wScan_27[0] , \wColumn_16[2] , 
        \wScan_24[3] , \wPDiag_9[3] , \wNDiag_9[23] , \wPDiag_23[4] , 
        \wNDiag_24[18] , \wPDiag_20[7] , \wPDiag_14[16] , \wNDiag_20[30] , 
        \wNDiag_20[29] , \wColumn_28[20] , \wColumn_28[13] , \wNDiag_28[7] , 
        \wColumn_31[7] , \wPDiag_22[13] , \wPDiag_14[25] , \wColumn_15[30] , 
        \wColumn_15[29] , \wPDiag_22[20] , \wColumn_29[5] , \wNDiag_30[5] , 
        \wPDiag_18[3] , \wColumn_6[11] , \wPDiag_12[21] , \wPDiag_24[24] , 
        \wPDiag_31[10] , \wScan_8[4] , \wPDiag_12[12] , \wColumn_25[31] , 
        \wColumn_25[28] , \wColumn_18[21] , \wPDiag_24[17] , \wPDiag_31[23] , 
        \wColumn_18[12] , \wColumn_28[8] , \wNDiag_10[31] , \wNDiag_10[28] , 
        \wColumn_12[2] , \wNDiag_31[8] , \wScan_20[3] , \wScan_23[0] , 
        \wColumn_2[20] , \wNDiag_4[18] , \wColumn_11[1] , \wNDiag_14[19] , 
        \wPDiag_24[7] , \wPDiag_27[4] , \wCall_5[0] , \wNDiag_13[0] , 
        \wPDiag_16[23] , \wColumn_6[3] , \wPDiag_20[26] , \wColumn_5[0] , 
        \wNDiag_10[3] , \wNDiag_29[23] , \wPDiag_20[15] , \wColumn_21[19] , 
        \wNDiag_1[23] , \wNDiag_1[6] , \wColumn_2[13] , \wPDiag_16[10] , 
        \wPDiag_22[9] , \wNDiag_2[5] , \wColumn_8[26] , \wNDiag_23[25] , 
        \wNDiag_29[10] , \wColumn_8[15] , \wNDiag_15[20] , \wNDiag_15[13] , 
        \wPDiag_29[2] , \wNDiag_23[16] , \wColumn_3[19] , \wNDiag_5[21] , 
        \wColumn_16[25] , \wColumn_20[20] , \wPDiag_31[0] , \wNDiag_5[12] , 
        \wColumn_8[5] , \wColumn_20[13] , \wColumn_16[16] , \wPDiag_17[30] , 
        \wNDiag_28[30] , \wNDiag_28[29] , \wPDiag_17[29] , \wColumn_19[9] , 
        \wNDiag_7[8] , \wScan_12[1] , \wPDiag_13[18] , \wPDiag_30[29] , 
        \wPDiag_30[30] , \wNDiag_1[10] , \wScan_11[2] , \wColumn_12[27] , 
        \wColumn_20[0] , \wColumn_23[3] , \wColumn_24[22] , \wColumn_31[16] , 
        \wPDiag_16[5] , \wColumn_3[23] , \wPDiag_3[5] , \wPDiag_4[23] , 
        \wPDiag_6[8] , \wColumn_7[31] , \wColumn_7[28] , \wNDiag_11[22] , 
        \wColumn_12[14] , \wPDiag_15[6] , \wColumn_31[25] , \wPDiag_18[27] , 
        \wNDiag_21[2] , \wColumn_24[11] , \wColumn_19[18] , \wNDiag_27[27] , 
        \wNDiag_22[1] , \wPDiag_4[10] , \wScan_5[1] , \wPDiag_18[14] , 
        \wReturn_29[0] , \wNDiag_4[2] , \wScan_6[2] , \wPDiag_13[8] , 
        \wNDiag_27[14] , \wNDiag_11[11] , \wScan_28[2] , \wNDiag_28[20] , 
        \wColumn_3[10] , \wNDiag_7[1] , \wPDiag_17[20] , \wColumn_19[0] , 
        \wPDiag_21[25] , \wNDiag_28[13] , \wPDiag_4[19] , \wNDiag_5[31] , 
        \wNDiag_5[28] , \wColumn_20[30] , \wPDiag_31[9] , \wColumn_20[29] , 
        \wReturn_10[0] , \wNDiag_15[30] , \wNDiag_15[29] , \wPDiag_17[13] , 
        \wNDiag_18[2] , \wPDiag_21[16] , \wScan_30[0] , \wPDiag_10[2] , 
        \wColumn_19[22] , \wNDiag_11[18] , \wPDiag_13[1] , \wScan_0[5] , 
        \wNDiag_1[19] , \wCall_12[0] , \wColumn_26[7] , \wScan_17[5] , 
        \wColumn_25[4] , \wColumn_19[11] , \wNDiag_22[8] , \wPDiag_5[2] , 
        \wPDiag_6[1] , \wPDiag_30[13] , \wPDiag_13[22] , \wPDiag_25[27] , 
        \wColumn_7[21] , \wPDiag_5[20] , \wColumn_7[12] , \wPDiag_13[11] , 
        \wColumn_24[18] , \wPDiag_25[14] , \wNDiag_27[5] , \wPDiag_30[20] , 
        \wColumn_20[9] , \wNDiag_24[6] , \wPDiag_5[13] , \wNDiag_10[21] , 
        \wNDiag_26[24] , \wColumn_28[1] , \wNDiag_10[12] , \wScan_19[3] , 
        \wPDiag_19[24] , \wNDiag_31[1] , \wColumn_18[31] , \wColumn_18[28] , 
        \wNDiag_26[17] , \wColumn_6[18] , \wPDiag_19[17] , \wColumn_13[24] , 
        \wColumn_25[21] , \wNDiag_29[3] , \wColumn_30[15] , \wColumn_30[3] , 
        \wPDiag_1[22] , \wColumn_2[30] , \wColumn_2[29] , \wNDiag_4[22] , 
        \wPDiag_8[7] , \wColumn_25[12] , \wPDiag_12[31] , \wPDiag_12[28] , 
        \wColumn_13[17] , \wColumn_30[26] , \wPDiag_31[19] , \wPDiag_16[19] , 
        \wPDiag_22[0] , \wNDiag_4[11] , \wColumn_14[5] , \wColumn_17[26] , 
        \wColumn_21[23] , \wPDiag_21[3] , \wNDiag_29[19] , \wColumn_5[9] , 
        \wNDiag_13[9] , \wScan_26[4] , \wNDiag_9[7] , \wColumn_9[25] , 
        \wNDiag_14[23] , \wColumn_17[15] , \wColumn_17[6] , \wColumn_21[10] , 
        \wNDiag_22[26] , \wPDiag_1[11] , \wNDiag_15[7] , \wNDiag_1[27] , 
        \wColumn_3[7] , \wPDiag_3[1] , \wPDiag_4[27] , \wColumn_9[16] , 
        \wNDiag_16[4] , \wColumn_11[8] , \wNDiag_14[10] , \wNDiag_22[15] , 
        \wNDiag_11[26] , \wNDiag_22[5] , \wColumn_25[9] , \wNDiag_27[23] , 
        \wNDiag_11[15] , \wPDiag_18[23] , \wNDiag_21[6] , \wNDiag_27[10] , 
        \wPDiag_4[14] , \wScan_5[5] , \wColumn_12[23] , \wPDiag_18[10] , 
        \wCall_17[0] , \wColumn_23[7] , \wColumn_24[26] , \wColumn_31[12] , 
        \wColumn_20[4] , \wNDiag_1[14] , \wReturn_8[0] , \wScan_12[5] , 
        \wPDiag_25[19] , \wColumn_12[10] , \wPDiag_15[2] , \wColumn_24[15] , 
        \wNDiag_27[8] , \wColumn_31[21] , \wNDiag_1[2] , \wNDiag_5[25] , 
        \wPDiag_16[1] , \wNDiag_5[16] , \wReturn_15[0] , \wColumn_16[21] , 
        \wColumn_20[24] , \wPDiag_31[4] , \wColumn_8[22] , \wColumn_8[1] , 
        \wColumn_16[12] , \wPDiag_21[31] , \wPDiag_21[28] , \wNDiag_15[24] , 
        \wColumn_20[17] , \wPDiag_29[6] , \wNDiag_23[21] , \wColumn_2[24] , 
        \wNDiag_2[1] , \wColumn_8[11] , \wColumn_5[4] , \wNDiag_15[17] , 
        \wNDiag_23[12] , \wColumn_17[18] , \wNDiag_10[7] , \wNDiag_29[27] , 
        \wColumn_2[17] , \wColumn_6[7] , \wPDiag_20[22] , \wNDiag_13[4] , 
        \wPDiag_16[27] , \wColumn_14[8] , \wNDiag_29[14] , \wPDiag_16[14] , 
        \wColumn_6[26] , \wScan_8[0] , \wColumn_9[31] , \wColumn_11[5] , 
        \wPDiag_20[11] , \wColumn_12[6] , \wNDiag_16[9] , \wNDiag_22[18] , 
        \wScan_23[4] , \wPDiag_27[0] , \wColumn_9[28] , \wPDiag_24[3] , 
        \wPDiag_12[25] , \wColumn_18[25] , \wColumn_18[16] , \wPDiag_19[30] , 
        \wPDiag_19[29] , \wNDiag_26[30] , \wNDiag_26[29] , \wPDiag_31[14] , 
        \wPDiag_24[20] , \wPDiag_12[16] , \wPDiag_18[7] , \wPDiag_24[13] , 
        \wPDiag_31[27] , \wColumn_13[30] , \wColumn_13[29] , \wColumn_30[18] , 
        \wCall_0[0] , \wPDiag_1[26] , \wColumn_6[15] , \wPDiag_1[15] , 
        \wColumn_9[21] , \wNDiag_22[22] , \wColumn_9[12] , \wNDiag_14[27] , 
        \wNDiag_14[14] , \wPDiag_27[9] , \wNDiag_22[11] , \wNDiag_16[0] , 
        \wColumn_3[3] , \wNDiag_4[26] , \wNDiag_15[3] , \wColumn_17[22] , 
        \wColumn_21[27] , \wPDiag_21[7] , \wNDiag_4[15] , \wNDiag_9[3] , 
        \wColumn_17[11] , \wColumn_17[2] , \wPDiag_20[18] , \wPDiag_22[4] , 
        \wColumn_21[14] , \wScan_25[3] , \wScan_26[0] , \wColumn_14[1] , 
        \wColumn_25[25] , \wColumn_30[7] , \wPDiag_8[3] , \wColumn_13[20] , 
        \wColumn_30[11] , \wColumn_13[13] , \wPDiag_24[30] , \wNDiag_29[7] , 
        \wPDiag_24[29] , \wColumn_30[22] , \wScan_0[1] , \wPDiag_5[24] , 
        \wNDiag_10[25] , \wPDiag_19[20] , \wColumn_25[16] , \wNDiag_31[5] , 
        \wNDiag_26[20] , \wColumn_28[5] , \wPDiag_5[17] , \wPDiag_19[13] , 
        \wNDiag_10[16] , \wNDiag_26[13] , \wColumn_12[19] , \wColumn_31[31] , 
        \wColumn_31[28] , \wScan_3[2] , \wPDiag_5[6] , \wColumn_7[25] , 
        \wPDiag_6[5] , \wPDiag_25[23] , \wPDiag_13[26] , \wPDiag_16[8] , 
        \wPDiag_30[17] , \wPDiag_3[8] , \wColumn_7[16] , \wPDiag_13[15] , 
        \wNDiag_24[2] , \wPDiag_13[5] , \wPDiag_25[10] , \wPDiag_30[24] , 
        \wNDiag_27[1] , \wColumn_19[26] , \wNDiag_27[19] , \wPDiag_10[6] , 
        \wScan_14[2] , \wScan_17[1] , \wPDiag_18[19] , \wColumn_19[15] , 
        \wColumn_25[0] , \wColumn_26[3] , \wScan_0[3] , \wNDiag_2[8] , 
        \wColumn_8[18] , \wNDiag_18[6] , \wScan_30[4] , \wScan_3[0] , 
        \wColumn_3[27] , \wNDiag_7[5] , \wNDiag_23[31] , \wNDiag_23[28] , 
        \wPDiag_17[24] , \wColumn_19[4] , \wPDiag_21[21] , \wColumn_3[14] , 
        \wNDiag_4[6] , \wColumn_8[8] , \wNDiag_28[24] , \wColumn_16[31] , 
        \wColumn_16[28] , \wPDiag_17[17] , \wPDiag_21[12] , \wNDiag_28[17] , 
        \wPDiag_5[4] , \wPDiag_6[7] , \wPDiag_13[24] , \wColumn_7[27] , 
        \wPDiag_25[21] , \wPDiag_30[15] , \wColumn_7[14] , \wColumn_12[31] , 
        \wColumn_12[28] , \wPDiag_13[17] , \wPDiag_15[9] , \wPDiag_25[12] , 
        \wNDiag_27[3] , \wPDiag_30[26] , \wColumn_31[19] , \wNDiag_24[0] , 
        \wPDiag_10[4] , \wPDiag_13[7] , \wColumn_19[24] , \wScan_14[0] , 
        \wPDiag_1[24] , \wNDiag_1[9] , \wScan_17[3] , \wPDiag_18[31] , 
        \wPDiag_18[28] , \wColumn_25[2] , \wColumn_26[1] , \wNDiag_27[31] , 
        \wNDiag_27[28] , \wColumn_19[17] , \wNDiag_23[19] , \wColumn_3[25] , 
        \wNDiag_4[4] , \wColumn_8[30] , \wColumn_8[29] , \wNDiag_18[4] , 
        \wColumn_16[19] , \wScan_28[4] , \wColumn_3[16] , \wNDiag_7[7] , 
        \wPDiag_17[26] , \wColumn_19[6] , \wPDiag_21[23] , \wNDiag_28[26] , 
        \wColumn_9[23] , \wNDiag_14[25] , \wPDiag_17[15] , \wNDiag_28[15] , 
        \wPDiag_21[10] , \wPDiag_24[8] , \wNDiag_22[20] , \wPDiag_1[17] , 
        \wColumn_3[1] , \wNDiag_15[1] , \wNDiag_4[24] , \wColumn_9[10] , 
        \wNDiag_16[2] , \wNDiag_22[13] , \wNDiag_14[16] , \wNDiag_4[17] , 
        \wColumn_14[3] , \wColumn_17[20] , \wColumn_21[25] , \wPDiag_21[5] , 
        \wPDiag_22[6] , \wNDiag_9[1] , \wPDiag_20[30] , \wPDiag_20[29] , 
        \wScan_26[2] , \wColumn_13[22] , \wColumn_17[13] , \wScan_25[1] , 
        \wColumn_17[0] , \wColumn_21[16] , \wNDiag_29[5] , \wColumn_30[13] , 
        \wPDiag_8[1] , \wPDiag_24[18] , \wColumn_25[27] , \wColumn_30[5] , 
        \wColumn_25[14] , \wColumn_2[26] , \wReturn_3[0] , \wPDiag_5[26] , 
        \wColumn_13[11] , \wColumn_30[20] , \wNDiag_10[27] , \wNDiag_26[22] , 
        \wColumn_28[7] , \wNDiag_10[14] , \wScan_19[5] , \wPDiag_19[22] , 
        \wNDiag_31[7] , \wPDiag_5[15] , \wNDiag_26[11] , \wColumn_6[5] , 
        \wNDiag_13[6] , \wPDiag_16[25] , \wPDiag_19[11] , \wNDiag_10[5] , 
        \wPDiag_20[20] , \wNDiag_29[25] , \wColumn_2[15] , \wColumn_5[6] , 
        \wNDiag_9[8] , \wPDiag_16[16] , \wColumn_17[9] , \wPDiag_20[13] , 
        \wColumn_17[30] , \wColumn_17[29] , \wNDiag_29[16] , \wColumn_3[8] , 
        \wColumn_12[4] , \wNDiag_15[8] , \wScan_20[5] , \wScan_8[2] , 
        \wColumn_9[19] , \wColumn_11[7] , \wCall_25[0] , \wColumn_18[27] , 
        \wNDiag_22[30] , \wNDiag_22[29] , \wPDiag_24[1] , \wNDiag_26[18] , 
        \wPDiag_27[2] , \wReturn_27[0] , \wPDiag_8[8] , \wColumn_13[18] , 
        \wColumn_18[14] , \wPDiag_19[18] , \wColumn_30[29] , \wColumn_30[30] , 
        \wColumn_6[24] , \wPDiag_18[5] , \wColumn_6[17] , \wPDiag_12[27] , 
        \wPDiag_24[22] , \wPDiag_31[16] , \wPDiag_12[14] , \wPDiag_31[25] , 
        \wNDiag_21[4] , \wPDiag_24[11] , \wNDiag_1[25] , \wPDiag_3[3] , 
        \wPDiag_4[25] , \wNDiag_11[24] , \wPDiag_18[21] , \wColumn_26[8] , 
        \wNDiag_27[21] , \wPDiag_4[16] , \wPDiag_18[12] , \wNDiag_22[7] , 
        \wScan_6[4] , \wNDiag_11[17] , \wNDiag_27[12] , \wColumn_20[6] , 
        \wNDiag_1[16] , \wScan_11[4] , \wColumn_12[21] , \wColumn_23[5] , 
        \wColumn_24[24] , \wNDiag_24[9] , \wColumn_31[10] , \wPDiag_16[3] , 
        \wNDiag_1[0] , \wNDiag_2[3] , \wNDiag_5[27] , \wColumn_12[12] , 
        \wPDiag_25[31] , \wPDiag_25[28] , \wPDiag_15[0] , \wColumn_16[23] , 
        \wColumn_24[17] , \wColumn_31[23] , \wColumn_20[26] , \wPDiag_31[6] , 
        \wNDiag_5[14] , \wColumn_8[3] , \wColumn_16[10] , \wColumn_20[15] , 
        \wPDiag_21[19] , \wColumn_8[20] , \wNDiag_15[26] , \wNDiag_23[23] , 
        \wNDiag_15[15] , \wPDiag_29[4] , \wColumn_8[13] , \wNDiag_23[10] , 
        \wPDiag_5[22] , \wNDiag_10[23] , \wScan_19[1] , \wPDiag_19[26] , 
        \wNDiag_31[3] , \wColumn_18[19] , \wNDiag_26[26] , \wColumn_28[3] , 
        \wPDiag_5[11] , \wPDiag_19[15] , \wNDiag_10[10] , \wNDiag_26[15] , 
        \wPDiag_12[19] , \wPDiag_31[31] , \wColumn_30[1] , \wPDiag_31[28] , 
        \wColumn_6[30] , \wColumn_6[29] , \wColumn_13[26] , \wColumn_25[23] , 
        \wNDiag_29[1] , \wPDiag_18[8] , \wReturn_22[0] , \wColumn_30[17] , 
        \wColumn_13[15] , \wColumn_25[10] , \wColumn_30[24] , \wPDiag_1[20] , 
        \wColumn_2[18] , \wPDiag_8[5] , \wNDiag_4[20] , \wColumn_17[24] , 
        \wColumn_21[21] , \wPDiag_21[1] , \wPDiag_22[2] , \wNDiag_4[13] , 
        \wColumn_6[8] , \wNDiag_9[5] , \wNDiag_10[8] , \wColumn_17[17] , 
        \wColumn_21[12] , \wColumn_17[4] , \wNDiag_29[31] , \wScan_25[5] , 
        \wNDiag_29[28] , \wPDiag_16[31] , \wPDiag_16[28] , \wColumn_14[7] , 
        \wCall_20[0] , \wPDiag_1[13] , \wColumn_3[5] , \wColumn_9[27] , 
        \wColumn_9[14] , \wNDiag_14[21] , \wNDiag_22[24] , \wNDiag_14[12] , 
        \wNDiag_16[6] , \wNDiag_22[17] , \wColumn_3[21] , \wNDiag_5[19] , 
        \wColumn_12[9] , \wNDiag_15[5] , \wNDiag_7[3] , \wPDiag_17[22] , 
        \wColumn_19[2] , \wPDiag_21[27] , \wNDiag_28[22] , \wColumn_3[12] , 
        \wNDiag_4[0] , \wColumn_20[18] , \wScan_28[0] , \wPDiag_17[11] , 
        \wPDiag_21[14] , \wNDiag_28[11] , \wPDiag_4[31] , \wPDiag_10[0] , 
        \wPDiag_13[3] , \wNDiag_15[18] , \wNDiag_18[0] , \wScan_30[2] , 
        \wPDiag_29[9] , \wColumn_19[20] , \wColumn_19[13] , \wPDiag_4[28] , 
        \wNDiag_11[30] , \wNDiag_11[29] , \wColumn_25[6] , \wColumn_26[5] , 
        \wPDiag_1[30] , \wPDiag_1[29] , \wNDiag_1[31] , \wNDiag_1[28] , 
        \wScan_3[4] , \wPDiag_5[0] , \wScan_14[4] , \wNDiag_21[9] , 
        \wPDiag_6[3] , \wColumn_7[23] , \wPDiag_13[20] , \wPDiag_25[25] , 
        \wPDiag_30[11] , \wColumn_7[10] , \wColumn_23[8] , \wNDiag_24[4] , 
        \wColumn_24[30] , \wColumn_24[29] , \wNDiag_1[21] , \wNDiag_1[4] , 
        \wColumn_8[24] , \wPDiag_13[13] , \wPDiag_30[22] , \wNDiag_15[22] , 
        \wPDiag_25[16] , \wNDiag_27[7] , \wPDiag_29[0] , \wNDiag_23[27] , 
        \wNDiag_2[7] , \wNDiag_18[9] , \wNDiag_23[14] , \wColumn_3[31] , 
        \wNDiag_5[23] , \wColumn_8[17] , \wNDiag_15[11] , \wPDiag_17[18] , 
        \wNDiag_5[10] , \wColumn_16[27] , \wColumn_20[22] , \wPDiag_31[2] , 
        \wNDiag_28[18] , \wColumn_3[28] , \wNDiag_4[9] , \wColumn_8[7] , 
        \wColumn_7[19] , \wScan_11[0] , \wColumn_16[14] , \wColumn_20[11] , 
        \wColumn_12[25] , \wColumn_31[14] , \wColumn_23[1] , \wColumn_24[20] , 
        \wNDiag_1[12] , \wPDiag_5[9] , \wScan_12[3] , \wColumn_20[2] , 
        \wColumn_12[16] , \wColumn_24[13] , \wReturn_31[0] , \wColumn_31[27] , 
        \wPDiag_15[4] , \wPDiag_13[30] , \wPDiag_13[29] , \wPDiag_30[18] , 
        \wPDiag_3[7] , \wPDiag_4[21] , \wPDiag_16[7] , \wNDiag_22[3] , 
        \wScan_6[0] , \wNDiag_11[20] , \wNDiag_27[25] , \wNDiag_11[13] , 
        \wPDiag_18[25] , \wNDiag_21[0] , \wColumn_19[30] , \wNDiag_27[16] , 
        \wPDiag_4[12] , \wColumn_19[29] , \wScan_5[3] , \wPDiag_5[18] , 
        \wReturn_6[0] , \wPDiag_10[9] , \wPDiag_18[16] , \wColumn_6[20] , 
        \wPDiag_12[23] , \wPDiag_24[26] , \wPDiag_31[12] , \wColumn_6[13] , 
        \wPDiag_12[10] , \wPDiag_18[1] , \wCall_19[0] , \wPDiag_24[15] , 
        \wColumn_25[19] , \wNDiag_29[8] , \wColumn_30[8] , \wPDiag_31[21] , 
        \wColumn_18[23] , \wNDiag_10[19] , \wColumn_11[3] , \wColumn_18[10] , 
        \wColumn_12[0] , \wScan_20[1] , \wScan_23[2] , \wColumn_2[22] , 
        \wColumn_5[2] , \wNDiag_14[31] , \wNDiag_14[28] , \wPDiag_27[6] , 
        \wPDiag_24[5] , \wColumn_2[11] , \wColumn_6[1] , \wNDiag_10[1] , 
        \wNDiag_29[21] , \wNDiag_13[2] , \wPDiag_16[21] , \wPDiag_20[24] , 
        \wNDiag_4[30] , \wColumn_21[31] , \wColumn_21[28] , \wNDiag_29[12] , 
        \wPDiag_21[8] , \wNDiag_4[29] , \wPDiag_16[12] , \wPDiag_20[17] ;
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_12 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_13[5] , \wScan_13[4] , \wScan_13[3] , 
        \wScan_13[2] , \wScan_13[1] , \wScan_13[0] }), .ScanOut({\wScan_12[5] , 
        \wScan_12[4] , \wScan_12[3] , \wScan_12[2] , \wScan_12[1] , 
        \wScan_12[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_12[0] ), .ReturnIn(\wReturn_13[0] ), 
        .ColIn({\wColumn_12[31] , \wColumn_12[30] , \wColumn_12[29] , 
        \wColumn_12[28] , \wColumn_12[27] , \wColumn_12[26] , \wColumn_12[25] , 
        \wColumn_12[24] , \wColumn_12[23] , \wColumn_12[22] , \wColumn_12[21] , 
        \wColumn_12[20] , \wColumn_12[19] , \wColumn_12[18] , \wColumn_12[17] , 
        \wColumn_12[16] , \wColumn_12[15] , \wColumn_12[14] , \wColumn_12[13] , 
        \wColumn_12[12] , \wColumn_12[11] , \wColumn_12[10] , \wColumn_12[9] , 
        \wColumn_12[8] , \wColumn_12[7] , \wColumn_12[6] , \wColumn_12[5] , 
        \wColumn_12[4] , \wColumn_12[3] , \wColumn_12[2] , \wColumn_12[1] , 
        \wColumn_12[0] }), .PDiagIn({\wPDiag_12[31] , \wPDiag_12[30] , 
        \wPDiag_12[29] , \wPDiag_12[28] , \wPDiag_12[27] , \wPDiag_12[26] , 
        \wPDiag_12[25] , \wPDiag_12[24] , \wPDiag_12[23] , \wPDiag_12[22] , 
        \wPDiag_12[21] , \wPDiag_12[20] , \wPDiag_12[19] , \wPDiag_12[18] , 
        \wPDiag_12[17] , \wPDiag_12[16] , \wPDiag_12[15] , \wPDiag_12[14] , 
        \wPDiag_12[13] , \wPDiag_12[12] , \wPDiag_12[11] , \wPDiag_12[10] , 
        \wPDiag_12[9] , \wPDiag_12[8] , \wPDiag_12[7] , \wPDiag_12[6] , 
        \wPDiag_12[5] , \wPDiag_12[4] , \wPDiag_12[3] , \wPDiag_12[2] , 
        \wPDiag_12[1] , \wPDiag_12[0] }), .NDiagIn({\wNDiag_12[31] , 
        \wNDiag_12[30] , \wNDiag_12[29] , \wNDiag_12[28] , \wNDiag_12[27] , 
        \wNDiag_12[26] , \wNDiag_12[25] , \wNDiag_12[24] , \wNDiag_12[23] , 
        \wNDiag_12[22] , \wNDiag_12[21] , \wNDiag_12[20] , \wNDiag_12[19] , 
        \wNDiag_12[18] , \wNDiag_12[17] , \wNDiag_12[16] , \wNDiag_12[15] , 
        \wNDiag_12[14] , \wNDiag_12[13] , \wNDiag_12[12] , \wNDiag_12[11] , 
        \wNDiag_12[10] , \wNDiag_12[9] , \wNDiag_12[8] , \wNDiag_12[7] , 
        \wNDiag_12[6] , \wNDiag_12[5] , \wNDiag_12[4] , \wNDiag_12[3] , 
        \wNDiag_12[2] , \wNDiag_12[1] , \wNDiag_12[0] }), .CallOut(
        \wCall_13[0] ), .ReturnOut(\wReturn_12[0] ), .ColOut({\wColumn_13[31] , 
        \wColumn_13[30] , \wColumn_13[29] , \wColumn_13[28] , \wColumn_13[27] , 
        \wColumn_13[26] , \wColumn_13[25] , \wColumn_13[24] , \wColumn_13[23] , 
        \wColumn_13[22] , \wColumn_13[21] , \wColumn_13[20] , \wColumn_13[19] , 
        \wColumn_13[18] , \wColumn_13[17] , \wColumn_13[16] , \wColumn_13[15] , 
        \wColumn_13[14] , \wColumn_13[13] , \wColumn_13[12] , \wColumn_13[11] , 
        \wColumn_13[10] , \wColumn_13[9] , \wColumn_13[8] , \wColumn_13[7] , 
        \wColumn_13[6] , \wColumn_13[5] , \wColumn_13[4] , \wColumn_13[3] , 
        \wColumn_13[2] , \wColumn_13[1] , \wColumn_13[0] }), .PDiagOut({
        \wPDiag_13[31] , \wPDiag_13[30] , \wPDiag_13[29] , \wPDiag_13[28] , 
        \wPDiag_13[27] , \wPDiag_13[26] , \wPDiag_13[25] , \wPDiag_13[24] , 
        \wPDiag_13[23] , \wPDiag_13[22] , \wPDiag_13[21] , \wPDiag_13[20] , 
        \wPDiag_13[19] , \wPDiag_13[18] , \wPDiag_13[17] , \wPDiag_13[16] , 
        \wPDiag_13[15] , \wPDiag_13[14] , \wPDiag_13[13] , \wPDiag_13[12] , 
        \wPDiag_13[11] , \wPDiag_13[10] , \wPDiag_13[9] , \wPDiag_13[8] , 
        \wPDiag_13[7] , \wPDiag_13[6] , \wPDiag_13[5] , \wPDiag_13[4] , 
        \wPDiag_13[3] , \wPDiag_13[2] , \wPDiag_13[1] , \wPDiag_13[0] }), 
        .NDiagOut({\wNDiag_13[31] , \wNDiag_13[30] , \wNDiag_13[29] , 
        \wNDiag_13[28] , \wNDiag_13[27] , \wNDiag_13[26] , \wNDiag_13[25] , 
        \wNDiag_13[24] , \wNDiag_13[23] , \wNDiag_13[22] , \wNDiag_13[21] , 
        \wNDiag_13[20] , \wNDiag_13[19] , \wNDiag_13[18] , \wNDiag_13[17] , 
        \wNDiag_13[16] , \wNDiag_13[15] , \wNDiag_13[14] , \wNDiag_13[13] , 
        \wNDiag_13[12] , \wNDiag_13[11] , \wNDiag_13[10] , \wNDiag_13[9] , 
        \wNDiag_13[8] , \wNDiag_13[7] , \wNDiag_13[6] , \wNDiag_13[5] , 
        \wNDiag_13[4] , \wNDiag_13[3] , \wNDiag_13[2] , \wNDiag_13[1] , 
        \wNDiag_13[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_0 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_1[5] , \wScan_1[4] , \wScan_1[3] , 
        \wScan_1[2] , \wScan_1[1] , \wScan_1[0] }), .ScanOut({\wScan_0[5] , 
        \wScan_0[4] , \wScan_0[3] , \wScan_0[2] , \wScan_0[1] , \wScan_0[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_0[0] ), .ReturnIn(\wReturn_1[0] ), .ColIn({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .PDiagIn({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .NDiagIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallOut(\wCall_1[0] ), .ReturnOut(\wReturn_0[0] ), 
        .ColOut({\wColumn_1[31] , \wColumn_1[30] , \wColumn_1[29] , 
        \wColumn_1[28] , \wColumn_1[27] , \wColumn_1[26] , \wColumn_1[25] , 
        \wColumn_1[24] , \wColumn_1[23] , \wColumn_1[22] , \wColumn_1[21] , 
        \wColumn_1[20] , \wColumn_1[19] , \wColumn_1[18] , \wColumn_1[17] , 
        \wColumn_1[16] , \wColumn_1[15] , \wColumn_1[14] , \wColumn_1[13] , 
        \wColumn_1[12] , \wColumn_1[11] , \wColumn_1[10] , \wColumn_1[9] , 
        \wColumn_1[8] , \wColumn_1[7] , \wColumn_1[6] , \wColumn_1[5] , 
        \wColumn_1[4] , \wColumn_1[3] , \wColumn_1[2] , \wColumn_1[1] , 
        \wColumn_1[0] }), .PDiagOut({\wPDiag_1[31] , \wPDiag_1[30] , 
        \wPDiag_1[29] , \wPDiag_1[28] , \wPDiag_1[27] , \wPDiag_1[26] , 
        \wPDiag_1[25] , \wPDiag_1[24] , \wPDiag_1[23] , \wPDiag_1[22] , 
        \wPDiag_1[21] , \wPDiag_1[20] , \wPDiag_1[19] , \wPDiag_1[18] , 
        \wPDiag_1[17] , \wPDiag_1[16] , \wPDiag_1[15] , \wPDiag_1[14] , 
        \wPDiag_1[13] , \wPDiag_1[12] , \wPDiag_1[11] , \wPDiag_1[10] , 
        \wPDiag_1[9] , \wPDiag_1[8] , \wPDiag_1[7] , \wPDiag_1[6] , 
        \wPDiag_1[5] , \wPDiag_1[4] , \wPDiag_1[3] , \wPDiag_1[2] , 
        \wPDiag_1[1] , \wPDiag_1[0] }), .NDiagOut({\wNDiag_1[31] , 
        \wNDiag_1[30] , \wNDiag_1[29] , \wNDiag_1[28] , \wNDiag_1[27] , 
        \wNDiag_1[26] , \wNDiag_1[25] , \wNDiag_1[24] , \wNDiag_1[23] , 
        \wNDiag_1[22] , \wNDiag_1[21] , \wNDiag_1[20] , \wNDiag_1[19] , 
        \wNDiag_1[18] , \wNDiag_1[17] , \wNDiag_1[16] , \wNDiag_1[15] , 
        \wNDiag_1[14] , \wNDiag_1[13] , \wNDiag_1[12] , \wNDiag_1[11] , 
        \wNDiag_1[10] , \wNDiag_1[9] , \wNDiag_1[8] , \wNDiag_1[7] , 
        \wNDiag_1[6] , \wNDiag_1[5] , \wNDiag_1[4] , \wNDiag_1[3] , 
        \wNDiag_1[2] , \wNDiag_1[1] , \wNDiag_1[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_2 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_3[5] , \wScan_3[4] , \wScan_3[3] , 
        \wScan_3[2] , \wScan_3[1] , \wScan_3[0] }), .ScanOut({\wScan_2[5] , 
        \wScan_2[4] , \wScan_2[3] , \wScan_2[2] , \wScan_2[1] , \wScan_2[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_2[0] ), .ReturnIn(\wReturn_3[0] ), .ColIn({
        \wColumn_2[31] , \wColumn_2[30] , \wColumn_2[29] , \wColumn_2[28] , 
        \wColumn_2[27] , \wColumn_2[26] , \wColumn_2[25] , \wColumn_2[24] , 
        \wColumn_2[23] , \wColumn_2[22] , \wColumn_2[21] , \wColumn_2[20] , 
        \wColumn_2[19] , \wColumn_2[18] , \wColumn_2[17] , \wColumn_2[16] , 
        \wColumn_2[15] , \wColumn_2[14] , \wColumn_2[13] , \wColumn_2[12] , 
        \wColumn_2[11] , \wColumn_2[10] , \wColumn_2[9] , \wColumn_2[8] , 
        \wColumn_2[7] , \wColumn_2[6] , \wColumn_2[5] , \wColumn_2[4] , 
        \wColumn_2[3] , \wColumn_2[2] , \wColumn_2[1] , \wColumn_2[0] }), 
        .PDiagIn({\wPDiag_2[31] , \wPDiag_2[30] , \wPDiag_2[29] , 
        \wPDiag_2[28] , \wPDiag_2[27] , \wPDiag_2[26] , \wPDiag_2[25] , 
        \wPDiag_2[24] , \wPDiag_2[23] , \wPDiag_2[22] , \wPDiag_2[21] , 
        \wPDiag_2[20] , \wPDiag_2[19] , \wPDiag_2[18] , \wPDiag_2[17] , 
        \wPDiag_2[16] , \wPDiag_2[15] , \wPDiag_2[14] , \wPDiag_2[13] , 
        \wPDiag_2[12] , \wPDiag_2[11] , \wPDiag_2[10] , \wPDiag_2[9] , 
        \wPDiag_2[8] , \wPDiag_2[7] , \wPDiag_2[6] , \wPDiag_2[5] , 
        \wPDiag_2[4] , \wPDiag_2[3] , \wPDiag_2[2] , \wPDiag_2[1] , 
        \wPDiag_2[0] }), .NDiagIn({\wNDiag_2[31] , \wNDiag_2[30] , 
        \wNDiag_2[29] , \wNDiag_2[28] , \wNDiag_2[27] , \wNDiag_2[26] , 
        \wNDiag_2[25] , \wNDiag_2[24] , \wNDiag_2[23] , \wNDiag_2[22] , 
        \wNDiag_2[21] , \wNDiag_2[20] , \wNDiag_2[19] , \wNDiag_2[18] , 
        \wNDiag_2[17] , \wNDiag_2[16] , \wNDiag_2[15] , \wNDiag_2[14] , 
        \wNDiag_2[13] , \wNDiag_2[12] , \wNDiag_2[11] , \wNDiag_2[10] , 
        \wNDiag_2[9] , \wNDiag_2[8] , \wNDiag_2[7] , \wNDiag_2[6] , 
        \wNDiag_2[5] , \wNDiag_2[4] , \wNDiag_2[3] , \wNDiag_2[2] , 
        \wNDiag_2[1] , \wNDiag_2[0] }), .CallOut(\wCall_3[0] ), .ReturnOut(
        \wReturn_2[0] ), .ColOut({\wColumn_3[31] , \wColumn_3[30] , 
        \wColumn_3[29] , \wColumn_3[28] , \wColumn_3[27] , \wColumn_3[26] , 
        \wColumn_3[25] , \wColumn_3[24] , \wColumn_3[23] , \wColumn_3[22] , 
        \wColumn_3[21] , \wColumn_3[20] , \wColumn_3[19] , \wColumn_3[18] , 
        \wColumn_3[17] , \wColumn_3[16] , \wColumn_3[15] , \wColumn_3[14] , 
        \wColumn_3[13] , \wColumn_3[12] , \wColumn_3[11] , \wColumn_3[10] , 
        \wColumn_3[9] , \wColumn_3[8] , \wColumn_3[7] , \wColumn_3[6] , 
        \wColumn_3[5] , \wColumn_3[4] , \wColumn_3[3] , \wColumn_3[2] , 
        \wColumn_3[1] , \wColumn_3[0] }), .PDiagOut({\wPDiag_3[31] , 
        \wPDiag_3[30] , \wPDiag_3[29] , \wPDiag_3[28] , \wPDiag_3[27] , 
        \wPDiag_3[26] , \wPDiag_3[25] , \wPDiag_3[24] , \wPDiag_3[23] , 
        \wPDiag_3[22] , \wPDiag_3[21] , \wPDiag_3[20] , \wPDiag_3[19] , 
        \wPDiag_3[18] , \wPDiag_3[17] , \wPDiag_3[16] , \wPDiag_3[15] , 
        \wPDiag_3[14] , \wPDiag_3[13] , \wPDiag_3[12] , \wPDiag_3[11] , 
        \wPDiag_3[10] , \wPDiag_3[9] , \wPDiag_3[8] , \wPDiag_3[7] , 
        \wPDiag_3[6] , \wPDiag_3[5] , \wPDiag_3[4] , \wPDiag_3[3] , 
        \wPDiag_3[2] , \wPDiag_3[1] , \wPDiag_3[0] }), .NDiagOut({
        \wNDiag_3[31] , \wNDiag_3[30] , \wNDiag_3[29] , \wNDiag_3[28] , 
        \wNDiag_3[27] , \wNDiag_3[26] , \wNDiag_3[25] , \wNDiag_3[24] , 
        \wNDiag_3[23] , \wNDiag_3[22] , \wNDiag_3[21] , \wNDiag_3[20] , 
        \wNDiag_3[19] , \wNDiag_3[18] , \wNDiag_3[17] , \wNDiag_3[16] , 
        \wNDiag_3[15] , \wNDiag_3[14] , \wNDiag_3[13] , \wNDiag_3[12] , 
        \wNDiag_3[11] , \wNDiag_3[10] , \wNDiag_3[9] , \wNDiag_3[8] , 
        \wNDiag_3[7] , \wNDiag_3[6] , \wNDiag_3[5] , \wNDiag_3[4] , 
        \wNDiag_3[3] , \wNDiag_3[2] , \wNDiag_3[1] , \wNDiag_3[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_3 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_4[5] , \wScan_4[4] , \wScan_4[3] , 
        \wScan_4[2] , \wScan_4[1] , \wScan_4[0] }), .ScanOut({\wScan_3[5] , 
        \wScan_3[4] , \wScan_3[3] , \wScan_3[2] , \wScan_3[1] , \wScan_3[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_3[0] ), .ReturnIn(\wReturn_4[0] ), .ColIn({
        \wColumn_3[31] , \wColumn_3[30] , \wColumn_3[29] , \wColumn_3[28] , 
        \wColumn_3[27] , \wColumn_3[26] , \wColumn_3[25] , \wColumn_3[24] , 
        \wColumn_3[23] , \wColumn_3[22] , \wColumn_3[21] , \wColumn_3[20] , 
        \wColumn_3[19] , \wColumn_3[18] , \wColumn_3[17] , \wColumn_3[16] , 
        \wColumn_3[15] , \wColumn_3[14] , \wColumn_3[13] , \wColumn_3[12] , 
        \wColumn_3[11] , \wColumn_3[10] , \wColumn_3[9] , \wColumn_3[8] , 
        \wColumn_3[7] , \wColumn_3[6] , \wColumn_3[5] , \wColumn_3[4] , 
        \wColumn_3[3] , \wColumn_3[2] , \wColumn_3[1] , \wColumn_3[0] }), 
        .PDiagIn({\wPDiag_3[31] , \wPDiag_3[30] , \wPDiag_3[29] , 
        \wPDiag_3[28] , \wPDiag_3[27] , \wPDiag_3[26] , \wPDiag_3[25] , 
        \wPDiag_3[24] , \wPDiag_3[23] , \wPDiag_3[22] , \wPDiag_3[21] , 
        \wPDiag_3[20] , \wPDiag_3[19] , \wPDiag_3[18] , \wPDiag_3[17] , 
        \wPDiag_3[16] , \wPDiag_3[15] , \wPDiag_3[14] , \wPDiag_3[13] , 
        \wPDiag_3[12] , \wPDiag_3[11] , \wPDiag_3[10] , \wPDiag_3[9] , 
        \wPDiag_3[8] , \wPDiag_3[7] , \wPDiag_3[6] , \wPDiag_3[5] , 
        \wPDiag_3[4] , \wPDiag_3[3] , \wPDiag_3[2] , \wPDiag_3[1] , 
        \wPDiag_3[0] }), .NDiagIn({\wNDiag_3[31] , \wNDiag_3[30] , 
        \wNDiag_3[29] , \wNDiag_3[28] , \wNDiag_3[27] , \wNDiag_3[26] , 
        \wNDiag_3[25] , \wNDiag_3[24] , \wNDiag_3[23] , \wNDiag_3[22] , 
        \wNDiag_3[21] , \wNDiag_3[20] , \wNDiag_3[19] , \wNDiag_3[18] , 
        \wNDiag_3[17] , \wNDiag_3[16] , \wNDiag_3[15] , \wNDiag_3[14] , 
        \wNDiag_3[13] , \wNDiag_3[12] , \wNDiag_3[11] , \wNDiag_3[10] , 
        \wNDiag_3[9] , \wNDiag_3[8] , \wNDiag_3[7] , \wNDiag_3[6] , 
        \wNDiag_3[5] , \wNDiag_3[4] , \wNDiag_3[3] , \wNDiag_3[2] , 
        \wNDiag_3[1] , \wNDiag_3[0] }), .CallOut(\wCall_4[0] ), .ReturnOut(
        \wReturn_3[0] ), .ColOut({\wColumn_4[31] , \wColumn_4[30] , 
        \wColumn_4[29] , \wColumn_4[28] , \wColumn_4[27] , \wColumn_4[26] , 
        \wColumn_4[25] , \wColumn_4[24] , \wColumn_4[23] , \wColumn_4[22] , 
        \wColumn_4[21] , \wColumn_4[20] , \wColumn_4[19] , \wColumn_4[18] , 
        \wColumn_4[17] , \wColumn_4[16] , \wColumn_4[15] , \wColumn_4[14] , 
        \wColumn_4[13] , \wColumn_4[12] , \wColumn_4[11] , \wColumn_4[10] , 
        \wColumn_4[9] , \wColumn_4[8] , \wColumn_4[7] , \wColumn_4[6] , 
        \wColumn_4[5] , \wColumn_4[4] , \wColumn_4[3] , \wColumn_4[2] , 
        \wColumn_4[1] , \wColumn_4[0] }), .PDiagOut({\wPDiag_4[31] , 
        \wPDiag_4[30] , \wPDiag_4[29] , \wPDiag_4[28] , \wPDiag_4[27] , 
        \wPDiag_4[26] , \wPDiag_4[25] , \wPDiag_4[24] , \wPDiag_4[23] , 
        \wPDiag_4[22] , \wPDiag_4[21] , \wPDiag_4[20] , \wPDiag_4[19] , 
        \wPDiag_4[18] , \wPDiag_4[17] , \wPDiag_4[16] , \wPDiag_4[15] , 
        \wPDiag_4[14] , \wPDiag_4[13] , \wPDiag_4[12] , \wPDiag_4[11] , 
        \wPDiag_4[10] , \wPDiag_4[9] , \wPDiag_4[8] , \wPDiag_4[7] , 
        \wPDiag_4[6] , \wPDiag_4[5] , \wPDiag_4[4] , \wPDiag_4[3] , 
        \wPDiag_4[2] , \wPDiag_4[1] , \wPDiag_4[0] }), .NDiagOut({
        \wNDiag_4[31] , \wNDiag_4[30] , \wNDiag_4[29] , \wNDiag_4[28] , 
        \wNDiag_4[27] , \wNDiag_4[26] , \wNDiag_4[25] , \wNDiag_4[24] , 
        \wNDiag_4[23] , \wNDiag_4[22] , \wNDiag_4[21] , \wNDiag_4[20] , 
        \wNDiag_4[19] , \wNDiag_4[18] , \wNDiag_4[17] , \wNDiag_4[16] , 
        \wNDiag_4[15] , \wNDiag_4[14] , \wNDiag_4[13] , \wNDiag_4[12] , 
        \wNDiag_4[11] , \wNDiag_4[10] , \wNDiag_4[9] , \wNDiag_4[8] , 
        \wNDiag_4[7] , \wNDiag_4[6] , \wNDiag_4[5] , \wNDiag_4[4] , 
        \wNDiag_4[3] , \wNDiag_4[2] , \wNDiag_4[1] , \wNDiag_4[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_27 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_28[5] , \wScan_28[4] , \wScan_28[3] , 
        \wScan_28[2] , \wScan_28[1] , \wScan_28[0] }), .ScanOut({\wScan_27[5] , 
        \wScan_27[4] , \wScan_27[3] , \wScan_27[2] , \wScan_27[1] , 
        \wScan_27[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_27[0] ), .ReturnIn(\wReturn_28[0] ), 
        .ColIn({\wColumn_27[31] , \wColumn_27[30] , \wColumn_27[29] , 
        \wColumn_27[28] , \wColumn_27[27] , \wColumn_27[26] , \wColumn_27[25] , 
        \wColumn_27[24] , \wColumn_27[23] , \wColumn_27[22] , \wColumn_27[21] , 
        \wColumn_27[20] , \wColumn_27[19] , \wColumn_27[18] , \wColumn_27[17] , 
        \wColumn_27[16] , \wColumn_27[15] , \wColumn_27[14] , \wColumn_27[13] , 
        \wColumn_27[12] , \wColumn_27[11] , \wColumn_27[10] , \wColumn_27[9] , 
        \wColumn_27[8] , \wColumn_27[7] , \wColumn_27[6] , \wColumn_27[5] , 
        \wColumn_27[4] , \wColumn_27[3] , \wColumn_27[2] , \wColumn_27[1] , 
        \wColumn_27[0] }), .PDiagIn({\wPDiag_27[31] , \wPDiag_27[30] , 
        \wPDiag_27[29] , \wPDiag_27[28] , \wPDiag_27[27] , \wPDiag_27[26] , 
        \wPDiag_27[25] , \wPDiag_27[24] , \wPDiag_27[23] , \wPDiag_27[22] , 
        \wPDiag_27[21] , \wPDiag_27[20] , \wPDiag_27[19] , \wPDiag_27[18] , 
        \wPDiag_27[17] , \wPDiag_27[16] , \wPDiag_27[15] , \wPDiag_27[14] , 
        \wPDiag_27[13] , \wPDiag_27[12] , \wPDiag_27[11] , \wPDiag_27[10] , 
        \wPDiag_27[9] , \wPDiag_27[8] , \wPDiag_27[7] , \wPDiag_27[6] , 
        \wPDiag_27[5] , \wPDiag_27[4] , \wPDiag_27[3] , \wPDiag_27[2] , 
        \wPDiag_27[1] , \wPDiag_27[0] }), .NDiagIn({\wNDiag_27[31] , 
        \wNDiag_27[30] , \wNDiag_27[29] , \wNDiag_27[28] , \wNDiag_27[27] , 
        \wNDiag_27[26] , \wNDiag_27[25] , \wNDiag_27[24] , \wNDiag_27[23] , 
        \wNDiag_27[22] , \wNDiag_27[21] , \wNDiag_27[20] , \wNDiag_27[19] , 
        \wNDiag_27[18] , \wNDiag_27[17] , \wNDiag_27[16] , \wNDiag_27[15] , 
        \wNDiag_27[14] , \wNDiag_27[13] , \wNDiag_27[12] , \wNDiag_27[11] , 
        \wNDiag_27[10] , \wNDiag_27[9] , \wNDiag_27[8] , \wNDiag_27[7] , 
        \wNDiag_27[6] , \wNDiag_27[5] , \wNDiag_27[4] , \wNDiag_27[3] , 
        \wNDiag_27[2] , \wNDiag_27[1] , \wNDiag_27[0] }), .CallOut(
        \wCall_28[0] ), .ReturnOut(\wReturn_27[0] ), .ColOut({\wColumn_28[31] , 
        \wColumn_28[30] , \wColumn_28[29] , \wColumn_28[28] , \wColumn_28[27] , 
        \wColumn_28[26] , \wColumn_28[25] , \wColumn_28[24] , \wColumn_28[23] , 
        \wColumn_28[22] , \wColumn_28[21] , \wColumn_28[20] , \wColumn_28[19] , 
        \wColumn_28[18] , \wColumn_28[17] , \wColumn_28[16] , \wColumn_28[15] , 
        \wColumn_28[14] , \wColumn_28[13] , \wColumn_28[12] , \wColumn_28[11] , 
        \wColumn_28[10] , \wColumn_28[9] , \wColumn_28[8] , \wColumn_28[7] , 
        \wColumn_28[6] , \wColumn_28[5] , \wColumn_28[4] , \wColumn_28[3] , 
        \wColumn_28[2] , \wColumn_28[1] , \wColumn_28[0] }), .PDiagOut({
        \wPDiag_28[31] , \wPDiag_28[30] , \wPDiag_28[29] , \wPDiag_28[28] , 
        \wPDiag_28[27] , \wPDiag_28[26] , \wPDiag_28[25] , \wPDiag_28[24] , 
        \wPDiag_28[23] , \wPDiag_28[22] , \wPDiag_28[21] , \wPDiag_28[20] , 
        \wPDiag_28[19] , \wPDiag_28[18] , \wPDiag_28[17] , \wPDiag_28[16] , 
        \wPDiag_28[15] , \wPDiag_28[14] , \wPDiag_28[13] , \wPDiag_28[12] , 
        \wPDiag_28[11] , \wPDiag_28[10] , \wPDiag_28[9] , \wPDiag_28[8] , 
        \wPDiag_28[7] , \wPDiag_28[6] , \wPDiag_28[5] , \wPDiag_28[4] , 
        \wPDiag_28[3] , \wPDiag_28[2] , \wPDiag_28[1] , \wPDiag_28[0] }), 
        .NDiagOut({\wNDiag_28[31] , \wNDiag_28[30] , \wNDiag_28[29] , 
        \wNDiag_28[28] , \wNDiag_28[27] , \wNDiag_28[26] , \wNDiag_28[25] , 
        \wNDiag_28[24] , \wNDiag_28[23] , \wNDiag_28[22] , \wNDiag_28[21] , 
        \wNDiag_28[20] , \wNDiag_28[19] , \wNDiag_28[18] , \wNDiag_28[17] , 
        \wNDiag_28[16] , \wNDiag_28[15] , \wNDiag_28[14] , \wNDiag_28[13] , 
        \wNDiag_28[12] , \wNDiag_28[11] , \wNDiag_28[10] , \wNDiag_28[9] , 
        \wNDiag_28[8] , \wNDiag_28[7] , \wNDiag_28[6] , \wNDiag_28[5] , 
        \wNDiag_28[4] , \wNDiag_28[3] , \wNDiag_28[2] , \wNDiag_28[1] , 
        \wNDiag_28[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_4 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_5[5] , \wScan_5[4] , \wScan_5[3] , 
        \wScan_5[2] , \wScan_5[1] , \wScan_5[0] }), .ScanOut({\wScan_4[5] , 
        \wScan_4[4] , \wScan_4[3] , \wScan_4[2] , \wScan_4[1] , \wScan_4[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_4[0] ), .ReturnIn(\wReturn_5[0] ), .ColIn({
        \wColumn_4[31] , \wColumn_4[30] , \wColumn_4[29] , \wColumn_4[28] , 
        \wColumn_4[27] , \wColumn_4[26] , \wColumn_4[25] , \wColumn_4[24] , 
        \wColumn_4[23] , \wColumn_4[22] , \wColumn_4[21] , \wColumn_4[20] , 
        \wColumn_4[19] , \wColumn_4[18] , \wColumn_4[17] , \wColumn_4[16] , 
        \wColumn_4[15] , \wColumn_4[14] , \wColumn_4[13] , \wColumn_4[12] , 
        \wColumn_4[11] , \wColumn_4[10] , \wColumn_4[9] , \wColumn_4[8] , 
        \wColumn_4[7] , \wColumn_4[6] , \wColumn_4[5] , \wColumn_4[4] , 
        \wColumn_4[3] , \wColumn_4[2] , \wColumn_4[1] , \wColumn_4[0] }), 
        .PDiagIn({\wPDiag_4[31] , \wPDiag_4[30] , \wPDiag_4[29] , 
        \wPDiag_4[28] , \wPDiag_4[27] , \wPDiag_4[26] , \wPDiag_4[25] , 
        \wPDiag_4[24] , \wPDiag_4[23] , \wPDiag_4[22] , \wPDiag_4[21] , 
        \wPDiag_4[20] , \wPDiag_4[19] , \wPDiag_4[18] , \wPDiag_4[17] , 
        \wPDiag_4[16] , \wPDiag_4[15] , \wPDiag_4[14] , \wPDiag_4[13] , 
        \wPDiag_4[12] , \wPDiag_4[11] , \wPDiag_4[10] , \wPDiag_4[9] , 
        \wPDiag_4[8] , \wPDiag_4[7] , \wPDiag_4[6] , \wPDiag_4[5] , 
        \wPDiag_4[4] , \wPDiag_4[3] , \wPDiag_4[2] , \wPDiag_4[1] , 
        \wPDiag_4[0] }), .NDiagIn({\wNDiag_4[31] , \wNDiag_4[30] , 
        \wNDiag_4[29] , \wNDiag_4[28] , \wNDiag_4[27] , \wNDiag_4[26] , 
        \wNDiag_4[25] , \wNDiag_4[24] , \wNDiag_4[23] , \wNDiag_4[22] , 
        \wNDiag_4[21] , \wNDiag_4[20] , \wNDiag_4[19] , \wNDiag_4[18] , 
        \wNDiag_4[17] , \wNDiag_4[16] , \wNDiag_4[15] , \wNDiag_4[14] , 
        \wNDiag_4[13] , \wNDiag_4[12] , \wNDiag_4[11] , \wNDiag_4[10] , 
        \wNDiag_4[9] , \wNDiag_4[8] , \wNDiag_4[7] , \wNDiag_4[6] , 
        \wNDiag_4[5] , \wNDiag_4[4] , \wNDiag_4[3] , \wNDiag_4[2] , 
        \wNDiag_4[1] , \wNDiag_4[0] }), .CallOut(\wCall_5[0] ), .ReturnOut(
        \wReturn_4[0] ), .ColOut({\wColumn_5[31] , \wColumn_5[30] , 
        \wColumn_5[29] , \wColumn_5[28] , \wColumn_5[27] , \wColumn_5[26] , 
        \wColumn_5[25] , \wColumn_5[24] , \wColumn_5[23] , \wColumn_5[22] , 
        \wColumn_5[21] , \wColumn_5[20] , \wColumn_5[19] , \wColumn_5[18] , 
        \wColumn_5[17] , \wColumn_5[16] , \wColumn_5[15] , \wColumn_5[14] , 
        \wColumn_5[13] , \wColumn_5[12] , \wColumn_5[11] , \wColumn_5[10] , 
        \wColumn_5[9] , \wColumn_5[8] , \wColumn_5[7] , \wColumn_5[6] , 
        \wColumn_5[5] , \wColumn_5[4] , \wColumn_5[3] , \wColumn_5[2] , 
        \wColumn_5[1] , \wColumn_5[0] }), .PDiagOut({\wPDiag_5[31] , 
        \wPDiag_5[30] , \wPDiag_5[29] , \wPDiag_5[28] , \wPDiag_5[27] , 
        \wPDiag_5[26] , \wPDiag_5[25] , \wPDiag_5[24] , \wPDiag_5[23] , 
        \wPDiag_5[22] , \wPDiag_5[21] , \wPDiag_5[20] , \wPDiag_5[19] , 
        \wPDiag_5[18] , \wPDiag_5[17] , \wPDiag_5[16] , \wPDiag_5[15] , 
        \wPDiag_5[14] , \wPDiag_5[13] , \wPDiag_5[12] , \wPDiag_5[11] , 
        \wPDiag_5[10] , \wPDiag_5[9] , \wPDiag_5[8] , \wPDiag_5[7] , 
        \wPDiag_5[6] , \wPDiag_5[5] , \wPDiag_5[4] , \wPDiag_5[3] , 
        \wPDiag_5[2] , \wPDiag_5[1] , \wPDiag_5[0] }), .NDiagOut({
        \wNDiag_5[31] , \wNDiag_5[30] , \wNDiag_5[29] , \wNDiag_5[28] , 
        \wNDiag_5[27] , \wNDiag_5[26] , \wNDiag_5[25] , \wNDiag_5[24] , 
        \wNDiag_5[23] , \wNDiag_5[22] , \wNDiag_5[21] , \wNDiag_5[20] , 
        \wNDiag_5[19] , \wNDiag_5[18] , \wNDiag_5[17] , \wNDiag_5[16] , 
        \wNDiag_5[15] , \wNDiag_5[14] , \wNDiag_5[13] , \wNDiag_5[12] , 
        \wNDiag_5[11] , \wNDiag_5[10] , \wNDiag_5[9] , \wNDiag_5[8] , 
        \wNDiag_5[7] , \wNDiag_5[6] , \wNDiag_5[5] , \wNDiag_5[4] , 
        \wNDiag_5[3] , \wNDiag_5[2] , \wNDiag_5[1] , \wNDiag_5[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_5 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_6[5] , \wScan_6[4] , \wScan_6[3] , 
        \wScan_6[2] , \wScan_6[1] , \wScan_6[0] }), .ScanOut({\wScan_5[5] , 
        \wScan_5[4] , \wScan_5[3] , \wScan_5[2] , \wScan_5[1] , \wScan_5[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_5[0] ), .ReturnIn(\wReturn_6[0] ), .ColIn({
        \wColumn_5[31] , \wColumn_5[30] , \wColumn_5[29] , \wColumn_5[28] , 
        \wColumn_5[27] , \wColumn_5[26] , \wColumn_5[25] , \wColumn_5[24] , 
        \wColumn_5[23] , \wColumn_5[22] , \wColumn_5[21] , \wColumn_5[20] , 
        \wColumn_5[19] , \wColumn_5[18] , \wColumn_5[17] , \wColumn_5[16] , 
        \wColumn_5[15] , \wColumn_5[14] , \wColumn_5[13] , \wColumn_5[12] , 
        \wColumn_5[11] , \wColumn_5[10] , \wColumn_5[9] , \wColumn_5[8] , 
        \wColumn_5[7] , \wColumn_5[6] , \wColumn_5[5] , \wColumn_5[4] , 
        \wColumn_5[3] , \wColumn_5[2] , \wColumn_5[1] , \wColumn_5[0] }), 
        .PDiagIn({\wPDiag_5[31] , \wPDiag_5[30] , \wPDiag_5[29] , 
        \wPDiag_5[28] , \wPDiag_5[27] , \wPDiag_5[26] , \wPDiag_5[25] , 
        \wPDiag_5[24] , \wPDiag_5[23] , \wPDiag_5[22] , \wPDiag_5[21] , 
        \wPDiag_5[20] , \wPDiag_5[19] , \wPDiag_5[18] , \wPDiag_5[17] , 
        \wPDiag_5[16] , \wPDiag_5[15] , \wPDiag_5[14] , \wPDiag_5[13] , 
        \wPDiag_5[12] , \wPDiag_5[11] , \wPDiag_5[10] , \wPDiag_5[9] , 
        \wPDiag_5[8] , \wPDiag_5[7] , \wPDiag_5[6] , \wPDiag_5[5] , 
        \wPDiag_5[4] , \wPDiag_5[3] , \wPDiag_5[2] , \wPDiag_5[1] , 
        \wPDiag_5[0] }), .NDiagIn({\wNDiag_5[31] , \wNDiag_5[30] , 
        \wNDiag_5[29] , \wNDiag_5[28] , \wNDiag_5[27] , \wNDiag_5[26] , 
        \wNDiag_5[25] , \wNDiag_5[24] , \wNDiag_5[23] , \wNDiag_5[22] , 
        \wNDiag_5[21] , \wNDiag_5[20] , \wNDiag_5[19] , \wNDiag_5[18] , 
        \wNDiag_5[17] , \wNDiag_5[16] , \wNDiag_5[15] , \wNDiag_5[14] , 
        \wNDiag_5[13] , \wNDiag_5[12] , \wNDiag_5[11] , \wNDiag_5[10] , 
        \wNDiag_5[9] , \wNDiag_5[8] , \wNDiag_5[7] , \wNDiag_5[6] , 
        \wNDiag_5[5] , \wNDiag_5[4] , \wNDiag_5[3] , \wNDiag_5[2] , 
        \wNDiag_5[1] , \wNDiag_5[0] }), .CallOut(\wCall_6[0] ), .ReturnOut(
        \wReturn_5[0] ), .ColOut({\wColumn_6[31] , \wColumn_6[30] , 
        \wColumn_6[29] , \wColumn_6[28] , \wColumn_6[27] , \wColumn_6[26] , 
        \wColumn_6[25] , \wColumn_6[24] , \wColumn_6[23] , \wColumn_6[22] , 
        \wColumn_6[21] , \wColumn_6[20] , \wColumn_6[19] , \wColumn_6[18] , 
        \wColumn_6[17] , \wColumn_6[16] , \wColumn_6[15] , \wColumn_6[14] , 
        \wColumn_6[13] , \wColumn_6[12] , \wColumn_6[11] , \wColumn_6[10] , 
        \wColumn_6[9] , \wColumn_6[8] , \wColumn_6[7] , \wColumn_6[6] , 
        \wColumn_6[5] , \wColumn_6[4] , \wColumn_6[3] , \wColumn_6[2] , 
        \wColumn_6[1] , \wColumn_6[0] }), .PDiagOut({\wPDiag_6[31] , 
        \wPDiag_6[30] , \wPDiag_6[29] , \wPDiag_6[28] , \wPDiag_6[27] , 
        \wPDiag_6[26] , \wPDiag_6[25] , \wPDiag_6[24] , \wPDiag_6[23] , 
        \wPDiag_6[22] , \wPDiag_6[21] , \wPDiag_6[20] , \wPDiag_6[19] , 
        \wPDiag_6[18] , \wPDiag_6[17] , \wPDiag_6[16] , \wPDiag_6[15] , 
        \wPDiag_6[14] , \wPDiag_6[13] , \wPDiag_6[12] , \wPDiag_6[11] , 
        \wPDiag_6[10] , \wPDiag_6[9] , \wPDiag_6[8] , \wPDiag_6[7] , 
        \wPDiag_6[6] , \wPDiag_6[5] , \wPDiag_6[4] , \wPDiag_6[3] , 
        \wPDiag_6[2] , \wPDiag_6[1] , \wPDiag_6[0] }), .NDiagOut({
        \wNDiag_6[31] , \wNDiag_6[30] , \wNDiag_6[29] , \wNDiag_6[28] , 
        \wNDiag_6[27] , \wNDiag_6[26] , \wNDiag_6[25] , \wNDiag_6[24] , 
        \wNDiag_6[23] , \wNDiag_6[22] , \wNDiag_6[21] , \wNDiag_6[20] , 
        \wNDiag_6[19] , \wNDiag_6[18] , \wNDiag_6[17] , \wNDiag_6[16] , 
        \wNDiag_6[15] , \wNDiag_6[14] , \wNDiag_6[13] , \wNDiag_6[12] , 
        \wNDiag_6[11] , \wNDiag_6[10] , \wNDiag_6[9] , \wNDiag_6[8] , 
        \wNDiag_6[7] , \wNDiag_6[6] , \wNDiag_6[5] , \wNDiag_6[4] , 
        \wNDiag_6[3] , \wNDiag_6[2] , \wNDiag_6[1] , \wNDiag_6[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_15 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_16[5] , \wScan_16[4] , \wScan_16[3] , 
        \wScan_16[2] , \wScan_16[1] , \wScan_16[0] }), .ScanOut({\wScan_15[5] , 
        \wScan_15[4] , \wScan_15[3] , \wScan_15[2] , \wScan_15[1] , 
        \wScan_15[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_15[0] ), .ReturnIn(\wReturn_16[0] ), 
        .ColIn({\wColumn_15[31] , \wColumn_15[30] , \wColumn_15[29] , 
        \wColumn_15[28] , \wColumn_15[27] , \wColumn_15[26] , \wColumn_15[25] , 
        \wColumn_15[24] , \wColumn_15[23] , \wColumn_15[22] , \wColumn_15[21] , 
        \wColumn_15[20] , \wColumn_15[19] , \wColumn_15[18] , \wColumn_15[17] , 
        \wColumn_15[16] , \wColumn_15[15] , \wColumn_15[14] , \wColumn_15[13] , 
        \wColumn_15[12] , \wColumn_15[11] , \wColumn_15[10] , \wColumn_15[9] , 
        \wColumn_15[8] , \wColumn_15[7] , \wColumn_15[6] , \wColumn_15[5] , 
        \wColumn_15[4] , \wColumn_15[3] , \wColumn_15[2] , \wColumn_15[1] , 
        \wColumn_15[0] }), .PDiagIn({\wPDiag_15[31] , \wPDiag_15[30] , 
        \wPDiag_15[29] , \wPDiag_15[28] , \wPDiag_15[27] , \wPDiag_15[26] , 
        \wPDiag_15[25] , \wPDiag_15[24] , \wPDiag_15[23] , \wPDiag_15[22] , 
        \wPDiag_15[21] , \wPDiag_15[20] , \wPDiag_15[19] , \wPDiag_15[18] , 
        \wPDiag_15[17] , \wPDiag_15[16] , \wPDiag_15[15] , \wPDiag_15[14] , 
        \wPDiag_15[13] , \wPDiag_15[12] , \wPDiag_15[11] , \wPDiag_15[10] , 
        \wPDiag_15[9] , \wPDiag_15[8] , \wPDiag_15[7] , \wPDiag_15[6] , 
        \wPDiag_15[5] , \wPDiag_15[4] , \wPDiag_15[3] , \wPDiag_15[2] , 
        \wPDiag_15[1] , \wPDiag_15[0] }), .NDiagIn({\wNDiag_15[31] , 
        \wNDiag_15[30] , \wNDiag_15[29] , \wNDiag_15[28] , \wNDiag_15[27] , 
        \wNDiag_15[26] , \wNDiag_15[25] , \wNDiag_15[24] , \wNDiag_15[23] , 
        \wNDiag_15[22] , \wNDiag_15[21] , \wNDiag_15[20] , \wNDiag_15[19] , 
        \wNDiag_15[18] , \wNDiag_15[17] , \wNDiag_15[16] , \wNDiag_15[15] , 
        \wNDiag_15[14] , \wNDiag_15[13] , \wNDiag_15[12] , \wNDiag_15[11] , 
        \wNDiag_15[10] , \wNDiag_15[9] , \wNDiag_15[8] , \wNDiag_15[7] , 
        \wNDiag_15[6] , \wNDiag_15[5] , \wNDiag_15[4] , \wNDiag_15[3] , 
        \wNDiag_15[2] , \wNDiag_15[1] , \wNDiag_15[0] }), .CallOut(
        \wCall_16[0] ), .ReturnOut(\wReturn_15[0] ), .ColOut({\wColumn_16[31] , 
        \wColumn_16[30] , \wColumn_16[29] , \wColumn_16[28] , \wColumn_16[27] , 
        \wColumn_16[26] , \wColumn_16[25] , \wColumn_16[24] , \wColumn_16[23] , 
        \wColumn_16[22] , \wColumn_16[21] , \wColumn_16[20] , \wColumn_16[19] , 
        \wColumn_16[18] , \wColumn_16[17] , \wColumn_16[16] , \wColumn_16[15] , 
        \wColumn_16[14] , \wColumn_16[13] , \wColumn_16[12] , \wColumn_16[11] , 
        \wColumn_16[10] , \wColumn_16[9] , \wColumn_16[8] , \wColumn_16[7] , 
        \wColumn_16[6] , \wColumn_16[5] , \wColumn_16[4] , \wColumn_16[3] , 
        \wColumn_16[2] , \wColumn_16[1] , \wColumn_16[0] }), .PDiagOut({
        \wPDiag_16[31] , \wPDiag_16[30] , \wPDiag_16[29] , \wPDiag_16[28] , 
        \wPDiag_16[27] , \wPDiag_16[26] , \wPDiag_16[25] , \wPDiag_16[24] , 
        \wPDiag_16[23] , \wPDiag_16[22] , \wPDiag_16[21] , \wPDiag_16[20] , 
        \wPDiag_16[19] , \wPDiag_16[18] , \wPDiag_16[17] , \wPDiag_16[16] , 
        \wPDiag_16[15] , \wPDiag_16[14] , \wPDiag_16[13] , \wPDiag_16[12] , 
        \wPDiag_16[11] , \wPDiag_16[10] , \wPDiag_16[9] , \wPDiag_16[8] , 
        \wPDiag_16[7] , \wPDiag_16[6] , \wPDiag_16[5] , \wPDiag_16[4] , 
        \wPDiag_16[3] , \wPDiag_16[2] , \wPDiag_16[1] , \wPDiag_16[0] }), 
        .NDiagOut({\wNDiag_16[31] , \wNDiag_16[30] , \wNDiag_16[29] , 
        \wNDiag_16[28] , \wNDiag_16[27] , \wNDiag_16[26] , \wNDiag_16[25] , 
        \wNDiag_16[24] , \wNDiag_16[23] , \wNDiag_16[22] , \wNDiag_16[21] , 
        \wNDiag_16[20] , \wNDiag_16[19] , \wNDiag_16[18] , \wNDiag_16[17] , 
        \wNDiag_16[16] , \wNDiag_16[15] , \wNDiag_16[14] , \wNDiag_16[13] , 
        \wNDiag_16[12] , \wNDiag_16[11] , \wNDiag_16[10] , \wNDiag_16[9] , 
        \wNDiag_16[8] , \wNDiag_16[7] , \wNDiag_16[6] , \wNDiag_16[5] , 
        \wNDiag_16[4] , \wNDiag_16[3] , \wNDiag_16[2] , \wNDiag_16[1] , 
        \wNDiag_16[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_20 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_21[5] , \wScan_21[4] , \wScan_21[3] , 
        \wScan_21[2] , \wScan_21[1] , \wScan_21[0] }), .ScanOut({\wScan_20[5] , 
        \wScan_20[4] , \wScan_20[3] , \wScan_20[2] , \wScan_20[1] , 
        \wScan_20[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_20[0] ), .ReturnIn(\wReturn_21[0] ), 
        .ColIn({\wColumn_20[31] , \wColumn_20[30] , \wColumn_20[29] , 
        \wColumn_20[28] , \wColumn_20[27] , \wColumn_20[26] , \wColumn_20[25] , 
        \wColumn_20[24] , \wColumn_20[23] , \wColumn_20[22] , \wColumn_20[21] , 
        \wColumn_20[20] , \wColumn_20[19] , \wColumn_20[18] , \wColumn_20[17] , 
        \wColumn_20[16] , \wColumn_20[15] , \wColumn_20[14] , \wColumn_20[13] , 
        \wColumn_20[12] , \wColumn_20[11] , \wColumn_20[10] , \wColumn_20[9] , 
        \wColumn_20[8] , \wColumn_20[7] , \wColumn_20[6] , \wColumn_20[5] , 
        \wColumn_20[4] , \wColumn_20[3] , \wColumn_20[2] , \wColumn_20[1] , 
        \wColumn_20[0] }), .PDiagIn({\wPDiag_20[31] , \wPDiag_20[30] , 
        \wPDiag_20[29] , \wPDiag_20[28] , \wPDiag_20[27] , \wPDiag_20[26] , 
        \wPDiag_20[25] , \wPDiag_20[24] , \wPDiag_20[23] , \wPDiag_20[22] , 
        \wPDiag_20[21] , \wPDiag_20[20] , \wPDiag_20[19] , \wPDiag_20[18] , 
        \wPDiag_20[17] , \wPDiag_20[16] , \wPDiag_20[15] , \wPDiag_20[14] , 
        \wPDiag_20[13] , \wPDiag_20[12] , \wPDiag_20[11] , \wPDiag_20[10] , 
        \wPDiag_20[9] , \wPDiag_20[8] , \wPDiag_20[7] , \wPDiag_20[6] , 
        \wPDiag_20[5] , \wPDiag_20[4] , \wPDiag_20[3] , \wPDiag_20[2] , 
        \wPDiag_20[1] , \wPDiag_20[0] }), .NDiagIn({\wNDiag_20[31] , 
        \wNDiag_20[30] , \wNDiag_20[29] , \wNDiag_20[28] , \wNDiag_20[27] , 
        \wNDiag_20[26] , \wNDiag_20[25] , \wNDiag_20[24] , \wNDiag_20[23] , 
        \wNDiag_20[22] , \wNDiag_20[21] , \wNDiag_20[20] , \wNDiag_20[19] , 
        \wNDiag_20[18] , \wNDiag_20[17] , \wNDiag_20[16] , \wNDiag_20[15] , 
        \wNDiag_20[14] , \wNDiag_20[13] , \wNDiag_20[12] , \wNDiag_20[11] , 
        \wNDiag_20[10] , \wNDiag_20[9] , \wNDiag_20[8] , \wNDiag_20[7] , 
        \wNDiag_20[6] , \wNDiag_20[5] , \wNDiag_20[4] , \wNDiag_20[3] , 
        \wNDiag_20[2] , \wNDiag_20[1] , \wNDiag_20[0] }), .CallOut(
        \wCall_21[0] ), .ReturnOut(\wReturn_20[0] ), .ColOut({\wColumn_21[31] , 
        \wColumn_21[30] , \wColumn_21[29] , \wColumn_21[28] , \wColumn_21[27] , 
        \wColumn_21[26] , \wColumn_21[25] , \wColumn_21[24] , \wColumn_21[23] , 
        \wColumn_21[22] , \wColumn_21[21] , \wColumn_21[20] , \wColumn_21[19] , 
        \wColumn_21[18] , \wColumn_21[17] , \wColumn_21[16] , \wColumn_21[15] , 
        \wColumn_21[14] , \wColumn_21[13] , \wColumn_21[12] , \wColumn_21[11] , 
        \wColumn_21[10] , \wColumn_21[9] , \wColumn_21[8] , \wColumn_21[7] , 
        \wColumn_21[6] , \wColumn_21[5] , \wColumn_21[4] , \wColumn_21[3] , 
        \wColumn_21[2] , \wColumn_21[1] , \wColumn_21[0] }), .PDiagOut({
        \wPDiag_21[31] , \wPDiag_21[30] , \wPDiag_21[29] , \wPDiag_21[28] , 
        \wPDiag_21[27] , \wPDiag_21[26] , \wPDiag_21[25] , \wPDiag_21[24] , 
        \wPDiag_21[23] , \wPDiag_21[22] , \wPDiag_21[21] , \wPDiag_21[20] , 
        \wPDiag_21[19] , \wPDiag_21[18] , \wPDiag_21[17] , \wPDiag_21[16] , 
        \wPDiag_21[15] , \wPDiag_21[14] , \wPDiag_21[13] , \wPDiag_21[12] , 
        \wPDiag_21[11] , \wPDiag_21[10] , \wPDiag_21[9] , \wPDiag_21[8] , 
        \wPDiag_21[7] , \wPDiag_21[6] , \wPDiag_21[5] , \wPDiag_21[4] , 
        \wPDiag_21[3] , \wPDiag_21[2] , \wPDiag_21[1] , \wPDiag_21[0] }), 
        .NDiagOut({\wNDiag_21[31] , \wNDiag_21[30] , \wNDiag_21[29] , 
        \wNDiag_21[28] , \wNDiag_21[27] , \wNDiag_21[26] , \wNDiag_21[25] , 
        \wNDiag_21[24] , \wNDiag_21[23] , \wNDiag_21[22] , \wNDiag_21[21] , 
        \wNDiag_21[20] , \wNDiag_21[19] , \wNDiag_21[18] , \wNDiag_21[17] , 
        \wNDiag_21[16] , \wNDiag_21[15] , \wNDiag_21[14] , \wNDiag_21[13] , 
        \wNDiag_21[12] , \wNDiag_21[11] , \wNDiag_21[10] , \wNDiag_21[9] , 
        \wNDiag_21[8] , \wNDiag_21[7] , \wNDiag_21[6] , \wNDiag_21[5] , 
        \wNDiag_21[4] , \wNDiag_21[3] , \wNDiag_21[2] , \wNDiag_21[1] , 
        \wNDiag_21[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_21 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_22[5] , \wScan_22[4] , \wScan_22[3] , 
        \wScan_22[2] , \wScan_22[1] , \wScan_22[0] }), .ScanOut({\wScan_21[5] , 
        \wScan_21[4] , \wScan_21[3] , \wScan_21[2] , \wScan_21[1] , 
        \wScan_21[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_21[0] ), .ReturnIn(\wReturn_22[0] ), 
        .ColIn({\wColumn_21[31] , \wColumn_21[30] , \wColumn_21[29] , 
        \wColumn_21[28] , \wColumn_21[27] , \wColumn_21[26] , \wColumn_21[25] , 
        \wColumn_21[24] , \wColumn_21[23] , \wColumn_21[22] , \wColumn_21[21] , 
        \wColumn_21[20] , \wColumn_21[19] , \wColumn_21[18] , \wColumn_21[17] , 
        \wColumn_21[16] , \wColumn_21[15] , \wColumn_21[14] , \wColumn_21[13] , 
        \wColumn_21[12] , \wColumn_21[11] , \wColumn_21[10] , \wColumn_21[9] , 
        \wColumn_21[8] , \wColumn_21[7] , \wColumn_21[6] , \wColumn_21[5] , 
        \wColumn_21[4] , \wColumn_21[3] , \wColumn_21[2] , \wColumn_21[1] , 
        \wColumn_21[0] }), .PDiagIn({\wPDiag_21[31] , \wPDiag_21[30] , 
        \wPDiag_21[29] , \wPDiag_21[28] , \wPDiag_21[27] , \wPDiag_21[26] , 
        \wPDiag_21[25] , \wPDiag_21[24] , \wPDiag_21[23] , \wPDiag_21[22] , 
        \wPDiag_21[21] , \wPDiag_21[20] , \wPDiag_21[19] , \wPDiag_21[18] , 
        \wPDiag_21[17] , \wPDiag_21[16] , \wPDiag_21[15] , \wPDiag_21[14] , 
        \wPDiag_21[13] , \wPDiag_21[12] , \wPDiag_21[11] , \wPDiag_21[10] , 
        \wPDiag_21[9] , \wPDiag_21[8] , \wPDiag_21[7] , \wPDiag_21[6] , 
        \wPDiag_21[5] , \wPDiag_21[4] , \wPDiag_21[3] , \wPDiag_21[2] , 
        \wPDiag_21[1] , \wPDiag_21[0] }), .NDiagIn({\wNDiag_21[31] , 
        \wNDiag_21[30] , \wNDiag_21[29] , \wNDiag_21[28] , \wNDiag_21[27] , 
        \wNDiag_21[26] , \wNDiag_21[25] , \wNDiag_21[24] , \wNDiag_21[23] , 
        \wNDiag_21[22] , \wNDiag_21[21] , \wNDiag_21[20] , \wNDiag_21[19] , 
        \wNDiag_21[18] , \wNDiag_21[17] , \wNDiag_21[16] , \wNDiag_21[15] , 
        \wNDiag_21[14] , \wNDiag_21[13] , \wNDiag_21[12] , \wNDiag_21[11] , 
        \wNDiag_21[10] , \wNDiag_21[9] , \wNDiag_21[8] , \wNDiag_21[7] , 
        \wNDiag_21[6] , \wNDiag_21[5] , \wNDiag_21[4] , \wNDiag_21[3] , 
        \wNDiag_21[2] , \wNDiag_21[1] , \wNDiag_21[0] }), .CallOut(
        \wCall_22[0] ), .ReturnOut(\wReturn_21[0] ), .ColOut({\wColumn_22[31] , 
        \wColumn_22[30] , \wColumn_22[29] , \wColumn_22[28] , \wColumn_22[27] , 
        \wColumn_22[26] , \wColumn_22[25] , \wColumn_22[24] , \wColumn_22[23] , 
        \wColumn_22[22] , \wColumn_22[21] , \wColumn_22[20] , \wColumn_22[19] , 
        \wColumn_22[18] , \wColumn_22[17] , \wColumn_22[16] , \wColumn_22[15] , 
        \wColumn_22[14] , \wColumn_22[13] , \wColumn_22[12] , \wColumn_22[11] , 
        \wColumn_22[10] , \wColumn_22[9] , \wColumn_22[8] , \wColumn_22[7] , 
        \wColumn_22[6] , \wColumn_22[5] , \wColumn_22[4] , \wColumn_22[3] , 
        \wColumn_22[2] , \wColumn_22[1] , \wColumn_22[0] }), .PDiagOut({
        \wPDiag_22[31] , \wPDiag_22[30] , \wPDiag_22[29] , \wPDiag_22[28] , 
        \wPDiag_22[27] , \wPDiag_22[26] , \wPDiag_22[25] , \wPDiag_22[24] , 
        \wPDiag_22[23] , \wPDiag_22[22] , \wPDiag_22[21] , \wPDiag_22[20] , 
        \wPDiag_22[19] , \wPDiag_22[18] , \wPDiag_22[17] , \wPDiag_22[16] , 
        \wPDiag_22[15] , \wPDiag_22[14] , \wPDiag_22[13] , \wPDiag_22[12] , 
        \wPDiag_22[11] , \wPDiag_22[10] , \wPDiag_22[9] , \wPDiag_22[8] , 
        \wPDiag_22[7] , \wPDiag_22[6] , \wPDiag_22[5] , \wPDiag_22[4] , 
        \wPDiag_22[3] , \wPDiag_22[2] , \wPDiag_22[1] , \wPDiag_22[0] }), 
        .NDiagOut({\wNDiag_22[31] , \wNDiag_22[30] , \wNDiag_22[29] , 
        \wNDiag_22[28] , \wNDiag_22[27] , \wNDiag_22[26] , \wNDiag_22[25] , 
        \wNDiag_22[24] , \wNDiag_22[23] , \wNDiag_22[22] , \wNDiag_22[21] , 
        \wNDiag_22[20] , \wNDiag_22[19] , \wNDiag_22[18] , \wNDiag_22[17] , 
        \wNDiag_22[16] , \wNDiag_22[15] , \wNDiag_22[14] , \wNDiag_22[13] , 
        \wNDiag_22[12] , \wNDiag_22[11] , \wNDiag_22[10] , \wNDiag_22[9] , 
        \wNDiag_22[8] , \wNDiag_22[7] , \wNDiag_22[6] , \wNDiag_22[5] , 
        \wNDiag_22[4] , \wNDiag_22[3] , \wNDiag_22[2] , \wNDiag_22[1] , 
        \wNDiag_22[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_29 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_30[5] , \wScan_30[4] , \wScan_30[3] , 
        \wScan_30[2] , \wScan_30[1] , \wScan_30[0] }), .ScanOut({\wScan_29[5] , 
        \wScan_29[4] , \wScan_29[3] , \wScan_29[2] , \wScan_29[1] , 
        \wScan_29[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_29[0] ), .ReturnIn(\wReturn_30[0] ), 
        .ColIn({\wColumn_29[31] , \wColumn_29[30] , \wColumn_29[29] , 
        \wColumn_29[28] , \wColumn_29[27] , \wColumn_29[26] , \wColumn_29[25] , 
        \wColumn_29[24] , \wColumn_29[23] , \wColumn_29[22] , \wColumn_29[21] , 
        \wColumn_29[20] , \wColumn_29[19] , \wColumn_29[18] , \wColumn_29[17] , 
        \wColumn_29[16] , \wColumn_29[15] , \wColumn_29[14] , \wColumn_29[13] , 
        \wColumn_29[12] , \wColumn_29[11] , \wColumn_29[10] , \wColumn_29[9] , 
        \wColumn_29[8] , \wColumn_29[7] , \wColumn_29[6] , \wColumn_29[5] , 
        \wColumn_29[4] , \wColumn_29[3] , \wColumn_29[2] , \wColumn_29[1] , 
        \wColumn_29[0] }), .PDiagIn({\wPDiag_29[31] , \wPDiag_29[30] , 
        \wPDiag_29[29] , \wPDiag_29[28] , \wPDiag_29[27] , \wPDiag_29[26] , 
        \wPDiag_29[25] , \wPDiag_29[24] , \wPDiag_29[23] , \wPDiag_29[22] , 
        \wPDiag_29[21] , \wPDiag_29[20] , \wPDiag_29[19] , \wPDiag_29[18] , 
        \wPDiag_29[17] , \wPDiag_29[16] , \wPDiag_29[15] , \wPDiag_29[14] , 
        \wPDiag_29[13] , \wPDiag_29[12] , \wPDiag_29[11] , \wPDiag_29[10] , 
        \wPDiag_29[9] , \wPDiag_29[8] , \wPDiag_29[7] , \wPDiag_29[6] , 
        \wPDiag_29[5] , \wPDiag_29[4] , \wPDiag_29[3] , \wPDiag_29[2] , 
        \wPDiag_29[1] , \wPDiag_29[0] }), .NDiagIn({\wNDiag_29[31] , 
        \wNDiag_29[30] , \wNDiag_29[29] , \wNDiag_29[28] , \wNDiag_29[27] , 
        \wNDiag_29[26] , \wNDiag_29[25] , \wNDiag_29[24] , \wNDiag_29[23] , 
        \wNDiag_29[22] , \wNDiag_29[21] , \wNDiag_29[20] , \wNDiag_29[19] , 
        \wNDiag_29[18] , \wNDiag_29[17] , \wNDiag_29[16] , \wNDiag_29[15] , 
        \wNDiag_29[14] , \wNDiag_29[13] , \wNDiag_29[12] , \wNDiag_29[11] , 
        \wNDiag_29[10] , \wNDiag_29[9] , \wNDiag_29[8] , \wNDiag_29[7] , 
        \wNDiag_29[6] , \wNDiag_29[5] , \wNDiag_29[4] , \wNDiag_29[3] , 
        \wNDiag_29[2] , \wNDiag_29[1] , \wNDiag_29[0] }), .CallOut(
        \wCall_30[0] ), .ReturnOut(\wReturn_29[0] ), .ColOut({\wColumn_30[31] , 
        \wColumn_30[30] , \wColumn_30[29] , \wColumn_30[28] , \wColumn_30[27] , 
        \wColumn_30[26] , \wColumn_30[25] , \wColumn_30[24] , \wColumn_30[23] , 
        \wColumn_30[22] , \wColumn_30[21] , \wColumn_30[20] , \wColumn_30[19] , 
        \wColumn_30[18] , \wColumn_30[17] , \wColumn_30[16] , \wColumn_30[15] , 
        \wColumn_30[14] , \wColumn_30[13] , \wColumn_30[12] , \wColumn_30[11] , 
        \wColumn_30[10] , \wColumn_30[9] , \wColumn_30[8] , \wColumn_30[7] , 
        \wColumn_30[6] , \wColumn_30[5] , \wColumn_30[4] , \wColumn_30[3] , 
        \wColumn_30[2] , \wColumn_30[1] , \wColumn_30[0] }), .PDiagOut({
        \wPDiag_30[31] , \wPDiag_30[30] , \wPDiag_30[29] , \wPDiag_30[28] , 
        \wPDiag_30[27] , \wPDiag_30[26] , \wPDiag_30[25] , \wPDiag_30[24] , 
        \wPDiag_30[23] , \wPDiag_30[22] , \wPDiag_30[21] , \wPDiag_30[20] , 
        \wPDiag_30[19] , \wPDiag_30[18] , \wPDiag_30[17] , \wPDiag_30[16] , 
        \wPDiag_30[15] , \wPDiag_30[14] , \wPDiag_30[13] , \wPDiag_30[12] , 
        \wPDiag_30[11] , \wPDiag_30[10] , \wPDiag_30[9] , \wPDiag_30[8] , 
        \wPDiag_30[7] , \wPDiag_30[6] , \wPDiag_30[5] , \wPDiag_30[4] , 
        \wPDiag_30[3] , \wPDiag_30[2] , \wPDiag_30[1] , \wPDiag_30[0] }), 
        .NDiagOut({\wNDiag_30[31] , \wNDiag_30[30] , \wNDiag_30[29] , 
        \wNDiag_30[28] , \wNDiag_30[27] , \wNDiag_30[26] , \wNDiag_30[25] , 
        \wNDiag_30[24] , \wNDiag_30[23] , \wNDiag_30[22] , \wNDiag_30[21] , 
        \wNDiag_30[20] , \wNDiag_30[19] , \wNDiag_30[18] , \wNDiag_30[17] , 
        \wNDiag_30[16] , \wNDiag_30[15] , \wNDiag_30[14] , \wNDiag_30[13] , 
        \wNDiag_30[12] , \wNDiag_30[11] , \wNDiag_30[10] , \wNDiag_30[9] , 
        \wNDiag_30[8] , \wNDiag_30[7] , \wNDiag_30[6] , \wNDiag_30[5] , 
        \wNDiag_30[4] , \wNDiag_30[3] , \wNDiag_30[2] , \wNDiag_30[1] , 
        \wNDiag_30[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_13 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_14[5] , \wScan_14[4] , \wScan_14[3] , 
        \wScan_14[2] , \wScan_14[1] , \wScan_14[0] }), .ScanOut({\wScan_13[5] , 
        \wScan_13[4] , \wScan_13[3] , \wScan_13[2] , \wScan_13[1] , 
        \wScan_13[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_13[0] ), .ReturnIn(\wReturn_14[0] ), 
        .ColIn({\wColumn_13[31] , \wColumn_13[30] , \wColumn_13[29] , 
        \wColumn_13[28] , \wColumn_13[27] , \wColumn_13[26] , \wColumn_13[25] , 
        \wColumn_13[24] , \wColumn_13[23] , \wColumn_13[22] , \wColumn_13[21] , 
        \wColumn_13[20] , \wColumn_13[19] , \wColumn_13[18] , \wColumn_13[17] , 
        \wColumn_13[16] , \wColumn_13[15] , \wColumn_13[14] , \wColumn_13[13] , 
        \wColumn_13[12] , \wColumn_13[11] , \wColumn_13[10] , \wColumn_13[9] , 
        \wColumn_13[8] , \wColumn_13[7] , \wColumn_13[6] , \wColumn_13[5] , 
        \wColumn_13[4] , \wColumn_13[3] , \wColumn_13[2] , \wColumn_13[1] , 
        \wColumn_13[0] }), .PDiagIn({\wPDiag_13[31] , \wPDiag_13[30] , 
        \wPDiag_13[29] , \wPDiag_13[28] , \wPDiag_13[27] , \wPDiag_13[26] , 
        \wPDiag_13[25] , \wPDiag_13[24] , \wPDiag_13[23] , \wPDiag_13[22] , 
        \wPDiag_13[21] , \wPDiag_13[20] , \wPDiag_13[19] , \wPDiag_13[18] , 
        \wPDiag_13[17] , \wPDiag_13[16] , \wPDiag_13[15] , \wPDiag_13[14] , 
        \wPDiag_13[13] , \wPDiag_13[12] , \wPDiag_13[11] , \wPDiag_13[10] , 
        \wPDiag_13[9] , \wPDiag_13[8] , \wPDiag_13[7] , \wPDiag_13[6] , 
        \wPDiag_13[5] , \wPDiag_13[4] , \wPDiag_13[3] , \wPDiag_13[2] , 
        \wPDiag_13[1] , \wPDiag_13[0] }), .NDiagIn({\wNDiag_13[31] , 
        \wNDiag_13[30] , \wNDiag_13[29] , \wNDiag_13[28] , \wNDiag_13[27] , 
        \wNDiag_13[26] , \wNDiag_13[25] , \wNDiag_13[24] , \wNDiag_13[23] , 
        \wNDiag_13[22] , \wNDiag_13[21] , \wNDiag_13[20] , \wNDiag_13[19] , 
        \wNDiag_13[18] , \wNDiag_13[17] , \wNDiag_13[16] , \wNDiag_13[15] , 
        \wNDiag_13[14] , \wNDiag_13[13] , \wNDiag_13[12] , \wNDiag_13[11] , 
        \wNDiag_13[10] , \wNDiag_13[9] , \wNDiag_13[8] , \wNDiag_13[7] , 
        \wNDiag_13[6] , \wNDiag_13[5] , \wNDiag_13[4] , \wNDiag_13[3] , 
        \wNDiag_13[2] , \wNDiag_13[1] , \wNDiag_13[0] }), .CallOut(
        \wCall_14[0] ), .ReturnOut(\wReturn_13[0] ), .ColOut({\wColumn_14[31] , 
        \wColumn_14[30] , \wColumn_14[29] , \wColumn_14[28] , \wColumn_14[27] , 
        \wColumn_14[26] , \wColumn_14[25] , \wColumn_14[24] , \wColumn_14[23] , 
        \wColumn_14[22] , \wColumn_14[21] , \wColumn_14[20] , \wColumn_14[19] , 
        \wColumn_14[18] , \wColumn_14[17] , \wColumn_14[16] , \wColumn_14[15] , 
        \wColumn_14[14] , \wColumn_14[13] , \wColumn_14[12] , \wColumn_14[11] , 
        \wColumn_14[10] , \wColumn_14[9] , \wColumn_14[8] , \wColumn_14[7] , 
        \wColumn_14[6] , \wColumn_14[5] , \wColumn_14[4] , \wColumn_14[3] , 
        \wColumn_14[2] , \wColumn_14[1] , \wColumn_14[0] }), .PDiagOut({
        \wPDiag_14[31] , \wPDiag_14[30] , \wPDiag_14[29] , \wPDiag_14[28] , 
        \wPDiag_14[27] , \wPDiag_14[26] , \wPDiag_14[25] , \wPDiag_14[24] , 
        \wPDiag_14[23] , \wPDiag_14[22] , \wPDiag_14[21] , \wPDiag_14[20] , 
        \wPDiag_14[19] , \wPDiag_14[18] , \wPDiag_14[17] , \wPDiag_14[16] , 
        \wPDiag_14[15] , \wPDiag_14[14] , \wPDiag_14[13] , \wPDiag_14[12] , 
        \wPDiag_14[11] , \wPDiag_14[10] , \wPDiag_14[9] , \wPDiag_14[8] , 
        \wPDiag_14[7] , \wPDiag_14[6] , \wPDiag_14[5] , \wPDiag_14[4] , 
        \wPDiag_14[3] , \wPDiag_14[2] , \wPDiag_14[1] , \wPDiag_14[0] }), 
        .NDiagOut({\wNDiag_14[31] , \wNDiag_14[30] , \wNDiag_14[29] , 
        \wNDiag_14[28] , \wNDiag_14[27] , \wNDiag_14[26] , \wNDiag_14[25] , 
        \wNDiag_14[24] , \wNDiag_14[23] , \wNDiag_14[22] , \wNDiag_14[21] , 
        \wNDiag_14[20] , \wNDiag_14[19] , \wNDiag_14[18] , \wNDiag_14[17] , 
        \wNDiag_14[16] , \wNDiag_14[15] , \wNDiag_14[14] , \wNDiag_14[13] , 
        \wNDiag_14[12] , \wNDiag_14[11] , \wNDiag_14[10] , \wNDiag_14[9] , 
        \wNDiag_14[8] , \wNDiag_14[7] , \wNDiag_14[6] , \wNDiag_14[5] , 
        \wNDiag_14[4] , \wNDiag_14[3] , \wNDiag_14[2] , \wNDiag_14[1] , 
        \wNDiag_14[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_14 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_15[5] , \wScan_15[4] , \wScan_15[3] , 
        \wScan_15[2] , \wScan_15[1] , \wScan_15[0] }), .ScanOut({\wScan_14[5] , 
        \wScan_14[4] , \wScan_14[3] , \wScan_14[2] , \wScan_14[1] , 
        \wScan_14[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_14[0] ), .ReturnIn(\wReturn_15[0] ), 
        .ColIn({\wColumn_14[31] , \wColumn_14[30] , \wColumn_14[29] , 
        \wColumn_14[28] , \wColumn_14[27] , \wColumn_14[26] , \wColumn_14[25] , 
        \wColumn_14[24] , \wColumn_14[23] , \wColumn_14[22] , \wColumn_14[21] , 
        \wColumn_14[20] , \wColumn_14[19] , \wColumn_14[18] , \wColumn_14[17] , 
        \wColumn_14[16] , \wColumn_14[15] , \wColumn_14[14] , \wColumn_14[13] , 
        \wColumn_14[12] , \wColumn_14[11] , \wColumn_14[10] , \wColumn_14[9] , 
        \wColumn_14[8] , \wColumn_14[7] , \wColumn_14[6] , \wColumn_14[5] , 
        \wColumn_14[4] , \wColumn_14[3] , \wColumn_14[2] , \wColumn_14[1] , 
        \wColumn_14[0] }), .PDiagIn({\wPDiag_14[31] , \wPDiag_14[30] , 
        \wPDiag_14[29] , \wPDiag_14[28] , \wPDiag_14[27] , \wPDiag_14[26] , 
        \wPDiag_14[25] , \wPDiag_14[24] , \wPDiag_14[23] , \wPDiag_14[22] , 
        \wPDiag_14[21] , \wPDiag_14[20] , \wPDiag_14[19] , \wPDiag_14[18] , 
        \wPDiag_14[17] , \wPDiag_14[16] , \wPDiag_14[15] , \wPDiag_14[14] , 
        \wPDiag_14[13] , \wPDiag_14[12] , \wPDiag_14[11] , \wPDiag_14[10] , 
        \wPDiag_14[9] , \wPDiag_14[8] , \wPDiag_14[7] , \wPDiag_14[6] , 
        \wPDiag_14[5] , \wPDiag_14[4] , \wPDiag_14[3] , \wPDiag_14[2] , 
        \wPDiag_14[1] , \wPDiag_14[0] }), .NDiagIn({\wNDiag_14[31] , 
        \wNDiag_14[30] , \wNDiag_14[29] , \wNDiag_14[28] , \wNDiag_14[27] , 
        \wNDiag_14[26] , \wNDiag_14[25] , \wNDiag_14[24] , \wNDiag_14[23] , 
        \wNDiag_14[22] , \wNDiag_14[21] , \wNDiag_14[20] , \wNDiag_14[19] , 
        \wNDiag_14[18] , \wNDiag_14[17] , \wNDiag_14[16] , \wNDiag_14[15] , 
        \wNDiag_14[14] , \wNDiag_14[13] , \wNDiag_14[12] , \wNDiag_14[11] , 
        \wNDiag_14[10] , \wNDiag_14[9] , \wNDiag_14[8] , \wNDiag_14[7] , 
        \wNDiag_14[6] , \wNDiag_14[5] , \wNDiag_14[4] , \wNDiag_14[3] , 
        \wNDiag_14[2] , \wNDiag_14[1] , \wNDiag_14[0] }), .CallOut(
        \wCall_15[0] ), .ReturnOut(\wReturn_14[0] ), .ColOut({\wColumn_15[31] , 
        \wColumn_15[30] , \wColumn_15[29] , \wColumn_15[28] , \wColumn_15[27] , 
        \wColumn_15[26] , \wColumn_15[25] , \wColumn_15[24] , \wColumn_15[23] , 
        \wColumn_15[22] , \wColumn_15[21] , \wColumn_15[20] , \wColumn_15[19] , 
        \wColumn_15[18] , \wColumn_15[17] , \wColumn_15[16] , \wColumn_15[15] , 
        \wColumn_15[14] , \wColumn_15[13] , \wColumn_15[12] , \wColumn_15[11] , 
        \wColumn_15[10] , \wColumn_15[9] , \wColumn_15[8] , \wColumn_15[7] , 
        \wColumn_15[6] , \wColumn_15[5] , \wColumn_15[4] , \wColumn_15[3] , 
        \wColumn_15[2] , \wColumn_15[1] , \wColumn_15[0] }), .PDiagOut({
        \wPDiag_15[31] , \wPDiag_15[30] , \wPDiag_15[29] , \wPDiag_15[28] , 
        \wPDiag_15[27] , \wPDiag_15[26] , \wPDiag_15[25] , \wPDiag_15[24] , 
        \wPDiag_15[23] , \wPDiag_15[22] , \wPDiag_15[21] , \wPDiag_15[20] , 
        \wPDiag_15[19] , \wPDiag_15[18] , \wPDiag_15[17] , \wPDiag_15[16] , 
        \wPDiag_15[15] , \wPDiag_15[14] , \wPDiag_15[13] , \wPDiag_15[12] , 
        \wPDiag_15[11] , \wPDiag_15[10] , \wPDiag_15[9] , \wPDiag_15[8] , 
        \wPDiag_15[7] , \wPDiag_15[6] , \wPDiag_15[5] , \wPDiag_15[4] , 
        \wPDiag_15[3] , \wPDiag_15[2] , \wPDiag_15[1] , \wPDiag_15[0] }), 
        .NDiagOut({\wNDiag_15[31] , \wNDiag_15[30] , \wNDiag_15[29] , 
        \wNDiag_15[28] , \wNDiag_15[27] , \wNDiag_15[26] , \wNDiag_15[25] , 
        \wNDiag_15[24] , \wNDiag_15[23] , \wNDiag_15[22] , \wNDiag_15[21] , 
        \wNDiag_15[20] , \wNDiag_15[19] , \wNDiag_15[18] , \wNDiag_15[17] , 
        \wNDiag_15[16] , \wNDiag_15[15] , \wNDiag_15[14] , \wNDiag_15[13] , 
        \wNDiag_15[12] , \wNDiag_15[11] , \wNDiag_15[10] , \wNDiag_15[9] , 
        \wNDiag_15[8] , \wNDiag_15[7] , \wNDiag_15[6] , \wNDiag_15[5] , 
        \wNDiag_15[4] , \wNDiag_15[3] , \wNDiag_15[2] , \wNDiag_15[1] , 
        \wNDiag_15[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_28 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_29[5] , \wScan_29[4] , \wScan_29[3] , 
        \wScan_29[2] , \wScan_29[1] , \wScan_29[0] }), .ScanOut({\wScan_28[5] , 
        \wScan_28[4] , \wScan_28[3] , \wScan_28[2] , \wScan_28[1] , 
        \wScan_28[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_28[0] ), .ReturnIn(\wReturn_29[0] ), 
        .ColIn({\wColumn_28[31] , \wColumn_28[30] , \wColumn_28[29] , 
        \wColumn_28[28] , \wColumn_28[27] , \wColumn_28[26] , \wColumn_28[25] , 
        \wColumn_28[24] , \wColumn_28[23] , \wColumn_28[22] , \wColumn_28[21] , 
        \wColumn_28[20] , \wColumn_28[19] , \wColumn_28[18] , \wColumn_28[17] , 
        \wColumn_28[16] , \wColumn_28[15] , \wColumn_28[14] , \wColumn_28[13] , 
        \wColumn_28[12] , \wColumn_28[11] , \wColumn_28[10] , \wColumn_28[9] , 
        \wColumn_28[8] , \wColumn_28[7] , \wColumn_28[6] , \wColumn_28[5] , 
        \wColumn_28[4] , \wColumn_28[3] , \wColumn_28[2] , \wColumn_28[1] , 
        \wColumn_28[0] }), .PDiagIn({\wPDiag_28[31] , \wPDiag_28[30] , 
        \wPDiag_28[29] , \wPDiag_28[28] , \wPDiag_28[27] , \wPDiag_28[26] , 
        \wPDiag_28[25] , \wPDiag_28[24] , \wPDiag_28[23] , \wPDiag_28[22] , 
        \wPDiag_28[21] , \wPDiag_28[20] , \wPDiag_28[19] , \wPDiag_28[18] , 
        \wPDiag_28[17] , \wPDiag_28[16] , \wPDiag_28[15] , \wPDiag_28[14] , 
        \wPDiag_28[13] , \wPDiag_28[12] , \wPDiag_28[11] , \wPDiag_28[10] , 
        \wPDiag_28[9] , \wPDiag_28[8] , \wPDiag_28[7] , \wPDiag_28[6] , 
        \wPDiag_28[5] , \wPDiag_28[4] , \wPDiag_28[3] , \wPDiag_28[2] , 
        \wPDiag_28[1] , \wPDiag_28[0] }), .NDiagIn({\wNDiag_28[31] , 
        \wNDiag_28[30] , \wNDiag_28[29] , \wNDiag_28[28] , \wNDiag_28[27] , 
        \wNDiag_28[26] , \wNDiag_28[25] , \wNDiag_28[24] , \wNDiag_28[23] , 
        \wNDiag_28[22] , \wNDiag_28[21] , \wNDiag_28[20] , \wNDiag_28[19] , 
        \wNDiag_28[18] , \wNDiag_28[17] , \wNDiag_28[16] , \wNDiag_28[15] , 
        \wNDiag_28[14] , \wNDiag_28[13] , \wNDiag_28[12] , \wNDiag_28[11] , 
        \wNDiag_28[10] , \wNDiag_28[9] , \wNDiag_28[8] , \wNDiag_28[7] , 
        \wNDiag_28[6] , \wNDiag_28[5] , \wNDiag_28[4] , \wNDiag_28[3] , 
        \wNDiag_28[2] , \wNDiag_28[1] , \wNDiag_28[0] }), .CallOut(
        \wCall_29[0] ), .ReturnOut(\wReturn_28[0] ), .ColOut({\wColumn_29[31] , 
        \wColumn_29[30] , \wColumn_29[29] , \wColumn_29[28] , \wColumn_29[27] , 
        \wColumn_29[26] , \wColumn_29[25] , \wColumn_29[24] , \wColumn_29[23] , 
        \wColumn_29[22] , \wColumn_29[21] , \wColumn_29[20] , \wColumn_29[19] , 
        \wColumn_29[18] , \wColumn_29[17] , \wColumn_29[16] , \wColumn_29[15] , 
        \wColumn_29[14] , \wColumn_29[13] , \wColumn_29[12] , \wColumn_29[11] , 
        \wColumn_29[10] , \wColumn_29[9] , \wColumn_29[8] , \wColumn_29[7] , 
        \wColumn_29[6] , \wColumn_29[5] , \wColumn_29[4] , \wColumn_29[3] , 
        \wColumn_29[2] , \wColumn_29[1] , \wColumn_29[0] }), .PDiagOut({
        \wPDiag_29[31] , \wPDiag_29[30] , \wPDiag_29[29] , \wPDiag_29[28] , 
        \wPDiag_29[27] , \wPDiag_29[26] , \wPDiag_29[25] , \wPDiag_29[24] , 
        \wPDiag_29[23] , \wPDiag_29[22] , \wPDiag_29[21] , \wPDiag_29[20] , 
        \wPDiag_29[19] , \wPDiag_29[18] , \wPDiag_29[17] , \wPDiag_29[16] , 
        \wPDiag_29[15] , \wPDiag_29[14] , \wPDiag_29[13] , \wPDiag_29[12] , 
        \wPDiag_29[11] , \wPDiag_29[10] , \wPDiag_29[9] , \wPDiag_29[8] , 
        \wPDiag_29[7] , \wPDiag_29[6] , \wPDiag_29[5] , \wPDiag_29[4] , 
        \wPDiag_29[3] , \wPDiag_29[2] , \wPDiag_29[1] , \wPDiag_29[0] }), 
        .NDiagOut({\wNDiag_29[31] , \wNDiag_29[30] , \wNDiag_29[29] , 
        \wNDiag_29[28] , \wNDiag_29[27] , \wNDiag_29[26] , \wNDiag_29[25] , 
        \wNDiag_29[24] , \wNDiag_29[23] , \wNDiag_29[22] , \wNDiag_29[21] , 
        \wNDiag_29[20] , \wNDiag_29[19] , \wNDiag_29[18] , \wNDiag_29[17] , 
        \wNDiag_29[16] , \wNDiag_29[15] , \wNDiag_29[14] , \wNDiag_29[13] , 
        \wNDiag_29[12] , \wNDiag_29[11] , \wNDiag_29[10] , \wNDiag_29[9] , 
        \wNDiag_29[8] , \wNDiag_29[7] , \wNDiag_29[6] , \wNDiag_29[5] , 
        \wNDiag_29[4] , \wNDiag_29[3] , \wNDiag_29[2] , \wNDiag_29[1] , 
        \wNDiag_29[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_9 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_10[5] , \wScan_10[4] , \wScan_10[3] , 
        \wScan_10[2] , \wScan_10[1] , \wScan_10[0] }), .ScanOut({\wScan_9[5] , 
        \wScan_9[4] , \wScan_9[3] , \wScan_9[2] , \wScan_9[1] , \wScan_9[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_9[0] ), .ReturnIn(\wReturn_10[0] ), .ColIn({
        \wColumn_9[31] , \wColumn_9[30] , \wColumn_9[29] , \wColumn_9[28] , 
        \wColumn_9[27] , \wColumn_9[26] , \wColumn_9[25] , \wColumn_9[24] , 
        \wColumn_9[23] , \wColumn_9[22] , \wColumn_9[21] , \wColumn_9[20] , 
        \wColumn_9[19] , \wColumn_9[18] , \wColumn_9[17] , \wColumn_9[16] , 
        \wColumn_9[15] , \wColumn_9[14] , \wColumn_9[13] , \wColumn_9[12] , 
        \wColumn_9[11] , \wColumn_9[10] , \wColumn_9[9] , \wColumn_9[8] , 
        \wColumn_9[7] , \wColumn_9[6] , \wColumn_9[5] , \wColumn_9[4] , 
        \wColumn_9[3] , \wColumn_9[2] , \wColumn_9[1] , \wColumn_9[0] }), 
        .PDiagIn({\wPDiag_9[31] , \wPDiag_9[30] , \wPDiag_9[29] , 
        \wPDiag_9[28] , \wPDiag_9[27] , \wPDiag_9[26] , \wPDiag_9[25] , 
        \wPDiag_9[24] , \wPDiag_9[23] , \wPDiag_9[22] , \wPDiag_9[21] , 
        \wPDiag_9[20] , \wPDiag_9[19] , \wPDiag_9[18] , \wPDiag_9[17] , 
        \wPDiag_9[16] , \wPDiag_9[15] , \wPDiag_9[14] , \wPDiag_9[13] , 
        \wPDiag_9[12] , \wPDiag_9[11] , \wPDiag_9[10] , \wPDiag_9[9] , 
        \wPDiag_9[8] , \wPDiag_9[7] , \wPDiag_9[6] , \wPDiag_9[5] , 
        \wPDiag_9[4] , \wPDiag_9[3] , \wPDiag_9[2] , \wPDiag_9[1] , 
        \wPDiag_9[0] }), .NDiagIn({\wNDiag_9[31] , \wNDiag_9[30] , 
        \wNDiag_9[29] , \wNDiag_9[28] , \wNDiag_9[27] , \wNDiag_9[26] , 
        \wNDiag_9[25] , \wNDiag_9[24] , \wNDiag_9[23] , \wNDiag_9[22] , 
        \wNDiag_9[21] , \wNDiag_9[20] , \wNDiag_9[19] , \wNDiag_9[18] , 
        \wNDiag_9[17] , \wNDiag_9[16] , \wNDiag_9[15] , \wNDiag_9[14] , 
        \wNDiag_9[13] , \wNDiag_9[12] , \wNDiag_9[11] , \wNDiag_9[10] , 
        \wNDiag_9[9] , \wNDiag_9[8] , \wNDiag_9[7] , \wNDiag_9[6] , 
        \wNDiag_9[5] , \wNDiag_9[4] , \wNDiag_9[3] , \wNDiag_9[2] , 
        \wNDiag_9[1] , \wNDiag_9[0] }), .CallOut(\wCall_10[0] ), .ReturnOut(
        \wReturn_9[0] ), .ColOut({\wColumn_10[31] , \wColumn_10[30] , 
        \wColumn_10[29] , \wColumn_10[28] , \wColumn_10[27] , \wColumn_10[26] , 
        \wColumn_10[25] , \wColumn_10[24] , \wColumn_10[23] , \wColumn_10[22] , 
        \wColumn_10[21] , \wColumn_10[20] , \wColumn_10[19] , \wColumn_10[18] , 
        \wColumn_10[17] , \wColumn_10[16] , \wColumn_10[15] , \wColumn_10[14] , 
        \wColumn_10[13] , \wColumn_10[12] , \wColumn_10[11] , \wColumn_10[10] , 
        \wColumn_10[9] , \wColumn_10[8] , \wColumn_10[7] , \wColumn_10[6] , 
        \wColumn_10[5] , \wColumn_10[4] , \wColumn_10[3] , \wColumn_10[2] , 
        \wColumn_10[1] , \wColumn_10[0] }), .PDiagOut({\wPDiag_10[31] , 
        \wPDiag_10[30] , \wPDiag_10[29] , \wPDiag_10[28] , \wPDiag_10[27] , 
        \wPDiag_10[26] , \wPDiag_10[25] , \wPDiag_10[24] , \wPDiag_10[23] , 
        \wPDiag_10[22] , \wPDiag_10[21] , \wPDiag_10[20] , \wPDiag_10[19] , 
        \wPDiag_10[18] , \wPDiag_10[17] , \wPDiag_10[16] , \wPDiag_10[15] , 
        \wPDiag_10[14] , \wPDiag_10[13] , \wPDiag_10[12] , \wPDiag_10[11] , 
        \wPDiag_10[10] , \wPDiag_10[9] , \wPDiag_10[8] , \wPDiag_10[7] , 
        \wPDiag_10[6] , \wPDiag_10[5] , \wPDiag_10[4] , \wPDiag_10[3] , 
        \wPDiag_10[2] , \wPDiag_10[1] , \wPDiag_10[0] }), .NDiagOut({
        \wNDiag_10[31] , \wNDiag_10[30] , \wNDiag_10[29] , \wNDiag_10[28] , 
        \wNDiag_10[27] , \wNDiag_10[26] , \wNDiag_10[25] , \wNDiag_10[24] , 
        \wNDiag_10[23] , \wNDiag_10[22] , \wNDiag_10[21] , \wNDiag_10[20] , 
        \wNDiag_10[19] , \wNDiag_10[18] , \wNDiag_10[17] , \wNDiag_10[16] , 
        \wNDiag_10[15] , \wNDiag_10[14] , \wNDiag_10[13] , \wNDiag_10[12] , 
        \wNDiag_10[11] , \wNDiag_10[10] , \wNDiag_10[9] , \wNDiag_10[8] , 
        \wNDiag_10[7] , \wNDiag_10[6] , \wNDiag_10[5] , \wNDiag_10[4] , 
        \wNDiag_10[3] , \wNDiag_10[2] , \wNDiag_10[1] , \wNDiag_10[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_26 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_27[5] , \wScan_27[4] , \wScan_27[3] , 
        \wScan_27[2] , \wScan_27[1] , \wScan_27[0] }), .ScanOut({\wScan_26[5] , 
        \wScan_26[4] , \wScan_26[3] , \wScan_26[2] , \wScan_26[1] , 
        \wScan_26[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_26[0] ), .ReturnIn(\wReturn_27[0] ), 
        .ColIn({\wColumn_26[31] , \wColumn_26[30] , \wColumn_26[29] , 
        \wColumn_26[28] , \wColumn_26[27] , \wColumn_26[26] , \wColumn_26[25] , 
        \wColumn_26[24] , \wColumn_26[23] , \wColumn_26[22] , \wColumn_26[21] , 
        \wColumn_26[20] , \wColumn_26[19] , \wColumn_26[18] , \wColumn_26[17] , 
        \wColumn_26[16] , \wColumn_26[15] , \wColumn_26[14] , \wColumn_26[13] , 
        \wColumn_26[12] , \wColumn_26[11] , \wColumn_26[10] , \wColumn_26[9] , 
        \wColumn_26[8] , \wColumn_26[7] , \wColumn_26[6] , \wColumn_26[5] , 
        \wColumn_26[4] , \wColumn_26[3] , \wColumn_26[2] , \wColumn_26[1] , 
        \wColumn_26[0] }), .PDiagIn({\wPDiag_26[31] , \wPDiag_26[30] , 
        \wPDiag_26[29] , \wPDiag_26[28] , \wPDiag_26[27] , \wPDiag_26[26] , 
        \wPDiag_26[25] , \wPDiag_26[24] , \wPDiag_26[23] , \wPDiag_26[22] , 
        \wPDiag_26[21] , \wPDiag_26[20] , \wPDiag_26[19] , \wPDiag_26[18] , 
        \wPDiag_26[17] , \wPDiag_26[16] , \wPDiag_26[15] , \wPDiag_26[14] , 
        \wPDiag_26[13] , \wPDiag_26[12] , \wPDiag_26[11] , \wPDiag_26[10] , 
        \wPDiag_26[9] , \wPDiag_26[8] , \wPDiag_26[7] , \wPDiag_26[6] , 
        \wPDiag_26[5] , \wPDiag_26[4] , \wPDiag_26[3] , \wPDiag_26[2] , 
        \wPDiag_26[1] , \wPDiag_26[0] }), .NDiagIn({\wNDiag_26[31] , 
        \wNDiag_26[30] , \wNDiag_26[29] , \wNDiag_26[28] , \wNDiag_26[27] , 
        \wNDiag_26[26] , \wNDiag_26[25] , \wNDiag_26[24] , \wNDiag_26[23] , 
        \wNDiag_26[22] , \wNDiag_26[21] , \wNDiag_26[20] , \wNDiag_26[19] , 
        \wNDiag_26[18] , \wNDiag_26[17] , \wNDiag_26[16] , \wNDiag_26[15] , 
        \wNDiag_26[14] , \wNDiag_26[13] , \wNDiag_26[12] , \wNDiag_26[11] , 
        \wNDiag_26[10] , \wNDiag_26[9] , \wNDiag_26[8] , \wNDiag_26[7] , 
        \wNDiag_26[6] , \wNDiag_26[5] , \wNDiag_26[4] , \wNDiag_26[3] , 
        \wNDiag_26[2] , \wNDiag_26[1] , \wNDiag_26[0] }), .CallOut(
        \wCall_27[0] ), .ReturnOut(\wReturn_26[0] ), .ColOut({\wColumn_27[31] , 
        \wColumn_27[30] , \wColumn_27[29] , \wColumn_27[28] , \wColumn_27[27] , 
        \wColumn_27[26] , \wColumn_27[25] , \wColumn_27[24] , \wColumn_27[23] , 
        \wColumn_27[22] , \wColumn_27[21] , \wColumn_27[20] , \wColumn_27[19] , 
        \wColumn_27[18] , \wColumn_27[17] , \wColumn_27[16] , \wColumn_27[15] , 
        \wColumn_27[14] , \wColumn_27[13] , \wColumn_27[12] , \wColumn_27[11] , 
        \wColumn_27[10] , \wColumn_27[9] , \wColumn_27[8] , \wColumn_27[7] , 
        \wColumn_27[6] , \wColumn_27[5] , \wColumn_27[4] , \wColumn_27[3] , 
        \wColumn_27[2] , \wColumn_27[1] , \wColumn_27[0] }), .PDiagOut({
        \wPDiag_27[31] , \wPDiag_27[30] , \wPDiag_27[29] , \wPDiag_27[28] , 
        \wPDiag_27[27] , \wPDiag_27[26] , \wPDiag_27[25] , \wPDiag_27[24] , 
        \wPDiag_27[23] , \wPDiag_27[22] , \wPDiag_27[21] , \wPDiag_27[20] , 
        \wPDiag_27[19] , \wPDiag_27[18] , \wPDiag_27[17] , \wPDiag_27[16] , 
        \wPDiag_27[15] , \wPDiag_27[14] , \wPDiag_27[13] , \wPDiag_27[12] , 
        \wPDiag_27[11] , \wPDiag_27[10] , \wPDiag_27[9] , \wPDiag_27[8] , 
        \wPDiag_27[7] , \wPDiag_27[6] , \wPDiag_27[5] , \wPDiag_27[4] , 
        \wPDiag_27[3] , \wPDiag_27[2] , \wPDiag_27[1] , \wPDiag_27[0] }), 
        .NDiagOut({\wNDiag_27[31] , \wNDiag_27[30] , \wNDiag_27[29] , 
        \wNDiag_27[28] , \wNDiag_27[27] , \wNDiag_27[26] , \wNDiag_27[25] , 
        \wNDiag_27[24] , \wNDiag_27[23] , \wNDiag_27[22] , \wNDiag_27[21] , 
        \wNDiag_27[20] , \wNDiag_27[19] , \wNDiag_27[18] , \wNDiag_27[17] , 
        \wNDiag_27[16] , \wNDiag_27[15] , \wNDiag_27[14] , \wNDiag_27[13] , 
        \wNDiag_27[12] , \wNDiag_27[11] , \wNDiag_27[10] , \wNDiag_27[9] , 
        \wNDiag_27[8] , \wNDiag_27[7] , \wNDiag_27[6] , \wNDiag_27[5] , 
        \wNDiag_27[4] , \wNDiag_27[3] , \wNDiag_27[2] , \wNDiag_27[1] , 
        \wNDiag_27[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_11 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_12[5] , \wScan_12[4] , \wScan_12[3] , 
        \wScan_12[2] , \wScan_12[1] , \wScan_12[0] }), .ScanOut({\wScan_11[5] , 
        \wScan_11[4] , \wScan_11[3] , \wScan_11[2] , \wScan_11[1] , 
        \wScan_11[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_11[0] ), .ReturnIn(\wReturn_12[0] ), 
        .ColIn({\wColumn_11[31] , \wColumn_11[30] , \wColumn_11[29] , 
        \wColumn_11[28] , \wColumn_11[27] , \wColumn_11[26] , \wColumn_11[25] , 
        \wColumn_11[24] , \wColumn_11[23] , \wColumn_11[22] , \wColumn_11[21] , 
        \wColumn_11[20] , \wColumn_11[19] , \wColumn_11[18] , \wColumn_11[17] , 
        \wColumn_11[16] , \wColumn_11[15] , \wColumn_11[14] , \wColumn_11[13] , 
        \wColumn_11[12] , \wColumn_11[11] , \wColumn_11[10] , \wColumn_11[9] , 
        \wColumn_11[8] , \wColumn_11[7] , \wColumn_11[6] , \wColumn_11[5] , 
        \wColumn_11[4] , \wColumn_11[3] , \wColumn_11[2] , \wColumn_11[1] , 
        \wColumn_11[0] }), .PDiagIn({\wPDiag_11[31] , \wPDiag_11[30] , 
        \wPDiag_11[29] , \wPDiag_11[28] , \wPDiag_11[27] , \wPDiag_11[26] , 
        \wPDiag_11[25] , \wPDiag_11[24] , \wPDiag_11[23] , \wPDiag_11[22] , 
        \wPDiag_11[21] , \wPDiag_11[20] , \wPDiag_11[19] , \wPDiag_11[18] , 
        \wPDiag_11[17] , \wPDiag_11[16] , \wPDiag_11[15] , \wPDiag_11[14] , 
        \wPDiag_11[13] , \wPDiag_11[12] , \wPDiag_11[11] , \wPDiag_11[10] , 
        \wPDiag_11[9] , \wPDiag_11[8] , \wPDiag_11[7] , \wPDiag_11[6] , 
        \wPDiag_11[5] , \wPDiag_11[4] , \wPDiag_11[3] , \wPDiag_11[2] , 
        \wPDiag_11[1] , \wPDiag_11[0] }), .NDiagIn({\wNDiag_11[31] , 
        \wNDiag_11[30] , \wNDiag_11[29] , \wNDiag_11[28] , \wNDiag_11[27] , 
        \wNDiag_11[26] , \wNDiag_11[25] , \wNDiag_11[24] , \wNDiag_11[23] , 
        \wNDiag_11[22] , \wNDiag_11[21] , \wNDiag_11[20] , \wNDiag_11[19] , 
        \wNDiag_11[18] , \wNDiag_11[17] , \wNDiag_11[16] , \wNDiag_11[15] , 
        \wNDiag_11[14] , \wNDiag_11[13] , \wNDiag_11[12] , \wNDiag_11[11] , 
        \wNDiag_11[10] , \wNDiag_11[9] , \wNDiag_11[8] , \wNDiag_11[7] , 
        \wNDiag_11[6] , \wNDiag_11[5] , \wNDiag_11[4] , \wNDiag_11[3] , 
        \wNDiag_11[2] , \wNDiag_11[1] , \wNDiag_11[0] }), .CallOut(
        \wCall_12[0] ), .ReturnOut(\wReturn_11[0] ), .ColOut({\wColumn_12[31] , 
        \wColumn_12[30] , \wColumn_12[29] , \wColumn_12[28] , \wColumn_12[27] , 
        \wColumn_12[26] , \wColumn_12[25] , \wColumn_12[24] , \wColumn_12[23] , 
        \wColumn_12[22] , \wColumn_12[21] , \wColumn_12[20] , \wColumn_12[19] , 
        \wColumn_12[18] , \wColumn_12[17] , \wColumn_12[16] , \wColumn_12[15] , 
        \wColumn_12[14] , \wColumn_12[13] , \wColumn_12[12] , \wColumn_12[11] , 
        \wColumn_12[10] , \wColumn_12[9] , \wColumn_12[8] , \wColumn_12[7] , 
        \wColumn_12[6] , \wColumn_12[5] , \wColumn_12[4] , \wColumn_12[3] , 
        \wColumn_12[2] , \wColumn_12[1] , \wColumn_12[0] }), .PDiagOut({
        \wPDiag_12[31] , \wPDiag_12[30] , \wPDiag_12[29] , \wPDiag_12[28] , 
        \wPDiag_12[27] , \wPDiag_12[26] , \wPDiag_12[25] , \wPDiag_12[24] , 
        \wPDiag_12[23] , \wPDiag_12[22] , \wPDiag_12[21] , \wPDiag_12[20] , 
        \wPDiag_12[19] , \wPDiag_12[18] , \wPDiag_12[17] , \wPDiag_12[16] , 
        \wPDiag_12[15] , \wPDiag_12[14] , \wPDiag_12[13] , \wPDiag_12[12] , 
        \wPDiag_12[11] , \wPDiag_12[10] , \wPDiag_12[9] , \wPDiag_12[8] , 
        \wPDiag_12[7] , \wPDiag_12[6] , \wPDiag_12[5] , \wPDiag_12[4] , 
        \wPDiag_12[3] , \wPDiag_12[2] , \wPDiag_12[1] , \wPDiag_12[0] }), 
        .NDiagOut({\wNDiag_12[31] , \wNDiag_12[30] , \wNDiag_12[29] , 
        \wNDiag_12[28] , \wNDiag_12[27] , \wNDiag_12[26] , \wNDiag_12[25] , 
        \wNDiag_12[24] , \wNDiag_12[23] , \wNDiag_12[22] , \wNDiag_12[21] , 
        \wNDiag_12[20] , \wNDiag_12[19] , \wNDiag_12[18] , \wNDiag_12[17] , 
        \wNDiag_12[16] , \wNDiag_12[15] , \wNDiag_12[14] , \wNDiag_12[13] , 
        \wNDiag_12[12] , \wNDiag_12[11] , \wNDiag_12[10] , \wNDiag_12[9] , 
        \wNDiag_12[8] , \wNDiag_12[7] , \wNDiag_12[6] , \wNDiag_12[5] , 
        \wNDiag_12[4] , \wNDiag_12[3] , \wNDiag_12[2] , \wNDiag_12[1] , 
        \wNDiag_12[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_24 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_25[5] , \wScan_25[4] , \wScan_25[3] , 
        \wScan_25[2] , \wScan_25[1] , \wScan_25[0] }), .ScanOut({\wScan_24[5] , 
        \wScan_24[4] , \wScan_24[3] , \wScan_24[2] , \wScan_24[1] , 
        \wScan_24[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_24[0] ), .ReturnIn(\wReturn_25[0] ), 
        .ColIn({\wColumn_24[31] , \wColumn_24[30] , \wColumn_24[29] , 
        \wColumn_24[28] , \wColumn_24[27] , \wColumn_24[26] , \wColumn_24[25] , 
        \wColumn_24[24] , \wColumn_24[23] , \wColumn_24[22] , \wColumn_24[21] , 
        \wColumn_24[20] , \wColumn_24[19] , \wColumn_24[18] , \wColumn_24[17] , 
        \wColumn_24[16] , \wColumn_24[15] , \wColumn_24[14] , \wColumn_24[13] , 
        \wColumn_24[12] , \wColumn_24[11] , \wColumn_24[10] , \wColumn_24[9] , 
        \wColumn_24[8] , \wColumn_24[7] , \wColumn_24[6] , \wColumn_24[5] , 
        \wColumn_24[4] , \wColumn_24[3] , \wColumn_24[2] , \wColumn_24[1] , 
        \wColumn_24[0] }), .PDiagIn({\wPDiag_24[31] , \wPDiag_24[30] , 
        \wPDiag_24[29] , \wPDiag_24[28] , \wPDiag_24[27] , \wPDiag_24[26] , 
        \wPDiag_24[25] , \wPDiag_24[24] , \wPDiag_24[23] , \wPDiag_24[22] , 
        \wPDiag_24[21] , \wPDiag_24[20] , \wPDiag_24[19] , \wPDiag_24[18] , 
        \wPDiag_24[17] , \wPDiag_24[16] , \wPDiag_24[15] , \wPDiag_24[14] , 
        \wPDiag_24[13] , \wPDiag_24[12] , \wPDiag_24[11] , \wPDiag_24[10] , 
        \wPDiag_24[9] , \wPDiag_24[8] , \wPDiag_24[7] , \wPDiag_24[6] , 
        \wPDiag_24[5] , \wPDiag_24[4] , \wPDiag_24[3] , \wPDiag_24[2] , 
        \wPDiag_24[1] , \wPDiag_24[0] }), .NDiagIn({\wNDiag_24[31] , 
        \wNDiag_24[30] , \wNDiag_24[29] , \wNDiag_24[28] , \wNDiag_24[27] , 
        \wNDiag_24[26] , \wNDiag_24[25] , \wNDiag_24[24] , \wNDiag_24[23] , 
        \wNDiag_24[22] , \wNDiag_24[21] , \wNDiag_24[20] , \wNDiag_24[19] , 
        \wNDiag_24[18] , \wNDiag_24[17] , \wNDiag_24[16] , \wNDiag_24[15] , 
        \wNDiag_24[14] , \wNDiag_24[13] , \wNDiag_24[12] , \wNDiag_24[11] , 
        \wNDiag_24[10] , \wNDiag_24[9] , \wNDiag_24[8] , \wNDiag_24[7] , 
        \wNDiag_24[6] , \wNDiag_24[5] , \wNDiag_24[4] , \wNDiag_24[3] , 
        \wNDiag_24[2] , \wNDiag_24[1] , \wNDiag_24[0] }), .CallOut(
        \wCall_25[0] ), .ReturnOut(\wReturn_24[0] ), .ColOut({\wColumn_25[31] , 
        \wColumn_25[30] , \wColumn_25[29] , \wColumn_25[28] , \wColumn_25[27] , 
        \wColumn_25[26] , \wColumn_25[25] , \wColumn_25[24] , \wColumn_25[23] , 
        \wColumn_25[22] , \wColumn_25[21] , \wColumn_25[20] , \wColumn_25[19] , 
        \wColumn_25[18] , \wColumn_25[17] , \wColumn_25[16] , \wColumn_25[15] , 
        \wColumn_25[14] , \wColumn_25[13] , \wColumn_25[12] , \wColumn_25[11] , 
        \wColumn_25[10] , \wColumn_25[9] , \wColumn_25[8] , \wColumn_25[7] , 
        \wColumn_25[6] , \wColumn_25[5] , \wColumn_25[4] , \wColumn_25[3] , 
        \wColumn_25[2] , \wColumn_25[1] , \wColumn_25[0] }), .PDiagOut({
        \wPDiag_25[31] , \wPDiag_25[30] , \wPDiag_25[29] , \wPDiag_25[28] , 
        \wPDiag_25[27] , \wPDiag_25[26] , \wPDiag_25[25] , \wPDiag_25[24] , 
        \wPDiag_25[23] , \wPDiag_25[22] , \wPDiag_25[21] , \wPDiag_25[20] , 
        \wPDiag_25[19] , \wPDiag_25[18] , \wPDiag_25[17] , \wPDiag_25[16] , 
        \wPDiag_25[15] , \wPDiag_25[14] , \wPDiag_25[13] , \wPDiag_25[12] , 
        \wPDiag_25[11] , \wPDiag_25[10] , \wPDiag_25[9] , \wPDiag_25[8] , 
        \wPDiag_25[7] , \wPDiag_25[6] , \wPDiag_25[5] , \wPDiag_25[4] , 
        \wPDiag_25[3] , \wPDiag_25[2] , \wPDiag_25[1] , \wPDiag_25[0] }), 
        .NDiagOut({\wNDiag_25[31] , \wNDiag_25[30] , \wNDiag_25[29] , 
        \wNDiag_25[28] , \wNDiag_25[27] , \wNDiag_25[26] , \wNDiag_25[25] , 
        \wNDiag_25[24] , \wNDiag_25[23] , \wNDiag_25[22] , \wNDiag_25[21] , 
        \wNDiag_25[20] , \wNDiag_25[19] , \wNDiag_25[18] , \wNDiag_25[17] , 
        \wNDiag_25[16] , \wNDiag_25[15] , \wNDiag_25[14] , \wNDiag_25[13] , 
        \wNDiag_25[12] , \wNDiag_25[11] , \wNDiag_25[10] , \wNDiag_25[9] , 
        \wNDiag_25[8] , \wNDiag_25[7] , \wNDiag_25[6] , \wNDiag_25[5] , 
        \wNDiag_25[4] , \wNDiag_25[3] , \wNDiag_25[2] , \wNDiag_25[1] , 
        \wNDiag_25[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_1 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_2[5] , \wScan_2[4] , \wScan_2[3] , 
        \wScan_2[2] , \wScan_2[1] , \wScan_2[0] }), .ScanOut({\wScan_1[5] , 
        \wScan_1[4] , \wScan_1[3] , \wScan_1[2] , \wScan_1[1] , \wScan_1[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_1[0] ), .ReturnIn(\wReturn_2[0] ), .ColIn({
        \wColumn_1[31] , \wColumn_1[30] , \wColumn_1[29] , \wColumn_1[28] , 
        \wColumn_1[27] , \wColumn_1[26] , \wColumn_1[25] , \wColumn_1[24] , 
        \wColumn_1[23] , \wColumn_1[22] , \wColumn_1[21] , \wColumn_1[20] , 
        \wColumn_1[19] , \wColumn_1[18] , \wColumn_1[17] , \wColumn_1[16] , 
        \wColumn_1[15] , \wColumn_1[14] , \wColumn_1[13] , \wColumn_1[12] , 
        \wColumn_1[11] , \wColumn_1[10] , \wColumn_1[9] , \wColumn_1[8] , 
        \wColumn_1[7] , \wColumn_1[6] , \wColumn_1[5] , \wColumn_1[4] , 
        \wColumn_1[3] , \wColumn_1[2] , \wColumn_1[1] , \wColumn_1[0] }), 
        .PDiagIn({\wPDiag_1[31] , \wPDiag_1[30] , \wPDiag_1[29] , 
        \wPDiag_1[28] , \wPDiag_1[27] , \wPDiag_1[26] , \wPDiag_1[25] , 
        \wPDiag_1[24] , \wPDiag_1[23] , \wPDiag_1[22] , \wPDiag_1[21] , 
        \wPDiag_1[20] , \wPDiag_1[19] , \wPDiag_1[18] , \wPDiag_1[17] , 
        \wPDiag_1[16] , \wPDiag_1[15] , \wPDiag_1[14] , \wPDiag_1[13] , 
        \wPDiag_1[12] , \wPDiag_1[11] , \wPDiag_1[10] , \wPDiag_1[9] , 
        \wPDiag_1[8] , \wPDiag_1[7] , \wPDiag_1[6] , \wPDiag_1[5] , 
        \wPDiag_1[4] , \wPDiag_1[3] , \wPDiag_1[2] , \wPDiag_1[1] , 
        \wPDiag_1[0] }), .NDiagIn({\wNDiag_1[31] , \wNDiag_1[30] , 
        \wNDiag_1[29] , \wNDiag_1[28] , \wNDiag_1[27] , \wNDiag_1[26] , 
        \wNDiag_1[25] , \wNDiag_1[24] , \wNDiag_1[23] , \wNDiag_1[22] , 
        \wNDiag_1[21] , \wNDiag_1[20] , \wNDiag_1[19] , \wNDiag_1[18] , 
        \wNDiag_1[17] , \wNDiag_1[16] , \wNDiag_1[15] , \wNDiag_1[14] , 
        \wNDiag_1[13] , \wNDiag_1[12] , \wNDiag_1[11] , \wNDiag_1[10] , 
        \wNDiag_1[9] , \wNDiag_1[8] , \wNDiag_1[7] , \wNDiag_1[6] , 
        \wNDiag_1[5] , \wNDiag_1[4] , \wNDiag_1[3] , \wNDiag_1[2] , 
        \wNDiag_1[1] , \wNDiag_1[0] }), .CallOut(\wCall_2[0] ), .ReturnOut(
        \wReturn_1[0] ), .ColOut({\wColumn_2[31] , \wColumn_2[30] , 
        \wColumn_2[29] , \wColumn_2[28] , \wColumn_2[27] , \wColumn_2[26] , 
        \wColumn_2[25] , \wColumn_2[24] , \wColumn_2[23] , \wColumn_2[22] , 
        \wColumn_2[21] , \wColumn_2[20] , \wColumn_2[19] , \wColumn_2[18] , 
        \wColumn_2[17] , \wColumn_2[16] , \wColumn_2[15] , \wColumn_2[14] , 
        \wColumn_2[13] , \wColumn_2[12] , \wColumn_2[11] , \wColumn_2[10] , 
        \wColumn_2[9] , \wColumn_2[8] , \wColumn_2[7] , \wColumn_2[6] , 
        \wColumn_2[5] , \wColumn_2[4] , \wColumn_2[3] , \wColumn_2[2] , 
        \wColumn_2[1] , \wColumn_2[0] }), .PDiagOut({\wPDiag_2[31] , 
        \wPDiag_2[30] , \wPDiag_2[29] , \wPDiag_2[28] , \wPDiag_2[27] , 
        \wPDiag_2[26] , \wPDiag_2[25] , \wPDiag_2[24] , \wPDiag_2[23] , 
        \wPDiag_2[22] , \wPDiag_2[21] , \wPDiag_2[20] , \wPDiag_2[19] , 
        \wPDiag_2[18] , \wPDiag_2[17] , \wPDiag_2[16] , \wPDiag_2[15] , 
        \wPDiag_2[14] , \wPDiag_2[13] , \wPDiag_2[12] , \wPDiag_2[11] , 
        \wPDiag_2[10] , \wPDiag_2[9] , \wPDiag_2[8] , \wPDiag_2[7] , 
        \wPDiag_2[6] , \wPDiag_2[5] , \wPDiag_2[4] , \wPDiag_2[3] , 
        \wPDiag_2[2] , \wPDiag_2[1] , \wPDiag_2[0] }), .NDiagOut({
        \wNDiag_2[31] , \wNDiag_2[30] , \wNDiag_2[29] , \wNDiag_2[28] , 
        \wNDiag_2[27] , \wNDiag_2[26] , \wNDiag_2[25] , \wNDiag_2[24] , 
        \wNDiag_2[23] , \wNDiag_2[22] , \wNDiag_2[21] , \wNDiag_2[20] , 
        \wNDiag_2[19] , \wNDiag_2[18] , \wNDiag_2[17] , \wNDiag_2[16] , 
        \wNDiag_2[15] , \wNDiag_2[14] , \wNDiag_2[13] , \wNDiag_2[12] , 
        \wNDiag_2[11] , \wNDiag_2[10] , \wNDiag_2[9] , \wNDiag_2[8] , 
        \wNDiag_2[7] , \wNDiag_2[6] , \wNDiag_2[5] , \wNDiag_2[4] , 
        \wNDiag_2[3] , \wNDiag_2[2] , \wNDiag_2[1] , \wNDiag_2[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_6 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_7[5] , \wScan_7[4] , \wScan_7[3] , 
        \wScan_7[2] , \wScan_7[1] , \wScan_7[0] }), .ScanOut({\wScan_6[5] , 
        \wScan_6[4] , \wScan_6[3] , \wScan_6[2] , \wScan_6[1] , \wScan_6[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_6[0] ), .ReturnIn(\wReturn_7[0] ), .ColIn({
        \wColumn_6[31] , \wColumn_6[30] , \wColumn_6[29] , \wColumn_6[28] , 
        \wColumn_6[27] , \wColumn_6[26] , \wColumn_6[25] , \wColumn_6[24] , 
        \wColumn_6[23] , \wColumn_6[22] , \wColumn_6[21] , \wColumn_6[20] , 
        \wColumn_6[19] , \wColumn_6[18] , \wColumn_6[17] , \wColumn_6[16] , 
        \wColumn_6[15] , \wColumn_6[14] , \wColumn_6[13] , \wColumn_6[12] , 
        \wColumn_6[11] , \wColumn_6[10] , \wColumn_6[9] , \wColumn_6[8] , 
        \wColumn_6[7] , \wColumn_6[6] , \wColumn_6[5] , \wColumn_6[4] , 
        \wColumn_6[3] , \wColumn_6[2] , \wColumn_6[1] , \wColumn_6[0] }), 
        .PDiagIn({\wPDiag_6[31] , \wPDiag_6[30] , \wPDiag_6[29] , 
        \wPDiag_6[28] , \wPDiag_6[27] , \wPDiag_6[26] , \wPDiag_6[25] , 
        \wPDiag_6[24] , \wPDiag_6[23] , \wPDiag_6[22] , \wPDiag_6[21] , 
        \wPDiag_6[20] , \wPDiag_6[19] , \wPDiag_6[18] , \wPDiag_6[17] , 
        \wPDiag_6[16] , \wPDiag_6[15] , \wPDiag_6[14] , \wPDiag_6[13] , 
        \wPDiag_6[12] , \wPDiag_6[11] , \wPDiag_6[10] , \wPDiag_6[9] , 
        \wPDiag_6[8] , \wPDiag_6[7] , \wPDiag_6[6] , \wPDiag_6[5] , 
        \wPDiag_6[4] , \wPDiag_6[3] , \wPDiag_6[2] , \wPDiag_6[1] , 
        \wPDiag_6[0] }), .NDiagIn({\wNDiag_6[31] , \wNDiag_6[30] , 
        \wNDiag_6[29] , \wNDiag_6[28] , \wNDiag_6[27] , \wNDiag_6[26] , 
        \wNDiag_6[25] , \wNDiag_6[24] , \wNDiag_6[23] , \wNDiag_6[22] , 
        \wNDiag_6[21] , \wNDiag_6[20] , \wNDiag_6[19] , \wNDiag_6[18] , 
        \wNDiag_6[17] , \wNDiag_6[16] , \wNDiag_6[15] , \wNDiag_6[14] , 
        \wNDiag_6[13] , \wNDiag_6[12] , \wNDiag_6[11] , \wNDiag_6[10] , 
        \wNDiag_6[9] , \wNDiag_6[8] , \wNDiag_6[7] , \wNDiag_6[6] , 
        \wNDiag_6[5] , \wNDiag_6[4] , \wNDiag_6[3] , \wNDiag_6[2] , 
        \wNDiag_6[1] , \wNDiag_6[0] }), .CallOut(\wCall_7[0] ), .ReturnOut(
        \wReturn_6[0] ), .ColOut({\wColumn_7[31] , \wColumn_7[30] , 
        \wColumn_7[29] , \wColumn_7[28] , \wColumn_7[27] , \wColumn_7[26] , 
        \wColumn_7[25] , \wColumn_7[24] , \wColumn_7[23] , \wColumn_7[22] , 
        \wColumn_7[21] , \wColumn_7[20] , \wColumn_7[19] , \wColumn_7[18] , 
        \wColumn_7[17] , \wColumn_7[16] , \wColumn_7[15] , \wColumn_7[14] , 
        \wColumn_7[13] , \wColumn_7[12] , \wColumn_7[11] , \wColumn_7[10] , 
        \wColumn_7[9] , \wColumn_7[8] , \wColumn_7[7] , \wColumn_7[6] , 
        \wColumn_7[5] , \wColumn_7[4] , \wColumn_7[3] , \wColumn_7[2] , 
        \wColumn_7[1] , \wColumn_7[0] }), .PDiagOut({\wPDiag_7[31] , 
        \wPDiag_7[30] , \wPDiag_7[29] , \wPDiag_7[28] , \wPDiag_7[27] , 
        \wPDiag_7[26] , \wPDiag_7[25] , \wPDiag_7[24] , \wPDiag_7[23] , 
        \wPDiag_7[22] , \wPDiag_7[21] , \wPDiag_7[20] , \wPDiag_7[19] , 
        \wPDiag_7[18] , \wPDiag_7[17] , \wPDiag_7[16] , \wPDiag_7[15] , 
        \wPDiag_7[14] , \wPDiag_7[13] , \wPDiag_7[12] , \wPDiag_7[11] , 
        \wPDiag_7[10] , \wPDiag_7[9] , \wPDiag_7[8] , \wPDiag_7[7] , 
        \wPDiag_7[6] , \wPDiag_7[5] , \wPDiag_7[4] , \wPDiag_7[3] , 
        \wPDiag_7[2] , \wPDiag_7[1] , \wPDiag_7[0] }), .NDiagOut({
        \wNDiag_7[31] , \wNDiag_7[30] , \wNDiag_7[29] , \wNDiag_7[28] , 
        \wNDiag_7[27] , \wNDiag_7[26] , \wNDiag_7[25] , \wNDiag_7[24] , 
        \wNDiag_7[23] , \wNDiag_7[22] , \wNDiag_7[21] , \wNDiag_7[20] , 
        \wNDiag_7[19] , \wNDiag_7[18] , \wNDiag_7[17] , \wNDiag_7[16] , 
        \wNDiag_7[15] , \wNDiag_7[14] , \wNDiag_7[13] , \wNDiag_7[12] , 
        \wNDiag_7[11] , \wNDiag_7[10] , \wNDiag_7[9] , \wNDiag_7[8] , 
        \wNDiag_7[7] , \wNDiag_7[6] , \wNDiag_7[5] , \wNDiag_7[4] , 
        \wNDiag_7[3] , \wNDiag_7[2] , \wNDiag_7[1] , \wNDiag_7[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_7 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_8[5] , \wScan_8[4] , \wScan_8[3] , 
        \wScan_8[2] , \wScan_8[1] , \wScan_8[0] }), .ScanOut({\wScan_7[5] , 
        \wScan_7[4] , \wScan_7[3] , \wScan_7[2] , \wScan_7[1] , \wScan_7[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_7[0] ), .ReturnIn(\wReturn_8[0] ), .ColIn({
        \wColumn_7[31] , \wColumn_7[30] , \wColumn_7[29] , \wColumn_7[28] , 
        \wColumn_7[27] , \wColumn_7[26] , \wColumn_7[25] , \wColumn_7[24] , 
        \wColumn_7[23] , \wColumn_7[22] , \wColumn_7[21] , \wColumn_7[20] , 
        \wColumn_7[19] , \wColumn_7[18] , \wColumn_7[17] , \wColumn_7[16] , 
        \wColumn_7[15] , \wColumn_7[14] , \wColumn_7[13] , \wColumn_7[12] , 
        \wColumn_7[11] , \wColumn_7[10] , \wColumn_7[9] , \wColumn_7[8] , 
        \wColumn_7[7] , \wColumn_7[6] , \wColumn_7[5] , \wColumn_7[4] , 
        \wColumn_7[3] , \wColumn_7[2] , \wColumn_7[1] , \wColumn_7[0] }), 
        .PDiagIn({\wPDiag_7[31] , \wPDiag_7[30] , \wPDiag_7[29] , 
        \wPDiag_7[28] , \wPDiag_7[27] , \wPDiag_7[26] , \wPDiag_7[25] , 
        \wPDiag_7[24] , \wPDiag_7[23] , \wPDiag_7[22] , \wPDiag_7[21] , 
        \wPDiag_7[20] , \wPDiag_7[19] , \wPDiag_7[18] , \wPDiag_7[17] , 
        \wPDiag_7[16] , \wPDiag_7[15] , \wPDiag_7[14] , \wPDiag_7[13] , 
        \wPDiag_7[12] , \wPDiag_7[11] , \wPDiag_7[10] , \wPDiag_7[9] , 
        \wPDiag_7[8] , \wPDiag_7[7] , \wPDiag_7[6] , \wPDiag_7[5] , 
        \wPDiag_7[4] , \wPDiag_7[3] , \wPDiag_7[2] , \wPDiag_7[1] , 
        \wPDiag_7[0] }), .NDiagIn({\wNDiag_7[31] , \wNDiag_7[30] , 
        \wNDiag_7[29] , \wNDiag_7[28] , \wNDiag_7[27] , \wNDiag_7[26] , 
        \wNDiag_7[25] , \wNDiag_7[24] , \wNDiag_7[23] , \wNDiag_7[22] , 
        \wNDiag_7[21] , \wNDiag_7[20] , \wNDiag_7[19] , \wNDiag_7[18] , 
        \wNDiag_7[17] , \wNDiag_7[16] , \wNDiag_7[15] , \wNDiag_7[14] , 
        \wNDiag_7[13] , \wNDiag_7[12] , \wNDiag_7[11] , \wNDiag_7[10] , 
        \wNDiag_7[9] , \wNDiag_7[8] , \wNDiag_7[7] , \wNDiag_7[6] , 
        \wNDiag_7[5] , \wNDiag_7[4] , \wNDiag_7[3] , \wNDiag_7[2] , 
        \wNDiag_7[1] , \wNDiag_7[0] }), .CallOut(\wCall_8[0] ), .ReturnOut(
        \wReturn_7[0] ), .ColOut({\wColumn_8[31] , \wColumn_8[30] , 
        \wColumn_8[29] , \wColumn_8[28] , \wColumn_8[27] , \wColumn_8[26] , 
        \wColumn_8[25] , \wColumn_8[24] , \wColumn_8[23] , \wColumn_8[22] , 
        \wColumn_8[21] , \wColumn_8[20] , \wColumn_8[19] , \wColumn_8[18] , 
        \wColumn_8[17] , \wColumn_8[16] , \wColumn_8[15] , \wColumn_8[14] , 
        \wColumn_8[13] , \wColumn_8[12] , \wColumn_8[11] , \wColumn_8[10] , 
        \wColumn_8[9] , \wColumn_8[8] , \wColumn_8[7] , \wColumn_8[6] , 
        \wColumn_8[5] , \wColumn_8[4] , \wColumn_8[3] , \wColumn_8[2] , 
        \wColumn_8[1] , \wColumn_8[0] }), .PDiagOut({\wPDiag_8[31] , 
        \wPDiag_8[30] , \wPDiag_8[29] , \wPDiag_8[28] , \wPDiag_8[27] , 
        \wPDiag_8[26] , \wPDiag_8[25] , \wPDiag_8[24] , \wPDiag_8[23] , 
        \wPDiag_8[22] , \wPDiag_8[21] , \wPDiag_8[20] , \wPDiag_8[19] , 
        \wPDiag_8[18] , \wPDiag_8[17] , \wPDiag_8[16] , \wPDiag_8[15] , 
        \wPDiag_8[14] , \wPDiag_8[13] , \wPDiag_8[12] , \wPDiag_8[11] , 
        \wPDiag_8[10] , \wPDiag_8[9] , \wPDiag_8[8] , \wPDiag_8[7] , 
        \wPDiag_8[6] , \wPDiag_8[5] , \wPDiag_8[4] , \wPDiag_8[3] , 
        \wPDiag_8[2] , \wPDiag_8[1] , \wPDiag_8[0] }), .NDiagOut({
        \wNDiag_8[31] , \wNDiag_8[30] , \wNDiag_8[29] , \wNDiag_8[28] , 
        \wNDiag_8[27] , \wNDiag_8[26] , \wNDiag_8[25] , \wNDiag_8[24] , 
        \wNDiag_8[23] , \wNDiag_8[22] , \wNDiag_8[21] , \wNDiag_8[20] , 
        \wNDiag_8[19] , \wNDiag_8[18] , \wNDiag_8[17] , \wNDiag_8[16] , 
        \wNDiag_8[15] , \wNDiag_8[14] , \wNDiag_8[13] , \wNDiag_8[12] , 
        \wNDiag_8[11] , \wNDiag_8[10] , \wNDiag_8[9] , \wNDiag_8[8] , 
        \wNDiag_8[7] , \wNDiag_8[6] , \wNDiag_8[5] , \wNDiag_8[4] , 
        \wNDiag_8[3] , \wNDiag_8[2] , \wNDiag_8[1] , \wNDiag_8[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_18 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_19[5] , \wScan_19[4] , \wScan_19[3] , 
        \wScan_19[2] , \wScan_19[1] , \wScan_19[0] }), .ScanOut({\wScan_18[5] , 
        \wScan_18[4] , \wScan_18[3] , \wScan_18[2] , \wScan_18[1] , 
        \wScan_18[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_18[0] ), .ReturnIn(\wReturn_19[0] ), 
        .ColIn({\wColumn_18[31] , \wColumn_18[30] , \wColumn_18[29] , 
        \wColumn_18[28] , \wColumn_18[27] , \wColumn_18[26] , \wColumn_18[25] , 
        \wColumn_18[24] , \wColumn_18[23] , \wColumn_18[22] , \wColumn_18[21] , 
        \wColumn_18[20] , \wColumn_18[19] , \wColumn_18[18] , \wColumn_18[17] , 
        \wColumn_18[16] , \wColumn_18[15] , \wColumn_18[14] , \wColumn_18[13] , 
        \wColumn_18[12] , \wColumn_18[11] , \wColumn_18[10] , \wColumn_18[9] , 
        \wColumn_18[8] , \wColumn_18[7] , \wColumn_18[6] , \wColumn_18[5] , 
        \wColumn_18[4] , \wColumn_18[3] , \wColumn_18[2] , \wColumn_18[1] , 
        \wColumn_18[0] }), .PDiagIn({\wPDiag_18[31] , \wPDiag_18[30] , 
        \wPDiag_18[29] , \wPDiag_18[28] , \wPDiag_18[27] , \wPDiag_18[26] , 
        \wPDiag_18[25] , \wPDiag_18[24] , \wPDiag_18[23] , \wPDiag_18[22] , 
        \wPDiag_18[21] , \wPDiag_18[20] , \wPDiag_18[19] , \wPDiag_18[18] , 
        \wPDiag_18[17] , \wPDiag_18[16] , \wPDiag_18[15] , \wPDiag_18[14] , 
        \wPDiag_18[13] , \wPDiag_18[12] , \wPDiag_18[11] , \wPDiag_18[10] , 
        \wPDiag_18[9] , \wPDiag_18[8] , \wPDiag_18[7] , \wPDiag_18[6] , 
        \wPDiag_18[5] , \wPDiag_18[4] , \wPDiag_18[3] , \wPDiag_18[2] , 
        \wPDiag_18[1] , \wPDiag_18[0] }), .NDiagIn({\wNDiag_18[31] , 
        \wNDiag_18[30] , \wNDiag_18[29] , \wNDiag_18[28] , \wNDiag_18[27] , 
        \wNDiag_18[26] , \wNDiag_18[25] , \wNDiag_18[24] , \wNDiag_18[23] , 
        \wNDiag_18[22] , \wNDiag_18[21] , \wNDiag_18[20] , \wNDiag_18[19] , 
        \wNDiag_18[18] , \wNDiag_18[17] , \wNDiag_18[16] , \wNDiag_18[15] , 
        \wNDiag_18[14] , \wNDiag_18[13] , \wNDiag_18[12] , \wNDiag_18[11] , 
        \wNDiag_18[10] , \wNDiag_18[9] , \wNDiag_18[8] , \wNDiag_18[7] , 
        \wNDiag_18[6] , \wNDiag_18[5] , \wNDiag_18[4] , \wNDiag_18[3] , 
        \wNDiag_18[2] , \wNDiag_18[1] , \wNDiag_18[0] }), .CallOut(
        \wCall_19[0] ), .ReturnOut(\wReturn_18[0] ), .ColOut({\wColumn_19[31] , 
        \wColumn_19[30] , \wColumn_19[29] , \wColumn_19[28] , \wColumn_19[27] , 
        \wColumn_19[26] , \wColumn_19[25] , \wColumn_19[24] , \wColumn_19[23] , 
        \wColumn_19[22] , \wColumn_19[21] , \wColumn_19[20] , \wColumn_19[19] , 
        \wColumn_19[18] , \wColumn_19[17] , \wColumn_19[16] , \wColumn_19[15] , 
        \wColumn_19[14] , \wColumn_19[13] , \wColumn_19[12] , \wColumn_19[11] , 
        \wColumn_19[10] , \wColumn_19[9] , \wColumn_19[8] , \wColumn_19[7] , 
        \wColumn_19[6] , \wColumn_19[5] , \wColumn_19[4] , \wColumn_19[3] , 
        \wColumn_19[2] , \wColumn_19[1] , \wColumn_19[0] }), .PDiagOut({
        \wPDiag_19[31] , \wPDiag_19[30] , \wPDiag_19[29] , \wPDiag_19[28] , 
        \wPDiag_19[27] , \wPDiag_19[26] , \wPDiag_19[25] , \wPDiag_19[24] , 
        \wPDiag_19[23] , \wPDiag_19[22] , \wPDiag_19[21] , \wPDiag_19[20] , 
        \wPDiag_19[19] , \wPDiag_19[18] , \wPDiag_19[17] , \wPDiag_19[16] , 
        \wPDiag_19[15] , \wPDiag_19[14] , \wPDiag_19[13] , \wPDiag_19[12] , 
        \wPDiag_19[11] , \wPDiag_19[10] , \wPDiag_19[9] , \wPDiag_19[8] , 
        \wPDiag_19[7] , \wPDiag_19[6] , \wPDiag_19[5] , \wPDiag_19[4] , 
        \wPDiag_19[3] , \wPDiag_19[2] , \wPDiag_19[1] , \wPDiag_19[0] }), 
        .NDiagOut({\wNDiag_19[31] , \wNDiag_19[30] , \wNDiag_19[29] , 
        \wNDiag_19[28] , \wNDiag_19[27] , \wNDiag_19[26] , \wNDiag_19[25] , 
        \wNDiag_19[24] , \wNDiag_19[23] , \wNDiag_19[22] , \wNDiag_19[21] , 
        \wNDiag_19[20] , \wNDiag_19[19] , \wNDiag_19[18] , \wNDiag_19[17] , 
        \wNDiag_19[16] , \wNDiag_19[15] , \wNDiag_19[14] , \wNDiag_19[13] , 
        \wNDiag_19[12] , \wNDiag_19[11] , \wNDiag_19[10] , \wNDiag_19[9] , 
        \wNDiag_19[8] , \wNDiag_19[7] , \wNDiag_19[6] , \wNDiag_19[5] , 
        \wNDiag_19[4] , \wNDiag_19[3] , \wNDiag_19[2] , \wNDiag_19[1] , 
        \wNDiag_19[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_16 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_17[5] , \wScan_17[4] , \wScan_17[3] , 
        \wScan_17[2] , \wScan_17[1] , \wScan_17[0] }), .ScanOut({\wScan_16[5] , 
        \wScan_16[4] , \wScan_16[3] , \wScan_16[2] , \wScan_16[1] , 
        \wScan_16[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_16[0] ), .ReturnIn(\wReturn_17[0] ), 
        .ColIn({\wColumn_16[31] , \wColumn_16[30] , \wColumn_16[29] , 
        \wColumn_16[28] , \wColumn_16[27] , \wColumn_16[26] , \wColumn_16[25] , 
        \wColumn_16[24] , \wColumn_16[23] , \wColumn_16[22] , \wColumn_16[21] , 
        \wColumn_16[20] , \wColumn_16[19] , \wColumn_16[18] , \wColumn_16[17] , 
        \wColumn_16[16] , \wColumn_16[15] , \wColumn_16[14] , \wColumn_16[13] , 
        \wColumn_16[12] , \wColumn_16[11] , \wColumn_16[10] , \wColumn_16[9] , 
        \wColumn_16[8] , \wColumn_16[7] , \wColumn_16[6] , \wColumn_16[5] , 
        \wColumn_16[4] , \wColumn_16[3] , \wColumn_16[2] , \wColumn_16[1] , 
        \wColumn_16[0] }), .PDiagIn({\wPDiag_16[31] , \wPDiag_16[30] , 
        \wPDiag_16[29] , \wPDiag_16[28] , \wPDiag_16[27] , \wPDiag_16[26] , 
        \wPDiag_16[25] , \wPDiag_16[24] , \wPDiag_16[23] , \wPDiag_16[22] , 
        \wPDiag_16[21] , \wPDiag_16[20] , \wPDiag_16[19] , \wPDiag_16[18] , 
        \wPDiag_16[17] , \wPDiag_16[16] , \wPDiag_16[15] , \wPDiag_16[14] , 
        \wPDiag_16[13] , \wPDiag_16[12] , \wPDiag_16[11] , \wPDiag_16[10] , 
        \wPDiag_16[9] , \wPDiag_16[8] , \wPDiag_16[7] , \wPDiag_16[6] , 
        \wPDiag_16[5] , \wPDiag_16[4] , \wPDiag_16[3] , \wPDiag_16[2] , 
        \wPDiag_16[1] , \wPDiag_16[0] }), .NDiagIn({\wNDiag_16[31] , 
        \wNDiag_16[30] , \wNDiag_16[29] , \wNDiag_16[28] , \wNDiag_16[27] , 
        \wNDiag_16[26] , \wNDiag_16[25] , \wNDiag_16[24] , \wNDiag_16[23] , 
        \wNDiag_16[22] , \wNDiag_16[21] , \wNDiag_16[20] , \wNDiag_16[19] , 
        \wNDiag_16[18] , \wNDiag_16[17] , \wNDiag_16[16] , \wNDiag_16[15] , 
        \wNDiag_16[14] , \wNDiag_16[13] , \wNDiag_16[12] , \wNDiag_16[11] , 
        \wNDiag_16[10] , \wNDiag_16[9] , \wNDiag_16[8] , \wNDiag_16[7] , 
        \wNDiag_16[6] , \wNDiag_16[5] , \wNDiag_16[4] , \wNDiag_16[3] , 
        \wNDiag_16[2] , \wNDiag_16[1] , \wNDiag_16[0] }), .CallOut(
        \wCall_17[0] ), .ReturnOut(\wReturn_16[0] ), .ColOut({\wColumn_17[31] , 
        \wColumn_17[30] , \wColumn_17[29] , \wColumn_17[28] , \wColumn_17[27] , 
        \wColumn_17[26] , \wColumn_17[25] , \wColumn_17[24] , \wColumn_17[23] , 
        \wColumn_17[22] , \wColumn_17[21] , \wColumn_17[20] , \wColumn_17[19] , 
        \wColumn_17[18] , \wColumn_17[17] , \wColumn_17[16] , \wColumn_17[15] , 
        \wColumn_17[14] , \wColumn_17[13] , \wColumn_17[12] , \wColumn_17[11] , 
        \wColumn_17[10] , \wColumn_17[9] , \wColumn_17[8] , \wColumn_17[7] , 
        \wColumn_17[6] , \wColumn_17[5] , \wColumn_17[4] , \wColumn_17[3] , 
        \wColumn_17[2] , \wColumn_17[1] , \wColumn_17[0] }), .PDiagOut({
        \wPDiag_17[31] , \wPDiag_17[30] , \wPDiag_17[29] , \wPDiag_17[28] , 
        \wPDiag_17[27] , \wPDiag_17[26] , \wPDiag_17[25] , \wPDiag_17[24] , 
        \wPDiag_17[23] , \wPDiag_17[22] , \wPDiag_17[21] , \wPDiag_17[20] , 
        \wPDiag_17[19] , \wPDiag_17[18] , \wPDiag_17[17] , \wPDiag_17[16] , 
        \wPDiag_17[15] , \wPDiag_17[14] , \wPDiag_17[13] , \wPDiag_17[12] , 
        \wPDiag_17[11] , \wPDiag_17[10] , \wPDiag_17[9] , \wPDiag_17[8] , 
        \wPDiag_17[7] , \wPDiag_17[6] , \wPDiag_17[5] , \wPDiag_17[4] , 
        \wPDiag_17[3] , \wPDiag_17[2] , \wPDiag_17[1] , \wPDiag_17[0] }), 
        .NDiagOut({\wNDiag_17[31] , \wNDiag_17[30] , \wNDiag_17[29] , 
        \wNDiag_17[28] , \wNDiag_17[27] , \wNDiag_17[26] , \wNDiag_17[25] , 
        \wNDiag_17[24] , \wNDiag_17[23] , \wNDiag_17[22] , \wNDiag_17[21] , 
        \wNDiag_17[20] , \wNDiag_17[19] , \wNDiag_17[18] , \wNDiag_17[17] , 
        \wNDiag_17[16] , \wNDiag_17[15] , \wNDiag_17[14] , \wNDiag_17[13] , 
        \wNDiag_17[12] , \wNDiag_17[11] , \wNDiag_17[10] , \wNDiag_17[9] , 
        \wNDiag_17[8] , \wNDiag_17[7] , \wNDiag_17[6] , \wNDiag_17[5] , 
        \wNDiag_17[4] , \wNDiag_17[3] , \wNDiag_17[2] , \wNDiag_17[1] , 
        \wNDiag_17[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_23 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_24[5] , \wScan_24[4] , \wScan_24[3] , 
        \wScan_24[2] , \wScan_24[1] , \wScan_24[0] }), .ScanOut({\wScan_23[5] , 
        \wScan_23[4] , \wScan_23[3] , \wScan_23[2] , \wScan_23[1] , 
        \wScan_23[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_23[0] ), .ReturnIn(\wReturn_24[0] ), 
        .ColIn({\wColumn_23[31] , \wColumn_23[30] , \wColumn_23[29] , 
        \wColumn_23[28] , \wColumn_23[27] , \wColumn_23[26] , \wColumn_23[25] , 
        \wColumn_23[24] , \wColumn_23[23] , \wColumn_23[22] , \wColumn_23[21] , 
        \wColumn_23[20] , \wColumn_23[19] , \wColumn_23[18] , \wColumn_23[17] , 
        \wColumn_23[16] , \wColumn_23[15] , \wColumn_23[14] , \wColumn_23[13] , 
        \wColumn_23[12] , \wColumn_23[11] , \wColumn_23[10] , \wColumn_23[9] , 
        \wColumn_23[8] , \wColumn_23[7] , \wColumn_23[6] , \wColumn_23[5] , 
        \wColumn_23[4] , \wColumn_23[3] , \wColumn_23[2] , \wColumn_23[1] , 
        \wColumn_23[0] }), .PDiagIn({\wPDiag_23[31] , \wPDiag_23[30] , 
        \wPDiag_23[29] , \wPDiag_23[28] , \wPDiag_23[27] , \wPDiag_23[26] , 
        \wPDiag_23[25] , \wPDiag_23[24] , \wPDiag_23[23] , \wPDiag_23[22] , 
        \wPDiag_23[21] , \wPDiag_23[20] , \wPDiag_23[19] , \wPDiag_23[18] , 
        \wPDiag_23[17] , \wPDiag_23[16] , \wPDiag_23[15] , \wPDiag_23[14] , 
        \wPDiag_23[13] , \wPDiag_23[12] , \wPDiag_23[11] , \wPDiag_23[10] , 
        \wPDiag_23[9] , \wPDiag_23[8] , \wPDiag_23[7] , \wPDiag_23[6] , 
        \wPDiag_23[5] , \wPDiag_23[4] , \wPDiag_23[3] , \wPDiag_23[2] , 
        \wPDiag_23[1] , \wPDiag_23[0] }), .NDiagIn({\wNDiag_23[31] , 
        \wNDiag_23[30] , \wNDiag_23[29] , \wNDiag_23[28] , \wNDiag_23[27] , 
        \wNDiag_23[26] , \wNDiag_23[25] , \wNDiag_23[24] , \wNDiag_23[23] , 
        \wNDiag_23[22] , \wNDiag_23[21] , \wNDiag_23[20] , \wNDiag_23[19] , 
        \wNDiag_23[18] , \wNDiag_23[17] , \wNDiag_23[16] , \wNDiag_23[15] , 
        \wNDiag_23[14] , \wNDiag_23[13] , \wNDiag_23[12] , \wNDiag_23[11] , 
        \wNDiag_23[10] , \wNDiag_23[9] , \wNDiag_23[8] , \wNDiag_23[7] , 
        \wNDiag_23[6] , \wNDiag_23[5] , \wNDiag_23[4] , \wNDiag_23[3] , 
        \wNDiag_23[2] , \wNDiag_23[1] , \wNDiag_23[0] }), .CallOut(
        \wCall_24[0] ), .ReturnOut(\wReturn_23[0] ), .ColOut({\wColumn_24[31] , 
        \wColumn_24[30] , \wColumn_24[29] , \wColumn_24[28] , \wColumn_24[27] , 
        \wColumn_24[26] , \wColumn_24[25] , \wColumn_24[24] , \wColumn_24[23] , 
        \wColumn_24[22] , \wColumn_24[21] , \wColumn_24[20] , \wColumn_24[19] , 
        \wColumn_24[18] , \wColumn_24[17] , \wColumn_24[16] , \wColumn_24[15] , 
        \wColumn_24[14] , \wColumn_24[13] , \wColumn_24[12] , \wColumn_24[11] , 
        \wColumn_24[10] , \wColumn_24[9] , \wColumn_24[8] , \wColumn_24[7] , 
        \wColumn_24[6] , \wColumn_24[5] , \wColumn_24[4] , \wColumn_24[3] , 
        \wColumn_24[2] , \wColumn_24[1] , \wColumn_24[0] }), .PDiagOut({
        \wPDiag_24[31] , \wPDiag_24[30] , \wPDiag_24[29] , \wPDiag_24[28] , 
        \wPDiag_24[27] , \wPDiag_24[26] , \wPDiag_24[25] , \wPDiag_24[24] , 
        \wPDiag_24[23] , \wPDiag_24[22] , \wPDiag_24[21] , \wPDiag_24[20] , 
        \wPDiag_24[19] , \wPDiag_24[18] , \wPDiag_24[17] , \wPDiag_24[16] , 
        \wPDiag_24[15] , \wPDiag_24[14] , \wPDiag_24[13] , \wPDiag_24[12] , 
        \wPDiag_24[11] , \wPDiag_24[10] , \wPDiag_24[9] , \wPDiag_24[8] , 
        \wPDiag_24[7] , \wPDiag_24[6] , \wPDiag_24[5] , \wPDiag_24[4] , 
        \wPDiag_24[3] , \wPDiag_24[2] , \wPDiag_24[1] , \wPDiag_24[0] }), 
        .NDiagOut({\wNDiag_24[31] , \wNDiag_24[30] , \wNDiag_24[29] , 
        \wNDiag_24[28] , \wNDiag_24[27] , \wNDiag_24[26] , \wNDiag_24[25] , 
        \wNDiag_24[24] , \wNDiag_24[23] , \wNDiag_24[22] , \wNDiag_24[21] , 
        \wNDiag_24[20] , \wNDiag_24[19] , \wNDiag_24[18] , \wNDiag_24[17] , 
        \wNDiag_24[16] , \wNDiag_24[15] , \wNDiag_24[14] , \wNDiag_24[13] , 
        \wNDiag_24[12] , \wNDiag_24[11] , \wNDiag_24[10] , \wNDiag_24[9] , 
        \wNDiag_24[8] , \wNDiag_24[7] , \wNDiag_24[6] , \wNDiag_24[5] , 
        \wNDiag_24[4] , \wNDiag_24[3] , \wNDiag_24[2] , \wNDiag_24[1] , 
        \wNDiag_24[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_31 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_32[5] , \wScan_32[4] , \wScan_32[3] , 
        \wScan_32[2] , \wScan_32[1] , \wScan_32[0] }), .ScanOut({\wScan_31[5] , 
        \wScan_31[4] , \wScan_31[3] , \wScan_31[2] , \wScan_31[1] , 
        \wScan_31[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_31[0] ), .ReturnIn(1'b0), .ColIn({
        \wColumn_31[31] , \wColumn_31[30] , \wColumn_31[29] , \wColumn_31[28] , 
        \wColumn_31[27] , \wColumn_31[26] , \wColumn_31[25] , \wColumn_31[24] , 
        \wColumn_31[23] , \wColumn_31[22] , \wColumn_31[21] , \wColumn_31[20] , 
        \wColumn_31[19] , \wColumn_31[18] , \wColumn_31[17] , \wColumn_31[16] , 
        \wColumn_31[15] , \wColumn_31[14] , \wColumn_31[13] , \wColumn_31[12] , 
        \wColumn_31[11] , \wColumn_31[10] , \wColumn_31[9] , \wColumn_31[8] , 
        \wColumn_31[7] , \wColumn_31[6] , \wColumn_31[5] , \wColumn_31[4] , 
        \wColumn_31[3] , \wColumn_31[2] , \wColumn_31[1] , \wColumn_31[0] }), 
        .PDiagIn({\wPDiag_31[31] , \wPDiag_31[30] , \wPDiag_31[29] , 
        \wPDiag_31[28] , \wPDiag_31[27] , \wPDiag_31[26] , \wPDiag_31[25] , 
        \wPDiag_31[24] , \wPDiag_31[23] , \wPDiag_31[22] , \wPDiag_31[21] , 
        \wPDiag_31[20] , \wPDiag_31[19] , \wPDiag_31[18] , \wPDiag_31[17] , 
        \wPDiag_31[16] , \wPDiag_31[15] , \wPDiag_31[14] , \wPDiag_31[13] , 
        \wPDiag_31[12] , \wPDiag_31[11] , \wPDiag_31[10] , \wPDiag_31[9] , 
        \wPDiag_31[8] , \wPDiag_31[7] , \wPDiag_31[6] , \wPDiag_31[5] , 
        \wPDiag_31[4] , \wPDiag_31[3] , \wPDiag_31[2] , \wPDiag_31[1] , 
        \wPDiag_31[0] }), .NDiagIn({\wNDiag_31[31] , \wNDiag_31[30] , 
        \wNDiag_31[29] , \wNDiag_31[28] , \wNDiag_31[27] , \wNDiag_31[26] , 
        \wNDiag_31[25] , \wNDiag_31[24] , \wNDiag_31[23] , \wNDiag_31[22] , 
        \wNDiag_31[21] , \wNDiag_31[20] , \wNDiag_31[19] , \wNDiag_31[18] , 
        \wNDiag_31[17] , \wNDiag_31[16] , \wNDiag_31[15] , \wNDiag_31[14] , 
        \wNDiag_31[13] , \wNDiag_31[12] , \wNDiag_31[11] , \wNDiag_31[10] , 
        \wNDiag_31[9] , \wNDiag_31[8] , \wNDiag_31[7] , \wNDiag_31[6] , 
        \wNDiag_31[5] , \wNDiag_31[4] , \wNDiag_31[3] , \wNDiag_31[2] , 
        \wNDiag_31[1] , \wNDiag_31[0] }), .CallOut(\wCall_32[0] ), .ReturnOut(
        \wReturn_31[0] ) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_22 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_23[5] , \wScan_23[4] , \wScan_23[3] , 
        \wScan_23[2] , \wScan_23[1] , \wScan_23[0] }), .ScanOut({\wScan_22[5] , 
        \wScan_22[4] , \wScan_22[3] , \wScan_22[2] , \wScan_22[1] , 
        \wScan_22[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_22[0] ), .ReturnIn(\wReturn_23[0] ), 
        .ColIn({\wColumn_22[31] , \wColumn_22[30] , \wColumn_22[29] , 
        \wColumn_22[28] , \wColumn_22[27] , \wColumn_22[26] , \wColumn_22[25] , 
        \wColumn_22[24] , \wColumn_22[23] , \wColumn_22[22] , \wColumn_22[21] , 
        \wColumn_22[20] , \wColumn_22[19] , \wColumn_22[18] , \wColumn_22[17] , 
        \wColumn_22[16] , \wColumn_22[15] , \wColumn_22[14] , \wColumn_22[13] , 
        \wColumn_22[12] , \wColumn_22[11] , \wColumn_22[10] , \wColumn_22[9] , 
        \wColumn_22[8] , \wColumn_22[7] , \wColumn_22[6] , \wColumn_22[5] , 
        \wColumn_22[4] , \wColumn_22[3] , \wColumn_22[2] , \wColumn_22[1] , 
        \wColumn_22[0] }), .PDiagIn({\wPDiag_22[31] , \wPDiag_22[30] , 
        \wPDiag_22[29] , \wPDiag_22[28] , \wPDiag_22[27] , \wPDiag_22[26] , 
        \wPDiag_22[25] , \wPDiag_22[24] , \wPDiag_22[23] , \wPDiag_22[22] , 
        \wPDiag_22[21] , \wPDiag_22[20] , \wPDiag_22[19] , \wPDiag_22[18] , 
        \wPDiag_22[17] , \wPDiag_22[16] , \wPDiag_22[15] , \wPDiag_22[14] , 
        \wPDiag_22[13] , \wPDiag_22[12] , \wPDiag_22[11] , \wPDiag_22[10] , 
        \wPDiag_22[9] , \wPDiag_22[8] , \wPDiag_22[7] , \wPDiag_22[6] , 
        \wPDiag_22[5] , \wPDiag_22[4] , \wPDiag_22[3] , \wPDiag_22[2] , 
        \wPDiag_22[1] , \wPDiag_22[0] }), .NDiagIn({\wNDiag_22[31] , 
        \wNDiag_22[30] , \wNDiag_22[29] , \wNDiag_22[28] , \wNDiag_22[27] , 
        \wNDiag_22[26] , \wNDiag_22[25] , \wNDiag_22[24] , \wNDiag_22[23] , 
        \wNDiag_22[22] , \wNDiag_22[21] , \wNDiag_22[20] , \wNDiag_22[19] , 
        \wNDiag_22[18] , \wNDiag_22[17] , \wNDiag_22[16] , \wNDiag_22[15] , 
        \wNDiag_22[14] , \wNDiag_22[13] , \wNDiag_22[12] , \wNDiag_22[11] , 
        \wNDiag_22[10] , \wNDiag_22[9] , \wNDiag_22[8] , \wNDiag_22[7] , 
        \wNDiag_22[6] , \wNDiag_22[5] , \wNDiag_22[4] , \wNDiag_22[3] , 
        \wNDiag_22[2] , \wNDiag_22[1] , \wNDiag_22[0] }), .CallOut(
        \wCall_23[0] ), .ReturnOut(\wReturn_22[0] ), .ColOut({\wColumn_23[31] , 
        \wColumn_23[30] , \wColumn_23[29] , \wColumn_23[28] , \wColumn_23[27] , 
        \wColumn_23[26] , \wColumn_23[25] , \wColumn_23[24] , \wColumn_23[23] , 
        \wColumn_23[22] , \wColumn_23[21] , \wColumn_23[20] , \wColumn_23[19] , 
        \wColumn_23[18] , \wColumn_23[17] , \wColumn_23[16] , \wColumn_23[15] , 
        \wColumn_23[14] , \wColumn_23[13] , \wColumn_23[12] , \wColumn_23[11] , 
        \wColumn_23[10] , \wColumn_23[9] , \wColumn_23[8] , \wColumn_23[7] , 
        \wColumn_23[6] , \wColumn_23[5] , \wColumn_23[4] , \wColumn_23[3] , 
        \wColumn_23[2] , \wColumn_23[1] , \wColumn_23[0] }), .PDiagOut({
        \wPDiag_23[31] , \wPDiag_23[30] , \wPDiag_23[29] , \wPDiag_23[28] , 
        \wPDiag_23[27] , \wPDiag_23[26] , \wPDiag_23[25] , \wPDiag_23[24] , 
        \wPDiag_23[23] , \wPDiag_23[22] , \wPDiag_23[21] , \wPDiag_23[20] , 
        \wPDiag_23[19] , \wPDiag_23[18] , \wPDiag_23[17] , \wPDiag_23[16] , 
        \wPDiag_23[15] , \wPDiag_23[14] , \wPDiag_23[13] , \wPDiag_23[12] , 
        \wPDiag_23[11] , \wPDiag_23[10] , \wPDiag_23[9] , \wPDiag_23[8] , 
        \wPDiag_23[7] , \wPDiag_23[6] , \wPDiag_23[5] , \wPDiag_23[4] , 
        \wPDiag_23[3] , \wPDiag_23[2] , \wPDiag_23[1] , \wPDiag_23[0] }), 
        .NDiagOut({\wNDiag_23[31] , \wNDiag_23[30] , \wNDiag_23[29] , 
        \wNDiag_23[28] , \wNDiag_23[27] , \wNDiag_23[26] , \wNDiag_23[25] , 
        \wNDiag_23[24] , \wNDiag_23[23] , \wNDiag_23[22] , \wNDiag_23[21] , 
        \wNDiag_23[20] , \wNDiag_23[19] , \wNDiag_23[18] , \wNDiag_23[17] , 
        \wNDiag_23[16] , \wNDiag_23[15] , \wNDiag_23[14] , \wNDiag_23[13] , 
        \wNDiag_23[12] , \wNDiag_23[11] , \wNDiag_23[10] , \wNDiag_23[9] , 
        \wNDiag_23[8] , \wNDiag_23[7] , \wNDiag_23[6] , \wNDiag_23[5] , 
        \wNDiag_23[4] , \wNDiag_23[3] , \wNDiag_23[2] , \wNDiag_23[1] , 
        \wNDiag_23[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_8 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_9[5] , \wScan_9[4] , \wScan_9[3] , 
        \wScan_9[2] , \wScan_9[1] , \wScan_9[0] }), .ScanOut({\wScan_8[5] , 
        \wScan_8[4] , \wScan_8[3] , \wScan_8[2] , \wScan_8[1] , \wScan_8[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0
        }), .CallIn(\wCall_8[0] ), .ReturnIn(\wReturn_9[0] ), .ColIn({
        \wColumn_8[31] , \wColumn_8[30] , \wColumn_8[29] , \wColumn_8[28] , 
        \wColumn_8[27] , \wColumn_8[26] , \wColumn_8[25] , \wColumn_8[24] , 
        \wColumn_8[23] , \wColumn_8[22] , \wColumn_8[21] , \wColumn_8[20] , 
        \wColumn_8[19] , \wColumn_8[18] , \wColumn_8[17] , \wColumn_8[16] , 
        \wColumn_8[15] , \wColumn_8[14] , \wColumn_8[13] , \wColumn_8[12] , 
        \wColumn_8[11] , \wColumn_8[10] , \wColumn_8[9] , \wColumn_8[8] , 
        \wColumn_8[7] , \wColumn_8[6] , \wColumn_8[5] , \wColumn_8[4] , 
        \wColumn_8[3] , \wColumn_8[2] , \wColumn_8[1] , \wColumn_8[0] }), 
        .PDiagIn({\wPDiag_8[31] , \wPDiag_8[30] , \wPDiag_8[29] , 
        \wPDiag_8[28] , \wPDiag_8[27] , \wPDiag_8[26] , \wPDiag_8[25] , 
        \wPDiag_8[24] , \wPDiag_8[23] , \wPDiag_8[22] , \wPDiag_8[21] , 
        \wPDiag_8[20] , \wPDiag_8[19] , \wPDiag_8[18] , \wPDiag_8[17] , 
        \wPDiag_8[16] , \wPDiag_8[15] , \wPDiag_8[14] , \wPDiag_8[13] , 
        \wPDiag_8[12] , \wPDiag_8[11] , \wPDiag_8[10] , \wPDiag_8[9] , 
        \wPDiag_8[8] , \wPDiag_8[7] , \wPDiag_8[6] , \wPDiag_8[5] , 
        \wPDiag_8[4] , \wPDiag_8[3] , \wPDiag_8[2] , \wPDiag_8[1] , 
        \wPDiag_8[0] }), .NDiagIn({\wNDiag_8[31] , \wNDiag_8[30] , 
        \wNDiag_8[29] , \wNDiag_8[28] , \wNDiag_8[27] , \wNDiag_8[26] , 
        \wNDiag_8[25] , \wNDiag_8[24] , \wNDiag_8[23] , \wNDiag_8[22] , 
        \wNDiag_8[21] , \wNDiag_8[20] , \wNDiag_8[19] , \wNDiag_8[18] , 
        \wNDiag_8[17] , \wNDiag_8[16] , \wNDiag_8[15] , \wNDiag_8[14] , 
        \wNDiag_8[13] , \wNDiag_8[12] , \wNDiag_8[11] , \wNDiag_8[10] , 
        \wNDiag_8[9] , \wNDiag_8[8] , \wNDiag_8[7] , \wNDiag_8[6] , 
        \wNDiag_8[5] , \wNDiag_8[4] , \wNDiag_8[3] , \wNDiag_8[2] , 
        \wNDiag_8[1] , \wNDiag_8[0] }), .CallOut(\wCall_9[0] ), .ReturnOut(
        \wReturn_8[0] ), .ColOut({\wColumn_9[31] , \wColumn_9[30] , 
        \wColumn_9[29] , \wColumn_9[28] , \wColumn_9[27] , \wColumn_9[26] , 
        \wColumn_9[25] , \wColumn_9[24] , \wColumn_9[23] , \wColumn_9[22] , 
        \wColumn_9[21] , \wColumn_9[20] , \wColumn_9[19] , \wColumn_9[18] , 
        \wColumn_9[17] , \wColumn_9[16] , \wColumn_9[15] , \wColumn_9[14] , 
        \wColumn_9[13] , \wColumn_9[12] , \wColumn_9[11] , \wColumn_9[10] , 
        \wColumn_9[9] , \wColumn_9[8] , \wColumn_9[7] , \wColumn_9[6] , 
        \wColumn_9[5] , \wColumn_9[4] , \wColumn_9[3] , \wColumn_9[2] , 
        \wColumn_9[1] , \wColumn_9[0] }), .PDiagOut({\wPDiag_9[31] , 
        \wPDiag_9[30] , \wPDiag_9[29] , \wPDiag_9[28] , \wPDiag_9[27] , 
        \wPDiag_9[26] , \wPDiag_9[25] , \wPDiag_9[24] , \wPDiag_9[23] , 
        \wPDiag_9[22] , \wPDiag_9[21] , \wPDiag_9[20] , \wPDiag_9[19] , 
        \wPDiag_9[18] , \wPDiag_9[17] , \wPDiag_9[16] , \wPDiag_9[15] , 
        \wPDiag_9[14] , \wPDiag_9[13] , \wPDiag_9[12] , \wPDiag_9[11] , 
        \wPDiag_9[10] , \wPDiag_9[9] , \wPDiag_9[8] , \wPDiag_9[7] , 
        \wPDiag_9[6] , \wPDiag_9[5] , \wPDiag_9[4] , \wPDiag_9[3] , 
        \wPDiag_9[2] , \wPDiag_9[1] , \wPDiag_9[0] }), .NDiagOut({
        \wNDiag_9[31] , \wNDiag_9[30] , \wNDiag_9[29] , \wNDiag_9[28] , 
        \wNDiag_9[27] , \wNDiag_9[26] , \wNDiag_9[25] , \wNDiag_9[24] , 
        \wNDiag_9[23] , \wNDiag_9[22] , \wNDiag_9[21] , \wNDiag_9[20] , 
        \wNDiag_9[19] , \wNDiag_9[18] , \wNDiag_9[17] , \wNDiag_9[16] , 
        \wNDiag_9[15] , \wNDiag_9[14] , \wNDiag_9[13] , \wNDiag_9[12] , 
        \wNDiag_9[11] , \wNDiag_9[10] , \wNDiag_9[9] , \wNDiag_9[8] , 
        \wNDiag_9[7] , \wNDiag_9[6] , \wNDiag_9[5] , \wNDiag_9[4] , 
        \wNDiag_9[3] , \wNDiag_9[2] , \wNDiag_9[1] , \wNDiag_9[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_10 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_11[5] , \wScan_11[4] , \wScan_11[3] , 
        \wScan_11[2] , \wScan_11[1] , \wScan_11[0] }), .ScanOut({\wScan_10[5] , 
        \wScan_10[4] , \wScan_10[3] , \wScan_10[2] , \wScan_10[1] , 
        \wScan_10[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_10[0] ), .ReturnIn(\wReturn_11[0] ), 
        .ColIn({\wColumn_10[31] , \wColumn_10[30] , \wColumn_10[29] , 
        \wColumn_10[28] , \wColumn_10[27] , \wColumn_10[26] , \wColumn_10[25] , 
        \wColumn_10[24] , \wColumn_10[23] , \wColumn_10[22] , \wColumn_10[21] , 
        \wColumn_10[20] , \wColumn_10[19] , \wColumn_10[18] , \wColumn_10[17] , 
        \wColumn_10[16] , \wColumn_10[15] , \wColumn_10[14] , \wColumn_10[13] , 
        \wColumn_10[12] , \wColumn_10[11] , \wColumn_10[10] , \wColumn_10[9] , 
        \wColumn_10[8] , \wColumn_10[7] , \wColumn_10[6] , \wColumn_10[5] , 
        \wColumn_10[4] , \wColumn_10[3] , \wColumn_10[2] , \wColumn_10[1] , 
        \wColumn_10[0] }), .PDiagIn({\wPDiag_10[31] , \wPDiag_10[30] , 
        \wPDiag_10[29] , \wPDiag_10[28] , \wPDiag_10[27] , \wPDiag_10[26] , 
        \wPDiag_10[25] , \wPDiag_10[24] , \wPDiag_10[23] , \wPDiag_10[22] , 
        \wPDiag_10[21] , \wPDiag_10[20] , \wPDiag_10[19] , \wPDiag_10[18] , 
        \wPDiag_10[17] , \wPDiag_10[16] , \wPDiag_10[15] , \wPDiag_10[14] , 
        \wPDiag_10[13] , \wPDiag_10[12] , \wPDiag_10[11] , \wPDiag_10[10] , 
        \wPDiag_10[9] , \wPDiag_10[8] , \wPDiag_10[7] , \wPDiag_10[6] , 
        \wPDiag_10[5] , \wPDiag_10[4] , \wPDiag_10[3] , \wPDiag_10[2] , 
        \wPDiag_10[1] , \wPDiag_10[0] }), .NDiagIn({\wNDiag_10[31] , 
        \wNDiag_10[30] , \wNDiag_10[29] , \wNDiag_10[28] , \wNDiag_10[27] , 
        \wNDiag_10[26] , \wNDiag_10[25] , \wNDiag_10[24] , \wNDiag_10[23] , 
        \wNDiag_10[22] , \wNDiag_10[21] , \wNDiag_10[20] , \wNDiag_10[19] , 
        \wNDiag_10[18] , \wNDiag_10[17] , \wNDiag_10[16] , \wNDiag_10[15] , 
        \wNDiag_10[14] , \wNDiag_10[13] , \wNDiag_10[12] , \wNDiag_10[11] , 
        \wNDiag_10[10] , \wNDiag_10[9] , \wNDiag_10[8] , \wNDiag_10[7] , 
        \wNDiag_10[6] , \wNDiag_10[5] , \wNDiag_10[4] , \wNDiag_10[3] , 
        \wNDiag_10[2] , \wNDiag_10[1] , \wNDiag_10[0] }), .CallOut(
        \wCall_11[0] ), .ReturnOut(\wReturn_10[0] ), .ColOut({\wColumn_11[31] , 
        \wColumn_11[30] , \wColumn_11[29] , \wColumn_11[28] , \wColumn_11[27] , 
        \wColumn_11[26] , \wColumn_11[25] , \wColumn_11[24] , \wColumn_11[23] , 
        \wColumn_11[22] , \wColumn_11[21] , \wColumn_11[20] , \wColumn_11[19] , 
        \wColumn_11[18] , \wColumn_11[17] , \wColumn_11[16] , \wColumn_11[15] , 
        \wColumn_11[14] , \wColumn_11[13] , \wColumn_11[12] , \wColumn_11[11] , 
        \wColumn_11[10] , \wColumn_11[9] , \wColumn_11[8] , \wColumn_11[7] , 
        \wColumn_11[6] , \wColumn_11[5] , \wColumn_11[4] , \wColumn_11[3] , 
        \wColumn_11[2] , \wColumn_11[1] , \wColumn_11[0] }), .PDiagOut({
        \wPDiag_11[31] , \wPDiag_11[30] , \wPDiag_11[29] , \wPDiag_11[28] , 
        \wPDiag_11[27] , \wPDiag_11[26] , \wPDiag_11[25] , \wPDiag_11[24] , 
        \wPDiag_11[23] , \wPDiag_11[22] , \wPDiag_11[21] , \wPDiag_11[20] , 
        \wPDiag_11[19] , \wPDiag_11[18] , \wPDiag_11[17] , \wPDiag_11[16] , 
        \wPDiag_11[15] , \wPDiag_11[14] , \wPDiag_11[13] , \wPDiag_11[12] , 
        \wPDiag_11[11] , \wPDiag_11[10] , \wPDiag_11[9] , \wPDiag_11[8] , 
        \wPDiag_11[7] , \wPDiag_11[6] , \wPDiag_11[5] , \wPDiag_11[4] , 
        \wPDiag_11[3] , \wPDiag_11[2] , \wPDiag_11[1] , \wPDiag_11[0] }), 
        .NDiagOut({\wNDiag_11[31] , \wNDiag_11[30] , \wNDiag_11[29] , 
        \wNDiag_11[28] , \wNDiag_11[27] , \wNDiag_11[26] , \wNDiag_11[25] , 
        \wNDiag_11[24] , \wNDiag_11[23] , \wNDiag_11[22] , \wNDiag_11[21] , 
        \wNDiag_11[20] , \wNDiag_11[19] , \wNDiag_11[18] , \wNDiag_11[17] , 
        \wNDiag_11[16] , \wNDiag_11[15] , \wNDiag_11[14] , \wNDiag_11[13] , 
        \wNDiag_11[12] , \wNDiag_11[11] , \wNDiag_11[10] , \wNDiag_11[9] , 
        \wNDiag_11[8] , \wNDiag_11[7] , \wNDiag_11[6] , \wNDiag_11[5] , 
        \wNDiag_11[4] , \wNDiag_11[3] , \wNDiag_11[2] , \wNDiag_11[1] , 
        \wNDiag_11[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_17 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_18[5] , \wScan_18[4] , \wScan_18[3] , 
        \wScan_18[2] , \wScan_18[1] , \wScan_18[0] }), .ScanOut({\wScan_17[5] , 
        \wScan_17[4] , \wScan_17[3] , \wScan_17[2] , \wScan_17[1] , 
        \wScan_17[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_17[0] ), .ReturnIn(\wReturn_18[0] ), 
        .ColIn({\wColumn_17[31] , \wColumn_17[30] , \wColumn_17[29] , 
        \wColumn_17[28] , \wColumn_17[27] , \wColumn_17[26] , \wColumn_17[25] , 
        \wColumn_17[24] , \wColumn_17[23] , \wColumn_17[22] , \wColumn_17[21] , 
        \wColumn_17[20] , \wColumn_17[19] , \wColumn_17[18] , \wColumn_17[17] , 
        \wColumn_17[16] , \wColumn_17[15] , \wColumn_17[14] , \wColumn_17[13] , 
        \wColumn_17[12] , \wColumn_17[11] , \wColumn_17[10] , \wColumn_17[9] , 
        \wColumn_17[8] , \wColumn_17[7] , \wColumn_17[6] , \wColumn_17[5] , 
        \wColumn_17[4] , \wColumn_17[3] , \wColumn_17[2] , \wColumn_17[1] , 
        \wColumn_17[0] }), .PDiagIn({\wPDiag_17[31] , \wPDiag_17[30] , 
        \wPDiag_17[29] , \wPDiag_17[28] , \wPDiag_17[27] , \wPDiag_17[26] , 
        \wPDiag_17[25] , \wPDiag_17[24] , \wPDiag_17[23] , \wPDiag_17[22] , 
        \wPDiag_17[21] , \wPDiag_17[20] , \wPDiag_17[19] , \wPDiag_17[18] , 
        \wPDiag_17[17] , \wPDiag_17[16] , \wPDiag_17[15] , \wPDiag_17[14] , 
        \wPDiag_17[13] , \wPDiag_17[12] , \wPDiag_17[11] , \wPDiag_17[10] , 
        \wPDiag_17[9] , \wPDiag_17[8] , \wPDiag_17[7] , \wPDiag_17[6] , 
        \wPDiag_17[5] , \wPDiag_17[4] , \wPDiag_17[3] , \wPDiag_17[2] , 
        \wPDiag_17[1] , \wPDiag_17[0] }), .NDiagIn({\wNDiag_17[31] , 
        \wNDiag_17[30] , \wNDiag_17[29] , \wNDiag_17[28] , \wNDiag_17[27] , 
        \wNDiag_17[26] , \wNDiag_17[25] , \wNDiag_17[24] , \wNDiag_17[23] , 
        \wNDiag_17[22] , \wNDiag_17[21] , \wNDiag_17[20] , \wNDiag_17[19] , 
        \wNDiag_17[18] , \wNDiag_17[17] , \wNDiag_17[16] , \wNDiag_17[15] , 
        \wNDiag_17[14] , \wNDiag_17[13] , \wNDiag_17[12] , \wNDiag_17[11] , 
        \wNDiag_17[10] , \wNDiag_17[9] , \wNDiag_17[8] , \wNDiag_17[7] , 
        \wNDiag_17[6] , \wNDiag_17[5] , \wNDiag_17[4] , \wNDiag_17[3] , 
        \wNDiag_17[2] , \wNDiag_17[1] , \wNDiag_17[0] }), .CallOut(
        \wCall_18[0] ), .ReturnOut(\wReturn_17[0] ), .ColOut({\wColumn_18[31] , 
        \wColumn_18[30] , \wColumn_18[29] , \wColumn_18[28] , \wColumn_18[27] , 
        \wColumn_18[26] , \wColumn_18[25] , \wColumn_18[24] , \wColumn_18[23] , 
        \wColumn_18[22] , \wColumn_18[21] , \wColumn_18[20] , \wColumn_18[19] , 
        \wColumn_18[18] , \wColumn_18[17] , \wColumn_18[16] , \wColumn_18[15] , 
        \wColumn_18[14] , \wColumn_18[13] , \wColumn_18[12] , \wColumn_18[11] , 
        \wColumn_18[10] , \wColumn_18[9] , \wColumn_18[8] , \wColumn_18[7] , 
        \wColumn_18[6] , \wColumn_18[5] , \wColumn_18[4] , \wColumn_18[3] , 
        \wColumn_18[2] , \wColumn_18[1] , \wColumn_18[0] }), .PDiagOut({
        \wPDiag_18[31] , \wPDiag_18[30] , \wPDiag_18[29] , \wPDiag_18[28] , 
        \wPDiag_18[27] , \wPDiag_18[26] , \wPDiag_18[25] , \wPDiag_18[24] , 
        \wPDiag_18[23] , \wPDiag_18[22] , \wPDiag_18[21] , \wPDiag_18[20] , 
        \wPDiag_18[19] , \wPDiag_18[18] , \wPDiag_18[17] , \wPDiag_18[16] , 
        \wPDiag_18[15] , \wPDiag_18[14] , \wPDiag_18[13] , \wPDiag_18[12] , 
        \wPDiag_18[11] , \wPDiag_18[10] , \wPDiag_18[9] , \wPDiag_18[8] , 
        \wPDiag_18[7] , \wPDiag_18[6] , \wPDiag_18[5] , \wPDiag_18[4] , 
        \wPDiag_18[3] , \wPDiag_18[2] , \wPDiag_18[1] , \wPDiag_18[0] }), 
        .NDiagOut({\wNDiag_18[31] , \wNDiag_18[30] , \wNDiag_18[29] , 
        \wNDiag_18[28] , \wNDiag_18[27] , \wNDiag_18[26] , \wNDiag_18[25] , 
        \wNDiag_18[24] , \wNDiag_18[23] , \wNDiag_18[22] , \wNDiag_18[21] , 
        \wNDiag_18[20] , \wNDiag_18[19] , \wNDiag_18[18] , \wNDiag_18[17] , 
        \wNDiag_18[16] , \wNDiag_18[15] , \wNDiag_18[14] , \wNDiag_18[13] , 
        \wNDiag_18[12] , \wNDiag_18[11] , \wNDiag_18[10] , \wNDiag_18[9] , 
        \wNDiag_18[8] , \wNDiag_18[7] , \wNDiag_18[6] , \wNDiag_18[5] , 
        \wNDiag_18[4] , \wNDiag_18[3] , \wNDiag_18[2] , \wNDiag_18[1] , 
        \wNDiag_18[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_30 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_31[5] , \wScan_31[4] , \wScan_31[3] , 
        \wScan_31[2] , \wScan_31[1] , \wScan_31[0] }), .ScanOut({\wScan_30[5] , 
        \wScan_30[4] , \wScan_30[3] , \wScan_30[2] , \wScan_30[1] , 
        \wScan_30[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_30[0] ), .ReturnIn(\wReturn_31[0] ), 
        .ColIn({\wColumn_30[31] , \wColumn_30[30] , \wColumn_30[29] , 
        \wColumn_30[28] , \wColumn_30[27] , \wColumn_30[26] , \wColumn_30[25] , 
        \wColumn_30[24] , \wColumn_30[23] , \wColumn_30[22] , \wColumn_30[21] , 
        \wColumn_30[20] , \wColumn_30[19] , \wColumn_30[18] , \wColumn_30[17] , 
        \wColumn_30[16] , \wColumn_30[15] , \wColumn_30[14] , \wColumn_30[13] , 
        \wColumn_30[12] , \wColumn_30[11] , \wColumn_30[10] , \wColumn_30[9] , 
        \wColumn_30[8] , \wColumn_30[7] , \wColumn_30[6] , \wColumn_30[5] , 
        \wColumn_30[4] , \wColumn_30[3] , \wColumn_30[2] , \wColumn_30[1] , 
        \wColumn_30[0] }), .PDiagIn({\wPDiag_30[31] , \wPDiag_30[30] , 
        \wPDiag_30[29] , \wPDiag_30[28] , \wPDiag_30[27] , \wPDiag_30[26] , 
        \wPDiag_30[25] , \wPDiag_30[24] , \wPDiag_30[23] , \wPDiag_30[22] , 
        \wPDiag_30[21] , \wPDiag_30[20] , \wPDiag_30[19] , \wPDiag_30[18] , 
        \wPDiag_30[17] , \wPDiag_30[16] , \wPDiag_30[15] , \wPDiag_30[14] , 
        \wPDiag_30[13] , \wPDiag_30[12] , \wPDiag_30[11] , \wPDiag_30[10] , 
        \wPDiag_30[9] , \wPDiag_30[8] , \wPDiag_30[7] , \wPDiag_30[6] , 
        \wPDiag_30[5] , \wPDiag_30[4] , \wPDiag_30[3] , \wPDiag_30[2] , 
        \wPDiag_30[1] , \wPDiag_30[0] }), .NDiagIn({\wNDiag_30[31] , 
        \wNDiag_30[30] , \wNDiag_30[29] , \wNDiag_30[28] , \wNDiag_30[27] , 
        \wNDiag_30[26] , \wNDiag_30[25] , \wNDiag_30[24] , \wNDiag_30[23] , 
        \wNDiag_30[22] , \wNDiag_30[21] , \wNDiag_30[20] , \wNDiag_30[19] , 
        \wNDiag_30[18] , \wNDiag_30[17] , \wNDiag_30[16] , \wNDiag_30[15] , 
        \wNDiag_30[14] , \wNDiag_30[13] , \wNDiag_30[12] , \wNDiag_30[11] , 
        \wNDiag_30[10] , \wNDiag_30[9] , \wNDiag_30[8] , \wNDiag_30[7] , 
        \wNDiag_30[6] , \wNDiag_30[5] , \wNDiag_30[4] , \wNDiag_30[3] , 
        \wNDiag_30[2] , \wNDiag_30[1] , \wNDiag_30[0] }), .CallOut(
        \wCall_31[0] ), .ReturnOut(\wReturn_30[0] ), .ColOut({\wColumn_31[31] , 
        \wColumn_31[30] , \wColumn_31[29] , \wColumn_31[28] , \wColumn_31[27] , 
        \wColumn_31[26] , \wColumn_31[25] , \wColumn_31[24] , \wColumn_31[23] , 
        \wColumn_31[22] , \wColumn_31[21] , \wColumn_31[20] , \wColumn_31[19] , 
        \wColumn_31[18] , \wColumn_31[17] , \wColumn_31[16] , \wColumn_31[15] , 
        \wColumn_31[14] , \wColumn_31[13] , \wColumn_31[12] , \wColumn_31[11] , 
        \wColumn_31[10] , \wColumn_31[9] , \wColumn_31[8] , \wColumn_31[7] , 
        \wColumn_31[6] , \wColumn_31[5] , \wColumn_31[4] , \wColumn_31[3] , 
        \wColumn_31[2] , \wColumn_31[1] , \wColumn_31[0] }), .PDiagOut({
        \wPDiag_31[31] , \wPDiag_31[30] , \wPDiag_31[29] , \wPDiag_31[28] , 
        \wPDiag_31[27] , \wPDiag_31[26] , \wPDiag_31[25] , \wPDiag_31[24] , 
        \wPDiag_31[23] , \wPDiag_31[22] , \wPDiag_31[21] , \wPDiag_31[20] , 
        \wPDiag_31[19] , \wPDiag_31[18] , \wPDiag_31[17] , \wPDiag_31[16] , 
        \wPDiag_31[15] , \wPDiag_31[14] , \wPDiag_31[13] , \wPDiag_31[12] , 
        \wPDiag_31[11] , \wPDiag_31[10] , \wPDiag_31[9] , \wPDiag_31[8] , 
        \wPDiag_31[7] , \wPDiag_31[6] , \wPDiag_31[5] , \wPDiag_31[4] , 
        \wPDiag_31[3] , \wPDiag_31[2] , \wPDiag_31[1] , \wPDiag_31[0] }), 
        .NDiagOut({\wNDiag_31[31] , \wNDiag_31[30] , \wNDiag_31[29] , 
        \wNDiag_31[28] , \wNDiag_31[27] , \wNDiag_31[26] , \wNDiag_31[25] , 
        \wNDiag_31[24] , \wNDiag_31[23] , \wNDiag_31[22] , \wNDiag_31[21] , 
        \wNDiag_31[20] , \wNDiag_31[19] , \wNDiag_31[18] , \wNDiag_31[17] , 
        \wNDiag_31[16] , \wNDiag_31[15] , \wNDiag_31[14] , \wNDiag_31[13] , 
        \wNDiag_31[12] , \wNDiag_31[11] , \wNDiag_31[10] , \wNDiag_31[9] , 
        \wNDiag_31[8] , \wNDiag_31[7] , \wNDiag_31[6] , \wNDiag_31[5] , 
        \wNDiag_31[4] , \wNDiag_31[3] , \wNDiag_31[2] , \wNDiag_31[1] , 
        \wNDiag_31[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_19 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_20[5] , \wScan_20[4] , \wScan_20[3] , 
        \wScan_20[2] , \wScan_20[1] , \wScan_20[0] }), .ScanOut({\wScan_19[5] , 
        \wScan_19[4] , \wScan_19[3] , \wScan_19[2] , \wScan_19[1] , 
        \wScan_19[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_19[0] ), .ReturnIn(\wReturn_20[0] ), 
        .ColIn({\wColumn_19[31] , \wColumn_19[30] , \wColumn_19[29] , 
        \wColumn_19[28] , \wColumn_19[27] , \wColumn_19[26] , \wColumn_19[25] , 
        \wColumn_19[24] , \wColumn_19[23] , \wColumn_19[22] , \wColumn_19[21] , 
        \wColumn_19[20] , \wColumn_19[19] , \wColumn_19[18] , \wColumn_19[17] , 
        \wColumn_19[16] , \wColumn_19[15] , \wColumn_19[14] , \wColumn_19[13] , 
        \wColumn_19[12] , \wColumn_19[11] , \wColumn_19[10] , \wColumn_19[9] , 
        \wColumn_19[8] , \wColumn_19[7] , \wColumn_19[6] , \wColumn_19[5] , 
        \wColumn_19[4] , \wColumn_19[3] , \wColumn_19[2] , \wColumn_19[1] , 
        \wColumn_19[0] }), .PDiagIn({\wPDiag_19[31] , \wPDiag_19[30] , 
        \wPDiag_19[29] , \wPDiag_19[28] , \wPDiag_19[27] , \wPDiag_19[26] , 
        \wPDiag_19[25] , \wPDiag_19[24] , \wPDiag_19[23] , \wPDiag_19[22] , 
        \wPDiag_19[21] , \wPDiag_19[20] , \wPDiag_19[19] , \wPDiag_19[18] , 
        \wPDiag_19[17] , \wPDiag_19[16] , \wPDiag_19[15] , \wPDiag_19[14] , 
        \wPDiag_19[13] , \wPDiag_19[12] , \wPDiag_19[11] , \wPDiag_19[10] , 
        \wPDiag_19[9] , \wPDiag_19[8] , \wPDiag_19[7] , \wPDiag_19[6] , 
        \wPDiag_19[5] , \wPDiag_19[4] , \wPDiag_19[3] , \wPDiag_19[2] , 
        \wPDiag_19[1] , \wPDiag_19[0] }), .NDiagIn({\wNDiag_19[31] , 
        \wNDiag_19[30] , \wNDiag_19[29] , \wNDiag_19[28] , \wNDiag_19[27] , 
        \wNDiag_19[26] , \wNDiag_19[25] , \wNDiag_19[24] , \wNDiag_19[23] , 
        \wNDiag_19[22] , \wNDiag_19[21] , \wNDiag_19[20] , \wNDiag_19[19] , 
        \wNDiag_19[18] , \wNDiag_19[17] , \wNDiag_19[16] , \wNDiag_19[15] , 
        \wNDiag_19[14] , \wNDiag_19[13] , \wNDiag_19[12] , \wNDiag_19[11] , 
        \wNDiag_19[10] , \wNDiag_19[9] , \wNDiag_19[8] , \wNDiag_19[7] , 
        \wNDiag_19[6] , \wNDiag_19[5] , \wNDiag_19[4] , \wNDiag_19[3] , 
        \wNDiag_19[2] , \wNDiag_19[1] , \wNDiag_19[0] }), .CallOut(
        \wCall_20[0] ), .ReturnOut(\wReturn_19[0] ), .ColOut({\wColumn_20[31] , 
        \wColumn_20[30] , \wColumn_20[29] , \wColumn_20[28] , \wColumn_20[27] , 
        \wColumn_20[26] , \wColumn_20[25] , \wColumn_20[24] , \wColumn_20[23] , 
        \wColumn_20[22] , \wColumn_20[21] , \wColumn_20[20] , \wColumn_20[19] , 
        \wColumn_20[18] , \wColumn_20[17] , \wColumn_20[16] , \wColumn_20[15] , 
        \wColumn_20[14] , \wColumn_20[13] , \wColumn_20[12] , \wColumn_20[11] , 
        \wColumn_20[10] , \wColumn_20[9] , \wColumn_20[8] , \wColumn_20[7] , 
        \wColumn_20[6] , \wColumn_20[5] , \wColumn_20[4] , \wColumn_20[3] , 
        \wColumn_20[2] , \wColumn_20[1] , \wColumn_20[0] }), .PDiagOut({
        \wPDiag_20[31] , \wPDiag_20[30] , \wPDiag_20[29] , \wPDiag_20[28] , 
        \wPDiag_20[27] , \wPDiag_20[26] , \wPDiag_20[25] , \wPDiag_20[24] , 
        \wPDiag_20[23] , \wPDiag_20[22] , \wPDiag_20[21] , \wPDiag_20[20] , 
        \wPDiag_20[19] , \wPDiag_20[18] , \wPDiag_20[17] , \wPDiag_20[16] , 
        \wPDiag_20[15] , \wPDiag_20[14] , \wPDiag_20[13] , \wPDiag_20[12] , 
        \wPDiag_20[11] , \wPDiag_20[10] , \wPDiag_20[9] , \wPDiag_20[8] , 
        \wPDiag_20[7] , \wPDiag_20[6] , \wPDiag_20[5] , \wPDiag_20[4] , 
        \wPDiag_20[3] , \wPDiag_20[2] , \wPDiag_20[1] , \wPDiag_20[0] }), 
        .NDiagOut({\wNDiag_20[31] , \wNDiag_20[30] , \wNDiag_20[29] , 
        \wNDiag_20[28] , \wNDiag_20[27] , \wNDiag_20[26] , \wNDiag_20[25] , 
        \wNDiag_20[24] , \wNDiag_20[23] , \wNDiag_20[22] , \wNDiag_20[21] , 
        \wNDiag_20[20] , \wNDiag_20[19] , \wNDiag_20[18] , \wNDiag_20[17] , 
        \wNDiag_20[16] , \wNDiag_20[15] , \wNDiag_20[14] , \wNDiag_20[13] , 
        \wNDiag_20[12] , \wNDiag_20[11] , \wNDiag_20[10] , \wNDiag_20[9] , 
        \wNDiag_20[8] , \wNDiag_20[7] , \wNDiag_20[6] , \wNDiag_20[5] , 
        \wNDiag_20[4] , \wNDiag_20[3] , \wNDiag_20[2] , \wNDiag_20[1] , 
        \wNDiag_20[0] }) );
    NQueens_Node_WIDTH32_IDWIDTH6_SCAN1 U_NQueens_Node_25 ( .Clk(Clk), .Reset(
        Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(
        DataOut), .ScanIn({\wScan_26[5] , \wScan_26[4] , \wScan_26[3] , 
        \wScan_26[2] , \wScan_26[1] , \wScan_26[0] }), .ScanOut({\wScan_25[5] , 
        \wScan_25[4] , \wScan_25[3] , \wScan_25[2] , \wScan_25[1] , 
        \wScan_25[0] }), .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CallIn(\wCall_25[0] ), .ReturnIn(\wReturn_26[0] ), 
        .ColIn({\wColumn_25[31] , \wColumn_25[30] , \wColumn_25[29] , 
        \wColumn_25[28] , \wColumn_25[27] , \wColumn_25[26] , \wColumn_25[25] , 
        \wColumn_25[24] , \wColumn_25[23] , \wColumn_25[22] , \wColumn_25[21] , 
        \wColumn_25[20] , \wColumn_25[19] , \wColumn_25[18] , \wColumn_25[17] , 
        \wColumn_25[16] , \wColumn_25[15] , \wColumn_25[14] , \wColumn_25[13] , 
        \wColumn_25[12] , \wColumn_25[11] , \wColumn_25[10] , \wColumn_25[9] , 
        \wColumn_25[8] , \wColumn_25[7] , \wColumn_25[6] , \wColumn_25[5] , 
        \wColumn_25[4] , \wColumn_25[3] , \wColumn_25[2] , \wColumn_25[1] , 
        \wColumn_25[0] }), .PDiagIn({\wPDiag_25[31] , \wPDiag_25[30] , 
        \wPDiag_25[29] , \wPDiag_25[28] , \wPDiag_25[27] , \wPDiag_25[26] , 
        \wPDiag_25[25] , \wPDiag_25[24] , \wPDiag_25[23] , \wPDiag_25[22] , 
        \wPDiag_25[21] , \wPDiag_25[20] , \wPDiag_25[19] , \wPDiag_25[18] , 
        \wPDiag_25[17] , \wPDiag_25[16] , \wPDiag_25[15] , \wPDiag_25[14] , 
        \wPDiag_25[13] , \wPDiag_25[12] , \wPDiag_25[11] , \wPDiag_25[10] , 
        \wPDiag_25[9] , \wPDiag_25[8] , \wPDiag_25[7] , \wPDiag_25[6] , 
        \wPDiag_25[5] , \wPDiag_25[4] , \wPDiag_25[3] , \wPDiag_25[2] , 
        \wPDiag_25[1] , \wPDiag_25[0] }), .NDiagIn({\wNDiag_25[31] , 
        \wNDiag_25[30] , \wNDiag_25[29] , \wNDiag_25[28] , \wNDiag_25[27] , 
        \wNDiag_25[26] , \wNDiag_25[25] , \wNDiag_25[24] , \wNDiag_25[23] , 
        \wNDiag_25[22] , \wNDiag_25[21] , \wNDiag_25[20] , \wNDiag_25[19] , 
        \wNDiag_25[18] , \wNDiag_25[17] , \wNDiag_25[16] , \wNDiag_25[15] , 
        \wNDiag_25[14] , \wNDiag_25[13] , \wNDiag_25[12] , \wNDiag_25[11] , 
        \wNDiag_25[10] , \wNDiag_25[9] , \wNDiag_25[8] , \wNDiag_25[7] , 
        \wNDiag_25[6] , \wNDiag_25[5] , \wNDiag_25[4] , \wNDiag_25[3] , 
        \wNDiag_25[2] , \wNDiag_25[1] , \wNDiag_25[0] }), .CallOut(
        \wCall_26[0] ), .ReturnOut(\wReturn_25[0] ), .ColOut({\wColumn_26[31] , 
        \wColumn_26[30] , \wColumn_26[29] , \wColumn_26[28] , \wColumn_26[27] , 
        \wColumn_26[26] , \wColumn_26[25] , \wColumn_26[24] , \wColumn_26[23] , 
        \wColumn_26[22] , \wColumn_26[21] , \wColumn_26[20] , \wColumn_26[19] , 
        \wColumn_26[18] , \wColumn_26[17] , \wColumn_26[16] , \wColumn_26[15] , 
        \wColumn_26[14] , \wColumn_26[13] , \wColumn_26[12] , \wColumn_26[11] , 
        \wColumn_26[10] , \wColumn_26[9] , \wColumn_26[8] , \wColumn_26[7] , 
        \wColumn_26[6] , \wColumn_26[5] , \wColumn_26[4] , \wColumn_26[3] , 
        \wColumn_26[2] , \wColumn_26[1] , \wColumn_26[0] }), .PDiagOut({
        \wPDiag_26[31] , \wPDiag_26[30] , \wPDiag_26[29] , \wPDiag_26[28] , 
        \wPDiag_26[27] , \wPDiag_26[26] , \wPDiag_26[25] , \wPDiag_26[24] , 
        \wPDiag_26[23] , \wPDiag_26[22] , \wPDiag_26[21] , \wPDiag_26[20] , 
        \wPDiag_26[19] , \wPDiag_26[18] , \wPDiag_26[17] , \wPDiag_26[16] , 
        \wPDiag_26[15] , \wPDiag_26[14] , \wPDiag_26[13] , \wPDiag_26[12] , 
        \wPDiag_26[11] , \wPDiag_26[10] , \wPDiag_26[9] , \wPDiag_26[8] , 
        \wPDiag_26[7] , \wPDiag_26[6] , \wPDiag_26[5] , \wPDiag_26[4] , 
        \wPDiag_26[3] , \wPDiag_26[2] , \wPDiag_26[1] , \wPDiag_26[0] }), 
        .NDiagOut({\wNDiag_26[31] , \wNDiag_26[30] , \wNDiag_26[29] , 
        \wNDiag_26[28] , \wNDiag_26[27] , \wNDiag_26[26] , \wNDiag_26[25] , 
        \wNDiag_26[24] , \wNDiag_26[23] , \wNDiag_26[22] , \wNDiag_26[21] , 
        \wNDiag_26[20] , \wNDiag_26[19] , \wNDiag_26[18] , \wNDiag_26[17] , 
        \wNDiag_26[16] , \wNDiag_26[15] , \wNDiag_26[14] , \wNDiag_26[13] , 
        \wNDiag_26[12] , \wNDiag_26[11] , \wNDiag_26[10] , \wNDiag_26[9] , 
        \wNDiag_26[8] , \wNDiag_26[7] , \wNDiag_26[6] , \wNDiag_26[5] , 
        \wNDiag_26[4] , \wNDiag_26[3] , \wNDiag_26[2] , \wNDiag_26[1] , 
        \wNDiag_26[0] }) );
    NQueens_Control_IDWIDTH6_SCAN1 U_NQueens_Control ( .Clk(Clk), .Reset(Reset
        ), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\wScan_0[5] , \wScan_0[4] , \wScan_0[3] , \wScan_0[2] , 
        \wScan_0[1] , \wScan_0[0] }), .ScanOut({\wScan_32[5] , \wScan_32[4] , 
        \wScan_32[3] , \wScan_32[2] , \wScan_32[1] , \wScan_32[0] }), 
        .ScanEnable(\wScanEnable[0] ), .Id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1
        }), .ScanId({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CallIn(
        \wCall_32[0] ), .ReturnIn(\wReturn_0[0] ), .CallOut(\wCall_0[0] ) );
endmodule

