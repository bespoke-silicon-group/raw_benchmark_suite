
module EdgeAux_DW01_add_16_0 ( A, B, CI, SUM, CO );
input  [15:0] A;
input  [15:0] B;
output [15:0] SUM;
input  CI;
output CO;
    wire \carry[15] , \carry[13] , \carry[9] , \carry[4] , \carry[6] , 
        \carry[2] , \carry[14] , \carry[11] , \carry[10] , \carry[12] , 
        \carry[8] , \carry[7] , \carry[3] , \carry[5] , \carry[1] , n1;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(
        \carry[9] ) );
    VMW_FADD U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(
        \carry[8] ) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(
        \carry[10] ) );
    VMW_FADD U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
    VMW_FADD U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
    VMW_FADD U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]) );
    VMW_FADD U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
    VMW_FADD U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
endmodule


module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [7:0] Eid;
input  [7:0] WeightAddr;
input  [15:0] InEdge;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire \Weight[11] , \Weight[6] , \Weight[15] , \Weight[2] , \Weight[0] , 
        \Weight[9] , \Weight[13] , \Weight[4] , \Weight[12] , \Weight[5] , 
        \Weight[1] , \Weight[8] , \Weight[14] , \Weight[3] , \Weight[10] , 
        \Weight[7] , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101, n102, n103;
    VMW_PULLDOWN U15 ( .Z(n103) );
    VMW_AO22 U16 ( .A(\Weight[9] ), .B(n76), .C(WeightData[9]), .D(n77), .Z(
        n93) );
    VMW_AO22 U17 ( .A(\Weight[8] ), .B(n76), .C(WeightData[8]), .D(n77), .Z(
        n94) );
    VMW_AO22 U18 ( .A(\Weight[7] ), .B(n76), .C(WeightData[7]), .D(n77), .Z(
        n95) );
    VMW_AO22 U19 ( .A(\Weight[6] ), .B(n76), .C(WeightData[6]), .D(n77), .Z(
        n96) );
    VMW_AO22 U20 ( .A(\Weight[5] ), .B(n76), .C(WeightData[5]), .D(n77), .Z(
        n97) );
    VMW_AO22 U21 ( .A(\Weight[4] ), .B(n76), .C(WeightData[4]), .D(n77), .Z(
        n98) );
    VMW_AO22 U22 ( .A(\Weight[3] ), .B(n76), .C(WeightData[3]), .D(n77), .Z(
        n99) );
    VMW_AO22 U23 ( .A(\Weight[2] ), .B(n76), .C(WeightData[2]), .D(n77), .Z(
        n100) );
    VMW_AO22 U24 ( .A(\Weight[1] ), .B(n76), .C(WeightData[1]), .D(n77), .Z(
        n101) );
    VMW_AO22 U25 ( .A(\Weight[15] ), .B(n76), .C(WeightData[15]), .D(n77), .Z(
        n87) );
    VMW_AO22 U26 ( .A(\Weight[14] ), .B(n76), .C(WeightData[14]), .D(n77), .Z(
        n88) );
    VMW_AO22 U27 ( .A(\Weight[13] ), .B(n76), .C(WeightData[13]), .D(n77), .Z(
        n89) );
    VMW_AO22 U28 ( .A(\Weight[12] ), .B(n76), .C(WeightData[12]), .D(n77), .Z(
        n90) );
    VMW_AO22 U29 ( .A(\Weight[11] ), .B(n76), .C(WeightData[11]), .D(n77), .Z(
        n91) );
    VMW_AO22 U30 ( .A(\Weight[10] ), .B(n76), .C(WeightData[10]), .D(n77), .Z(
        n92) );
    VMW_AO22 U31 ( .A(\Weight[0] ), .B(n76), .C(WeightData[0]), .D(n77), .Z(
        n102) );
    VMW_AND4 U32 ( .A(n79), .B(n80), .C(n81), .D(n82), .Z(n78) );
    VMW_AND5 U33 ( .A(n83), .B(n84), .C(n85), .D(n86), .E(n78), .Z(n77) );
    VMW_XNOR2 U34 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n82) );
    VMW_XNOR2 U35 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n81) );
    VMW_XNOR2 U36 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n80) );
    VMW_XNOR2 U37 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n79) );
    VMW_XNOR2 U38 ( .A(WeightAddr[6]), .B(Eid[6]), .Z(n86) );
    VMW_XNOR2 U39 ( .A(WeightAddr[7]), .B(Eid[7]), .Z(n85) );
    VMW_XNOR2 U40 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n84) );
    VMW_XNOR2 U41 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n83) );
    VMW_INV U42 ( .A(n77), .Z(n76) );
    VMW_FD \Weight_reg[15]  ( .D(n87), .CP(Clk), .Q(\Weight[15] ) );
    VMW_FD \Weight_reg[14]  ( .D(n88), .CP(Clk), .Q(\Weight[14] ) );
    VMW_FD \Weight_reg[13]  ( .D(n89), .CP(Clk), .Q(\Weight[13] ) );
    VMW_FD \Weight_reg[12]  ( .D(n90), .CP(Clk), .Q(\Weight[12] ) );
    VMW_FD \Weight_reg[11]  ( .D(n91), .CP(Clk), .Q(\Weight[11] ) );
    VMW_FD \Weight_reg[10]  ( .D(n92), .CP(Clk), .Q(\Weight[10] ) );
    VMW_FD \Weight_reg[9]  ( .D(n93), .CP(Clk), .Q(\Weight[9] ) );
    VMW_FD \Weight_reg[8]  ( .D(n94), .CP(Clk), .Q(\Weight[8] ) );
    VMW_FD \Weight_reg[7]  ( .D(n95), .CP(Clk), .Q(\Weight[7] ) );
    VMW_FD \Weight_reg[6]  ( .D(n96), .CP(Clk), .Q(\Weight[6] ) );
    VMW_FD \Weight_reg[5]  ( .D(n97), .CP(Clk), .Q(\Weight[5] ) );
    VMW_FD \Weight_reg[4]  ( .D(n98), .CP(Clk), .Q(\Weight[4] ) );
    VMW_FD \Weight_reg[3]  ( .D(n99), .CP(Clk), .Q(\Weight[3] ) );
    VMW_FD \Weight_reg[2]  ( .D(n100), .CP(Clk), .Q(\Weight[2] ) );
    VMW_FD \Weight_reg[1]  ( .D(n101), .CP(Clk), .Q(\Weight[1] ) );
    VMW_FD \Weight_reg[0]  ( .D(n102), .CP(Clk), .Q(\Weight[0] ) );
    EdgeAux_DW01_add_16_0 add_92 ( .A({\Weight[15] , \Weight[14] , 
        \Weight[13] , \Weight[12] , \Weight[11] , \Weight[10] , \Weight[9] , 
        \Weight[8] , \Weight[7] , \Weight[6] , \Weight[5] , \Weight[4] , 
        \Weight[3] , \Weight[2] , \Weight[1] , \Weight[0] }), .B(InEdge), .CI(
        n103), .SUM(OutEdge) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, 
        n107, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n91), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, 
        n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n131), .D(n129), .Z(n133) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n167), .C(n166), .D(n161), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n156) );
    VMW_INV U34 ( .A(B[7]), .Z(n145) );
    VMW_INV U35 ( .A(A[7]), .Z(n148) );
    VMW_INV U36 ( .A(A[3]), .Z(n134) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n150) );
    VMW_INV U39 ( .A(B[9]), .Z(n152) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n162) );
    VMW_INV U43 ( .A(B[11]), .Z(n158) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n167) );
    VMW_INV U48 ( .A(B[13]), .Z(n164) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216;
    VMW_OAI21 U3 ( .A(B[15]), .B(n168), .C(n169), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n171), .B(B[2]), .Z(n170) );
    VMW_AO22 U5 ( .A(n173), .B(B[0]), .C(n174), .D(B[1]), .Z(n172) );
    VMW_OR2 U6 ( .A(B[2]), .B(n171), .Z(n175) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n174), .C(n175), .D(n172), .Z(n176) );
    VMW_NAND2 U8 ( .A(n178), .B(B[4]), .Z(n177) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n180), .C(n176), .D(n170), .Z(n179) );
    VMW_OR2 U10 ( .A(B[4]), .B(n178), .Z(n181) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n183), .C(n181), .D(n179), .Z(n182) );
    VMW_NAND2 U12 ( .A(n185), .B(B[6]), .Z(n184) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n187), .C(n182), .D(n177), .Z(n186) );
    VMW_OR2 U14 ( .A(B[6]), .B(n185), .Z(n188) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n190), .C(n188), .D(n186), .Z(n189) );
    VMW_NAND2 U16 ( .A(n192), .B(B[8]), .Z(n191) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n194), .C(n189), .D(n184), .Z(n193) );
    VMW_OR2 U18 ( .A(B[8]), .B(n192), .Z(n195) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n197), .C(n195), .D(n193), .Z(n196) );
    VMW_NAND2 U20 ( .A(n199), .B(B[10]), .Z(n198) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n201), .C(n196), .D(n191), .Z(n200) );
    VMW_NAND2 U22 ( .A(n201), .B(A[9]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n199), .C(n202), .D(n200), .Z(n203) );
    VMW_NAND2 U24 ( .A(n205), .B(B[12]), .Z(n204) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n207), .C(n203), .D(n198), .Z(n206) );
    VMW_NAND2 U26 ( .A(n207), .B(A[11]), .Z(n208) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n205), .C(n208), .D(n206), .Z(n209) );
    VMW_NAND2 U28 ( .A(n211), .B(B[14]), .Z(n210) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n213), .C(n209), .D(n204), .Z(n212) );
    VMW_NAND2 U30 ( .A(n213), .B(A[13]), .Z(n214) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n211), .C(n214), .D(n212), .Z(n215) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n216), .C(n215), .D(n210), .Z(n169) );
    VMW_INV U33 ( .A(A[12]), .Z(n205) );
    VMW_INV U34 ( .A(B[7]), .Z(n194) );
    VMW_INV U35 ( .A(A[7]), .Z(n197) );
    VMW_INV U36 ( .A(A[3]), .Z(n183) );
    VMW_INV U37 ( .A(B[3]), .Z(n180) );
    VMW_INV U38 ( .A(A[10]), .Z(n199) );
    VMW_INV U39 ( .A(B[9]), .Z(n201) );
    VMW_INV U40 ( .A(A[4]), .Z(n178) );
    VMW_INV U41 ( .A(A[8]), .Z(n192) );
    VMW_INV U42 ( .A(A[14]), .Z(n211) );
    VMW_INV U43 ( .A(B[11]), .Z(n207) );
    VMW_INV U44 ( .A(A[5]), .Z(n190) );
    VMW_INV U45 ( .A(B[5]), .Z(n187) );
    VMW_INV U46 ( .A(A[1]), .Z(n174) );
    VMW_INV U47 ( .A(B[15]), .Z(n216) );
    VMW_INV U48 ( .A(B[13]), .Z(n213) );
    VMW_INV U49 ( .A(A[6]), .Z(n185) );
    VMW_INV U50 ( .A(A[2]), .Z(n171) );
    VMW_INV U51 ( .A(A[0]), .Z(n173) );
    VMW_INV U52 ( .A(A[15]), .Z(n168) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265;
    VMW_OAI21 U3 ( .A(B[15]), .B(n217), .C(n218), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n220), .B(B[2]), .Z(n219) );
    VMW_AO22 U5 ( .A(n222), .B(B[0]), .C(n223), .D(B[1]), .Z(n221) );
    VMW_OR2 U6 ( .A(B[2]), .B(n220), .Z(n224) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n223), .C(n224), .D(n221), .Z(n225) );
    VMW_NAND2 U8 ( .A(n227), .B(B[4]), .Z(n226) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n229), .C(n225), .D(n219), .Z(n228) );
    VMW_OR2 U10 ( .A(B[4]), .B(n227), .Z(n230) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n232), .C(n230), .D(n228), .Z(n231) );
    VMW_NAND2 U12 ( .A(n234), .B(B[6]), .Z(n233) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n236), .C(n231), .D(n226), .Z(n235) );
    VMW_OR2 U14 ( .A(B[6]), .B(n234), .Z(n237) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n239), .C(n237), .D(n235), .Z(n238) );
    VMW_NAND2 U16 ( .A(n241), .B(B[8]), .Z(n240) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n243), .C(n238), .D(n233), .Z(n242) );
    VMW_OR2 U18 ( .A(B[8]), .B(n241), .Z(n244) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n246), .C(n244), .D(n242), .Z(n245) );
    VMW_NAND2 U20 ( .A(n248), .B(B[10]), .Z(n247) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n250), .C(n245), .D(n240), .Z(n249) );
    VMW_NAND2 U22 ( .A(n250), .B(A[9]), .Z(n251) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n248), .C(n251), .D(n249), .Z(n252) );
    VMW_NAND2 U24 ( .A(n254), .B(B[12]), .Z(n253) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n256), .C(n252), .D(n247), .Z(n255) );
    VMW_NAND2 U26 ( .A(n256), .B(A[11]), .Z(n257) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n254), .C(n257), .D(n255), .Z(n258) );
    VMW_NAND2 U28 ( .A(n260), .B(B[14]), .Z(n259) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n262), .C(n258), .D(n253), .Z(n261) );
    VMW_NAND2 U30 ( .A(n262), .B(A[13]), .Z(n263) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n260), .C(n263), .D(n261), .Z(n264) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n265), .C(n264), .D(n259), .Z(n218) );
    VMW_INV U33 ( .A(A[12]), .Z(n254) );
    VMW_INV U34 ( .A(B[7]), .Z(n243) );
    VMW_INV U35 ( .A(A[7]), .Z(n246) );
    VMW_INV U36 ( .A(A[3]), .Z(n232) );
    VMW_INV U37 ( .A(B[3]), .Z(n229) );
    VMW_INV U38 ( .A(A[10]), .Z(n248) );
    VMW_INV U39 ( .A(B[9]), .Z(n250) );
    VMW_INV U40 ( .A(A[4]), .Z(n227) );
    VMW_INV U41 ( .A(A[8]), .Z(n241) );
    VMW_INV U42 ( .A(A[14]), .Z(n260) );
    VMW_INV U43 ( .A(B[11]), .Z(n256) );
    VMW_INV U44 ( .A(A[5]), .Z(n239) );
    VMW_INV U45 ( .A(B[5]), .Z(n236) );
    VMW_INV U46 ( .A(A[1]), .Z(n223) );
    VMW_INV U47 ( .A(B[15]), .Z(n265) );
    VMW_INV U48 ( .A(B[13]), .Z(n262) );
    VMW_INV U49 ( .A(A[6]), .Z(n234) );
    VMW_INV U50 ( .A(A[2]), .Z(n220) );
    VMW_INV U51 ( .A(A[0]), .Z(n222) );
    VMW_INV U52 ( .A(A[15]), .Z(n217) );
endmodule


module NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314;
    VMW_OAI21 U3 ( .A(B[15]), .B(n266), .C(n267), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n269), .B(B[2]), .Z(n268) );
    VMW_AO22 U5 ( .A(n271), .B(B[0]), .C(n272), .D(B[1]), .Z(n270) );
    VMW_OR2 U6 ( .A(B[2]), .B(n269), .Z(n273) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n272), .C(n273), .D(n270), .Z(n274) );
    VMW_NAND2 U8 ( .A(n276), .B(B[4]), .Z(n275) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n278), .C(n274), .D(n268), .Z(n277) );
    VMW_OR2 U10 ( .A(B[4]), .B(n276), .Z(n279) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n281), .C(n279), .D(n277), .Z(n280) );
    VMW_NAND2 U12 ( .A(n283), .B(B[6]), .Z(n282) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n285), .C(n280), .D(n275), .Z(n284) );
    VMW_OR2 U14 ( .A(B[6]), .B(n283), .Z(n286) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n288), .C(n286), .D(n284), .Z(n287) );
    VMW_NAND2 U16 ( .A(n290), .B(B[8]), .Z(n289) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n292), .C(n287), .D(n282), .Z(n291) );
    VMW_OR2 U18 ( .A(B[8]), .B(n290), .Z(n293) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n295), .C(n293), .D(n291), .Z(n294) );
    VMW_NAND2 U20 ( .A(n297), .B(B[10]), .Z(n296) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n299), .C(n294), .D(n289), .Z(n298) );
    VMW_NAND2 U22 ( .A(n299), .B(A[9]), .Z(n300) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n297), .C(n300), .D(n298), .Z(n301) );
    VMW_NAND2 U24 ( .A(n303), .B(B[12]), .Z(n302) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n305), .C(n301), .D(n296), .Z(n304) );
    VMW_NAND2 U26 ( .A(n305), .B(A[11]), .Z(n306) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n303), .C(n306), .D(n304), .Z(n307) );
    VMW_NAND2 U28 ( .A(n309), .B(B[14]), .Z(n308) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n311), .C(n307), .D(n302), .Z(n310) );
    VMW_NAND2 U30 ( .A(n311), .B(A[13]), .Z(n312) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n309), .C(n312), .D(n310), .Z(n313) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n314), .C(n313), .D(n308), .Z(n267) );
    VMW_INV U33 ( .A(A[12]), .Z(n303) );
    VMW_INV U34 ( .A(B[7]), .Z(n292) );
    VMW_INV U35 ( .A(A[7]), .Z(n295) );
    VMW_INV U36 ( .A(A[3]), .Z(n281) );
    VMW_INV U37 ( .A(B[3]), .Z(n278) );
    VMW_INV U38 ( .A(A[10]), .Z(n297) );
    VMW_INV U39 ( .A(B[9]), .Z(n299) );
    VMW_INV U40 ( .A(A[4]), .Z(n276) );
    VMW_INV U41 ( .A(A[8]), .Z(n290) );
    VMW_INV U42 ( .A(A[14]), .Z(n309) );
    VMW_INV U43 ( .A(B[11]), .Z(n305) );
    VMW_INV U44 ( .A(A[5]), .Z(n288) );
    VMW_INV U45 ( .A(B[5]), .Z(n285) );
    VMW_INV U46 ( .A(A[1]), .Z(n272) );
    VMW_INV U47 ( .A(B[15]), .Z(n314) );
    VMW_INV U48 ( .A(B[13]), .Z(n311) );
    VMW_INV U49 ( .A(A[6]), .Z(n283) );
    VMW_INV U50 ( .A(A[2]), .Z(n269) );
    VMW_INV U51 ( .A(A[0]), .Z(n271) );
    VMW_INV U52 ( .A(A[15]), .Z(n266) );
endmodule


module NodeAux_INDEGREE6_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp494[7] , \temp584[2] , n100, \OutEdge146[7] , \temp314[15] , 
        \OutEdge146[12] , \temp314[11] , \OutEdge146[3] , \temp494[3] , 
        \temp584[6] , \path[2] , \path[0] , \temp314[13] , \temp494[1] , 
        \OutEdge146[1] , \temp584[4] , \OutEdge146[8] , \temp494[8] , n132, 
        \OutEdge146[10] , \temp584[0] , \OutEdge146[5] , \temp494[5] , 
        \OutEdge146[14] , \temp584[9] , \temp220[10] , \temp220[4] , 
        \temp314[7] , \temp494[11] , \temp404[6] , \temp584[13] , 
        \temp404[11] , \temp404[2] , \temp220[0] , \temp314[3] , \temp494[15] , 
        \temp220[14] , \temp404[15] , \temp220[9] , \temp404[9] , \temp314[8] , 
        \temp220[2] , \temp404[0] , \temp314[1] , \temp584[15] , n108, 
        \temp404[13] , \temp584[11] , \temp220[12] , \temp220[6] , 
        \temp314[5] , \temp404[4] , \temp494[13] , \temp404[12] , 
        \temp584[10] , \temp220[7] , \temp314[4] , n124, \temp494[12] , 
        \temp220[13] , \temp404[5] , \temp404[8] , \temp314[9] , \temp404[1] , 
        \temp220[3] , \temp314[0] , \temp584[14] , \temp404[3] , \temp220[15] , 
        \temp220[1] , \temp314[2] , \temp494[14] , \temp220[8] , \temp404[14] , 
        n116, \temp220[5] , \temp314[6] , \temp494[10] , \temp220[11] , 
        \temp404[7] , \temp584[12] , \temp404[10] , \temp584[1] , 
        \OutEdge146[4] , \temp494[4] , \OutEdge146[15] , \temp584[8] , 
        \path[1] , \temp494[0] , \OutEdge146[0] , \temp314[12] , n92, 
        \temp584[5] , \OutEdge146[9] , \temp494[9] , \OutEdge146[11] , 
        \OutEdge146[13] , \temp494[2] , \OutEdge146[2] , \temp314[10] , 
        \path[3] , \temp584[7] , \temp584[3] , \temp314[14] , \temp494[6] , 
        \OutEdge146[6] , n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
        n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
        n800, n801, n802;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U91 ( .Z(n801) );
    VMW_PULLDOWN U92 ( .Z(n800) );
    VMW_PULLDOWN U93 ( .Z(n799) );
    VMW_PULLDOWN U94 ( .Z(n798) );
    VMW_PULLDOWN U95 ( .Z(n802) );
    VMW_PULLDOWN U96 ( .Z(n797) );
    VMW_AO22 U97 ( .A(n767), .B(\temp584[15] ), .C(InEdges[95]), .D(n768), .Z(
        \OutEdge146[15] ) );
    VMW_AO22 U98 ( .A(n767), .B(\temp584[14] ), .C(InEdges[94]), .D(n768), .Z(
        \OutEdge146[14] ) );
    VMW_AO22 U99 ( .A(n767), .B(\temp584[13] ), .C(InEdges[93]), .D(n768), .Z(
        \OutEdge146[13] ) );
    VMW_AO22 U100 ( .A(n767), .B(\temp584[12] ), .C(InEdges[92]), .D(n768), 
        .Z(\OutEdge146[12] ) );
    VMW_AO22 U101 ( .A(n767), .B(\temp584[11] ), .C(InEdges[91]), .D(n768), 
        .Z(\OutEdge146[11] ) );
    VMW_AO22 U102 ( .A(n767), .B(\temp584[10] ), .C(InEdges[90]), .D(n768), 
        .Z(\OutEdge146[10] ) );
    VMW_AO22 U103 ( .A(n767), .B(\temp584[9] ), .C(InEdges[89]), .D(n768), .Z(
        \OutEdge146[9] ) );
    VMW_AO22 U104 ( .A(n767), .B(\temp584[8] ), .C(InEdges[88]), .D(n768), .Z(
        \OutEdge146[8] ) );
    VMW_AO22 U105 ( .A(n767), .B(\temp584[7] ), .C(InEdges[87]), .D(n768), .Z(
        \OutEdge146[7] ) );
    VMW_AO22 U106 ( .A(n767), .B(\temp584[6] ), .C(InEdges[86]), .D(n768), .Z(
        \OutEdge146[6] ) );
    VMW_AO22 U107 ( .A(n767), .B(\temp584[5] ), .C(InEdges[85]), .D(n768), .Z(
        \OutEdge146[5] ) );
    VMW_AO22 U108 ( .A(n767), .B(\temp584[4] ), .C(InEdges[84]), .D(n768), .Z(
        \OutEdge146[4] ) );
    VMW_AO22 U109 ( .A(n767), .B(\temp584[3] ), .C(InEdges[83]), .D(n768), .Z(
        \OutEdge146[3] ) );
    VMW_AO22 U110 ( .A(n767), .B(\temp584[2] ), .C(InEdges[82]), .D(n768), .Z(
        \OutEdge146[2] ) );
    VMW_AO22 U111 ( .A(n767), .B(\temp584[1] ), .C(InEdges[81]), .D(n768), .Z(
        \OutEdge146[1] ) );
    VMW_AO22 U112 ( .A(n767), .B(\temp584[0] ), .C(InEdges[80]), .D(n768), .Z(
        \OutEdge146[0] ) );
    VMW_AO21 U113 ( .A(Start), .B(\path[1] ), .C(n769), .Z(n796) );
    VMW_AO22 U114 ( .A(\path[3] ), .B(Start), .C(n767), .D(n770), .Z(n795) );
    VMW_OR2 U115 ( .A(n771), .B(n768), .Z(n794) );
    VMW_NAND2 U116 ( .A(n772), .B(n773), .Z(n793) );
    VMW_AO22 U117 ( .A(InEdges[73]), .B(n124), .C(\temp494[9] ), .D(n774), .Z(
        \temp584[9] ) );
    VMW_AO22 U118 ( .A(InEdges[72]), .B(n124), .C(\temp494[8] ), .D(n774), .Z(
        \temp584[8] ) );
    VMW_AO22 U119 ( .A(InEdges[71]), .B(n124), .C(\temp494[7] ), .D(n774), .Z(
        \temp584[7] ) );
    VMW_AO22 U120 ( .A(InEdges[70]), .B(n124), .C(\temp494[6] ), .D(n774), .Z(
        \temp584[6] ) );
    VMW_AO22 U121 ( .A(InEdges[69]), .B(n124), .C(\temp494[5] ), .D(n774), .Z(
        \temp584[5] ) );
    VMW_AO22 U122 ( .A(InEdges[68]), .B(n124), .C(\temp494[4] ), .D(n774), .Z(
        \temp584[4] ) );
    VMW_AO22 U123 ( .A(InEdges[67]), .B(n124), .C(\temp494[3] ), .D(n774), .Z(
        \temp584[3] ) );
    VMW_AO22 U124 ( .A(InEdges[66]), .B(n124), .C(\temp494[2] ), .D(n774), .Z(
        \temp584[2] ) );
    VMW_AO22 U125 ( .A(InEdges[65]), .B(n124), .C(\temp494[1] ), .D(n774), .Z(
        \temp584[1] ) );
    VMW_AO22 U126 ( .A(InEdges[79]), .B(n124), .C(\temp494[15] ), .D(n774), 
        .Z(\temp584[15] ) );
    VMW_AO22 U127 ( .A(InEdges[78]), .B(n124), .C(\temp494[14] ), .D(n774), 
        .Z(\temp584[14] ) );
    VMW_AO22 U128 ( .A(InEdges[77]), .B(n124), .C(\temp494[13] ), .D(n774), 
        .Z(\temp584[13] ) );
    VMW_AO22 U129 ( .A(InEdges[76]), .B(n124), .C(\temp494[12] ), .D(n774), 
        .Z(\temp584[12] ) );
    VMW_AO22 U130 ( .A(InEdges[75]), .B(n124), .C(\temp494[11] ), .D(n774), 
        .Z(\temp584[11] ) );
    VMW_AO22 U131 ( .A(InEdges[74]), .B(n124), .C(\temp494[10] ), .D(n774), 
        .Z(\temp584[10] ) );
    VMW_AO22 U132 ( .A(InEdges[64]), .B(n124), .C(\temp494[0] ), .D(n774), .Z(
        \temp584[0] ) );
    VMW_AND4 U133 ( .A(n776), .B(n777), .C(n778), .D(n779), .Z(n775) );
    VMW_NOR2 U134 ( .A(Start), .B(n132), .Z(n767) );
    VMW_AND2 U135 ( .A(n132), .B(n780), .Z(n768) );
    VMW_OR2 U136 ( .A(n775), .B(n124), .Z(n781) );
    VMW_OAI22 U137 ( .A(\path[0] ), .B(n780), .C(n782), .D(Start), .Z(n773) );
    VMW_AND2 U138 ( .A(n774), .B(n775), .Z(n770) );
    VMW_AND3 U139 ( .A(n784), .B(n785), .C(n786), .Z(n783) );
    VMW_INV U140 ( .A(n116), .Z(n779) );
    VMW_INV U141 ( .A(n108), .Z(n777) );
    VMW_INV U142 ( .A(n124), .Z(n774) );
    VMW_OAI211 U143 ( .A(n92), .B(n100), .C(n777), .D(n779), .Z(n787) );
    VMW_AND3 U144 ( .A(n787), .B(n774), .C(n767), .Z(n769) );
    VMW_AO21 U145 ( .A(n776), .B(n92), .C(n108), .Z(n788) );
    VMW_AND4 U146 ( .A(n789), .B(n790), .C(n791), .D(n783), .Z(n792) );
    VMW_XNOR2 U147 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n785) );
    VMW_XNOR2 U148 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n784) );
    VMW_XNOR2 U149 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n786) );
    VMW_XNOR2 U150 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n790) );
    VMW_XNOR2 U151 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n789) );
    VMW_XNOR2 U152 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n791) );
    VMW_AO22 U153 ( .A(InEdges[9]), .B(n92), .C(OutEdge[9]), .D(n778), .Z(
        \temp220[9] ) );
    VMW_AO22 U154 ( .A(\temp220[9] ), .B(n776), .C(InEdges[25]), .D(n100), .Z(
        \temp314[9] ) );
    VMW_AO22 U155 ( .A(InEdges[41]), .B(n108), .C(\temp314[9] ), .D(n777), .Z(
        \temp404[9] ) );
    VMW_AO22 U156 ( .A(InEdges[57]), .B(n116), .C(\temp404[9] ), .D(n779), .Z(
        \temp494[9] ) );
    VMW_AO22 U157 ( .A(InEdges[8]), .B(n92), .C(OutEdge[8]), .D(n778), .Z(
        \temp220[8] ) );
    VMW_AO22 U158 ( .A(\temp220[8] ), .B(n776), .C(InEdges[24]), .D(n100), .Z(
        \temp314[8] ) );
    VMW_AO22 U159 ( .A(InEdges[40]), .B(n108), .C(\temp314[8] ), .D(n777), .Z(
        \temp404[8] ) );
    VMW_AO22 U160 ( .A(InEdges[56]), .B(n116), .C(\temp404[8] ), .D(n779), .Z(
        \temp494[8] ) );
    VMW_AO22 U161 ( .A(InEdges[7]), .B(n92), .C(OutEdge[7]), .D(n778), .Z(
        \temp220[7] ) );
    VMW_AO22 U162 ( .A(\temp220[7] ), .B(n776), .C(InEdges[23]), .D(n100), .Z(
        \temp314[7] ) );
    VMW_AO22 U163 ( .A(InEdges[39]), .B(n108), .C(\temp314[7] ), .D(n777), .Z(
        \temp404[7] ) );
    VMW_AO22 U164 ( .A(InEdges[55]), .B(n116), .C(\temp404[7] ), .D(n779), .Z(
        \temp494[7] ) );
    VMW_AO22 U165 ( .A(InEdges[6]), .B(n92), .C(OutEdge[6]), .D(n778), .Z(
        \temp220[6] ) );
    VMW_AO22 U166 ( .A(\temp220[6] ), .B(n776), .C(InEdges[22]), .D(n100), .Z(
        \temp314[6] ) );
    VMW_AO22 U167 ( .A(InEdges[38]), .B(n108), .C(\temp314[6] ), .D(n777), .Z(
        \temp404[6] ) );
    VMW_AO22 U168 ( .A(InEdges[54]), .B(n116), .C(\temp404[6] ), .D(n779), .Z(
        \temp494[6] ) );
    VMW_AO22 U169 ( .A(InEdges[5]), .B(n92), .C(OutEdge[5]), .D(n778), .Z(
        \temp220[5] ) );
    VMW_AO22 U170 ( .A(\temp220[5] ), .B(n776), .C(InEdges[21]), .D(n100), .Z(
        \temp314[5] ) );
    VMW_AO22 U171 ( .A(InEdges[37]), .B(n108), .C(\temp314[5] ), .D(n777), .Z(
        \temp404[5] ) );
    VMW_AO22 U172 ( .A(InEdges[53]), .B(n116), .C(\temp404[5] ), .D(n779), .Z(
        \temp494[5] ) );
    VMW_AO22 U173 ( .A(InEdges[4]), .B(n92), .C(OutEdge[4]), .D(n778), .Z(
        \temp220[4] ) );
    VMW_AO22 U174 ( .A(\temp220[4] ), .B(n776), .C(InEdges[20]), .D(n100), .Z(
        \temp314[4] ) );
    VMW_AO22 U175 ( .A(InEdges[36]), .B(n108), .C(\temp314[4] ), .D(n777), .Z(
        \temp404[4] ) );
    VMW_AO22 U176 ( .A(InEdges[52]), .B(n116), .C(\temp404[4] ), .D(n779), .Z(
        \temp494[4] ) );
    VMW_AO22 U177 ( .A(InEdges[3]), .B(n92), .C(OutEdge[3]), .D(n778), .Z(
        \temp220[3] ) );
    VMW_AO22 U178 ( .A(\temp220[3] ), .B(n776), .C(InEdges[19]), .D(n100), .Z(
        \temp314[3] ) );
    VMW_AO22 U179 ( .A(InEdges[35]), .B(n108), .C(\temp314[3] ), .D(n777), .Z(
        \temp404[3] ) );
    VMW_AO22 U180 ( .A(InEdges[51]), .B(n116), .C(\temp404[3] ), .D(n779), .Z(
        \temp494[3] ) );
    VMW_AO22 U181 ( .A(InEdges[2]), .B(n92), .C(OutEdge[2]), .D(n778), .Z(
        \temp220[2] ) );
    VMW_AO22 U182 ( .A(\temp220[2] ), .B(n776), .C(InEdges[18]), .D(n100), .Z(
        \temp314[2] ) );
    VMW_AO22 U183 ( .A(InEdges[34]), .B(n108), .C(\temp314[2] ), .D(n777), .Z(
        \temp404[2] ) );
    VMW_AO22 U184 ( .A(InEdges[50]), .B(n116), .C(\temp404[2] ), .D(n779), .Z(
        \temp494[2] ) );
    VMW_AO22 U185 ( .A(InEdges[1]), .B(n92), .C(OutEdge[1]), .D(n778), .Z(
        \temp220[1] ) );
    VMW_AO22 U186 ( .A(\temp220[1] ), .B(n776), .C(InEdges[17]), .D(n100), .Z(
        \temp314[1] ) );
    VMW_AO22 U187 ( .A(InEdges[33]), .B(n108), .C(\temp314[1] ), .D(n777), .Z(
        \temp404[1] ) );
    VMW_AO22 U188 ( .A(InEdges[49]), .B(n116), .C(\temp404[1] ), .D(n779), .Z(
        \temp494[1] ) );
    VMW_AO22 U189 ( .A(InEdges[15]), .B(n92), .C(OutEdge[15]), .D(n778), .Z(
        \temp220[15] ) );
    VMW_AO22 U190 ( .A(\temp220[15] ), .B(n776), .C(InEdges[31]), .D(n100), 
        .Z(\temp314[15] ) );
    VMW_AO22 U191 ( .A(InEdges[47]), .B(n108), .C(\temp314[15] ), .D(n777), 
        .Z(\temp404[15] ) );
    VMW_AO22 U192 ( .A(InEdges[63]), .B(n116), .C(\temp404[15] ), .D(n779), 
        .Z(\temp494[15] ) );
    VMW_AO22 U193 ( .A(InEdges[14]), .B(n92), .C(OutEdge[14]), .D(n778), .Z(
        \temp220[14] ) );
    VMW_AO22 U194 ( .A(\temp220[14] ), .B(n776), .C(InEdges[30]), .D(n100), 
        .Z(\temp314[14] ) );
    VMW_AO22 U195 ( .A(InEdges[46]), .B(n108), .C(\temp314[14] ), .D(n777), 
        .Z(\temp404[14] ) );
    VMW_AO22 U196 ( .A(InEdges[62]), .B(n116), .C(\temp404[14] ), .D(n779), 
        .Z(\temp494[14] ) );
    VMW_AO22 U197 ( .A(InEdges[13]), .B(n92), .C(OutEdge[13]), .D(n778), .Z(
        \temp220[13] ) );
    VMW_AO22 U198 ( .A(\temp220[13] ), .B(n776), .C(InEdges[29]), .D(n100), 
        .Z(\temp314[13] ) );
    VMW_AO22 U199 ( .A(InEdges[45]), .B(n108), .C(\temp314[13] ), .D(n777), 
        .Z(\temp404[13] ) );
    VMW_AO22 U200 ( .A(InEdges[61]), .B(n116), .C(\temp404[13] ), .D(n779), 
        .Z(\temp494[13] ) );
    VMW_AO22 U201 ( .A(InEdges[12]), .B(n92), .C(OutEdge[12]), .D(n778), .Z(
        \temp220[12] ) );
    VMW_AO22 U202 ( .A(\temp220[12] ), .B(n776), .C(InEdges[28]), .D(n100), 
        .Z(\temp314[12] ) );
    VMW_AO22 U203 ( .A(InEdges[44]), .B(n108), .C(\temp314[12] ), .D(n777), 
        .Z(\temp404[12] ) );
    VMW_AO22 U204 ( .A(InEdges[60]), .B(n116), .C(\temp404[12] ), .D(n779), 
        .Z(\temp494[12] ) );
    VMW_AO22 U205 ( .A(InEdges[11]), .B(n92), .C(OutEdge[11]), .D(n778), .Z(
        \temp220[11] ) );
    VMW_AO22 U206 ( .A(\temp220[11] ), .B(n776), .C(InEdges[27]), .D(n100), 
        .Z(\temp314[11] ) );
    VMW_AO22 U207 ( .A(InEdges[43]), .B(n108), .C(\temp314[11] ), .D(n777), 
        .Z(\temp404[11] ) );
    VMW_AO22 U208 ( .A(InEdges[59]), .B(n116), .C(\temp404[11] ), .D(n779), 
        .Z(\temp494[11] ) );
    VMW_AO22 U209 ( .A(InEdges[10]), .B(n92), .C(OutEdge[10]), .D(n778), .Z(
        \temp220[10] ) );
    VMW_AO22 U210 ( .A(\temp220[10] ), .B(n776), .C(InEdges[26]), .D(n100), 
        .Z(\temp314[10] ) );
    VMW_AO22 U211 ( .A(InEdges[42]), .B(n108), .C(\temp314[10] ), .D(n777), 
        .Z(\temp404[10] ) );
    VMW_AO22 U212 ( .A(InEdges[58]), .B(n116), .C(\temp404[10] ), .D(n779), 
        .Z(\temp494[10] ) );
    VMW_AO22 U213 ( .A(InEdges[0]), .B(n92), .C(OutEdge[0]), .D(n778), .Z(
        \temp220[0] ) );
    VMW_AO22 U214 ( .A(\temp220[0] ), .B(n776), .C(InEdges[16]), .D(n100), .Z(
        \temp314[0] ) );
    VMW_AO22 U215 ( .A(InEdges[32]), .B(n108), .C(\temp314[0] ), .D(n777), .Z(
        \temp404[0] ) );
    VMW_AO22 U216 ( .A(InEdges[48]), .B(n116), .C(\temp404[0] ), .D(n779), .Z(
        \temp494[0] ) );
    VMW_AO22 U217 ( .A(n781), .B(n780), .C(\path[2] ), .D(Start), .Z(n771) );
    VMW_AOI21 U218 ( .A(n779), .B(n788), .C(n124), .Z(n782) );
    VMW_INV U219 ( .A(n92), .Z(n778) );
    VMW_INV U220 ( .A(Start), .Z(n780) );
    VMW_INV U221 ( .A(n100), .Z(n776) );
    VMW_INV U222 ( .A(n768), .Z(n772) );
    VMW_BUFIZ U223 ( .A(\path[3] ), .E(n792), .Z(\PathData[3] ) );
    VMW_BUFIZ U224 ( .A(\path[1] ), .E(n792), .Z(\PathData[1] ) );
    VMW_BUFIZ U225 ( .A(\path[0] ), .E(n792), .Z(\PathData[0] ) );
    VMW_BUFIZ U226 ( .A(\path[2] ), .E(n792), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n793), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n794), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n795), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n796), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge146[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge146[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge146[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge146[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge146[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge146[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge146[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge146[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge146[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge146[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge146[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge146[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge146[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge146[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge146[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge146[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_5 lte_55_1 ( .A({\temp220[15] , 
        \temp220[14] , \temp220[13] , \temp220[12] , \temp220[11] , 
        \temp220[10] , \temp220[9] , \temp220[8] , \temp220[7] , \temp220[6] , 
        \temp220[5] , \temp220[4] , \temp220[3] , \temp220[2] , \temp220[1] , 
        \temp220[0] }), .B(InEdges[31:16]), .LEQ(n802), .TC(n802), .GE_GT(n100
        ) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_4 lte_55_5 ( .A({\temp584[15] , 
        \temp584[14] , \temp584[13] , \temp584[12] , \temp584[11] , 
        \temp584[10] , \temp584[9] , \temp584[8] , \temp584[7] , \temp584[6] , 
        \temp584[5] , \temp584[4] , \temp584[3] , \temp584[2] , \temp584[1] , 
        \temp584[0] }), .B(InEdges[95:80]), .LEQ(n801), .TC(n801), .GE_GT(n132
        ) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_3 lte_55_4 ( .A({\temp494[15] , 
        \temp494[14] , \temp494[13] , \temp494[12] , \temp494[11] , 
        \temp494[10] , \temp494[9] , \temp494[8] , \temp494[7] , \temp494[6] , 
        \temp494[5] , \temp494[4] , \temp494[3] , \temp494[2] , \temp494[1] , 
        \temp494[0] }), .B(InEdges[79:64]), .LEQ(n800), .TC(n800), .GE_GT(n124
        ) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_2 lte_55_3 ( .A({\temp404[15] , 
        \temp404[14] , \temp404[13] , \temp404[12] , \temp404[11] , 
        \temp404[10] , \temp404[9] , \temp404[8] , \temp404[7] , \temp404[6] , 
        \temp404[5] , \temp404[4] , \temp404[3] , \temp404[2] , \temp404[1] , 
        \temp404[0] }), .B(InEdges[63:48]), .LEQ(n799), .TC(n799), .GE_GT(n116
        ) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_1 lte_55_2 ( .A({\temp314[15] , 
        \temp314[14] , \temp314[13] , \temp314[12] , \temp314[11] , 
        \temp314[10] , \temp314[9] , \temp314[8] , \temp314[7] , \temp314[6] , 
        \temp314[5] , \temp314[4] , \temp314[3] , \temp314[2] , \temp314[1] , 
        \temp314[0] }), .B(InEdges[47:32]), .LEQ(n798), .TC(n798), .GE_GT(n108
        ) );
    NodeAux_INDEGREE6_SOURCE1_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n797), .TC(n797), .GE_GT(n92) );
endmodule


module NodeAux_INDEGREE0_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [-1:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge86[6] , \OutEdge86[2] , \OutEdge86[13] , 
        \OutEdge86[11] , \OutEdge86[9] , \OutEdge86[0] , \OutEdge86[15] , 
        \OutEdge86[4] , \OutEdge86[14] , \OutEdge86[5] , \OutEdge86[10] , 
        \OutEdge86[8] , \OutEdge86[1] , \OutEdge86[3] , \OutEdge86[12] , 
        \OutEdge86[7] , \path[1] , \path[3] , n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_AND2 U29 ( .A(OutEdge[15]), .B(n122), .Z(\OutEdge86[15] ) );
    VMW_OR2 U30 ( .A(OutEdge[14]), .B(Start), .Z(\OutEdge86[14] ) );
    VMW_OR2 U31 ( .A(OutEdge[13]), .B(Start), .Z(\OutEdge86[13] ) );
    VMW_OR2 U32 ( .A(OutEdge[12]), .B(Start), .Z(\OutEdge86[12] ) );
    VMW_OR2 U33 ( .A(OutEdge[11]), .B(Start), .Z(\OutEdge86[11] ) );
    VMW_OR2 U34 ( .A(OutEdge[10]), .B(Start), .Z(\OutEdge86[10] ) );
    VMW_OR2 U35 ( .A(OutEdge[9]), .B(Start), .Z(\OutEdge86[9] ) );
    VMW_OR2 U36 ( .A(OutEdge[8]), .B(Start), .Z(\OutEdge86[8] ) );
    VMW_OR2 U37 ( .A(OutEdge[7]), .B(Start), .Z(\OutEdge86[7] ) );
    VMW_OR2 U38 ( .A(OutEdge[6]), .B(Start), .Z(\OutEdge86[6] ) );
    VMW_OR2 U39 ( .A(OutEdge[5]), .B(Start), .Z(\OutEdge86[5] ) );
    VMW_OR2 U40 ( .A(OutEdge[4]), .B(Start), .Z(\OutEdge86[4] ) );
    VMW_OR2 U41 ( .A(OutEdge[3]), .B(Start), .Z(\OutEdge86[3] ) );
    VMW_OR2 U42 ( .A(OutEdge[2]), .B(Start), .Z(\OutEdge86[2] ) );
    VMW_OR2 U43 ( .A(OutEdge[1]), .B(Start), .Z(\OutEdge86[1] ) );
    VMW_OR2 U44 ( .A(OutEdge[0]), .B(Start), .Z(\OutEdge86[0] ) );
    VMW_OR2 U45 ( .A(n122), .B(\path[1] ), .Z(n134) );
    VMW_OR2 U46 ( .A(n122), .B(\path[3] ), .Z(n133) );
    VMW_OR2 U47 ( .A(n122), .B(\path[2] ), .Z(n132) );
    VMW_OR2 U48 ( .A(n122), .B(\path[0] ), .Z(n131) );
    VMW_AND3 U49 ( .A(n124), .B(n125), .C(n126), .Z(n123) );
    VMW_AND4 U50 ( .A(n127), .B(n128), .C(n129), .D(n123), .Z(n130) );
    VMW_XNOR2 U51 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n125) );
    VMW_XNOR2 U52 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n124) );
    VMW_XNOR2 U53 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n126) );
    VMW_XNOR2 U54 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n128) );
    VMW_XNOR2 U55 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n127) );
    VMW_XNOR2 U56 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n129) );
    VMW_INV U57 ( .A(Start), .Z(n122) );
    VMW_BUFIZ U58 ( .A(\path[3] ), .E(n130), .Z(\PathData[3] ) );
    VMW_BUFIZ U59 ( .A(\path[1] ), .E(n130), .Z(\PathData[1] ) );
    VMW_BUFIZ U60 ( .A(\path[0] ), .E(n130), .Z(\PathData[0] ) );
    VMW_BUFIZ U61 ( .A(\path[2] ), .E(n130), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n131), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n132), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n133), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n134), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge86[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge86[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge86[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge86[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge86[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge86[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge86[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge86[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge86[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge86[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge86[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge86[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge86[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge86[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge86[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge86[0] ), .CP(Clk), .Q(OutEdge[0]) );
endmodule


module NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , \path[3] , n267, n268, 
        n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
        n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
        n293, n294, n295, n296, n297;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n297) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(n268), .D(InEdges[15]), .Z(
        \OutEdge96[15] ) );
    VMW_OR2 U48 ( .A(n269), .B(Start), .Z(\OutEdge96[14] ) );
    VMW_OR2 U49 ( .A(n270), .B(Start), .Z(\OutEdge96[13] ) );
    VMW_OR2 U50 ( .A(n271), .B(Start), .Z(\OutEdge96[12] ) );
    VMW_OR2 U51 ( .A(n272), .B(Start), .Z(\OutEdge96[11] ) );
    VMW_OR2 U52 ( .A(n273), .B(Start), .Z(\OutEdge96[10] ) );
    VMW_OR2 U53 ( .A(n274), .B(Start), .Z(\OutEdge96[9] ) );
    VMW_OR2 U54 ( .A(n275), .B(Start), .Z(\OutEdge96[8] ) );
    VMW_OR2 U55 ( .A(n276), .B(Start), .Z(\OutEdge96[7] ) );
    VMW_OR2 U56 ( .A(n277), .B(Start), .Z(\OutEdge96[6] ) );
    VMW_OR2 U57 ( .A(n278), .B(Start), .Z(\OutEdge96[5] ) );
    VMW_OR2 U58 ( .A(n279), .B(Start), .Z(\OutEdge96[4] ) );
    VMW_OR2 U59 ( .A(n280), .B(Start), .Z(\OutEdge96[3] ) );
    VMW_OR2 U60 ( .A(n281), .B(Start), .Z(\OutEdge96[2] ) );
    VMW_OR2 U61 ( .A(n282), .B(Start), .Z(\OutEdge96[1] ) );
    VMW_OR2 U62 ( .A(n283), .B(Start), .Z(\OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(\path[1] ), .B(Start), .C(n267), .Z(n296) );
    VMW_AO21 U64 ( .A(Start), .B(\path[3] ), .C(n267), .Z(n295) );
    VMW_AO21 U65 ( .A(\path[2] ), .B(Start), .C(n267), .Z(n294) );
    VMW_AO21 U66 ( .A(\path[0] ), .B(Start), .C(n267), .Z(n293) );
    VMW_INV U67 ( .A(n82), .Z(n284) );
    VMW_NOR2 U68 ( .A(Start), .B(n82), .Z(n267) );
    VMW_AND3 U69 ( .A(n286), .B(n287), .C(n288), .Z(n285) );
    VMW_NOR2 U70 ( .A(Start), .B(n284), .Z(n268) );
    VMW_AND4 U71 ( .A(n289), .B(n290), .C(n291), .D(n285), .Z(n292) );
    VMW_XNOR2 U72 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n287) );
    VMW_XNOR2 U73 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n286) );
    VMW_XNOR2 U74 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n288) );
    VMW_XNOR2 U75 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n290) );
    VMW_XNOR2 U76 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n289) );
    VMW_XNOR2 U77 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n291) );
    VMW_AO22 U78 ( .A(InEdges[9]), .B(n82), .C(OutEdge[9]), .D(n284), .Z(n274)
         );
    VMW_AO22 U79 ( .A(InEdges[8]), .B(n82), .C(OutEdge[8]), .D(n284), .Z(n275)
         );
    VMW_AO22 U80 ( .A(InEdges[7]), .B(n82), .C(OutEdge[7]), .D(n284), .Z(n276)
         );
    VMW_AO22 U81 ( .A(InEdges[6]), .B(n82), .C(OutEdge[6]), .D(n284), .Z(n277)
         );
    VMW_AO22 U82 ( .A(InEdges[5]), .B(n82), .C(OutEdge[5]), .D(n284), .Z(n278)
         );
    VMW_AO22 U83 ( .A(InEdges[4]), .B(n82), .C(OutEdge[4]), .D(n284), .Z(n279)
         );
    VMW_AO22 U84 ( .A(InEdges[3]), .B(n82), .C(OutEdge[3]), .D(n284), .Z(n280)
         );
    VMW_AO22 U85 ( .A(InEdges[2]), .B(n82), .C(OutEdge[2]), .D(n284), .Z(n281)
         );
    VMW_AO22 U86 ( .A(InEdges[1]), .B(n82), .C(OutEdge[1]), .D(n284), .Z(n282)
         );
    VMW_AO22 U87 ( .A(InEdges[14]), .B(n82), .C(OutEdge[14]), .D(n284), .Z(
        n269) );
    VMW_AO22 U88 ( .A(InEdges[13]), .B(n82), .C(OutEdge[13]), .D(n284), .Z(
        n270) );
    VMW_AO22 U89 ( .A(InEdges[12]), .B(n82), .C(OutEdge[12]), .D(n284), .Z(
        n271) );
    VMW_AO22 U90 ( .A(InEdges[11]), .B(n82), .C(OutEdge[11]), .D(n284), .Z(
        n272) );
    VMW_AO22 U91 ( .A(InEdges[10]), .B(n82), .C(OutEdge[10]), .D(n284), .Z(
        n273) );
    VMW_AO22 U92 ( .A(InEdges[0]), .B(n82), .C(OutEdge[0]), .D(n284), .Z(n283)
         );
    VMW_BUFIZ U93 ( .A(\path[3] ), .E(n292), .Z(\PathData[3] ) );
    VMW_BUFIZ U94 ( .A(\path[1] ), .E(n292), .Z(\PathData[1] ) );
    VMW_BUFIZ U95 ( .A(\path[0] ), .E(n292), .Z(\PathData[0] ) );
    VMW_BUFIZ U96 ( .A(\path[2] ), .E(n292), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n293), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n294), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n295), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n296), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n297), .TC(n297), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \path[3] , 
        \OutEdge106[0] , \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, 
        n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
        n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
        n392, n393, n394, n395, n396, n397, n398, n399, n400, n401;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n400) );
    VMW_PULLDOWN U56 ( .Z(n401) );
    VMW_NOR2 U57 ( .A(Start), .B(n367), .Z(\OutEdge106[15] ) );
    VMW_NAND2 U58 ( .A(n368), .B(n369), .Z(\OutEdge106[14] ) );
    VMW_NAND2 U59 ( .A(n370), .B(n369), .Z(\OutEdge106[13] ) );
    VMW_NAND2 U60 ( .A(n371), .B(n369), .Z(\OutEdge106[12] ) );
    VMW_NAND2 U61 ( .A(n372), .B(n369), .Z(\OutEdge106[11] ) );
    VMW_NAND2 U62 ( .A(n373), .B(n369), .Z(\OutEdge106[10] ) );
    VMW_NAND2 U63 ( .A(n374), .B(n369), .Z(\OutEdge106[9] ) );
    VMW_NAND2 U64 ( .A(n375), .B(n369), .Z(\OutEdge106[8] ) );
    VMW_NAND2 U65 ( .A(n376), .B(n369), .Z(\OutEdge106[7] ) );
    VMW_NAND2 U66 ( .A(n377), .B(n369), .Z(\OutEdge106[6] ) );
    VMW_NAND2 U67 ( .A(n378), .B(n369), .Z(\OutEdge106[5] ) );
    VMW_NAND2 U68 ( .A(n379), .B(n369), .Z(\OutEdge106[4] ) );
    VMW_NAND2 U69 ( .A(n380), .B(n369), .Z(\OutEdge106[3] ) );
    VMW_NAND2 U70 ( .A(n381), .B(n369), .Z(\OutEdge106[2] ) );
    VMW_NAND2 U71 ( .A(n382), .B(n369), .Z(\OutEdge106[1] ) );
    VMW_NAND2 U72 ( .A(n383), .B(n369), .Z(\OutEdge106[0] ) );
    VMW_AO21 U73 ( .A(Start), .B(\path[1] ), .C(n384), .Z(n399) );
    VMW_AO21 U74 ( .A(\path[3] ), .B(Start), .C(n384), .Z(n398) );
    VMW_AO21 U75 ( .A(Start), .B(\path[2] ), .C(n384), .Z(n397) );
    VMW_OR2 U76 ( .A(n386), .B(n92), .Z(n385) );
    VMW_AO22 U77 ( .A(OutEdge[15]), .B(n386), .C(InEdges[15]), .D(n84), .Z(
        \temp180[15] ) );
    VMW_OAI22 U78 ( .A(\path[0] ), .B(n369), .C(n385), .D(Start), .Z(n387) );
    VMW_MUX2I U79 ( .A(\temp180[15] ), .B(InEdges[31]), .S(n92), .Z(n367) );
    VMW_AND3 U80 ( .A(n389), .B(n390), .C(n391), .Z(n388) );
    VMW_NOR3 U81 ( .A(Start), .B(n84), .C(n92), .Z(n384) );
    VMW_AND4 U82 ( .A(n392), .B(n393), .C(n394), .D(n388), .Z(n395) );
    VMW_XNOR2 U83 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n390) );
    VMW_XNOR2 U84 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n389) );
    VMW_XNOR2 U85 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n391) );
    VMW_XNOR2 U86 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n393) );
    VMW_XNOR2 U87 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n392) );
    VMW_XNOR2 U88 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n394) );
    VMW_AO22 U89 ( .A(OutEdge[9]), .B(n386), .C(InEdges[9]), .D(n84), .Z(
        \temp180[9] ) );
    VMW_AO22 U90 ( .A(OutEdge[8]), .B(n386), .C(InEdges[8]), .D(n84), .Z(
        \temp180[8] ) );
    VMW_AO22 U91 ( .A(OutEdge[7]), .B(n386), .C(InEdges[7]), .D(n84), .Z(
        \temp180[7] ) );
    VMW_AO22 U92 ( .A(OutEdge[6]), .B(n386), .C(InEdges[6]), .D(n84), .Z(
        \temp180[6] ) );
    VMW_AO22 U93 ( .A(OutEdge[5]), .B(n386), .C(InEdges[5]), .D(n84), .Z(
        \temp180[5] ) );
    VMW_AO22 U94 ( .A(OutEdge[4]), .B(n386), .C(InEdges[4]), .D(n84), .Z(
        \temp180[4] ) );
    VMW_AO22 U95 ( .A(OutEdge[3]), .B(n386), .C(InEdges[3]), .D(n84), .Z(
        \temp180[3] ) );
    VMW_AO22 U96 ( .A(OutEdge[2]), .B(n386), .C(InEdges[2]), .D(n84), .Z(
        \temp180[2] ) );
    VMW_AO22 U97 ( .A(OutEdge[1]), .B(n386), .C(InEdges[1]), .D(n84), .Z(
        \temp180[1] ) );
    VMW_AO22 U98 ( .A(OutEdge[14]), .B(n386), .C(InEdges[14]), .D(n84), .Z(
        \temp180[14] ) );
    VMW_AO22 U99 ( .A(OutEdge[13]), .B(n386), .C(InEdges[13]), .D(n84), .Z(
        \temp180[13] ) );
    VMW_AO22 U100 ( .A(OutEdge[12]), .B(n386), .C(InEdges[12]), .D(n84), .Z(
        \temp180[12] ) );
    VMW_AO22 U101 ( .A(OutEdge[11]), .B(n386), .C(InEdges[11]), .D(n84), .Z(
        \temp180[11] ) );
    VMW_AO22 U102 ( .A(OutEdge[10]), .B(n386), .C(InEdges[10]), .D(n84), .Z(
        \temp180[10] ) );
    VMW_AO22 U103 ( .A(OutEdge[0]), .B(n386), .C(InEdges[0]), .D(n84), .Z(
        \temp180[0] ) );
    VMW_MUX2I U104 ( .A(\temp180[9] ), .B(InEdges[25]), .S(n92), .Z(n374) );
    VMW_MUX2I U105 ( .A(\temp180[8] ), .B(InEdges[24]), .S(n92), .Z(n375) );
    VMW_MUX2I U106 ( .A(\temp180[7] ), .B(InEdges[23]), .S(n92), .Z(n376) );
    VMW_MUX2I U107 ( .A(\temp180[6] ), .B(InEdges[22]), .S(n92), .Z(n377) );
    VMW_MUX2I U108 ( .A(\temp180[5] ), .B(InEdges[21]), .S(n92), .Z(n378) );
    VMW_MUX2I U109 ( .A(\temp180[4] ), .B(InEdges[20]), .S(n92), .Z(n379) );
    VMW_MUX2I U110 ( .A(\temp180[3] ), .B(InEdges[19]), .S(n92), .Z(n380) );
    VMW_MUX2I U111 ( .A(\temp180[2] ), .B(InEdges[18]), .S(n92), .Z(n381) );
    VMW_MUX2I U112 ( .A(\temp180[1] ), .B(InEdges[17]), .S(n92), .Z(n382) );
    VMW_MUX2I U113 ( .A(\temp180[14] ), .B(InEdges[30]), .S(n92), .Z(n368) );
    VMW_MUX2I U114 ( .A(\temp180[13] ), .B(InEdges[29]), .S(n92), .Z(n370) );
    VMW_MUX2I U115 ( .A(\temp180[12] ), .B(InEdges[28]), .S(n92), .Z(n371) );
    VMW_MUX2I U116 ( .A(\temp180[11] ), .B(InEdges[27]), .S(n92), .Z(n372) );
    VMW_MUX2I U117 ( .A(\temp180[10] ), .B(InEdges[26]), .S(n92), .Z(n373) );
    VMW_MUX2I U118 ( .A(\temp180[0] ), .B(InEdges[16]), .S(n92), .Z(n383) );
    VMW_INV U119 ( .A(n84), .Z(n386) );
    VMW_INV U120 ( .A(Start), .Z(n369) );
    VMW_INV U121 ( .A(n387), .Z(n396) );
    VMW_BUFIZ U122 ( .A(\path[3] ), .E(n395), .Z(\PathData[3] ) );
    VMW_BUFIZ U123 ( .A(\path[1] ), .E(n395), .Z(\PathData[1] ) );
    VMW_BUFIZ U124 ( .A(\path[0] ), .E(n395), .Z(\PathData[0] ) );
    VMW_BUFIZ U125 ( .A(\path[2] ), .E(n395), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n396), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n397), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n398), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n399), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n401), .TC(n401), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n400), .TC(n400), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, 
        n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n104), .B(B[12]), .Z(n103) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n96), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n104), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n103), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n104) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n121), .B(B[0]), .C(n122), .D(B[1]), .Z(n120) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n123) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n122), .C(n123), .D(n120), .Z(n124) );
    VMW_NAND2 U8 ( .A(n126), .B(B[4]), .Z(n125) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n128), .C(n124), .D(n118), .Z(n127) );
    VMW_OR2 U10 ( .A(B[4]), .B(n126), .Z(n129) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n131), .C(n129), .D(n127), .Z(n130) );
    VMW_NAND2 U12 ( .A(n133), .B(B[6]), .Z(n132) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n135), .C(n130), .D(n125), .Z(n134) );
    VMW_OR2 U14 ( .A(B[6]), .B(n133), .Z(n136) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n138), .C(n136), .D(n134), .Z(n137) );
    VMW_NAND2 U16 ( .A(n140), .B(B[8]), .Z(n139) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n142), .C(n137), .D(n132), .Z(n141) );
    VMW_OR2 U18 ( .A(B[8]), .B(n140), .Z(n143) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n145), .C(n143), .D(n141), .Z(n144) );
    VMW_NAND2 U20 ( .A(n147), .B(B[10]), .Z(n146) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n149), .C(n144), .D(n139), .Z(n148) );
    VMW_NAND2 U22 ( .A(n149), .B(A[9]), .Z(n150) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n147), .C(n150), .D(n148), .Z(n151) );
    VMW_NAND2 U24 ( .A(n153), .B(B[12]), .Z(n152) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n155), .C(n151), .D(n146), .Z(n154) );
    VMW_NAND2 U26 ( .A(n155), .B(A[11]), .Z(n156) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n153), .C(n156), .D(n154), .Z(n157) );
    VMW_NAND2 U28 ( .A(n159), .B(B[14]), .Z(n158) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n161), .C(n157), .D(n152), .Z(n160) );
    VMW_NAND2 U30 ( .A(n161), .B(A[13]), .Z(n162) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n159), .C(n162), .D(n160), .Z(n163) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n164), .C(n163), .D(n158), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n153) );
    VMW_INV U34 ( .A(B[7]), .Z(n142) );
    VMW_INV U35 ( .A(A[7]), .Z(n145) );
    VMW_INV U36 ( .A(A[3]), .Z(n131) );
    VMW_INV U37 ( .A(B[3]), .Z(n128) );
    VMW_INV U38 ( .A(A[10]), .Z(n147) );
    VMW_INV U39 ( .A(B[9]), .Z(n149) );
    VMW_INV U40 ( .A(A[4]), .Z(n126) );
    VMW_INV U41 ( .A(A[8]), .Z(n140) );
    VMW_INV U42 ( .A(A[14]), .Z(n159) );
    VMW_INV U43 ( .A(B[11]), .Z(n155) );
    VMW_INV U44 ( .A(A[5]), .Z(n138) );
    VMW_INV U45 ( .A(B[5]), .Z(n135) );
    VMW_INV U46 ( .A(A[1]), .Z(n122) );
    VMW_INV U47 ( .A(B[15]), .Z(n164) );
    VMW_INV U48 ( .A(B[13]), .Z(n161) );
    VMW_INV U49 ( .A(A[6]), .Z(n133) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n121) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp284[0] , \OutEdge116[6] , \temp284[9] , \temp284[11] , 
        \temp190[2] , \OutEdge116[2] , \temp284[4] , \temp190[6] , 
        \temp284[15] , \path[2] , \OutEdge116[9] , \path[0] , \temp190[4] , 
        \OutEdge116[0] , \temp284[6] , \temp284[13] , \temp190[0] , 
        \temp284[2] , \OutEdge116[4] , \temp190[9] , \temp190[10] , 
        \OutEdge116[11] , \OutEdge116[15] , \temp190[14] , \OutEdge116[13] , 
        \temp190[12] , n94, \OutEdge116[12] , \temp190[13] , n86, 
        \OutEdge116[14] , \temp190[15] , \temp190[11] , \OutEdge116[10] , 
        \temp284[12] , \temp190[1] , \temp284[3] , \OutEdge116[5] , 
        \temp190[8] , \path[1] , \OutEdge116[8] , \temp190[5] , 
        \OutEdge116[1] , \temp284[7] , n102, \OutEdge116[3] , \temp284[5] , 
        \temp190[7] , \temp284[14] , \path[3] , \temp284[1] , \OutEdge116[7] , 
        \temp284[8] , \temp284[10] , \temp190[3] , n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U64 ( .Z(n504) );
    VMW_PULLDOWN U65 ( .Z(n506) );
    VMW_PULLDOWN U66 ( .Z(n505) );
    VMW_NOR2 U67 ( .A(Start), .B(n467), .Z(\OutEdge116[15] ) );
    VMW_NAND2 U68 ( .A(n468), .B(n469), .Z(\OutEdge116[14] ) );
    VMW_NAND2 U69 ( .A(n470), .B(n469), .Z(\OutEdge116[13] ) );
    VMW_NAND2 U70 ( .A(n471), .B(n469), .Z(\OutEdge116[12] ) );
    VMW_NAND2 U71 ( .A(n472), .B(n469), .Z(\OutEdge116[11] ) );
    VMW_NAND2 U72 ( .A(n473), .B(n469), .Z(\OutEdge116[10] ) );
    VMW_NAND2 U73 ( .A(n474), .B(n469), .Z(\OutEdge116[9] ) );
    VMW_NAND2 U74 ( .A(n475), .B(n469), .Z(\OutEdge116[8] ) );
    VMW_NAND2 U75 ( .A(n476), .B(n469), .Z(\OutEdge116[7] ) );
    VMW_NAND2 U76 ( .A(n477), .B(n469), .Z(\OutEdge116[6] ) );
    VMW_NAND2 U77 ( .A(n478), .B(n469), .Z(\OutEdge116[5] ) );
    VMW_NAND2 U78 ( .A(n479), .B(n469), .Z(\OutEdge116[4] ) );
    VMW_NAND2 U79 ( .A(n480), .B(n469), .Z(\OutEdge116[3] ) );
    VMW_NAND2 U80 ( .A(n481), .B(n469), .Z(\OutEdge116[2] ) );
    VMW_NAND2 U81 ( .A(n482), .B(n469), .Z(\OutEdge116[1] ) );
    VMW_NAND2 U82 ( .A(n483), .B(n469), .Z(\OutEdge116[0] ) );
    VMW_OR2 U83 ( .A(n484), .B(n485), .Z(n503) );
    VMW_AO21 U84 ( .A(\path[3] ), .B(Start), .C(n486), .Z(n502) );
    VMW_AO21 U85 ( .A(Start), .B(\path[2] ), .C(n486), .Z(n501) );
    VMW_AO22 U86 ( .A(InEdges[31]), .B(n94), .C(\temp190[15] ), .D(n487), .Z(
        \temp284[15] ) );
    VMW_INV U87 ( .A(Start), .Z(n469) );
    VMW_AND3 U88 ( .A(n469), .B(n488), .C(n487), .Z(n485) );
    VMW_OAI22 U89 ( .A(\path[0] ), .B(n469), .C(n490), .D(Start), .Z(n489) );
    VMW_MUX2I U90 ( .A(\temp284[15] ), .B(InEdges[47]), .S(n102), .Z(n467) );
    VMW_AND3 U91 ( .A(n492), .B(n493), .C(n494), .Z(n491) );
    VMW_NOR2 U92 ( .A(n102), .B(n495), .Z(n486) );
    VMW_AND4 U93 ( .A(n496), .B(n497), .C(n498), .D(n491), .Z(n499) );
    VMW_XNOR2 U94 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n493) );
    VMW_XNOR2 U95 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n492) );
    VMW_XNOR2 U96 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n494) );
    VMW_XNOR2 U97 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n497) );
    VMW_XNOR2 U98 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n496) );
    VMW_XNOR2 U99 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n498) );
    VMW_AO22 U100 ( .A(OutEdge[9]), .B(n488), .C(InEdges[9]), .D(n86), .Z(
        \temp190[9] ) );
    VMW_AO22 U101 ( .A(InEdges[25]), .B(n94), .C(\temp190[9] ), .D(n487), .Z(
        \temp284[9] ) );
    VMW_AO22 U102 ( .A(OutEdge[8]), .B(n488), .C(InEdges[8]), .D(n86), .Z(
        \temp190[8] ) );
    VMW_AO22 U103 ( .A(InEdges[24]), .B(n94), .C(\temp190[8] ), .D(n487), .Z(
        \temp284[8] ) );
    VMW_AO22 U104 ( .A(OutEdge[7]), .B(n488), .C(InEdges[7]), .D(n86), .Z(
        \temp190[7] ) );
    VMW_AO22 U105 ( .A(InEdges[23]), .B(n94), .C(\temp190[7] ), .D(n487), .Z(
        \temp284[7] ) );
    VMW_AO22 U106 ( .A(OutEdge[6]), .B(n488), .C(InEdges[6]), .D(n86), .Z(
        \temp190[6] ) );
    VMW_AO22 U107 ( .A(InEdges[22]), .B(n94), .C(\temp190[6] ), .D(n487), .Z(
        \temp284[6] ) );
    VMW_AO22 U108 ( .A(OutEdge[5]), .B(n488), .C(InEdges[5]), .D(n86), .Z(
        \temp190[5] ) );
    VMW_AO22 U109 ( .A(InEdges[21]), .B(n94), .C(\temp190[5] ), .D(n487), .Z(
        \temp284[5] ) );
    VMW_AO22 U110 ( .A(OutEdge[4]), .B(n488), .C(InEdges[4]), .D(n86), .Z(
        \temp190[4] ) );
    VMW_AO22 U111 ( .A(InEdges[20]), .B(n94), .C(\temp190[4] ), .D(n487), .Z(
        \temp284[4] ) );
    VMW_AO22 U112 ( .A(OutEdge[3]), .B(n488), .C(InEdges[3]), .D(n86), .Z(
        \temp190[3] ) );
    VMW_AO22 U113 ( .A(InEdges[19]), .B(n94), .C(\temp190[3] ), .D(n487), .Z(
        \temp284[3] ) );
    VMW_AO22 U114 ( .A(OutEdge[2]), .B(n488), .C(InEdges[2]), .D(n86), .Z(
        \temp190[2] ) );
    VMW_AO22 U115 ( .A(InEdges[18]), .B(n94), .C(\temp190[2] ), .D(n487), .Z(
        \temp284[2] ) );
    VMW_AO22 U116 ( .A(OutEdge[1]), .B(n488), .C(InEdges[1]), .D(n86), .Z(
        \temp190[1] ) );
    VMW_AO22 U117 ( .A(InEdges[17]), .B(n94), .C(\temp190[1] ), .D(n487), .Z(
        \temp284[1] ) );
    VMW_AO22 U118 ( .A(OutEdge[15]), .B(n488), .C(InEdges[15]), .D(n86), .Z(
        \temp190[15] ) );
    VMW_AO22 U119 ( .A(OutEdge[14]), .B(n488), .C(InEdges[14]), .D(n86), .Z(
        \temp190[14] ) );
    VMW_AO22 U120 ( .A(InEdges[30]), .B(n94), .C(\temp190[14] ), .D(n487), .Z(
        \temp284[14] ) );
    VMW_AO22 U121 ( .A(OutEdge[13]), .B(n488), .C(InEdges[13]), .D(n86), .Z(
        \temp190[13] ) );
    VMW_AO22 U122 ( .A(InEdges[29]), .B(n94), .C(\temp190[13] ), .D(n487), .Z(
        \temp284[13] ) );
    VMW_AO22 U123 ( .A(OutEdge[12]), .B(n488), .C(InEdges[12]), .D(n86), .Z(
        \temp190[12] ) );
    VMW_AO22 U124 ( .A(InEdges[28]), .B(n94), .C(\temp190[12] ), .D(n487), .Z(
        \temp284[12] ) );
    VMW_AO22 U125 ( .A(OutEdge[11]), .B(n488), .C(InEdges[11]), .D(n86), .Z(
        \temp190[11] ) );
    VMW_AO22 U126 ( .A(InEdges[27]), .B(n94), .C(\temp190[11] ), .D(n487), .Z(
        \temp284[11] ) );
    VMW_AO22 U127 ( .A(OutEdge[10]), .B(n488), .C(InEdges[10]), .D(n86), .Z(
        \temp190[10] ) );
    VMW_AO22 U128 ( .A(InEdges[26]), .B(n94), .C(\temp190[10] ), .D(n487), .Z(
        \temp284[10] ) );
    VMW_AO22 U129 ( .A(OutEdge[0]), .B(n488), .C(InEdges[0]), .D(n86), .Z(
        \temp190[0] ) );
    VMW_AO22 U130 ( .A(InEdges[16]), .B(n94), .C(\temp190[0] ), .D(n487), .Z(
        \temp284[0] ) );
    VMW_AO22 U131 ( .A(\path[1] ), .B(Start), .C(n102), .D(n469), .Z(n484) );
    VMW_AOI21 U132 ( .A(n487), .B(n86), .C(n102), .Z(n490) );
    VMW_MUX2I U133 ( .A(\temp284[9] ), .B(InEdges[41]), .S(n102), .Z(n474) );
    VMW_MUX2I U134 ( .A(\temp284[8] ), .B(InEdges[40]), .S(n102), .Z(n475) );
    VMW_MUX2I U135 ( .A(\temp284[7] ), .B(InEdges[39]), .S(n102), .Z(n476) );
    VMW_MUX2I U136 ( .A(\temp284[6] ), .B(InEdges[38]), .S(n102), .Z(n477) );
    VMW_MUX2I U137 ( .A(\temp284[5] ), .B(InEdges[37]), .S(n102), .Z(n478) );
    VMW_MUX2I U138 ( .A(\temp284[4] ), .B(InEdges[36]), .S(n102), .Z(n479) );
    VMW_MUX2I U139 ( .A(\temp284[3] ), .B(InEdges[35]), .S(n102), .Z(n480) );
    VMW_MUX2I U140 ( .A(\temp284[2] ), .B(InEdges[34]), .S(n102), .Z(n481) );
    VMW_MUX2I U141 ( .A(\temp284[1] ), .B(InEdges[33]), .S(n102), .Z(n482) );
    VMW_MUX2I U142 ( .A(\temp284[14] ), .B(InEdges[46]), .S(n102), .Z(n468) );
    VMW_MUX2I U143 ( .A(\temp284[13] ), .B(InEdges[45]), .S(n102), .Z(n470) );
    VMW_MUX2I U144 ( .A(\temp284[12] ), .B(InEdges[44]), .S(n102), .Z(n471) );
    VMW_MUX2I U145 ( .A(\temp284[11] ), .B(InEdges[43]), .S(n102), .Z(n472) );
    VMW_MUX2I U146 ( .A(\temp284[10] ), .B(InEdges[42]), .S(n102), .Z(n473) );
    VMW_MUX2I U147 ( .A(\temp284[0] ), .B(InEdges[32]), .S(n102), .Z(n483) );
    VMW_INV U148 ( .A(n94), .Z(n487) );
    VMW_INV U149 ( .A(n86), .Z(n488) );
    VMW_INV U150 ( .A(n485), .Z(n495) );
    VMW_INV U151 ( .A(n489), .Z(n500) );
    VMW_BUFIZ U152 ( .A(\path[3] ), .E(n499), .Z(\PathData[3] ) );
    VMW_BUFIZ U153 ( .A(\path[1] ), .E(n499), .Z(\PathData[1] ) );
    VMW_BUFIZ U154 ( .A(\path[0] ), .E(n499), .Z(\PathData[0] ) );
    VMW_BUFIZ U155 ( .A(\path[2] ), .E(n499), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n500), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n501), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n502), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n503), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge116[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge116[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge116[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge116[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge116[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge116[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge116[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge116[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge116[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge116[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge116[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge116[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge116[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge116[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge116[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge116[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp190[15] , 
        \temp190[14] , \temp190[13] , \temp190[12] , \temp190[11] , 
        \temp190[10] , \temp190[9] , \temp190[8] , \temp190[7] , \temp190[6] , 
        \temp190[5] , \temp190[4] , \temp190[3] , \temp190[2] , \temp190[1] , 
        \temp190[0] }), .B(InEdges[31:16]), .LEQ(n506), .TC(n506), .GE_GT(n94)
         );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n505), .TC(n505), .GE_GT(n86) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 lte_55_2 ( .A({\temp284[15] , 
        \temp284[14] , \temp284[13] , \temp284[12] , \temp284[11] , 
        \temp284[10] , \temp284[9] , \temp284[8] , \temp284[7] , \temp284[6] , 
        \temp284[5] , \temp284[4] , \temp284[3] , \temp284[2] , \temp284[1] , 
        \temp284[0] }), .B(InEdges[47:32]), .LEQ(n504), .TC(n504), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, 
        n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, 
        n108, n109, n110, n111, n113, n114, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n95), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n113), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n113), .B(A[13]), .Z(n114) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n114), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n113) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n129), .C(n125), .D(n119), .Z(n128) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n130) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n132), .C(n130), .D(n128), .Z(n131) );
    VMW_NAND2 U12 ( .A(n134), .B(B[6]), .Z(n133) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n136), .C(n131), .D(n126), .Z(n135) );
    VMW_OR2 U14 ( .A(B[6]), .B(n134), .Z(n137) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n139), .C(n137), .D(n135), .Z(n138) );
    VMW_NAND2 U16 ( .A(n141), .B(B[8]), .Z(n140) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n143), .C(n138), .D(n133), .Z(n142) );
    VMW_OR2 U18 ( .A(B[8]), .B(n141), .Z(n144) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n146), .C(n144), .D(n142), .Z(n145) );
    VMW_NAND2 U20 ( .A(n148), .B(B[10]), .Z(n147) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n150), .C(n145), .D(n140), .Z(n149) );
    VMW_NAND2 U22 ( .A(n150), .B(A[9]), .Z(n151) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n148), .C(n151), .D(n149), .Z(n152) );
    VMW_NAND2 U24 ( .A(n154), .B(B[12]), .Z(n153) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n156), .C(n152), .D(n147), .Z(n155) );
    VMW_NAND2 U26 ( .A(n156), .B(A[11]), .Z(n157) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n154), .C(n157), .D(n155), .Z(n158) );
    VMW_NAND2 U28 ( .A(n160), .B(B[14]), .Z(n159) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n162), .C(n158), .D(n153), .Z(n161) );
    VMW_NAND2 U30 ( .A(n162), .B(A[13]), .Z(n163) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n160), .C(n163), .D(n161), .Z(n164) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n165), .C(n164), .D(n159), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n154) );
    VMW_INV U34 ( .A(B[7]), .Z(n143) );
    VMW_INV U35 ( .A(A[7]), .Z(n146) );
    VMW_INV U36 ( .A(A[3]), .Z(n132) );
    VMW_INV U37 ( .A(B[3]), .Z(n129) );
    VMW_INV U38 ( .A(A[10]), .Z(n148) );
    VMW_INV U39 ( .A(B[9]), .Z(n150) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n141) );
    VMW_INV U42 ( .A(A[14]), .Z(n160) );
    VMW_INV U43 ( .A(B[11]), .Z(n156) );
    VMW_INV U44 ( .A(A[5]), .Z(n139) );
    VMW_INV U45 ( .A(B[5]), .Z(n136) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n165) );
    VMW_INV U48 ( .A(B[13]), .Z(n162) );
    VMW_INV U49 ( .A(A[6]), .Z(n134) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
        n213, n214;
    VMW_OAI21 U3 ( .A(B[15]), .B(n166), .C(n167), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n169), .B(B[2]), .Z(n168) );
    VMW_AO22 U5 ( .A(n171), .B(B[0]), .C(n172), .D(B[1]), .Z(n170) );
    VMW_OR2 U6 ( .A(B[2]), .B(n169), .Z(n173) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n172), .C(n173), .D(n170), .Z(n174) );
    VMW_NAND2 U8 ( .A(n176), .B(B[4]), .Z(n175) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n178), .C(n174), .D(n168), .Z(n177) );
    VMW_OR2 U10 ( .A(B[4]), .B(n176), .Z(n179) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n181), .C(n179), .D(n177), .Z(n180) );
    VMW_NAND2 U12 ( .A(n183), .B(B[6]), .Z(n182) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n185), .C(n180), .D(n175), .Z(n184) );
    VMW_OR2 U14 ( .A(B[6]), .B(n183), .Z(n186) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n188), .C(n186), .D(n184), .Z(n187) );
    VMW_NAND2 U16 ( .A(n190), .B(B[8]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n192), .C(n187), .D(n182), .Z(n191) );
    VMW_OR2 U18 ( .A(B[8]), .B(n190), .Z(n193) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n195), .C(n193), .D(n191), .Z(n194) );
    VMW_NAND2 U20 ( .A(n197), .B(B[10]), .Z(n196) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n199), .C(n194), .D(n189), .Z(n198) );
    VMW_NAND2 U22 ( .A(n199), .B(A[9]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n197), .C(n200), .D(n198), .Z(n201) );
    VMW_NAND2 U24 ( .A(n203), .B(B[12]), .Z(n202) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n205), .C(n201), .D(n196), .Z(n204) );
    VMW_NAND2 U26 ( .A(n205), .B(A[11]), .Z(n206) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n203), .C(n206), .D(n204), .Z(n207) );
    VMW_NAND2 U28 ( .A(n209), .B(B[14]), .Z(n208) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n211), .C(n207), .D(n202), .Z(n210) );
    VMW_NAND2 U30 ( .A(n211), .B(A[13]), .Z(n212) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n209), .C(n212), .D(n210), .Z(n213) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n214), .C(n213), .D(n208), .Z(n167) );
    VMW_INV U33 ( .A(A[12]), .Z(n203) );
    VMW_INV U34 ( .A(B[7]), .Z(n192) );
    VMW_INV U35 ( .A(A[7]), .Z(n195) );
    VMW_INV U36 ( .A(A[3]), .Z(n181) );
    VMW_INV U37 ( .A(B[3]), .Z(n178) );
    VMW_INV U38 ( .A(A[10]), .Z(n197) );
    VMW_INV U39 ( .A(B[9]), .Z(n199) );
    VMW_INV U40 ( .A(A[4]), .Z(n176) );
    VMW_INV U41 ( .A(A[8]), .Z(n190) );
    VMW_INV U42 ( .A(A[14]), .Z(n209) );
    VMW_INV U43 ( .A(B[11]), .Z(n205) );
    VMW_INV U44 ( .A(A[5]), .Z(n188) );
    VMW_INV U45 ( .A(B[5]), .Z(n185) );
    VMW_INV U46 ( .A(A[1]), .Z(n172) );
    VMW_INV U47 ( .A(B[15]), .Z(n214) );
    VMW_INV U48 ( .A(B[13]), .Z(n211) );
    VMW_INV U49 ( .A(A[6]), .Z(n183) );
    VMW_INV U50 ( .A(A[2]), .Z(n169) );
    VMW_INV U51 ( .A(A[0]), .Z(n171) );
    VMW_INV U52 ( .A(A[15]), .Z(n166) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp200[0] , \temp384[15] , \OutEdge126[12] , \temp200[15] , 
        \temp200[9] , \temp384[6] , \temp294[3] , n112, \temp294[13] , 
        \temp384[11] , \temp200[4] , \temp294[7] , \temp384[2] , \path[2] , 
        \temp200[11] , \temp200[13] , \path[0] , \temp294[5] , \temp384[0] , 
        \temp384[13] , \temp200[6] , \temp384[9] , \OutEdge126[14] , 
        \temp294[11] , \temp384[4] , \temp294[1] , \OutEdge126[10] , 
        \temp294[15] , \temp200[2] , \temp294[8] , \OutEdge126[8] , 
        \OutEdge126[1] , \OutEdge126[5] , n96, \OutEdge126[7] , 
        \OutEdge126[3] , \OutEdge126[2] , \OutEdge126[6] , \OutEdge126[4] , 
        n104, \OutEdge126[9] , n88, \OutEdge126[0] , \temp384[5] , 
        \temp294[0] , \OutEdge126[11] , \temp294[14] , \temp200[3] , 
        \temp294[9] , \path[1] , \temp200[12] , \temp294[4] , \temp384[1] , 
        \temp384[12] , \temp384[8] , \temp200[7] , \OutEdge126[15] , 
        \temp294[10] , \temp294[12] , \temp384[10] , \temp200[5] , 
        \temp294[6] , \path[3] , \temp384[3] , \temp200[10] , \temp200[1] , 
        \temp384[14] , \OutEdge126[13] , \temp200[14] , \temp384[7] , 
        \temp200[8] , \temp294[2] , n567, n568, n569, n570, n571, n572, n573, 
        n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
        n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
        n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U73 ( .Z(n606) );
    VMW_PULLDOWN U74 ( .Z(n607) );
    VMW_PULLDOWN U75 ( .Z(n608) );
    VMW_PULLDOWN U76 ( .Z(n609) );
    VMW_NOR2 U77 ( .A(Start), .B(n567), .Z(\OutEdge126[15] ) );
    VMW_NAND2 U78 ( .A(n568), .B(n569), .Z(\OutEdge126[14] ) );
    VMW_NAND2 U79 ( .A(n570), .B(n569), .Z(\OutEdge126[13] ) );
    VMW_NAND2 U80 ( .A(n571), .B(n569), .Z(\OutEdge126[12] ) );
    VMW_NAND2 U81 ( .A(n572), .B(n569), .Z(\OutEdge126[11] ) );
    VMW_NAND2 U82 ( .A(n573), .B(n569), .Z(\OutEdge126[10] ) );
    VMW_NAND2 U83 ( .A(n574), .B(n569), .Z(\OutEdge126[9] ) );
    VMW_NAND2 U84 ( .A(n575), .B(n569), .Z(\OutEdge126[8] ) );
    VMW_NAND2 U85 ( .A(n576), .B(n569), .Z(\OutEdge126[7] ) );
    VMW_NAND2 U86 ( .A(n577), .B(n569), .Z(\OutEdge126[6] ) );
    VMW_NAND2 U87 ( .A(n578), .B(n569), .Z(\OutEdge126[5] ) );
    VMW_NAND2 U88 ( .A(n579), .B(n569), .Z(\OutEdge126[4] ) );
    VMW_NAND2 U89 ( .A(n580), .B(n569), .Z(\OutEdge126[3] ) );
    VMW_NAND2 U90 ( .A(n581), .B(n569), .Z(\OutEdge126[2] ) );
    VMW_NAND2 U91 ( .A(n582), .B(n569), .Z(\OutEdge126[1] ) );
    VMW_NAND2 U92 ( .A(n583), .B(n569), .Z(\OutEdge126[0] ) );
    VMW_AO21 U93 ( .A(Start), .B(\path[3] ), .C(n584), .Z(n604) );
    VMW_AO21 U94 ( .A(\path[2] ), .B(Start), .C(n584), .Z(n603) );
    VMW_OAI211 U95 ( .A(n96), .B(n88), .C(n586), .D(n587), .Z(n585) );
    VMW_NAND2 U96 ( .A(n586), .B(n589), .Z(n588) );
    VMW_AO22 U97 ( .A(\temp294[15] ), .B(n587), .C(InEdges[47]), .D(n104), .Z(
        \temp384[15] ) );
    VMW_INV U98 ( .A(n88), .Z(n590) );
    VMW_INV U99 ( .A(Start), .Z(n569) );
    VMW_OAI22 U100 ( .A(n585), .B(Start), .C(\path[1] ), .D(n569), .Z(n591) );
    VMW_OAI22 U101 ( .A(n588), .B(Start), .C(\path[0] ), .D(n569), .Z(n592) );
    VMW_MUX2I U102 ( .A(\temp384[15] ), .B(InEdges[63]), .S(n112), .Z(n567) );
    VMW_AND3 U103 ( .A(n594), .B(n595), .C(n596), .Z(n593) );
    VMW_INV U104 ( .A(n96), .Z(n597) );
    VMW_AND5 U105 ( .A(n590), .B(n569), .C(n586), .D(n587), .E(n597), .Z(n584)
         );
    VMW_OAI21 U106 ( .A(n96), .B(n590), .C(n587), .Z(n589) );
    VMW_AND4 U107 ( .A(n598), .B(n599), .C(n600), .D(n593), .Z(n601) );
    VMW_XNOR2 U108 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n595) );
    VMW_XNOR2 U109 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n594) );
    VMW_XNOR2 U110 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n596) );
    VMW_XNOR2 U111 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n599) );
    VMW_XNOR2 U112 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n598) );
    VMW_XNOR2 U113 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n600) );
    VMW_AO22 U114 ( .A(InEdges[9]), .B(n88), .C(OutEdge[9]), .D(n590), .Z(
        \temp200[9] ) );
    VMW_AO22 U115 ( .A(InEdges[25]), .B(n96), .C(\temp200[9] ), .D(n597), .Z(
        \temp294[9] ) );
    VMW_AO22 U116 ( .A(\temp294[9] ), .B(n587), .C(InEdges[41]), .D(n104), .Z(
        \temp384[9] ) );
    VMW_AO22 U117 ( .A(InEdges[8]), .B(n88), .C(OutEdge[8]), .D(n590), .Z(
        \temp200[8] ) );
    VMW_AO22 U118 ( .A(InEdges[24]), .B(n96), .C(\temp200[8] ), .D(n597), .Z(
        \temp294[8] ) );
    VMW_AO22 U119 ( .A(\temp294[8] ), .B(n587), .C(InEdges[40]), .D(n104), .Z(
        \temp384[8] ) );
    VMW_AO22 U120 ( .A(InEdges[7]), .B(n88), .C(OutEdge[7]), .D(n590), .Z(
        \temp200[7] ) );
    VMW_AO22 U121 ( .A(InEdges[23]), .B(n96), .C(\temp200[7] ), .D(n597), .Z(
        \temp294[7] ) );
    VMW_AO22 U122 ( .A(\temp294[7] ), .B(n587), .C(InEdges[39]), .D(n104), .Z(
        \temp384[7] ) );
    VMW_AO22 U123 ( .A(InEdges[6]), .B(n88), .C(OutEdge[6]), .D(n590), .Z(
        \temp200[6] ) );
    VMW_AO22 U124 ( .A(InEdges[22]), .B(n96), .C(\temp200[6] ), .D(n597), .Z(
        \temp294[6] ) );
    VMW_AO22 U125 ( .A(\temp294[6] ), .B(n587), .C(InEdges[38]), .D(n104), .Z(
        \temp384[6] ) );
    VMW_AO22 U126 ( .A(InEdges[5]), .B(n88), .C(OutEdge[5]), .D(n590), .Z(
        \temp200[5] ) );
    VMW_AO22 U127 ( .A(InEdges[21]), .B(n96), .C(\temp200[5] ), .D(n597), .Z(
        \temp294[5] ) );
    VMW_AO22 U128 ( .A(\temp294[5] ), .B(n587), .C(InEdges[37]), .D(n104), .Z(
        \temp384[5] ) );
    VMW_AO22 U129 ( .A(InEdges[4]), .B(n88), .C(OutEdge[4]), .D(n590), .Z(
        \temp200[4] ) );
    VMW_AO22 U130 ( .A(InEdges[20]), .B(n96), .C(\temp200[4] ), .D(n597), .Z(
        \temp294[4] ) );
    VMW_AO22 U131 ( .A(\temp294[4] ), .B(n587), .C(InEdges[36]), .D(n104), .Z(
        \temp384[4] ) );
    VMW_AO22 U132 ( .A(InEdges[3]), .B(n88), .C(OutEdge[3]), .D(n590), .Z(
        \temp200[3] ) );
    VMW_AO22 U133 ( .A(InEdges[19]), .B(n96), .C(\temp200[3] ), .D(n597), .Z(
        \temp294[3] ) );
    VMW_AO22 U134 ( .A(\temp294[3] ), .B(n587), .C(InEdges[35]), .D(n104), .Z(
        \temp384[3] ) );
    VMW_AO22 U135 ( .A(InEdges[2]), .B(n88), .C(OutEdge[2]), .D(n590), .Z(
        \temp200[2] ) );
    VMW_AO22 U136 ( .A(InEdges[18]), .B(n96), .C(\temp200[2] ), .D(n597), .Z(
        \temp294[2] ) );
    VMW_AO22 U137 ( .A(\temp294[2] ), .B(n587), .C(InEdges[34]), .D(n104), .Z(
        \temp384[2] ) );
    VMW_AO22 U138 ( .A(InEdges[1]), .B(n88), .C(OutEdge[1]), .D(n590), .Z(
        \temp200[1] ) );
    VMW_AO22 U139 ( .A(InEdges[17]), .B(n96), .C(\temp200[1] ), .D(n597), .Z(
        \temp294[1] ) );
    VMW_AO22 U140 ( .A(\temp294[1] ), .B(n587), .C(InEdges[33]), .D(n104), .Z(
        \temp384[1] ) );
    VMW_AO22 U141 ( .A(InEdges[15]), .B(n88), .C(OutEdge[15]), .D(n590), .Z(
        \temp200[15] ) );
    VMW_AO22 U142 ( .A(InEdges[31]), .B(n96), .C(\temp200[15] ), .D(n597), .Z(
        \temp294[15] ) );
    VMW_AO22 U143 ( .A(InEdges[14]), .B(n88), .C(OutEdge[14]), .D(n590), .Z(
        \temp200[14] ) );
    VMW_AO22 U144 ( .A(InEdges[30]), .B(n96), .C(\temp200[14] ), .D(n597), .Z(
        \temp294[14] ) );
    VMW_AO22 U145 ( .A(\temp294[14] ), .B(n587), .C(InEdges[46]), .D(n104), 
        .Z(\temp384[14] ) );
    VMW_AO22 U146 ( .A(InEdges[13]), .B(n88), .C(OutEdge[13]), .D(n590), .Z(
        \temp200[13] ) );
    VMW_AO22 U147 ( .A(InEdges[29]), .B(n96), .C(\temp200[13] ), .D(n597), .Z(
        \temp294[13] ) );
    VMW_AO22 U148 ( .A(\temp294[13] ), .B(n587), .C(InEdges[45]), .D(n104), 
        .Z(\temp384[13] ) );
    VMW_AO22 U149 ( .A(InEdges[12]), .B(n88), .C(OutEdge[12]), .D(n590), .Z(
        \temp200[12] ) );
    VMW_AO22 U150 ( .A(InEdges[28]), .B(n96), .C(\temp200[12] ), .D(n597), .Z(
        \temp294[12] ) );
    VMW_AO22 U151 ( .A(\temp294[12] ), .B(n587), .C(InEdges[44]), .D(n104), 
        .Z(\temp384[12] ) );
    VMW_AO22 U152 ( .A(InEdges[11]), .B(n88), .C(OutEdge[11]), .D(n590), .Z(
        \temp200[11] ) );
    VMW_AO22 U153 ( .A(InEdges[27]), .B(n96), .C(\temp200[11] ), .D(n597), .Z(
        \temp294[11] ) );
    VMW_AO22 U154 ( .A(\temp294[11] ), .B(n587), .C(InEdges[43]), .D(n104), 
        .Z(\temp384[11] ) );
    VMW_AO22 U155 ( .A(InEdges[10]), .B(n88), .C(OutEdge[10]), .D(n590), .Z(
        \temp200[10] ) );
    VMW_AO22 U156 ( .A(InEdges[26]), .B(n96), .C(\temp200[10] ), .D(n597), .Z(
        \temp294[10] ) );
    VMW_AO22 U157 ( .A(\temp294[10] ), .B(n587), .C(InEdges[42]), .D(n104), 
        .Z(\temp384[10] ) );
    VMW_AO22 U158 ( .A(InEdges[0]), .B(n88), .C(OutEdge[0]), .D(n590), .Z(
        \temp200[0] ) );
    VMW_AO22 U159 ( .A(InEdges[16]), .B(n96), .C(\temp200[0] ), .D(n597), .Z(
        \temp294[0] ) );
    VMW_AO22 U160 ( .A(\temp294[0] ), .B(n587), .C(InEdges[32]), .D(n104), .Z(
        \temp384[0] ) );
    VMW_MUX2I U161 ( .A(\temp384[9] ), .B(InEdges[57]), .S(n112), .Z(n574) );
    VMW_MUX2I U162 ( .A(\temp384[8] ), .B(InEdges[56]), .S(n112), .Z(n575) );
    VMW_MUX2I U163 ( .A(\temp384[7] ), .B(InEdges[55]), .S(n112), .Z(n576) );
    VMW_MUX2I U164 ( .A(\temp384[6] ), .B(InEdges[54]), .S(n112), .Z(n577) );
    VMW_MUX2I U165 ( .A(\temp384[5] ), .B(InEdges[53]), .S(n112), .Z(n578) );
    VMW_MUX2I U166 ( .A(\temp384[4] ), .B(InEdges[52]), .S(n112), .Z(n579) );
    VMW_MUX2I U167 ( .A(\temp384[3] ), .B(InEdges[51]), .S(n112), .Z(n580) );
    VMW_MUX2I U168 ( .A(\temp384[2] ), .B(InEdges[50]), .S(n112), .Z(n581) );
    VMW_MUX2I U169 ( .A(\temp384[1] ), .B(InEdges[49]), .S(n112), .Z(n582) );
    VMW_MUX2I U170 ( .A(\temp384[14] ), .B(InEdges[62]), .S(n112), .Z(n568) );
    VMW_MUX2I U171 ( .A(\temp384[13] ), .B(InEdges[61]), .S(n112), .Z(n570) );
    VMW_MUX2I U172 ( .A(\temp384[12] ), .B(InEdges[60]), .S(n112), .Z(n571) );
    VMW_MUX2I U173 ( .A(\temp384[11] ), .B(InEdges[59]), .S(n112), .Z(n572) );
    VMW_MUX2I U174 ( .A(\temp384[10] ), .B(InEdges[58]), .S(n112), .Z(n573) );
    VMW_MUX2I U175 ( .A(\temp384[0] ), .B(InEdges[48]), .S(n112), .Z(n583) );
    VMW_INV U176 ( .A(n104), .Z(n587) );
    VMW_INV U177 ( .A(n112), .Z(n586) );
    VMW_INV U178 ( .A(n591), .Z(n605) );
    VMW_INV U179 ( .A(n592), .Z(n602) );
    VMW_BUFIZ U180 ( .A(\path[3] ), .E(n601), .Z(\PathData[3] ) );
    VMW_BUFIZ U181 ( .A(\path[1] ), .E(n601), .Z(\PathData[1] ) );
    VMW_BUFIZ U182 ( .A(\path[0] ), .E(n601), .Z(\PathData[0] ) );
    VMW_BUFIZ U183 ( .A(\path[2] ), .E(n601), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n602), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n603), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n604), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n605), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge126[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge126[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge126[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge126[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge126[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge126[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge126[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge126[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge126[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge126[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge126[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge126[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge126[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge126[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge126[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge126[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n609), .TC(n609), .GE_GT(n88) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp200[15] , 
        \temp200[14] , \temp200[13] , \temp200[12] , \temp200[11] , 
        \temp200[10] , \temp200[9] , \temp200[8] , \temp200[7] , \temp200[6] , 
        \temp200[5] , \temp200[4] , \temp200[3] , \temp200[2] , \temp200[1] , 
        \temp200[0] }), .B(InEdges[31:16]), .LEQ(n608), .TC(n608), .GE_GT(n96)
         );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp294[15] , 
        \temp294[14] , \temp294[13] , \temp294[12] , \temp294[11] , 
        \temp294[10] , \temp294[9] , \temp294[8] , \temp294[7] , \temp294[6] , 
        \temp294[5] , \temp294[4] , \temp294[3] , \temp294[2] , \temp294[1] , 
        \temp294[0] }), .B(InEdges[47:32]), .LEQ(n607), .TC(n607), .GE_GT(n104
        ) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp384[15] , 
        \temp384[14] , \temp384[13] , \temp384[12] , \temp384[11] , 
        \temp384[10] , \temp384[9] , \temp384[8] , \temp384[7] , \temp384[6] , 
        \temp384[5] , \temp384[4] , \temp384[3] , \temp384[2] , \temp384[1] , 
        \temp384[0] }), .B(InEdges[63:48]), .LEQ(n606), .TC(n606), .GE_GT(n112
        ) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, 
        n93, n94, n95, n96, n97, n99, n100, n101, n102, n103, n104, n105, n107, 
        n108, n109, n110, n111, n112, n113, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n100), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n104), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n123), .B(B[0]), .C(n124), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n124), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n137), .C(n132), .D(n127), .Z(n136) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n138) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n140), .C(n138), .D(n136), .Z(n139) );
    VMW_NAND2 U16 ( .A(n142), .B(B[8]), .Z(n141) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n144), .C(n139), .D(n134), .Z(n143) );
    VMW_OR2 U18 ( .A(B[8]), .B(n142), .Z(n145) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n147), .C(n145), .D(n143), .Z(n146) );
    VMW_NAND2 U20 ( .A(n149), .B(B[10]), .Z(n148) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n151), .C(n146), .D(n141), .Z(n150) );
    VMW_NAND2 U22 ( .A(n151), .B(A[9]), .Z(n152) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n149), .C(n152), .D(n150), .Z(n153) );
    VMW_NAND2 U24 ( .A(n155), .B(B[12]), .Z(n154) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n157), .C(n153), .D(n148), .Z(n156) );
    VMW_NAND2 U26 ( .A(n157), .B(A[11]), .Z(n158) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n155), .C(n158), .D(n156), .Z(n159) );
    VMW_NAND2 U28 ( .A(n161), .B(B[14]), .Z(n160) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n163), .C(n159), .D(n154), .Z(n162) );
    VMW_NAND2 U30 ( .A(n163), .B(A[13]), .Z(n164) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n161), .C(n164), .D(n162), .Z(n165) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n166), .C(n165), .D(n160), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n155) );
    VMW_INV U34 ( .A(B[7]), .Z(n144) );
    VMW_INV U35 ( .A(A[7]), .Z(n147) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n149) );
    VMW_INV U39 ( .A(B[9]), .Z(n151) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n142) );
    VMW_INV U42 ( .A(A[14]), .Z(n161) );
    VMW_INV U43 ( .A(B[11]), .Z(n157) );
    VMW_INV U44 ( .A(A[5]), .Z(n140) );
    VMW_INV U45 ( .A(B[5]), .Z(n137) );
    VMW_INV U46 ( .A(A[1]), .Z(n124) );
    VMW_INV U47 ( .A(B[15]), .Z(n166) );
    VMW_INV U48 ( .A(B[13]), .Z(n163) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n123) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
        n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
        n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
        n214, n215;
    VMW_OAI21 U3 ( .A(B[15]), .B(n167), .C(n168), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n170), .B(B[2]), .Z(n169) );
    VMW_AO22 U5 ( .A(n172), .B(B[0]), .C(n173), .D(B[1]), .Z(n171) );
    VMW_OR2 U6 ( .A(B[2]), .B(n170), .Z(n174) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n173), .C(n174), .D(n171), .Z(n175) );
    VMW_NAND2 U8 ( .A(n177), .B(B[4]), .Z(n176) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n179), .C(n175), .D(n169), .Z(n178) );
    VMW_OR2 U10 ( .A(B[4]), .B(n177), .Z(n180) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n182), .C(n180), .D(n178), .Z(n181) );
    VMW_NAND2 U12 ( .A(n184), .B(B[6]), .Z(n183) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n186), .C(n181), .D(n176), .Z(n185) );
    VMW_OR2 U14 ( .A(B[6]), .B(n184), .Z(n187) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n189), .C(n187), .D(n185), .Z(n188) );
    VMW_NAND2 U16 ( .A(n191), .B(B[8]), .Z(n190) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n193), .C(n188), .D(n183), .Z(n192) );
    VMW_OR2 U18 ( .A(B[8]), .B(n191), .Z(n194) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n196), .C(n194), .D(n192), .Z(n195) );
    VMW_NAND2 U20 ( .A(n198), .B(B[10]), .Z(n197) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n200), .C(n195), .D(n190), .Z(n199) );
    VMW_NAND2 U22 ( .A(n200), .B(A[9]), .Z(n201) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n198), .C(n201), .D(n199), .Z(n202) );
    VMW_NAND2 U24 ( .A(n204), .B(B[12]), .Z(n203) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n206), .C(n202), .D(n197), .Z(n205) );
    VMW_NAND2 U26 ( .A(n206), .B(A[11]), .Z(n207) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n204), .C(n207), .D(n205), .Z(n208) );
    VMW_NAND2 U28 ( .A(n210), .B(B[14]), .Z(n209) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n212), .C(n208), .D(n203), .Z(n211) );
    VMW_NAND2 U30 ( .A(n212), .B(A[13]), .Z(n213) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n210), .C(n213), .D(n211), .Z(n214) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n215), .C(n214), .D(n209), .Z(n168) );
    VMW_INV U33 ( .A(A[12]), .Z(n204) );
    VMW_INV U34 ( .A(B[7]), .Z(n193) );
    VMW_INV U35 ( .A(A[7]), .Z(n196) );
    VMW_INV U36 ( .A(A[3]), .Z(n182) );
    VMW_INV U37 ( .A(B[3]), .Z(n179) );
    VMW_INV U38 ( .A(A[10]), .Z(n198) );
    VMW_INV U39 ( .A(B[9]), .Z(n200) );
    VMW_INV U40 ( .A(A[4]), .Z(n177) );
    VMW_INV U41 ( .A(A[8]), .Z(n191) );
    VMW_INV U42 ( .A(A[14]), .Z(n210) );
    VMW_INV U43 ( .A(B[11]), .Z(n206) );
    VMW_INV U44 ( .A(A[5]), .Z(n189) );
    VMW_INV U45 ( .A(B[5]), .Z(n186) );
    VMW_INV U46 ( .A(A[1]), .Z(n173) );
    VMW_INV U47 ( .A(B[15]), .Z(n215) );
    VMW_INV U48 ( .A(B[13]), .Z(n212) );
    VMW_INV U49 ( .A(A[6]), .Z(n184) );
    VMW_INV U50 ( .A(A[2]), .Z(n170) );
    VMW_INV U51 ( .A(A[0]), .Z(n172) );
    VMW_INV U52 ( .A(A[15]), .Z(n167) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264;
    VMW_OAI21 U3 ( .A(B[15]), .B(n216), .C(n217), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n219), .B(B[2]), .Z(n218) );
    VMW_AO22 U5 ( .A(n221), .B(B[0]), .C(n222), .D(B[1]), .Z(n220) );
    VMW_OR2 U6 ( .A(B[2]), .B(n219), .Z(n223) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n222), .C(n223), .D(n220), .Z(n224) );
    VMW_NAND2 U8 ( .A(n226), .B(B[4]), .Z(n225) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n228), .C(n224), .D(n218), .Z(n227) );
    VMW_OR2 U10 ( .A(B[4]), .B(n226), .Z(n229) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n231), .C(n229), .D(n227), .Z(n230) );
    VMW_NAND2 U12 ( .A(n233), .B(B[6]), .Z(n232) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n235), .C(n230), .D(n225), .Z(n234) );
    VMW_OR2 U14 ( .A(B[6]), .B(n233), .Z(n236) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n238), .C(n236), .D(n234), .Z(n237) );
    VMW_NAND2 U16 ( .A(n240), .B(B[8]), .Z(n239) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n242), .C(n237), .D(n232), .Z(n241) );
    VMW_OR2 U18 ( .A(B[8]), .B(n240), .Z(n243) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n245), .C(n243), .D(n241), .Z(n244) );
    VMW_NAND2 U20 ( .A(n247), .B(B[10]), .Z(n246) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n249), .C(n244), .D(n239), .Z(n248) );
    VMW_NAND2 U22 ( .A(n249), .B(A[9]), .Z(n250) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n247), .C(n250), .D(n248), .Z(n251) );
    VMW_NAND2 U24 ( .A(n253), .B(B[12]), .Z(n252) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n255), .C(n251), .D(n246), .Z(n254) );
    VMW_NAND2 U26 ( .A(n255), .B(A[11]), .Z(n256) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n253), .C(n256), .D(n254), .Z(n257) );
    VMW_NAND2 U28 ( .A(n259), .B(B[14]), .Z(n258) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n261), .C(n257), .D(n252), .Z(n260) );
    VMW_NAND2 U30 ( .A(n261), .B(A[13]), .Z(n262) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n259), .C(n262), .D(n260), .Z(n263) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n264), .C(n263), .D(n258), .Z(n217) );
    VMW_INV U33 ( .A(A[12]), .Z(n253) );
    VMW_INV U34 ( .A(B[7]), .Z(n242) );
    VMW_INV U35 ( .A(A[7]), .Z(n245) );
    VMW_INV U36 ( .A(A[3]), .Z(n231) );
    VMW_INV U37 ( .A(B[3]), .Z(n228) );
    VMW_INV U38 ( .A(A[10]), .Z(n247) );
    VMW_INV U39 ( .A(B[9]), .Z(n249) );
    VMW_INV U40 ( .A(A[4]), .Z(n226) );
    VMW_INV U41 ( .A(A[8]), .Z(n240) );
    VMW_INV U42 ( .A(A[14]), .Z(n259) );
    VMW_INV U43 ( .A(B[11]), .Z(n255) );
    VMW_INV U44 ( .A(A[5]), .Z(n238) );
    VMW_INV U45 ( .A(B[5]), .Z(n235) );
    VMW_INV U46 ( .A(A[1]), .Z(n222) );
    VMW_INV U47 ( .A(B[15]), .Z(n264) );
    VMW_INV U48 ( .A(B[13]), .Z(n261) );
    VMW_INV U49 ( .A(A[6]), .Z(n233) );
    VMW_INV U50 ( .A(A[2]), .Z(n219) );
    VMW_INV U51 ( .A(A[0]), .Z(n221) );
    VMW_INV U52 ( .A(A[15]), .Z(n216) );
endmodule


module NodeAux_INDEGREE5_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp210[13] , \temp484[4] , \temp394[5] , \temp304[13] , 
        \temp210[3] , \temp394[13] , \OutEdge136[14] , \temp394[1] , 
        \temp484[0] , \OutEdge136[10] , \path[2] , \temp394[8] , \temp210[7] , 
        \temp484[9] , \temp394[15] , \path[0] , \temp210[5] , \OutEdge136[12] , 
        \temp210[15] , \temp304[15] , \temp394[3] , \temp484[2] , \temp210[1] , 
        n90, \temp394[11] , \temp484[6] , \temp394[7] , \temp210[8] , 
        \temp304[11] , \temp210[11] , n98, n114, \OutEdge136[2] , \temp304[4] , 
        \OutEdge136[6] , \temp304[9] , \temp304[0] , \temp484[13] , n106, 
        \temp304[2] , \temp484[11] , \OutEdge136[4] , \temp484[15] , 
        \temp304[6] , \OutEdge136[9] , \OutEdge136[0] , \temp484[14] , 
        \OutEdge136[8] , \temp304[7] , \OutEdge136[1] , \temp304[3] , 
        \temp484[10] , \OutEdge136[5] , \OutEdge136[7] , \temp304[8] , 
        \temp304[1] , \temp484[12] , \OutEdge136[3] , \temp304[5] , 
        \temp394[10] , \temp210[0] , \temp484[7] , \temp210[9] , \temp304[10] , 
        \temp394[6] , \temp210[10] , \temp210[4] , \path[1] , \temp394[14] , 
        \OutEdge136[13] , \temp210[14] , n122, \temp394[2] , \temp304[14] , 
        \temp484[3] , \temp394[0] , \temp484[1] , \path[3] , \OutEdge136[11] , 
        \temp210[6] , \temp394[9] , \temp484[8] , \temp210[12] , \temp484[5] , 
        \temp304[12] , \temp394[4] , \OutEdge136[15] , \temp394[12] , 
        \temp210[2] , n667, n668, n669, n670, n671, n672, n673, n674, n675, 
        n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
        n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
        n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
        n712;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U82 ( .Z(n711) );
    VMW_PULLDOWN U83 ( .Z(n708) );
    VMW_PULLDOWN U84 ( .Z(n710) );
    VMW_PULLDOWN U85 ( .Z(n709) );
    VMW_PULLDOWN U86 ( .Z(n712) );
    VMW_AO21 U87 ( .A(\temp484[15] ), .B(n667), .C(n668), .Z(\OutEdge136[15] )
         );
    VMW_OR2 U88 ( .A(n669), .B(Start), .Z(\OutEdge136[14] ) );
    VMW_OR2 U89 ( .A(n670), .B(Start), .Z(\OutEdge136[13] ) );
    VMW_OR2 U90 ( .A(n671), .B(Start), .Z(\OutEdge136[12] ) );
    VMW_OR2 U91 ( .A(n672), .B(Start), .Z(\OutEdge136[11] ) );
    VMW_OR2 U92 ( .A(n673), .B(Start), .Z(\OutEdge136[10] ) );
    VMW_OR2 U93 ( .A(n674), .B(Start), .Z(\OutEdge136[9] ) );
    VMW_OR2 U94 ( .A(n675), .B(Start), .Z(\OutEdge136[8] ) );
    VMW_OR2 U95 ( .A(n676), .B(Start), .Z(\OutEdge136[7] ) );
    VMW_OR2 U96 ( .A(n677), .B(Start), .Z(\OutEdge136[6] ) );
    VMW_OR2 U97 ( .A(n678), .B(Start), .Z(\OutEdge136[5] ) );
    VMW_OR2 U98 ( .A(n679), .B(Start), .Z(\OutEdge136[4] ) );
    VMW_OR2 U99 ( .A(n680), .B(Start), .Z(\OutEdge136[3] ) );
    VMW_OR2 U100 ( .A(n681), .B(Start), .Z(\OutEdge136[2] ) );
    VMW_OR2 U101 ( .A(n682), .B(Start), .Z(\OutEdge136[1] ) );
    VMW_OR2 U102 ( .A(n683), .B(Start), .Z(\OutEdge136[0] ) );
    VMW_AO22 U103 ( .A(\path[1] ), .B(Start), .C(n667), .D(n684), .Z(n707) );
    VMW_AO22 U104 ( .A(Start), .B(\path[3] ), .C(n685), .D(n686), .Z(n706) );
    VMW_OR2 U105 ( .A(n685), .B(n687), .Z(n705) );
    VMW_AO21 U106 ( .A(Start), .B(\path[0] ), .C(n688), .Z(n704) );
    VMW_AO22 U107 ( .A(\temp394[15] ), .B(n689), .C(InEdges[63]), .D(n114), 
        .Z(\temp484[15] ) );
    VMW_NOR5 U108 ( .A(n90), .B(Start), .C(n114), .D(n106), .E(n98), .Z(n685)
         );
    VMW_INV U109 ( .A(Start), .Z(n690) );
    VMW_INV U110 ( .A(n122), .Z(n686) );
    VMW_AND2 U111 ( .A(n690), .B(n686), .Z(n667) );
    VMW_AO22 U112 ( .A(\path[2] ), .B(Start), .C(n122), .D(n690), .Z(n687) );
    VMW_AND3 U113 ( .A(n692), .B(n693), .C(n694), .Z(n691) );
    VMW_INV U114 ( .A(n114), .Z(n689) );
    VMW_INV U115 ( .A(n106), .Z(n695) );
    VMW_OAI211 U116 ( .A(n90), .B(n98), .C(n695), .D(n689), .Z(n684) );
    VMW_OAI21 U117 ( .A(n98), .B(n697), .C(n695), .Z(n696) );
    VMW_AOI21 U118 ( .A(n689), .B(n696), .C(n698), .Z(n688) );
    VMW_AND4 U119 ( .A(n699), .B(n700), .C(n701), .D(n691), .Z(n703) );
    VMW_AND3 U120 ( .A(n122), .B(n690), .C(InEdges[79]), .Z(n668) );
    VMW_XNOR2 U121 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n693) );
    VMW_XNOR2 U122 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n692) );
    VMW_XNOR2 U123 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n694) );
    VMW_XNOR2 U124 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n700) );
    VMW_XNOR2 U125 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n699) );
    VMW_XNOR2 U126 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n701) );
    VMW_AO22 U127 ( .A(OutEdge[9]), .B(n697), .C(InEdges[9]), .D(n90), .Z(
        \temp210[9] ) );
    VMW_AO22 U128 ( .A(\temp210[9] ), .B(n702), .C(InEdges[25]), .D(n98), .Z(
        \temp304[9] ) );
    VMW_AO22 U129 ( .A(InEdges[41]), .B(n106), .C(\temp304[9] ), .D(n695), .Z(
        \temp394[9] ) );
    VMW_AO22 U130 ( .A(InEdges[57]), .B(n114), .C(\temp394[9] ), .D(n689), .Z(
        \temp484[9] ) );
    VMW_AO22 U131 ( .A(OutEdge[8]), .B(n697), .C(InEdges[8]), .D(n90), .Z(
        \temp210[8] ) );
    VMW_AO22 U132 ( .A(\temp210[8] ), .B(n702), .C(InEdges[24]), .D(n98), .Z(
        \temp304[8] ) );
    VMW_AO22 U133 ( .A(InEdges[40]), .B(n106), .C(\temp304[8] ), .D(n695), .Z(
        \temp394[8] ) );
    VMW_AO22 U134 ( .A(InEdges[56]), .B(n114), .C(\temp394[8] ), .D(n689), .Z(
        \temp484[8] ) );
    VMW_AO22 U135 ( .A(OutEdge[7]), .B(n697), .C(InEdges[7]), .D(n90), .Z(
        \temp210[7] ) );
    VMW_AO22 U136 ( .A(\temp210[7] ), .B(n702), .C(InEdges[23]), .D(n98), .Z(
        \temp304[7] ) );
    VMW_AO22 U137 ( .A(InEdges[39]), .B(n106), .C(\temp304[7] ), .D(n695), .Z(
        \temp394[7] ) );
    VMW_AO22 U138 ( .A(InEdges[55]), .B(n114), .C(\temp394[7] ), .D(n689), .Z(
        \temp484[7] ) );
    VMW_AO22 U139 ( .A(OutEdge[6]), .B(n697), .C(InEdges[6]), .D(n90), .Z(
        \temp210[6] ) );
    VMW_AO22 U140 ( .A(\temp210[6] ), .B(n702), .C(InEdges[22]), .D(n98), .Z(
        \temp304[6] ) );
    VMW_AO22 U141 ( .A(InEdges[38]), .B(n106), .C(\temp304[6] ), .D(n695), .Z(
        \temp394[6] ) );
    VMW_AO22 U142 ( .A(InEdges[54]), .B(n114), .C(\temp394[6] ), .D(n689), .Z(
        \temp484[6] ) );
    VMW_AO22 U143 ( .A(OutEdge[5]), .B(n697), .C(InEdges[5]), .D(n90), .Z(
        \temp210[5] ) );
    VMW_AO22 U144 ( .A(\temp210[5] ), .B(n702), .C(InEdges[21]), .D(n98), .Z(
        \temp304[5] ) );
    VMW_AO22 U145 ( .A(InEdges[37]), .B(n106), .C(\temp304[5] ), .D(n695), .Z(
        \temp394[5] ) );
    VMW_AO22 U146 ( .A(InEdges[53]), .B(n114), .C(\temp394[5] ), .D(n689), .Z(
        \temp484[5] ) );
    VMW_AO22 U147 ( .A(OutEdge[4]), .B(n697), .C(InEdges[4]), .D(n90), .Z(
        \temp210[4] ) );
    VMW_AO22 U148 ( .A(\temp210[4] ), .B(n702), .C(InEdges[20]), .D(n98), .Z(
        \temp304[4] ) );
    VMW_AO22 U149 ( .A(InEdges[36]), .B(n106), .C(\temp304[4] ), .D(n695), .Z(
        \temp394[4] ) );
    VMW_AO22 U150 ( .A(InEdges[52]), .B(n114), .C(\temp394[4] ), .D(n689), .Z(
        \temp484[4] ) );
    VMW_AO22 U151 ( .A(OutEdge[3]), .B(n697), .C(InEdges[3]), .D(n90), .Z(
        \temp210[3] ) );
    VMW_AO22 U152 ( .A(\temp210[3] ), .B(n702), .C(InEdges[19]), .D(n98), .Z(
        \temp304[3] ) );
    VMW_AO22 U153 ( .A(InEdges[35]), .B(n106), .C(\temp304[3] ), .D(n695), .Z(
        \temp394[3] ) );
    VMW_AO22 U154 ( .A(InEdges[51]), .B(n114), .C(\temp394[3] ), .D(n689), .Z(
        \temp484[3] ) );
    VMW_AO22 U155 ( .A(OutEdge[2]), .B(n697), .C(InEdges[2]), .D(n90), .Z(
        \temp210[2] ) );
    VMW_AO22 U156 ( .A(\temp210[2] ), .B(n702), .C(InEdges[18]), .D(n98), .Z(
        \temp304[2] ) );
    VMW_AO22 U157 ( .A(InEdges[34]), .B(n106), .C(\temp304[2] ), .D(n695), .Z(
        \temp394[2] ) );
    VMW_AO22 U158 ( .A(InEdges[50]), .B(n114), .C(\temp394[2] ), .D(n689), .Z(
        \temp484[2] ) );
    VMW_AO22 U159 ( .A(OutEdge[1]), .B(n697), .C(InEdges[1]), .D(n90), .Z(
        \temp210[1] ) );
    VMW_AO22 U160 ( .A(\temp210[1] ), .B(n702), .C(InEdges[17]), .D(n98), .Z(
        \temp304[1] ) );
    VMW_AO22 U161 ( .A(InEdges[33]), .B(n106), .C(\temp304[1] ), .D(n695), .Z(
        \temp394[1] ) );
    VMW_AO22 U162 ( .A(InEdges[49]), .B(n114), .C(\temp394[1] ), .D(n689), .Z(
        \temp484[1] ) );
    VMW_AO22 U163 ( .A(OutEdge[15]), .B(n697), .C(InEdges[15]), .D(n90), .Z(
        \temp210[15] ) );
    VMW_AO22 U164 ( .A(\temp210[15] ), .B(n702), .C(InEdges[31]), .D(n98), .Z(
        \temp304[15] ) );
    VMW_AO22 U165 ( .A(InEdges[47]), .B(n106), .C(\temp304[15] ), .D(n695), 
        .Z(\temp394[15] ) );
    VMW_AO22 U166 ( .A(OutEdge[14]), .B(n697), .C(InEdges[14]), .D(n90), .Z(
        \temp210[14] ) );
    VMW_AO22 U167 ( .A(\temp210[14] ), .B(n702), .C(InEdges[30]), .D(n98), .Z(
        \temp304[14] ) );
    VMW_AO22 U168 ( .A(InEdges[46]), .B(n106), .C(\temp304[14] ), .D(n695), 
        .Z(\temp394[14] ) );
    VMW_AO22 U169 ( .A(InEdges[62]), .B(n114), .C(\temp394[14] ), .D(n689), 
        .Z(\temp484[14] ) );
    VMW_AO22 U170 ( .A(OutEdge[13]), .B(n697), .C(InEdges[13]), .D(n90), .Z(
        \temp210[13] ) );
    VMW_AO22 U171 ( .A(\temp210[13] ), .B(n702), .C(InEdges[29]), .D(n98), .Z(
        \temp304[13] ) );
    VMW_AO22 U172 ( .A(InEdges[45]), .B(n106), .C(\temp304[13] ), .D(n695), 
        .Z(\temp394[13] ) );
    VMW_AO22 U173 ( .A(InEdges[61]), .B(n114), .C(\temp394[13] ), .D(n689), 
        .Z(\temp484[13] ) );
    VMW_AO22 U174 ( .A(OutEdge[12]), .B(n697), .C(InEdges[12]), .D(n90), .Z(
        \temp210[12] ) );
    VMW_AO22 U175 ( .A(\temp210[12] ), .B(n702), .C(InEdges[28]), .D(n98), .Z(
        \temp304[12] ) );
    VMW_AO22 U176 ( .A(InEdges[44]), .B(n106), .C(\temp304[12] ), .D(n695), 
        .Z(\temp394[12] ) );
    VMW_AO22 U177 ( .A(InEdges[60]), .B(n114), .C(\temp394[12] ), .D(n689), 
        .Z(\temp484[12] ) );
    VMW_AO22 U178 ( .A(OutEdge[11]), .B(n697), .C(InEdges[11]), .D(n90), .Z(
        \temp210[11] ) );
    VMW_AO22 U179 ( .A(\temp210[11] ), .B(n702), .C(InEdges[27]), .D(n98), .Z(
        \temp304[11] ) );
    VMW_AO22 U180 ( .A(InEdges[43]), .B(n106), .C(\temp304[11] ), .D(n695), 
        .Z(\temp394[11] ) );
    VMW_AO22 U181 ( .A(InEdges[59]), .B(n114), .C(\temp394[11] ), .D(n689), 
        .Z(\temp484[11] ) );
    VMW_AO22 U182 ( .A(OutEdge[10]), .B(n697), .C(InEdges[10]), .D(n90), .Z(
        \temp210[10] ) );
    VMW_AO22 U183 ( .A(\temp210[10] ), .B(n702), .C(InEdges[26]), .D(n98), .Z(
        \temp304[10] ) );
    VMW_AO22 U184 ( .A(InEdges[42]), .B(n106), .C(\temp304[10] ), .D(n695), 
        .Z(\temp394[10] ) );
    VMW_AO22 U185 ( .A(InEdges[58]), .B(n114), .C(\temp394[10] ), .D(n689), 
        .Z(\temp484[10] ) );
    VMW_AO22 U186 ( .A(OutEdge[0]), .B(n697), .C(InEdges[0]), .D(n90), .Z(
        \temp210[0] ) );
    VMW_AO22 U187 ( .A(\temp210[0] ), .B(n702), .C(InEdges[16]), .D(n98), .Z(
        \temp304[0] ) );
    VMW_AO22 U188 ( .A(InEdges[32]), .B(n106), .C(\temp304[0] ), .D(n695), .Z(
        \temp394[0] ) );
    VMW_AO22 U189 ( .A(InEdges[48]), .B(n114), .C(\temp394[0] ), .D(n689), .Z(
        \temp484[0] ) );
    VMW_AO22 U190 ( .A(\temp484[9] ), .B(n686), .C(InEdges[73]), .D(n122), .Z(
        n674) );
    VMW_AO22 U191 ( .A(\temp484[8] ), .B(n686), .C(InEdges[72]), .D(n122), .Z(
        n675) );
    VMW_AO22 U192 ( .A(\temp484[7] ), .B(n686), .C(InEdges[71]), .D(n122), .Z(
        n676) );
    VMW_AO22 U193 ( .A(\temp484[6] ), .B(n686), .C(InEdges[70]), .D(n122), .Z(
        n677) );
    VMW_AO22 U194 ( .A(\temp484[5] ), .B(n686), .C(InEdges[69]), .D(n122), .Z(
        n678) );
    VMW_AO22 U195 ( .A(\temp484[4] ), .B(n686), .C(InEdges[68]), .D(n122), .Z(
        n679) );
    VMW_AO22 U196 ( .A(\temp484[3] ), .B(n686), .C(InEdges[67]), .D(n122), .Z(
        n680) );
    VMW_AO22 U197 ( .A(\temp484[2] ), .B(n686), .C(InEdges[66]), .D(n122), .Z(
        n681) );
    VMW_AO22 U198 ( .A(\temp484[1] ), .B(n686), .C(InEdges[65]), .D(n122), .Z(
        n682) );
    VMW_AO22 U199 ( .A(\temp484[14] ), .B(n686), .C(InEdges[78]), .D(n122), 
        .Z(n669) );
    VMW_AO22 U200 ( .A(\temp484[13] ), .B(n686), .C(InEdges[77]), .D(n122), 
        .Z(n670) );
    VMW_AO22 U201 ( .A(\temp484[12] ), .B(n686), .C(InEdges[76]), .D(n122), 
        .Z(n671) );
    VMW_AO22 U202 ( .A(\temp484[11] ), .B(n686), .C(InEdges[75]), .D(n122), 
        .Z(n672) );
    VMW_AO22 U203 ( .A(\temp484[10] ), .B(n686), .C(InEdges[74]), .D(n122), 
        .Z(n673) );
    VMW_AO22 U204 ( .A(\temp484[0] ), .B(n686), .C(InEdges[64]), .D(n122), .Z(
        n683) );
    VMW_INV U205 ( .A(n90), .Z(n697) );
    VMW_INV U206 ( .A(n98), .Z(n702) );
    VMW_INV U207 ( .A(n667), .Z(n698) );
    VMW_BUFIZ U208 ( .A(\path[3] ), .E(n703), .Z(\PathData[3] ) );
    VMW_BUFIZ U209 ( .A(\path[1] ), .E(n703), .Z(\PathData[1] ) );
    VMW_BUFIZ U210 ( .A(\path[0] ), .E(n703), .Z(\PathData[0] ) );
    VMW_BUFIZ U211 ( .A(\path[2] ), .E(n703), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n704), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n705), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n706), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n707), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge136[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge136[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge136[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge136[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge136[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge136[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge136[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge136[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge136[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge136[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge136[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge136[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge136[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge136[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge136[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge136[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n712), .TC(n712), .GE_GT(n90) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp484[15] , 
        \temp484[14] , \temp484[13] , \temp484[12] , \temp484[11] , 
        \temp484[10] , \temp484[9] , \temp484[8] , \temp484[7] , \temp484[6] , 
        \temp484[5] , \temp484[4] , \temp484[3] , \temp484[2] , \temp484[1] , 
        \temp484[0] }), .B(InEdges[79:64]), .LEQ(n711), .TC(n711), .GE_GT(n122
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 lte_55_2 ( .A({\temp304[15] , 
        \temp304[14] , \temp304[13] , \temp304[12] , \temp304[11] , 
        \temp304[10] , \temp304[9] , \temp304[8] , \temp304[7] , \temp304[6] , 
        \temp304[5] , \temp304[4] , \temp304[3] , \temp304[2] , \temp304[1] , 
        \temp304[0] }), .B(InEdges[47:32]), .LEQ(n710), .TC(n710), .GE_GT(n106
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 lte_55_1 ( .A({\temp210[15] , 
        \temp210[14] , \temp210[13] , \temp210[12] , \temp210[11] , 
        \temp210[10] , \temp210[9] , \temp210[8] , \temp210[7] , \temp210[6] , 
        \temp210[5] , \temp210[4] , \temp210[3] , \temp210[2] , \temp210[1] , 
        \temp210[0] }), .B(InEdges[31:16]), .LEQ(n709), .TC(n709), .GE_GT(n98)
         );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp394[15] , 
        \temp394[14] , \temp394[13] , \temp394[12] , \temp394[11] , 
        \temp394[10] , \temp394[9] , \temp394[8] , \temp394[7] , \temp394[6] , 
        \temp394[5] , \temp394[4] , \temp394[3] , \temp394[2] , \temp394[1] , 
        \temp394[0] }), .B(InEdges[63:48]), .LEQ(n708), .TC(n708), .GE_GT(n114
        ) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, 
        n107, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n91), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, 
        n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n131), .D(n129), .Z(n133) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n167), .C(n166), .D(n161), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n156) );
    VMW_INV U34 ( .A(B[7]), .Z(n145) );
    VMW_INV U35 ( .A(A[7]), .Z(n148) );
    VMW_INV U36 ( .A(A[3]), .Z(n134) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n150) );
    VMW_INV U39 ( .A(B[9]), .Z(n152) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n162) );
    VMW_INV U43 ( .A(B[11]), .Z(n158) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n167) );
    VMW_INV U48 ( .A(B[13]), .Z(n164) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216;
    VMW_OAI21 U3 ( .A(B[15]), .B(n168), .C(n169), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n171), .B(B[2]), .Z(n170) );
    VMW_AO22 U5 ( .A(n173), .B(B[0]), .C(n174), .D(B[1]), .Z(n172) );
    VMW_OR2 U6 ( .A(B[2]), .B(n171), .Z(n175) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n174), .C(n175), .D(n172), .Z(n176) );
    VMW_NAND2 U8 ( .A(n178), .B(B[4]), .Z(n177) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n180), .C(n176), .D(n170), .Z(n179) );
    VMW_OR2 U10 ( .A(B[4]), .B(n178), .Z(n181) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n183), .C(n181), .D(n179), .Z(n182) );
    VMW_NAND2 U12 ( .A(n185), .B(B[6]), .Z(n184) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n187), .C(n182), .D(n177), .Z(n186) );
    VMW_OR2 U14 ( .A(B[6]), .B(n185), .Z(n188) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n190), .C(n188), .D(n186), .Z(n189) );
    VMW_NAND2 U16 ( .A(n192), .B(B[8]), .Z(n191) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n194), .C(n189), .D(n184), .Z(n193) );
    VMW_OR2 U18 ( .A(B[8]), .B(n192), .Z(n195) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n197), .C(n195), .D(n193), .Z(n196) );
    VMW_NAND2 U20 ( .A(n199), .B(B[10]), .Z(n198) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n201), .C(n196), .D(n191), .Z(n200) );
    VMW_NAND2 U22 ( .A(n201), .B(A[9]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n199), .C(n202), .D(n200), .Z(n203) );
    VMW_NAND2 U24 ( .A(n205), .B(B[12]), .Z(n204) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n207), .C(n203), .D(n198), .Z(n206) );
    VMW_NAND2 U26 ( .A(n207), .B(A[11]), .Z(n208) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n205), .C(n208), .D(n206), .Z(n209) );
    VMW_NAND2 U28 ( .A(n211), .B(B[14]), .Z(n210) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n213), .C(n209), .D(n204), .Z(n212) );
    VMW_NAND2 U30 ( .A(n213), .B(A[13]), .Z(n214) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n211), .C(n214), .D(n212), .Z(n215) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n216), .C(n215), .D(n210), .Z(n169) );
    VMW_INV U33 ( .A(A[12]), .Z(n205) );
    VMW_INV U34 ( .A(B[7]), .Z(n194) );
    VMW_INV U35 ( .A(A[7]), .Z(n197) );
    VMW_INV U36 ( .A(A[3]), .Z(n183) );
    VMW_INV U37 ( .A(B[3]), .Z(n180) );
    VMW_INV U38 ( .A(A[10]), .Z(n199) );
    VMW_INV U39 ( .A(B[9]), .Z(n201) );
    VMW_INV U40 ( .A(A[4]), .Z(n178) );
    VMW_INV U41 ( .A(A[8]), .Z(n192) );
    VMW_INV U42 ( .A(A[14]), .Z(n211) );
    VMW_INV U43 ( .A(B[11]), .Z(n207) );
    VMW_INV U44 ( .A(A[5]), .Z(n190) );
    VMW_INV U45 ( .A(B[5]), .Z(n187) );
    VMW_INV U46 ( .A(A[1]), .Z(n174) );
    VMW_INV U47 ( .A(B[15]), .Z(n216) );
    VMW_INV U48 ( .A(B[13]), .Z(n213) );
    VMW_INV U49 ( .A(A[6]), .Z(n185) );
    VMW_INV U50 ( .A(A[2]), .Z(n171) );
    VMW_INV U51 ( .A(A[0]), .Z(n173) );
    VMW_INV U52 ( .A(A[15]), .Z(n168) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265;
    VMW_OAI21 U3 ( .A(B[15]), .B(n217), .C(n218), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n220), .B(B[2]), .Z(n219) );
    VMW_AO22 U5 ( .A(n222), .B(B[0]), .C(n223), .D(B[1]), .Z(n221) );
    VMW_OR2 U6 ( .A(B[2]), .B(n220), .Z(n224) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n223), .C(n224), .D(n221), .Z(n225) );
    VMW_NAND2 U8 ( .A(n227), .B(B[4]), .Z(n226) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n229), .C(n225), .D(n219), .Z(n228) );
    VMW_OR2 U10 ( .A(B[4]), .B(n227), .Z(n230) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n232), .C(n230), .D(n228), .Z(n231) );
    VMW_NAND2 U12 ( .A(n234), .B(B[6]), .Z(n233) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n236), .C(n231), .D(n226), .Z(n235) );
    VMW_OR2 U14 ( .A(B[6]), .B(n234), .Z(n237) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n239), .C(n237), .D(n235), .Z(n238) );
    VMW_NAND2 U16 ( .A(n241), .B(B[8]), .Z(n240) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n243), .C(n238), .D(n233), .Z(n242) );
    VMW_OR2 U18 ( .A(B[8]), .B(n241), .Z(n244) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n246), .C(n244), .D(n242), .Z(n245) );
    VMW_NAND2 U20 ( .A(n248), .B(B[10]), .Z(n247) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n250), .C(n245), .D(n240), .Z(n249) );
    VMW_NAND2 U22 ( .A(n250), .B(A[9]), .Z(n251) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n248), .C(n251), .D(n249), .Z(n252) );
    VMW_NAND2 U24 ( .A(n254), .B(B[12]), .Z(n253) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n256), .C(n252), .D(n247), .Z(n255) );
    VMW_NAND2 U26 ( .A(n256), .B(A[11]), .Z(n257) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n254), .C(n257), .D(n255), .Z(n258) );
    VMW_NAND2 U28 ( .A(n260), .B(B[14]), .Z(n259) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n262), .C(n258), .D(n253), .Z(n261) );
    VMW_NAND2 U30 ( .A(n262), .B(A[13]), .Z(n263) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n260), .C(n263), .D(n261), .Z(n264) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n265), .C(n264), .D(n259), .Z(n218) );
    VMW_INV U33 ( .A(A[12]), .Z(n254) );
    VMW_INV U34 ( .A(B[7]), .Z(n243) );
    VMW_INV U35 ( .A(A[7]), .Z(n246) );
    VMW_INV U36 ( .A(A[3]), .Z(n232) );
    VMW_INV U37 ( .A(B[3]), .Z(n229) );
    VMW_INV U38 ( .A(A[10]), .Z(n248) );
    VMW_INV U39 ( .A(B[9]), .Z(n250) );
    VMW_INV U40 ( .A(A[4]), .Z(n227) );
    VMW_INV U41 ( .A(A[8]), .Z(n241) );
    VMW_INV U42 ( .A(A[14]), .Z(n260) );
    VMW_INV U43 ( .A(B[11]), .Z(n256) );
    VMW_INV U44 ( .A(A[5]), .Z(n239) );
    VMW_INV U45 ( .A(B[5]), .Z(n236) );
    VMW_INV U46 ( .A(A[1]), .Z(n223) );
    VMW_INV U47 ( .A(B[15]), .Z(n265) );
    VMW_INV U48 ( .A(B[13]), .Z(n262) );
    VMW_INV U49 ( .A(A[6]), .Z(n234) );
    VMW_INV U50 ( .A(A[2]), .Z(n220) );
    VMW_INV U51 ( .A(A[0]), .Z(n222) );
    VMW_INV U52 ( .A(A[15]), .Z(n217) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314;
    VMW_OAI21 U3 ( .A(B[15]), .B(n266), .C(n267), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n269), .B(B[2]), .Z(n268) );
    VMW_AO22 U5 ( .A(n271), .B(B[0]), .C(n272), .D(B[1]), .Z(n270) );
    VMW_OR2 U6 ( .A(B[2]), .B(n269), .Z(n273) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n272), .C(n273), .D(n270), .Z(n274) );
    VMW_NAND2 U8 ( .A(n276), .B(B[4]), .Z(n275) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n278), .C(n274), .D(n268), .Z(n277) );
    VMW_OR2 U10 ( .A(B[4]), .B(n276), .Z(n279) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n281), .C(n279), .D(n277), .Z(n280) );
    VMW_NAND2 U12 ( .A(n283), .B(B[6]), .Z(n282) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n285), .C(n280), .D(n275), .Z(n284) );
    VMW_OR2 U14 ( .A(B[6]), .B(n283), .Z(n286) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n288), .C(n286), .D(n284), .Z(n287) );
    VMW_NAND2 U16 ( .A(n290), .B(B[8]), .Z(n289) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n292), .C(n287), .D(n282), .Z(n291) );
    VMW_OR2 U18 ( .A(B[8]), .B(n290), .Z(n293) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n295), .C(n293), .D(n291), .Z(n294) );
    VMW_NAND2 U20 ( .A(n297), .B(B[10]), .Z(n296) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n299), .C(n294), .D(n289), .Z(n298) );
    VMW_NAND2 U22 ( .A(n299), .B(A[9]), .Z(n300) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n297), .C(n300), .D(n298), .Z(n301) );
    VMW_NAND2 U24 ( .A(n303), .B(B[12]), .Z(n302) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n305), .C(n301), .D(n296), .Z(n304) );
    VMW_NAND2 U26 ( .A(n305), .B(A[11]), .Z(n306) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n303), .C(n306), .D(n304), .Z(n307) );
    VMW_NAND2 U28 ( .A(n309), .B(B[14]), .Z(n308) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n311), .C(n307), .D(n302), .Z(n310) );
    VMW_NAND2 U30 ( .A(n311), .B(A[13]), .Z(n312) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n309), .C(n312), .D(n310), .Z(n313) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n314), .C(n313), .D(n308), .Z(n267) );
    VMW_INV U33 ( .A(A[12]), .Z(n303) );
    VMW_INV U34 ( .A(B[7]), .Z(n292) );
    VMW_INV U35 ( .A(A[7]), .Z(n295) );
    VMW_INV U36 ( .A(A[3]), .Z(n281) );
    VMW_INV U37 ( .A(B[3]), .Z(n278) );
    VMW_INV U38 ( .A(A[10]), .Z(n297) );
    VMW_INV U39 ( .A(B[9]), .Z(n299) );
    VMW_INV U40 ( .A(A[4]), .Z(n276) );
    VMW_INV U41 ( .A(A[8]), .Z(n290) );
    VMW_INV U42 ( .A(A[14]), .Z(n309) );
    VMW_INV U43 ( .A(B[11]), .Z(n305) );
    VMW_INV U44 ( .A(A[5]), .Z(n288) );
    VMW_INV U45 ( .A(B[5]), .Z(n285) );
    VMW_INV U46 ( .A(A[1]), .Z(n272) );
    VMW_INV U47 ( .A(B[15]), .Z(n314) );
    VMW_INV U48 ( .A(B[13]), .Z(n311) );
    VMW_INV U49 ( .A(A[6]), .Z(n283) );
    VMW_INV U50 ( .A(A[2]), .Z(n269) );
    VMW_INV U51 ( .A(A[0]), .Z(n271) );
    VMW_INV U52 ( .A(A[15]), .Z(n266) );
endmodule


module NodeAux_INDEGREE6_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp494[7] , \temp584[2] , n100, \OutEdge146[7] , \temp314[15] , 
        \OutEdge146[12] , \temp314[11] , \OutEdge146[3] , \temp494[3] , 
        \temp584[6] , \path[2] , \path[0] , \temp314[13] , \temp494[1] , 
        \OutEdge146[1] , \temp584[4] , \OutEdge146[8] , \temp494[8] , n132, 
        \OutEdge146[10] , \temp584[0] , \OutEdge146[5] , \temp494[5] , 
        \OutEdge146[14] , \temp584[9] , \temp220[10] , \temp220[4] , 
        \temp314[7] , \temp494[11] , \temp404[6] , \temp584[13] , 
        \temp404[11] , \temp404[2] , \temp220[0] , \temp314[3] , \temp494[15] , 
        \temp220[14] , \temp404[15] , \temp220[9] , \temp404[9] , \temp314[8] , 
        \temp220[2] , \temp404[0] , \temp314[1] , \temp584[15] , n108, 
        \temp404[13] , \temp584[11] , \temp220[12] , \temp220[6] , 
        \temp314[5] , \temp404[4] , \temp494[13] , \temp404[12] , 
        \temp584[10] , \temp220[7] , \temp314[4] , n124, \temp494[12] , 
        \temp220[13] , \temp404[5] , \temp404[8] , \temp314[9] , \temp404[1] , 
        \temp220[3] , \temp314[0] , \temp584[14] , \temp404[3] , \temp220[15] , 
        \temp220[1] , \temp314[2] , \temp494[14] , \temp220[8] , \temp404[14] , 
        n116, \temp220[5] , \temp314[6] , \temp494[10] , \temp220[11] , 
        \temp404[7] , \temp584[12] , \temp404[10] , \temp584[1] , 
        \OutEdge146[4] , \temp494[4] , \OutEdge146[15] , \temp584[8] , 
        \path[1] , \temp494[0] , \OutEdge146[0] , \temp314[12] , n92, 
        \temp584[5] , \OutEdge146[9] , \temp494[9] , \OutEdge146[11] , 
        \OutEdge146[13] , \temp494[2] , \OutEdge146[2] , \temp314[10] , 
        \path[3] , \temp584[7] , \temp584[3] , \temp314[14] , \temp494[6] , 
        \OutEdge146[6] , n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
        n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
        n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
        n812, n813, n814, n815, n816;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U91 ( .Z(n815) );
    VMW_PULLDOWN U92 ( .Z(n814) );
    VMW_PULLDOWN U93 ( .Z(n813) );
    VMW_PULLDOWN U94 ( .Z(n812) );
    VMW_PULLDOWN U95 ( .Z(n816) );
    VMW_PULLDOWN U96 ( .Z(n811) );
    VMW_NOR2 U97 ( .A(Start), .B(n767), .Z(\OutEdge146[15] ) );
    VMW_NAND2 U98 ( .A(n768), .B(n769), .Z(\OutEdge146[14] ) );
    VMW_NAND2 U99 ( .A(n770), .B(n769), .Z(\OutEdge146[13] ) );
    VMW_NAND2 U100 ( .A(n771), .B(n769), .Z(\OutEdge146[12] ) );
    VMW_NAND2 U101 ( .A(n772), .B(n769), .Z(\OutEdge146[11] ) );
    VMW_NAND2 U102 ( .A(n773), .B(n769), .Z(\OutEdge146[10] ) );
    VMW_NAND2 U103 ( .A(n774), .B(n769), .Z(\OutEdge146[9] ) );
    VMW_NAND2 U104 ( .A(n775), .B(n769), .Z(\OutEdge146[8] ) );
    VMW_NAND2 U105 ( .A(n776), .B(n769), .Z(\OutEdge146[7] ) );
    VMW_NAND2 U106 ( .A(n777), .B(n769), .Z(\OutEdge146[6] ) );
    VMW_NAND2 U107 ( .A(n778), .B(n769), .Z(\OutEdge146[5] ) );
    VMW_NAND2 U108 ( .A(n779), .B(n769), .Z(\OutEdge146[4] ) );
    VMW_NAND2 U109 ( .A(n780), .B(n769), .Z(\OutEdge146[3] ) );
    VMW_NAND2 U110 ( .A(n781), .B(n769), .Z(\OutEdge146[2] ) );
    VMW_NAND2 U111 ( .A(n782), .B(n769), .Z(\OutEdge146[1] ) );
    VMW_NAND2 U112 ( .A(n783), .B(n769), .Z(\OutEdge146[0] ) );
    VMW_AO21 U113 ( .A(Start), .B(\path[1] ), .C(n784), .Z(n810) );
    VMW_AO22 U114 ( .A(\path[3] ), .B(Start), .C(n785), .D(n786), .Z(n809) );
    VMW_OR2 U115 ( .A(n787), .B(n788), .Z(n807) );
    VMW_OR3 U116 ( .A(n785), .B(n124), .C(n132), .Z(n789) );
    VMW_AO22 U117 ( .A(\temp494[15] ), .B(n790), .C(InEdges[79]), .D(n124), 
        .Z(\temp584[15] ) );
    VMW_NAND2 U118 ( .A(n769), .B(n790), .Z(n791) );
    VMW_AND4 U119 ( .A(n792), .B(n793), .C(n794), .D(n795), .Z(n785) );
    VMW_INV U120 ( .A(Start), .Z(n769) );
    VMW_OAI22 U121 ( .A(n789), .B(Start), .C(\path[2] ), .D(n769), .Z(n796) );
    VMW_MUX2I U122 ( .A(\temp584[15] ), .B(InEdges[95]), .S(n132), .Z(n767) );
    VMW_NOR2 U123 ( .A(n132), .B(n791), .Z(n786) );
    VMW_AND3 U124 ( .A(n798), .B(n799), .C(n800), .Z(n797) );
    VMW_INV U125 ( .A(n116), .Z(n795) );
    VMW_AOI211 U126 ( .A(n794), .B(n792), .C(n108), .D(n116), .Z(n801) );
    VMW_NOR3 U127 ( .A(n801), .B(n132), .C(n791), .Z(n784) );
    VMW_OAI21 U128 ( .A(n100), .B(n794), .C(n793), .Z(n802) );
    VMW_AOI21 U129 ( .A(n795), .B(n802), .C(n791), .Z(n788) );
    VMW_AND4 U130 ( .A(n803), .B(n804), .C(n805), .D(n797), .Z(n806) );
    VMW_XNOR2 U131 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n799) );
    VMW_XNOR2 U132 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n798) );
    VMW_XNOR2 U133 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n800) );
    VMW_XNOR2 U134 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n804) );
    VMW_XNOR2 U135 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n803) );
    VMW_XNOR2 U136 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n805) );
    VMW_AO22 U137 ( .A(InEdges[9]), .B(n92), .C(OutEdge[9]), .D(n794), .Z(
        \temp220[9] ) );
    VMW_AO22 U138 ( .A(InEdges[25]), .B(n100), .C(\temp220[9] ), .D(n792), .Z(
        \temp314[9] ) );
    VMW_AO22 U139 ( .A(\temp314[9] ), .B(n793), .C(InEdges[41]), .D(n108), .Z(
        \temp404[9] ) );
    VMW_AO22 U140 ( .A(InEdges[57]), .B(n116), .C(\temp404[9] ), .D(n795), .Z(
        \temp494[9] ) );
    VMW_AO22 U141 ( .A(\temp494[9] ), .B(n790), .C(InEdges[73]), .D(n124), .Z(
        \temp584[9] ) );
    VMW_AO22 U142 ( .A(InEdges[8]), .B(n92), .C(OutEdge[8]), .D(n794), .Z(
        \temp220[8] ) );
    VMW_AO22 U143 ( .A(InEdges[24]), .B(n100), .C(\temp220[8] ), .D(n792), .Z(
        \temp314[8] ) );
    VMW_AO22 U144 ( .A(\temp314[8] ), .B(n793), .C(InEdges[40]), .D(n108), .Z(
        \temp404[8] ) );
    VMW_AO22 U145 ( .A(InEdges[56]), .B(n116), .C(\temp404[8] ), .D(n795), .Z(
        \temp494[8] ) );
    VMW_AO22 U146 ( .A(\temp494[8] ), .B(n790), .C(InEdges[72]), .D(n124), .Z(
        \temp584[8] ) );
    VMW_AO22 U147 ( .A(InEdges[7]), .B(n92), .C(OutEdge[7]), .D(n794), .Z(
        \temp220[7] ) );
    VMW_AO22 U148 ( .A(InEdges[23]), .B(n100), .C(\temp220[7] ), .D(n792), .Z(
        \temp314[7] ) );
    VMW_AO22 U149 ( .A(\temp314[7] ), .B(n793), .C(InEdges[39]), .D(n108), .Z(
        \temp404[7] ) );
    VMW_AO22 U150 ( .A(InEdges[55]), .B(n116), .C(\temp404[7] ), .D(n795), .Z(
        \temp494[7] ) );
    VMW_AO22 U151 ( .A(\temp494[7] ), .B(n790), .C(InEdges[71]), .D(n124), .Z(
        \temp584[7] ) );
    VMW_AO22 U152 ( .A(InEdges[6]), .B(n92), .C(OutEdge[6]), .D(n794), .Z(
        \temp220[6] ) );
    VMW_AO22 U153 ( .A(InEdges[22]), .B(n100), .C(\temp220[6] ), .D(n792), .Z(
        \temp314[6] ) );
    VMW_AO22 U154 ( .A(\temp314[6] ), .B(n793), .C(InEdges[38]), .D(n108), .Z(
        \temp404[6] ) );
    VMW_AO22 U155 ( .A(InEdges[54]), .B(n116), .C(\temp404[6] ), .D(n795), .Z(
        \temp494[6] ) );
    VMW_AO22 U156 ( .A(\temp494[6] ), .B(n790), .C(InEdges[70]), .D(n124), .Z(
        \temp584[6] ) );
    VMW_AO22 U157 ( .A(InEdges[5]), .B(n92), .C(OutEdge[5]), .D(n794), .Z(
        \temp220[5] ) );
    VMW_AO22 U158 ( .A(InEdges[21]), .B(n100), .C(\temp220[5] ), .D(n792), .Z(
        \temp314[5] ) );
    VMW_AO22 U159 ( .A(\temp314[5] ), .B(n793), .C(InEdges[37]), .D(n108), .Z(
        \temp404[5] ) );
    VMW_AO22 U160 ( .A(InEdges[53]), .B(n116), .C(\temp404[5] ), .D(n795), .Z(
        \temp494[5] ) );
    VMW_AO22 U161 ( .A(\temp494[5] ), .B(n790), .C(InEdges[69]), .D(n124), .Z(
        \temp584[5] ) );
    VMW_AO22 U162 ( .A(InEdges[4]), .B(n92), .C(OutEdge[4]), .D(n794), .Z(
        \temp220[4] ) );
    VMW_AO22 U163 ( .A(InEdges[20]), .B(n100), .C(\temp220[4] ), .D(n792), .Z(
        \temp314[4] ) );
    VMW_AO22 U164 ( .A(\temp314[4] ), .B(n793), .C(InEdges[36]), .D(n108), .Z(
        \temp404[4] ) );
    VMW_AO22 U165 ( .A(InEdges[52]), .B(n116), .C(\temp404[4] ), .D(n795), .Z(
        \temp494[4] ) );
    VMW_AO22 U166 ( .A(\temp494[4] ), .B(n790), .C(InEdges[68]), .D(n124), .Z(
        \temp584[4] ) );
    VMW_AO22 U167 ( .A(InEdges[3]), .B(n92), .C(OutEdge[3]), .D(n794), .Z(
        \temp220[3] ) );
    VMW_AO22 U168 ( .A(InEdges[19]), .B(n100), .C(\temp220[3] ), .D(n792), .Z(
        \temp314[3] ) );
    VMW_AO22 U169 ( .A(\temp314[3] ), .B(n793), .C(InEdges[35]), .D(n108), .Z(
        \temp404[3] ) );
    VMW_AO22 U170 ( .A(InEdges[51]), .B(n116), .C(\temp404[3] ), .D(n795), .Z(
        \temp494[3] ) );
    VMW_AO22 U171 ( .A(\temp494[3] ), .B(n790), .C(InEdges[67]), .D(n124), .Z(
        \temp584[3] ) );
    VMW_AO22 U172 ( .A(InEdges[2]), .B(n92), .C(OutEdge[2]), .D(n794), .Z(
        \temp220[2] ) );
    VMW_AO22 U173 ( .A(InEdges[18]), .B(n100), .C(\temp220[2] ), .D(n792), .Z(
        \temp314[2] ) );
    VMW_AO22 U174 ( .A(\temp314[2] ), .B(n793), .C(InEdges[34]), .D(n108), .Z(
        \temp404[2] ) );
    VMW_AO22 U175 ( .A(InEdges[50]), .B(n116), .C(\temp404[2] ), .D(n795), .Z(
        \temp494[2] ) );
    VMW_AO22 U176 ( .A(\temp494[2] ), .B(n790), .C(InEdges[66]), .D(n124), .Z(
        \temp584[2] ) );
    VMW_AO22 U177 ( .A(InEdges[1]), .B(n92), .C(OutEdge[1]), .D(n794), .Z(
        \temp220[1] ) );
    VMW_AO22 U178 ( .A(InEdges[17]), .B(n100), .C(\temp220[1] ), .D(n792), .Z(
        \temp314[1] ) );
    VMW_AO22 U179 ( .A(\temp314[1] ), .B(n793), .C(InEdges[33]), .D(n108), .Z(
        \temp404[1] ) );
    VMW_AO22 U180 ( .A(InEdges[49]), .B(n116), .C(\temp404[1] ), .D(n795), .Z(
        \temp494[1] ) );
    VMW_AO22 U181 ( .A(\temp494[1] ), .B(n790), .C(InEdges[65]), .D(n124), .Z(
        \temp584[1] ) );
    VMW_AO22 U182 ( .A(InEdges[15]), .B(n92), .C(OutEdge[15]), .D(n794), .Z(
        \temp220[15] ) );
    VMW_AO22 U183 ( .A(InEdges[31]), .B(n100), .C(\temp220[15] ), .D(n792), 
        .Z(\temp314[15] ) );
    VMW_AO22 U184 ( .A(\temp314[15] ), .B(n793), .C(InEdges[47]), .D(n108), 
        .Z(\temp404[15] ) );
    VMW_AO22 U185 ( .A(InEdges[63]), .B(n116), .C(\temp404[15] ), .D(n795), 
        .Z(\temp494[15] ) );
    VMW_AO22 U186 ( .A(InEdges[14]), .B(n92), .C(OutEdge[14]), .D(n794), .Z(
        \temp220[14] ) );
    VMW_AO22 U187 ( .A(InEdges[30]), .B(n100), .C(\temp220[14] ), .D(n792), 
        .Z(\temp314[14] ) );
    VMW_AO22 U188 ( .A(\temp314[14] ), .B(n793), .C(InEdges[46]), .D(n108), 
        .Z(\temp404[14] ) );
    VMW_AO22 U189 ( .A(InEdges[62]), .B(n116), .C(\temp404[14] ), .D(n795), 
        .Z(\temp494[14] ) );
    VMW_AO22 U190 ( .A(\temp494[14] ), .B(n790), .C(InEdges[78]), .D(n124), 
        .Z(\temp584[14] ) );
    VMW_AO22 U191 ( .A(InEdges[13]), .B(n92), .C(OutEdge[13]), .D(n794), .Z(
        \temp220[13] ) );
    VMW_AO22 U192 ( .A(InEdges[29]), .B(n100), .C(\temp220[13] ), .D(n792), 
        .Z(\temp314[13] ) );
    VMW_AO22 U193 ( .A(\temp314[13] ), .B(n793), .C(InEdges[45]), .D(n108), 
        .Z(\temp404[13] ) );
    VMW_AO22 U194 ( .A(InEdges[61]), .B(n116), .C(\temp404[13] ), .D(n795), 
        .Z(\temp494[13] ) );
    VMW_AO22 U195 ( .A(\temp494[13] ), .B(n790), .C(InEdges[77]), .D(n124), 
        .Z(\temp584[13] ) );
    VMW_AO22 U196 ( .A(InEdges[12]), .B(n92), .C(OutEdge[12]), .D(n794), .Z(
        \temp220[12] ) );
    VMW_AO22 U197 ( .A(InEdges[28]), .B(n100), .C(\temp220[12] ), .D(n792), 
        .Z(\temp314[12] ) );
    VMW_AO22 U198 ( .A(\temp314[12] ), .B(n793), .C(InEdges[44]), .D(n108), 
        .Z(\temp404[12] ) );
    VMW_AO22 U199 ( .A(InEdges[60]), .B(n116), .C(\temp404[12] ), .D(n795), 
        .Z(\temp494[12] ) );
    VMW_AO22 U200 ( .A(\temp494[12] ), .B(n790), .C(InEdges[76]), .D(n124), 
        .Z(\temp584[12] ) );
    VMW_AO22 U201 ( .A(InEdges[11]), .B(n92), .C(OutEdge[11]), .D(n794), .Z(
        \temp220[11] ) );
    VMW_AO22 U202 ( .A(InEdges[27]), .B(n100), .C(\temp220[11] ), .D(n792), 
        .Z(\temp314[11] ) );
    VMW_AO22 U203 ( .A(\temp314[11] ), .B(n793), .C(InEdges[43]), .D(n108), 
        .Z(\temp404[11] ) );
    VMW_AO22 U204 ( .A(InEdges[59]), .B(n116), .C(\temp404[11] ), .D(n795), 
        .Z(\temp494[11] ) );
    VMW_AO22 U205 ( .A(\temp494[11] ), .B(n790), .C(InEdges[75]), .D(n124), 
        .Z(\temp584[11] ) );
    VMW_AO22 U206 ( .A(InEdges[10]), .B(n92), .C(OutEdge[10]), .D(n794), .Z(
        \temp220[10] ) );
    VMW_AO22 U207 ( .A(InEdges[26]), .B(n100), .C(\temp220[10] ), .D(n792), 
        .Z(\temp314[10] ) );
    VMW_AO22 U208 ( .A(\temp314[10] ), .B(n793), .C(InEdges[42]), .D(n108), 
        .Z(\temp404[10] ) );
    VMW_AO22 U209 ( .A(InEdges[58]), .B(n116), .C(\temp404[10] ), .D(n795), 
        .Z(\temp494[10] ) );
    VMW_AO22 U210 ( .A(\temp494[10] ), .B(n790), .C(InEdges[74]), .D(n124), 
        .Z(\temp584[10] ) );
    VMW_AO22 U211 ( .A(InEdges[0]), .B(n92), .C(OutEdge[0]), .D(n794), .Z(
        \temp220[0] ) );
    VMW_AO22 U212 ( .A(InEdges[16]), .B(n100), .C(\temp220[0] ), .D(n792), .Z(
        \temp314[0] ) );
    VMW_AO22 U213 ( .A(\temp314[0] ), .B(n793), .C(InEdges[32]), .D(n108), .Z(
        \temp404[0] ) );
    VMW_AO22 U214 ( .A(InEdges[48]), .B(n116), .C(\temp404[0] ), .D(n795), .Z(
        \temp494[0] ) );
    VMW_AO22 U215 ( .A(\temp494[0] ), .B(n790), .C(InEdges[64]), .D(n124), .Z(
        \temp584[0] ) );
    VMW_AO22 U216 ( .A(n132), .B(n769), .C(\path[0] ), .D(Start), .Z(n787) );
    VMW_MUX2I U217 ( .A(\temp584[9] ), .B(InEdges[89]), .S(n132), .Z(n774) );
    VMW_MUX2I U218 ( .A(\temp584[8] ), .B(InEdges[88]), .S(n132), .Z(n775) );
    VMW_MUX2I U219 ( .A(\temp584[7] ), .B(InEdges[87]), .S(n132), .Z(n776) );
    VMW_MUX2I U220 ( .A(\temp584[6] ), .B(InEdges[86]), .S(n132), .Z(n777) );
    VMW_MUX2I U221 ( .A(\temp584[5] ), .B(InEdges[85]), .S(n132), .Z(n778) );
    VMW_MUX2I U222 ( .A(\temp584[4] ), .B(InEdges[84]), .S(n132), .Z(n779) );
    VMW_MUX2I U223 ( .A(\temp584[3] ), .B(InEdges[83]), .S(n132), .Z(n780) );
    VMW_MUX2I U224 ( .A(\temp584[2] ), .B(InEdges[82]), .S(n132), .Z(n781) );
    VMW_MUX2I U225 ( .A(\temp584[1] ), .B(InEdges[81]), .S(n132), .Z(n782) );
    VMW_MUX2I U226 ( .A(\temp584[14] ), .B(InEdges[94]), .S(n132), .Z(n768) );
    VMW_MUX2I U227 ( .A(\temp584[13] ), .B(InEdges[93]), .S(n132), .Z(n770) );
    VMW_MUX2I U228 ( .A(\temp584[12] ), .B(InEdges[92]), .S(n132), .Z(n771) );
    VMW_MUX2I U229 ( .A(\temp584[11] ), .B(InEdges[91]), .S(n132), .Z(n772) );
    VMW_MUX2I U230 ( .A(\temp584[10] ), .B(InEdges[90]), .S(n132), .Z(n773) );
    VMW_MUX2I U231 ( .A(\temp584[0] ), .B(InEdges[80]), .S(n132), .Z(n783) );
    VMW_INV U232 ( .A(n100), .Z(n792) );
    VMW_INV U233 ( .A(n92), .Z(n794) );
    VMW_INV U234 ( .A(n108), .Z(n793) );
    VMW_INV U235 ( .A(n124), .Z(n790) );
    VMW_INV U236 ( .A(n796), .Z(n808) );
    VMW_BUFIZ U237 ( .A(\path[3] ), .E(n806), .Z(\PathData[3] ) );
    VMW_BUFIZ U238 ( .A(\path[1] ), .E(n806), .Z(\PathData[1] ) );
    VMW_BUFIZ U239 ( .A(\path[0] ), .E(n806), .Z(\PathData[0] ) );
    VMW_BUFIZ U240 ( .A(\path[2] ), .E(n806), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n807), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n808), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n809), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n810), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge146[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge146[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge146[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge146[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge146[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge146[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge146[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge146[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge146[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge146[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge146[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge146[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge146[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge146[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge146[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge146[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 lte_55_1 ( .A({\temp220[15] , 
        \temp220[14] , \temp220[13] , \temp220[12] , \temp220[11] , 
        \temp220[10] , \temp220[9] , \temp220[8] , \temp220[7] , \temp220[6] , 
        \temp220[5] , \temp220[4] , \temp220[3] , \temp220[2] , \temp220[1] , 
        \temp220[0] }), .B(InEdges[31:16]), .LEQ(n816), .TC(n816), .GE_GT(n100
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp584[15] , 
        \temp584[14] , \temp584[13] , \temp584[12] , \temp584[11] , 
        \temp584[10] , \temp584[9] , \temp584[8] , \temp584[7] , \temp584[6] , 
        \temp584[5] , \temp584[4] , \temp584[3] , \temp584[2] , \temp584[1] , 
        \temp584[0] }), .B(InEdges[95:80]), .LEQ(n815), .TC(n815), .GE_GT(n132
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp494[15] , 
        \temp494[14] , \temp494[13] , \temp494[12] , \temp494[11] , 
        \temp494[10] , \temp494[9] , \temp494[8] , \temp494[7] , \temp494[6] , 
        \temp494[5] , \temp494[4] , \temp494[3] , \temp494[2] , \temp494[1] , 
        \temp494[0] }), .B(InEdges[79:64]), .LEQ(n814), .TC(n814), .GE_GT(n124
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 lte_55_3 ( .A({\temp404[15] , 
        \temp404[14] , \temp404[13] , \temp404[12] , \temp404[11] , 
        \temp404[10] , \temp404[9] , \temp404[8] , \temp404[7] , \temp404[6] , 
        \temp404[5] , \temp404[4] , \temp404[3] , \temp404[2] , \temp404[1] , 
        \temp404[0] }), .B(InEdges[63:48]), .LEQ(n813), .TC(n813), .GE_GT(n116
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp314[15] , 
        \temp314[14] , \temp314[13] , \temp314[12] , \temp314[11] , 
        \temp314[10] , \temp314[9] , \temp314[8] , \temp314[7] , \temp314[6] , 
        \temp314[5] , \temp314[4] , \temp314[3] , \temp314[2] , \temp314[1] , 
        \temp314[0] }), .B(InEdges[47:32]), .LEQ(n812), .TC(n812), .GE_GT(n108
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n811), .TC(n811), .GE_GT(n92) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, 
        n107, n108, n109, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n101), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n119, n120, n121, n122, n123, n124, n125, n127, n128, 
        n129, n130, n131, n132, n133, n135, n136, n137, n138, n139, n140, n141, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n144), .B(B[8]), .Z(n143) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n135), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n144), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n153), .C(n148), .D(n143), .Z(n152) );
    VMW_NAND2 U22 ( .A(n153), .B(A[9]), .Z(n154) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U24 ( .A(n157), .B(B[12]), .Z(n156) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_NAND2 U26 ( .A(n159), .B(A[11]), .Z(n160) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_NAND2 U28 ( .A(n163), .B(B[14]), .Z(n162) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_NAND2 U30 ( .A(n165), .B(A[13]), .Z(n166) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n163), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n168), .C(n167), .D(n162), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n157) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n153) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n144) );
    VMW_INV U42 ( .A(A[14]), .Z(n163) );
    VMW_INV U43 ( .A(B[11]), .Z(n159) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n168) );
    VMW_INV U48 ( .A(B[13]), .Z(n165) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
        n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
        n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
        n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
        n216, n217;
    VMW_OAI21 U3 ( .A(B[15]), .B(n169), .C(n170), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n172), .B(B[2]), .Z(n171) );
    VMW_AO22 U5 ( .A(n174), .B(B[0]), .C(n175), .D(B[1]), .Z(n173) );
    VMW_OR2 U6 ( .A(B[2]), .B(n172), .Z(n176) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n175), .C(n176), .D(n173), .Z(n177) );
    VMW_NAND2 U8 ( .A(n179), .B(B[4]), .Z(n178) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n181), .C(n177), .D(n171), .Z(n180) );
    VMW_OR2 U10 ( .A(B[4]), .B(n179), .Z(n182) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n184), .C(n182), .D(n180), .Z(n183) );
    VMW_NAND2 U12 ( .A(n186), .B(B[6]), .Z(n185) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n188), .C(n183), .D(n178), .Z(n187) );
    VMW_OR2 U14 ( .A(B[6]), .B(n186), .Z(n189) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n191), .C(n189), .D(n187), .Z(n190) );
    VMW_NAND2 U16 ( .A(n193), .B(B[8]), .Z(n192) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n195), .C(n190), .D(n185), .Z(n194) );
    VMW_OR2 U18 ( .A(B[8]), .B(n193), .Z(n196) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n198), .C(n196), .D(n194), .Z(n197) );
    VMW_NAND2 U20 ( .A(n200), .B(B[10]), .Z(n199) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n202), .C(n197), .D(n192), .Z(n201) );
    VMW_NAND2 U22 ( .A(n202), .B(A[9]), .Z(n203) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n200), .C(n203), .D(n201), .Z(n204) );
    VMW_NAND2 U24 ( .A(n206), .B(B[12]), .Z(n205) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n208), .C(n204), .D(n199), .Z(n207) );
    VMW_NAND2 U26 ( .A(n208), .B(A[11]), .Z(n209) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n206), .C(n209), .D(n207), .Z(n210) );
    VMW_NAND2 U28 ( .A(n212), .B(B[14]), .Z(n211) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n214), .C(n210), .D(n205), .Z(n213) );
    VMW_NAND2 U30 ( .A(n214), .B(A[13]), .Z(n215) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n212), .C(n215), .D(n213), .Z(n216) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n217), .C(n216), .D(n211), .Z(n170) );
    VMW_INV U33 ( .A(A[12]), .Z(n206) );
    VMW_INV U34 ( .A(B[7]), .Z(n195) );
    VMW_INV U35 ( .A(A[7]), .Z(n198) );
    VMW_INV U36 ( .A(A[3]), .Z(n184) );
    VMW_INV U37 ( .A(B[3]), .Z(n181) );
    VMW_INV U38 ( .A(A[10]), .Z(n200) );
    VMW_INV U39 ( .A(B[9]), .Z(n202) );
    VMW_INV U40 ( .A(A[4]), .Z(n179) );
    VMW_INV U41 ( .A(A[8]), .Z(n193) );
    VMW_INV U42 ( .A(A[14]), .Z(n212) );
    VMW_INV U43 ( .A(B[11]), .Z(n208) );
    VMW_INV U44 ( .A(A[5]), .Z(n191) );
    VMW_INV U45 ( .A(B[5]), .Z(n188) );
    VMW_INV U46 ( .A(A[1]), .Z(n175) );
    VMW_INV U47 ( .A(B[15]), .Z(n217) );
    VMW_INV U48 ( .A(B[13]), .Z(n214) );
    VMW_INV U49 ( .A(A[6]), .Z(n186) );
    VMW_INV U50 ( .A(A[2]), .Z(n172) );
    VMW_INV U51 ( .A(A[0]), .Z(n174) );
    VMW_INV U52 ( .A(A[15]), .Z(n169) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266;
    VMW_OAI21 U3 ( .A(B[15]), .B(n218), .C(n219), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n221), .B(B[2]), .Z(n220) );
    VMW_AO22 U5 ( .A(n223), .B(B[0]), .C(n224), .D(B[1]), .Z(n222) );
    VMW_OR2 U6 ( .A(B[2]), .B(n221), .Z(n225) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n224), .C(n225), .D(n222), .Z(n226) );
    VMW_NAND2 U8 ( .A(n228), .B(B[4]), .Z(n227) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n230), .C(n226), .D(n220), .Z(n229) );
    VMW_OR2 U10 ( .A(B[4]), .B(n228), .Z(n231) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n233), .C(n231), .D(n229), .Z(n232) );
    VMW_NAND2 U12 ( .A(n235), .B(B[6]), .Z(n234) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n237), .C(n232), .D(n227), .Z(n236) );
    VMW_OR2 U14 ( .A(B[6]), .B(n235), .Z(n238) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n240), .C(n238), .D(n236), .Z(n239) );
    VMW_NAND2 U16 ( .A(n242), .B(B[8]), .Z(n241) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n244), .C(n239), .D(n234), .Z(n243) );
    VMW_OR2 U18 ( .A(B[8]), .B(n242), .Z(n245) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n247), .C(n245), .D(n243), .Z(n246) );
    VMW_NAND2 U20 ( .A(n249), .B(B[10]), .Z(n248) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n251), .C(n246), .D(n241), .Z(n250) );
    VMW_NAND2 U22 ( .A(n251), .B(A[9]), .Z(n252) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n249), .C(n252), .D(n250), .Z(n253) );
    VMW_NAND2 U24 ( .A(n255), .B(B[12]), .Z(n254) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n257), .C(n253), .D(n248), .Z(n256) );
    VMW_NAND2 U26 ( .A(n257), .B(A[11]), .Z(n258) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n255), .C(n258), .D(n256), .Z(n259) );
    VMW_NAND2 U28 ( .A(n261), .B(B[14]), .Z(n260) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n263), .C(n259), .D(n254), .Z(n262) );
    VMW_NAND2 U30 ( .A(n263), .B(A[13]), .Z(n264) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n261), .C(n264), .D(n262), .Z(n265) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n266), .C(n265), .D(n260), .Z(n219) );
    VMW_INV U33 ( .A(A[12]), .Z(n255) );
    VMW_INV U34 ( .A(B[7]), .Z(n244) );
    VMW_INV U35 ( .A(A[7]), .Z(n247) );
    VMW_INV U36 ( .A(A[3]), .Z(n233) );
    VMW_INV U37 ( .A(B[3]), .Z(n230) );
    VMW_INV U38 ( .A(A[10]), .Z(n249) );
    VMW_INV U39 ( .A(B[9]), .Z(n251) );
    VMW_INV U40 ( .A(A[4]), .Z(n228) );
    VMW_INV U41 ( .A(A[8]), .Z(n242) );
    VMW_INV U42 ( .A(A[14]), .Z(n261) );
    VMW_INV U43 ( .A(B[11]), .Z(n257) );
    VMW_INV U44 ( .A(A[5]), .Z(n240) );
    VMW_INV U45 ( .A(B[5]), .Z(n237) );
    VMW_INV U46 ( .A(A[1]), .Z(n224) );
    VMW_INV U47 ( .A(B[15]), .Z(n266) );
    VMW_INV U48 ( .A(B[13]), .Z(n263) );
    VMW_INV U49 ( .A(A[6]), .Z(n235) );
    VMW_INV U50 ( .A(A[2]), .Z(n221) );
    VMW_INV U51 ( .A(A[0]), .Z(n223) );
    VMW_INV U52 ( .A(A[15]), .Z(n218) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315;
    VMW_OAI21 U3 ( .A(B[15]), .B(n267), .C(n268), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n270), .B(B[2]), .Z(n269) );
    VMW_AO22 U5 ( .A(n272), .B(B[0]), .C(n273), .D(B[1]), .Z(n271) );
    VMW_OR2 U6 ( .A(B[2]), .B(n270), .Z(n274) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n273), .C(n274), .D(n271), .Z(n275) );
    VMW_NAND2 U8 ( .A(n277), .B(B[4]), .Z(n276) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n279), .C(n275), .D(n269), .Z(n278) );
    VMW_OR2 U10 ( .A(B[4]), .B(n277), .Z(n280) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n282), .C(n280), .D(n278), .Z(n281) );
    VMW_NAND2 U12 ( .A(n284), .B(B[6]), .Z(n283) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n286), .C(n281), .D(n276), .Z(n285) );
    VMW_OR2 U14 ( .A(B[6]), .B(n284), .Z(n287) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n289), .C(n287), .D(n285), .Z(n288) );
    VMW_NAND2 U16 ( .A(n291), .B(B[8]), .Z(n290) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n293), .C(n288), .D(n283), .Z(n292) );
    VMW_OR2 U18 ( .A(B[8]), .B(n291), .Z(n294) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n296), .C(n294), .D(n292), .Z(n295) );
    VMW_NAND2 U20 ( .A(n298), .B(B[10]), .Z(n297) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n300), .C(n295), .D(n290), .Z(n299) );
    VMW_NAND2 U22 ( .A(n300), .B(A[9]), .Z(n301) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n298), .C(n301), .D(n299), .Z(n302) );
    VMW_NAND2 U24 ( .A(n304), .B(B[12]), .Z(n303) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n306), .C(n302), .D(n297), .Z(n305) );
    VMW_NAND2 U26 ( .A(n306), .B(A[11]), .Z(n307) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n304), .C(n307), .D(n305), .Z(n308) );
    VMW_NAND2 U28 ( .A(n310), .B(B[14]), .Z(n309) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n312), .C(n308), .D(n303), .Z(n311) );
    VMW_NAND2 U30 ( .A(n312), .B(A[13]), .Z(n313) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n310), .C(n313), .D(n311), .Z(n314) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n315), .C(n314), .D(n309), .Z(n268) );
    VMW_INV U33 ( .A(A[12]), .Z(n304) );
    VMW_INV U34 ( .A(B[7]), .Z(n293) );
    VMW_INV U35 ( .A(A[7]), .Z(n296) );
    VMW_INV U36 ( .A(A[3]), .Z(n282) );
    VMW_INV U37 ( .A(B[3]), .Z(n279) );
    VMW_INV U38 ( .A(A[10]), .Z(n298) );
    VMW_INV U39 ( .A(B[9]), .Z(n300) );
    VMW_INV U40 ( .A(A[4]), .Z(n277) );
    VMW_INV U41 ( .A(A[8]), .Z(n291) );
    VMW_INV U42 ( .A(A[14]), .Z(n310) );
    VMW_INV U43 ( .A(B[11]), .Z(n306) );
    VMW_INV U44 ( .A(A[5]), .Z(n289) );
    VMW_INV U45 ( .A(B[5]), .Z(n286) );
    VMW_INV U46 ( .A(A[1]), .Z(n273) );
    VMW_INV U47 ( .A(B[15]), .Z(n315) );
    VMW_INV U48 ( .A(B[13]), .Z(n312) );
    VMW_INV U49 ( .A(A[6]), .Z(n284) );
    VMW_INV U50 ( .A(A[2]), .Z(n270) );
    VMW_INV U51 ( .A(A[0]), .Z(n272) );
    VMW_INV U52 ( .A(A[15]), .Z(n267) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
        n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
        n363, n364;
    VMW_OAI21 U3 ( .A(B[15]), .B(n316), .C(n317), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n319), .B(B[2]), .Z(n318) );
    VMW_AO22 U5 ( .A(n321), .B(B[0]), .C(n322), .D(B[1]), .Z(n320) );
    VMW_OR2 U6 ( .A(B[2]), .B(n319), .Z(n323) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n322), .C(n323), .D(n320), .Z(n324) );
    VMW_NAND2 U8 ( .A(n326), .B(B[4]), .Z(n325) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n328), .C(n324), .D(n318), .Z(n327) );
    VMW_OR2 U10 ( .A(B[4]), .B(n326), .Z(n329) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n331), .C(n329), .D(n327), .Z(n330) );
    VMW_NAND2 U12 ( .A(n333), .B(B[6]), .Z(n332) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n335), .C(n330), .D(n325), .Z(n334) );
    VMW_OR2 U14 ( .A(B[6]), .B(n333), .Z(n336) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n338), .C(n336), .D(n334), .Z(n337) );
    VMW_NAND2 U16 ( .A(n340), .B(B[8]), .Z(n339) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n342), .C(n337), .D(n332), .Z(n341) );
    VMW_OR2 U18 ( .A(B[8]), .B(n340), .Z(n343) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n345), .C(n343), .D(n341), .Z(n344) );
    VMW_NAND2 U20 ( .A(n347), .B(B[10]), .Z(n346) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n349), .C(n344), .D(n339), .Z(n348) );
    VMW_NAND2 U22 ( .A(n349), .B(A[9]), .Z(n350) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n347), .C(n350), .D(n348), .Z(n351) );
    VMW_NAND2 U24 ( .A(n353), .B(B[12]), .Z(n352) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n355), .C(n351), .D(n346), .Z(n354) );
    VMW_NAND2 U26 ( .A(n355), .B(A[11]), .Z(n356) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n353), .C(n356), .D(n354), .Z(n357) );
    VMW_NAND2 U28 ( .A(n359), .B(B[14]), .Z(n358) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n361), .C(n357), .D(n352), .Z(n360) );
    VMW_NAND2 U30 ( .A(n361), .B(A[13]), .Z(n362) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n359), .C(n362), .D(n360), .Z(n363) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n364), .C(n363), .D(n358), .Z(n317) );
    VMW_INV U33 ( .A(A[12]), .Z(n353) );
    VMW_INV U34 ( .A(B[7]), .Z(n342) );
    VMW_INV U35 ( .A(A[7]), .Z(n345) );
    VMW_INV U36 ( .A(A[3]), .Z(n331) );
    VMW_INV U37 ( .A(B[3]), .Z(n328) );
    VMW_INV U38 ( .A(A[10]), .Z(n347) );
    VMW_INV U39 ( .A(B[9]), .Z(n349) );
    VMW_INV U40 ( .A(A[4]), .Z(n326) );
    VMW_INV U41 ( .A(A[8]), .Z(n340) );
    VMW_INV U42 ( .A(A[14]), .Z(n359) );
    VMW_INV U43 ( .A(B[11]), .Z(n355) );
    VMW_INV U44 ( .A(A[5]), .Z(n338) );
    VMW_INV U45 ( .A(B[5]), .Z(n335) );
    VMW_INV U46 ( .A(A[1]), .Z(n322) );
    VMW_INV U47 ( .A(B[15]), .Z(n364) );
    VMW_INV U48 ( .A(B[13]), .Z(n361) );
    VMW_INV U49 ( .A(A[6]), .Z(n333) );
    VMW_INV U50 ( .A(A[2]), .Z(n319) );
    VMW_INV U51 ( .A(A[0]), .Z(n321) );
    VMW_INV U52 ( .A(A[15]), .Z(n316) );
endmodule


module NodeAux_INDEGREE7_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \OutEdge156[4] , \temp324[9] , \temp594[1] , \temp324[0] , 
        \temp594[8] , \OutEdge156[10] , \OutEdge156[0] , \temp594[5] , 
        \temp684[12] , \OutEdge156[14] , \path[2] , \OutEdge156[9] , 
        \temp324[4] , \path[0] , \temp324[6] , \temp684[10] , \temp594[7] , 
        \OutEdge156[2] , \OutEdge156[12] , \temp324[2] , \OutEdge156[6] , 
        \temp594[3] , \temp684[14] , \temp504[15] , \temp684[8] , \temp504[9] , 
        \temp414[5] , \temp230[7] , \temp504[0] , \temp594[15] , \temp684[1] , 
        \temp414[13] , \temp414[8] , \temp504[11] , \temp684[5] , 
        \temp594[11] , \temp324[12] , \temp230[3] , \temp504[4] , \temp414[1] , 
        \temp230[12] , \temp230[1] , \temp504[6] , \temp414[3] , \temp230[10] , 
        n126, \temp594[13] , \temp684[7] , \temp324[10] , \temp504[13] , 
        \temp230[8] , \temp414[11] , \temp324[14] , \temp684[3] , 
        \temp230[14] , \temp414[7] , \temp230[5] , \temp504[2] , \temp414[15] , 
        n134, \temp324[15] , n118, \temp684[2] , \temp414[6] , \temp230[15] , 
        n94, \temp504[3] , \temp230[4] , \temp414[14] , \temp230[0] , 
        \temp504[7] , \temp230[11] , \temp414[2] , \temp684[6] , \temp594[12] , 
        \temp324[11] , \temp504[12] , \temp230[9] , \temp414[10] , 
        \temp414[9] , \temp414[12] , \temp504[10] , \temp684[4] , 
        \temp594[10] , \temp324[13] , \temp230[2] , \temp504[5] , 
        \temp230[13] , \temp414[0] , \temp504[14] , \temp684[9] , \temp504[8] , 
        \temp414[4] , \temp230[6] , \temp504[1] , \temp684[0] , \temp594[14] , 
        \OutEdge156[13] , \temp324[3] , \OutEdge156[7] , \temp594[2] , 
        \temp684[15] , \temp324[7] , \path[1] , \temp684[11] , \temp594[6] , 
        \OutEdge156[3] , n102, \temp594[4] , \OutEdge156[1] , \temp684[13] , 
        \path[3] , \OutEdge156[15] , \temp324[5] , \OutEdge156[8] , 
        \OutEdge156[5] , n142, \temp324[8] , \temp594[0] , \OutEdge156[11] , 
        \temp594[9] , \temp324[1] , n110, n867, n868, n869, n870, n871, n872, 
        n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
        n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
        n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
        n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U100 ( .Z(n916) );
    VMW_PULLDOWN U101 ( .Z(n920) );
    VMW_PULLDOWN U102 ( .Z(n918) );
    VMW_PULLDOWN U103 ( .Z(n919) );
    VMW_PULLDOWN U104 ( .Z(n915) );
    VMW_PULLDOWN U105 ( .Z(n914) );
    VMW_PULLDOWN U106 ( .Z(n917) );
    VMW_AO21 U107 ( .A(\temp684[15] ), .B(n867), .C(n868), .Z(\OutEdge156[15] 
        ) );
    VMW_NAND2 U108 ( .A(n869), .B(n870), .Z(\OutEdge156[14] ) );
    VMW_NAND2 U109 ( .A(n871), .B(n870), .Z(\OutEdge156[13] ) );
    VMW_NAND2 U110 ( .A(n872), .B(n870), .Z(\OutEdge156[12] ) );
    VMW_NAND2 U111 ( .A(n873), .B(n870), .Z(\OutEdge156[11] ) );
    VMW_NAND2 U112 ( .A(n874), .B(n870), .Z(\OutEdge156[10] ) );
    VMW_NAND2 U113 ( .A(n875), .B(n870), .Z(\OutEdge156[9] ) );
    VMW_NAND2 U114 ( .A(n876), .B(n870), .Z(\OutEdge156[8] ) );
    VMW_NAND2 U115 ( .A(n877), .B(n870), .Z(\OutEdge156[7] ) );
    VMW_NAND2 U116 ( .A(n878), .B(n870), .Z(\OutEdge156[6] ) );
    VMW_NAND2 U117 ( .A(n879), .B(n870), .Z(\OutEdge156[5] ) );
    VMW_NAND2 U118 ( .A(n880), .B(n870), .Z(\OutEdge156[4] ) );
    VMW_NAND2 U119 ( .A(n881), .B(n870), .Z(\OutEdge156[3] ) );
    VMW_NAND2 U120 ( .A(n882), .B(n870), .Z(\OutEdge156[2] ) );
    VMW_NAND2 U121 ( .A(n883), .B(n870), .Z(\OutEdge156[1] ) );
    VMW_NAND2 U122 ( .A(n884), .B(n870), .Z(\OutEdge156[0] ) );
    VMW_AO21 U123 ( .A(Start), .B(\path[3] ), .C(n885), .Z(n912) );
    VMW_AO22 U124 ( .A(\path[0] ), .B(Start), .C(n867), .D(n886), .Z(n910) );
    VMW_AND4 U125 ( .A(n887), .B(n888), .C(n867), .D(n889), .Z(n885) );
    VMW_OR4 U126 ( .A(n142), .B(n126), .C(n134), .D(n889), .Z(n890) );
    VMW_AND3 U127 ( .A(n888), .B(n887), .C(n892), .Z(n891) );
    VMW_OR2 U128 ( .A(n891), .B(n142), .Z(n893) );
    VMW_AO22 U129 ( .A(\temp594[15] ), .B(n888), .C(InEdges[95]), .D(n134), 
        .Z(\temp684[15] ) );
    VMW_NOR2 U130 ( .A(Start), .B(n142), .Z(n867) );
    VMW_AND4 U131 ( .A(n894), .B(n895), .C(n896), .D(n897), .Z(n889) );
    VMW_INV U132 ( .A(Start), .Z(n870) );
    VMW_OAI22 U133 ( .A(\path[2] ), .B(n870), .C(n890), .D(Start), .Z(n898) );
    VMW_OAI22 U134 ( .A(\path[1] ), .B(n870), .C(n893), .D(Start), .Z(n899) );
    VMW_AND3 U135 ( .A(n901), .B(n902), .C(n903), .Z(n900) );
    VMW_INV U136 ( .A(n118), .Z(n897) );
    VMW_INV U137 ( .A(n110), .Z(n895) );
    VMW_INV U138 ( .A(n126), .Z(n887) );
    VMW_INV U139 ( .A(n134), .Z(n888) );
    VMW_OAI211 U140 ( .A(n94), .B(n102), .C(n895), .D(n897), .Z(n892) );
    VMW_AO21 U141 ( .A(n894), .B(n94), .C(n110), .Z(n904) );
    VMW_AO21 U142 ( .A(n897), .B(n904), .C(n126), .Z(n905) );
    VMW_NAND2 U143 ( .A(n888), .B(n905), .Z(n886) );
    VMW_AND4 U144 ( .A(n906), .B(n907), .C(n908), .D(n900), .Z(n909) );
    VMW_AND3 U145 ( .A(n142), .B(n870), .C(InEdges[111]), .Z(n868) );
    VMW_XNOR2 U146 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n902) );
    VMW_XNOR2 U147 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n901) );
    VMW_XNOR2 U148 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n903) );
    VMW_XNOR2 U149 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n907) );
    VMW_XNOR2 U150 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n906) );
    VMW_XNOR2 U151 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n908) );
    VMW_AO22 U152 ( .A(OutEdge[9]), .B(n896), .C(InEdges[9]), .D(n94), .Z(
        \temp230[9] ) );
    VMW_AO22 U153 ( .A(\temp230[9] ), .B(n894), .C(InEdges[25]), .D(n102), .Z(
        \temp324[9] ) );
    VMW_AO22 U154 ( .A(\temp324[9] ), .B(n895), .C(InEdges[41]), .D(n110), .Z(
        \temp414[9] ) );
    VMW_AO22 U155 ( .A(\temp414[9] ), .B(n897), .C(InEdges[57]), .D(n118), .Z(
        \temp504[9] ) );
    VMW_AO22 U156 ( .A(\temp504[9] ), .B(n887), .C(InEdges[73]), .D(n126), .Z(
        \temp594[9] ) );
    VMW_AO22 U157 ( .A(\temp594[9] ), .B(n888), .C(InEdges[89]), .D(n134), .Z(
        \temp684[9] ) );
    VMW_AO22 U158 ( .A(OutEdge[8]), .B(n896), .C(InEdges[8]), .D(n94), .Z(
        \temp230[8] ) );
    VMW_AO22 U159 ( .A(\temp230[8] ), .B(n894), .C(InEdges[24]), .D(n102), .Z(
        \temp324[8] ) );
    VMW_AO22 U160 ( .A(\temp324[8] ), .B(n895), .C(InEdges[40]), .D(n110), .Z(
        \temp414[8] ) );
    VMW_AO22 U161 ( .A(\temp414[8] ), .B(n897), .C(InEdges[56]), .D(n118), .Z(
        \temp504[8] ) );
    VMW_AO22 U162 ( .A(\temp504[8] ), .B(n887), .C(InEdges[72]), .D(n126), .Z(
        \temp594[8] ) );
    VMW_AO22 U163 ( .A(\temp594[8] ), .B(n888), .C(InEdges[88]), .D(n134), .Z(
        \temp684[8] ) );
    VMW_AO22 U164 ( .A(OutEdge[7]), .B(n896), .C(InEdges[7]), .D(n94), .Z(
        \temp230[7] ) );
    VMW_AO22 U165 ( .A(\temp230[7] ), .B(n894), .C(InEdges[23]), .D(n102), .Z(
        \temp324[7] ) );
    VMW_AO22 U166 ( .A(\temp324[7] ), .B(n895), .C(InEdges[39]), .D(n110), .Z(
        \temp414[7] ) );
    VMW_AO22 U167 ( .A(\temp414[7] ), .B(n897), .C(InEdges[55]), .D(n118), .Z(
        \temp504[7] ) );
    VMW_AO22 U168 ( .A(\temp504[7] ), .B(n887), .C(InEdges[71]), .D(n126), .Z(
        \temp594[7] ) );
    VMW_AO22 U169 ( .A(\temp594[7] ), .B(n888), .C(InEdges[87]), .D(n134), .Z(
        \temp684[7] ) );
    VMW_AO22 U170 ( .A(OutEdge[6]), .B(n896), .C(InEdges[6]), .D(n94), .Z(
        \temp230[6] ) );
    VMW_AO22 U171 ( .A(\temp230[6] ), .B(n894), .C(InEdges[22]), .D(n102), .Z(
        \temp324[6] ) );
    VMW_AO22 U172 ( .A(\temp324[6] ), .B(n895), .C(InEdges[38]), .D(n110), .Z(
        \temp414[6] ) );
    VMW_AO22 U173 ( .A(\temp414[6] ), .B(n897), .C(InEdges[54]), .D(n118), .Z(
        \temp504[6] ) );
    VMW_AO22 U174 ( .A(\temp504[6] ), .B(n887), .C(InEdges[70]), .D(n126), .Z(
        \temp594[6] ) );
    VMW_AO22 U175 ( .A(\temp594[6] ), .B(n888), .C(InEdges[86]), .D(n134), .Z(
        \temp684[6] ) );
    VMW_AO22 U176 ( .A(OutEdge[5]), .B(n896), .C(InEdges[5]), .D(n94), .Z(
        \temp230[5] ) );
    VMW_AO22 U177 ( .A(\temp230[5] ), .B(n894), .C(InEdges[21]), .D(n102), .Z(
        \temp324[5] ) );
    VMW_AO22 U178 ( .A(\temp324[5] ), .B(n895), .C(InEdges[37]), .D(n110), .Z(
        \temp414[5] ) );
    VMW_AO22 U179 ( .A(\temp414[5] ), .B(n897), .C(InEdges[53]), .D(n118), .Z(
        \temp504[5] ) );
    VMW_AO22 U180 ( .A(\temp504[5] ), .B(n887), .C(InEdges[69]), .D(n126), .Z(
        \temp594[5] ) );
    VMW_AO22 U181 ( .A(\temp594[5] ), .B(n888), .C(InEdges[85]), .D(n134), .Z(
        \temp684[5] ) );
    VMW_AO22 U182 ( .A(OutEdge[4]), .B(n896), .C(InEdges[4]), .D(n94), .Z(
        \temp230[4] ) );
    VMW_AO22 U183 ( .A(\temp230[4] ), .B(n894), .C(InEdges[20]), .D(n102), .Z(
        \temp324[4] ) );
    VMW_AO22 U184 ( .A(\temp324[4] ), .B(n895), .C(InEdges[36]), .D(n110), .Z(
        \temp414[4] ) );
    VMW_AO22 U185 ( .A(\temp414[4] ), .B(n897), .C(InEdges[52]), .D(n118), .Z(
        \temp504[4] ) );
    VMW_AO22 U186 ( .A(\temp504[4] ), .B(n887), .C(InEdges[68]), .D(n126), .Z(
        \temp594[4] ) );
    VMW_AO22 U187 ( .A(\temp594[4] ), .B(n888), .C(InEdges[84]), .D(n134), .Z(
        \temp684[4] ) );
    VMW_AO22 U188 ( .A(OutEdge[3]), .B(n896), .C(InEdges[3]), .D(n94), .Z(
        \temp230[3] ) );
    VMW_AO22 U189 ( .A(\temp230[3] ), .B(n894), .C(InEdges[19]), .D(n102), .Z(
        \temp324[3] ) );
    VMW_AO22 U190 ( .A(\temp324[3] ), .B(n895), .C(InEdges[35]), .D(n110), .Z(
        \temp414[3] ) );
    VMW_AO22 U191 ( .A(\temp414[3] ), .B(n897), .C(InEdges[51]), .D(n118), .Z(
        \temp504[3] ) );
    VMW_AO22 U192 ( .A(\temp504[3] ), .B(n887), .C(InEdges[67]), .D(n126), .Z(
        \temp594[3] ) );
    VMW_AO22 U193 ( .A(\temp594[3] ), .B(n888), .C(InEdges[83]), .D(n134), .Z(
        \temp684[3] ) );
    VMW_AO22 U194 ( .A(OutEdge[2]), .B(n896), .C(InEdges[2]), .D(n94), .Z(
        \temp230[2] ) );
    VMW_AO22 U195 ( .A(\temp230[2] ), .B(n894), .C(InEdges[18]), .D(n102), .Z(
        \temp324[2] ) );
    VMW_AO22 U196 ( .A(\temp324[2] ), .B(n895), .C(InEdges[34]), .D(n110), .Z(
        \temp414[2] ) );
    VMW_AO22 U197 ( .A(\temp414[2] ), .B(n897), .C(InEdges[50]), .D(n118), .Z(
        \temp504[2] ) );
    VMW_AO22 U198 ( .A(\temp504[2] ), .B(n887), .C(InEdges[66]), .D(n126), .Z(
        \temp594[2] ) );
    VMW_AO22 U199 ( .A(\temp594[2] ), .B(n888), .C(InEdges[82]), .D(n134), .Z(
        \temp684[2] ) );
    VMW_AO22 U200 ( .A(OutEdge[1]), .B(n896), .C(InEdges[1]), .D(n94), .Z(
        \temp230[1] ) );
    VMW_AO22 U201 ( .A(\temp230[1] ), .B(n894), .C(InEdges[17]), .D(n102), .Z(
        \temp324[1] ) );
    VMW_AO22 U202 ( .A(\temp324[1] ), .B(n895), .C(InEdges[33]), .D(n110), .Z(
        \temp414[1] ) );
    VMW_AO22 U203 ( .A(\temp414[1] ), .B(n897), .C(InEdges[49]), .D(n118), .Z(
        \temp504[1] ) );
    VMW_AO22 U204 ( .A(\temp504[1] ), .B(n887), .C(InEdges[65]), .D(n126), .Z(
        \temp594[1] ) );
    VMW_AO22 U205 ( .A(\temp594[1] ), .B(n888), .C(InEdges[81]), .D(n134), .Z(
        \temp684[1] ) );
    VMW_AO22 U206 ( .A(OutEdge[15]), .B(n896), .C(InEdges[15]), .D(n94), .Z(
        \temp230[15] ) );
    VMW_AO22 U207 ( .A(\temp230[15] ), .B(n894), .C(InEdges[31]), .D(n102), 
        .Z(\temp324[15] ) );
    VMW_AO22 U208 ( .A(\temp324[15] ), .B(n895), .C(InEdges[47]), .D(n110), 
        .Z(\temp414[15] ) );
    VMW_AO22 U209 ( .A(\temp414[15] ), .B(n897), .C(InEdges[63]), .D(n118), 
        .Z(\temp504[15] ) );
    VMW_AO22 U210 ( .A(\temp504[15] ), .B(n887), .C(InEdges[79]), .D(n126), 
        .Z(\temp594[15] ) );
    VMW_AO22 U211 ( .A(OutEdge[14]), .B(n896), .C(InEdges[14]), .D(n94), .Z(
        \temp230[14] ) );
    VMW_AO22 U212 ( .A(\temp230[14] ), .B(n894), .C(InEdges[30]), .D(n102), 
        .Z(\temp324[14] ) );
    VMW_AO22 U213 ( .A(\temp324[14] ), .B(n895), .C(InEdges[46]), .D(n110), 
        .Z(\temp414[14] ) );
    VMW_AO22 U214 ( .A(\temp414[14] ), .B(n897), .C(InEdges[62]), .D(n118), 
        .Z(\temp504[14] ) );
    VMW_AO22 U215 ( .A(\temp504[14] ), .B(n887), .C(InEdges[78]), .D(n126), 
        .Z(\temp594[14] ) );
    VMW_AO22 U216 ( .A(\temp594[14] ), .B(n888), .C(InEdges[94]), .D(n134), 
        .Z(\temp684[14] ) );
    VMW_AO22 U217 ( .A(OutEdge[13]), .B(n896), .C(InEdges[13]), .D(n94), .Z(
        \temp230[13] ) );
    VMW_AO22 U218 ( .A(\temp230[13] ), .B(n894), .C(InEdges[29]), .D(n102), 
        .Z(\temp324[13] ) );
    VMW_AO22 U219 ( .A(\temp324[13] ), .B(n895), .C(InEdges[45]), .D(n110), 
        .Z(\temp414[13] ) );
    VMW_AO22 U220 ( .A(\temp414[13] ), .B(n897), .C(InEdges[61]), .D(n118), 
        .Z(\temp504[13] ) );
    VMW_AO22 U221 ( .A(\temp504[13] ), .B(n887), .C(InEdges[77]), .D(n126), 
        .Z(\temp594[13] ) );
    VMW_AO22 U222 ( .A(\temp594[13] ), .B(n888), .C(InEdges[93]), .D(n134), 
        .Z(\temp684[13] ) );
    VMW_AO22 U223 ( .A(OutEdge[12]), .B(n896), .C(InEdges[12]), .D(n94), .Z(
        \temp230[12] ) );
    VMW_AO22 U224 ( .A(\temp230[12] ), .B(n894), .C(InEdges[28]), .D(n102), 
        .Z(\temp324[12] ) );
    VMW_AO22 U225 ( .A(\temp324[12] ), .B(n895), .C(InEdges[44]), .D(n110), 
        .Z(\temp414[12] ) );
    VMW_AO22 U226 ( .A(\temp414[12] ), .B(n897), .C(InEdges[60]), .D(n118), 
        .Z(\temp504[12] ) );
    VMW_AO22 U227 ( .A(\temp504[12] ), .B(n887), .C(InEdges[76]), .D(n126), 
        .Z(\temp594[12] ) );
    VMW_AO22 U228 ( .A(\temp594[12] ), .B(n888), .C(InEdges[92]), .D(n134), 
        .Z(\temp684[12] ) );
    VMW_AO22 U229 ( .A(OutEdge[11]), .B(n896), .C(InEdges[11]), .D(n94), .Z(
        \temp230[11] ) );
    VMW_AO22 U230 ( .A(\temp230[11] ), .B(n894), .C(InEdges[27]), .D(n102), 
        .Z(\temp324[11] ) );
    VMW_AO22 U231 ( .A(\temp324[11] ), .B(n895), .C(InEdges[43]), .D(n110), 
        .Z(\temp414[11] ) );
    VMW_AO22 U232 ( .A(\temp414[11] ), .B(n897), .C(InEdges[59]), .D(n118), 
        .Z(\temp504[11] ) );
    VMW_AO22 U233 ( .A(\temp504[11] ), .B(n887), .C(InEdges[75]), .D(n126), 
        .Z(\temp594[11] ) );
    VMW_AO22 U234 ( .A(\temp594[11] ), .B(n888), .C(InEdges[91]), .D(n134), 
        .Z(\temp684[11] ) );
    VMW_AO22 U235 ( .A(OutEdge[10]), .B(n896), .C(InEdges[10]), .D(n94), .Z(
        \temp230[10] ) );
    VMW_AO22 U236 ( .A(\temp230[10] ), .B(n894), .C(InEdges[26]), .D(n102), 
        .Z(\temp324[10] ) );
    VMW_AO22 U237 ( .A(\temp324[10] ), .B(n895), .C(InEdges[42]), .D(n110), 
        .Z(\temp414[10] ) );
    VMW_AO22 U238 ( .A(\temp414[10] ), .B(n897), .C(InEdges[58]), .D(n118), 
        .Z(\temp504[10] ) );
    VMW_AO22 U239 ( .A(\temp504[10] ), .B(n887), .C(InEdges[74]), .D(n126), 
        .Z(\temp594[10] ) );
    VMW_AO22 U240 ( .A(\temp594[10] ), .B(n888), .C(InEdges[90]), .D(n134), 
        .Z(\temp684[10] ) );
    VMW_AO22 U241 ( .A(OutEdge[0]), .B(n896), .C(InEdges[0]), .D(n94), .Z(
        \temp230[0] ) );
    VMW_AO22 U242 ( .A(\temp230[0] ), .B(n894), .C(InEdges[16]), .D(n102), .Z(
        \temp324[0] ) );
    VMW_AO22 U243 ( .A(\temp324[0] ), .B(n895), .C(InEdges[32]), .D(n110), .Z(
        \temp414[0] ) );
    VMW_AO22 U244 ( .A(\temp414[0] ), .B(n897), .C(InEdges[48]), .D(n118), .Z(
        \temp504[0] ) );
    VMW_AO22 U245 ( .A(\temp504[0] ), .B(n887), .C(InEdges[64]), .D(n126), .Z(
        \temp594[0] ) );
    VMW_AO22 U246 ( .A(\temp594[0] ), .B(n888), .C(InEdges[80]), .D(n134), .Z(
        \temp684[0] ) );
    VMW_MUX2I U247 ( .A(\temp684[9] ), .B(InEdges[105]), .S(n142), .Z(n875) );
    VMW_MUX2I U248 ( .A(\temp684[8] ), .B(InEdges[104]), .S(n142), .Z(n876) );
    VMW_MUX2I U249 ( .A(\temp684[7] ), .B(InEdges[103]), .S(n142), .Z(n877) );
    VMW_MUX2I U250 ( .A(\temp684[6] ), .B(InEdges[102]), .S(n142), .Z(n878) );
    VMW_MUX2I U251 ( .A(\temp684[5] ), .B(InEdges[101]), .S(n142), .Z(n879) );
    VMW_MUX2I U252 ( .A(\temp684[4] ), .B(InEdges[100]), .S(n142), .Z(n880) );
    VMW_MUX2I U253 ( .A(\temp684[3] ), .B(InEdges[99]), .S(n142), .Z(n881) );
    VMW_MUX2I U254 ( .A(\temp684[2] ), .B(InEdges[98]), .S(n142), .Z(n882) );
    VMW_MUX2I U255 ( .A(\temp684[1] ), .B(InEdges[97]), .S(n142), .Z(n883) );
    VMW_MUX2I U256 ( .A(\temp684[14] ), .B(InEdges[110]), .S(n142), .Z(n869)
         );
    VMW_MUX2I U257 ( .A(\temp684[13] ), .B(InEdges[109]), .S(n142), .Z(n871)
         );
    VMW_MUX2I U258 ( .A(\temp684[12] ), .B(InEdges[108]), .S(n142), .Z(n872)
         );
    VMW_MUX2I U259 ( .A(\temp684[11] ), .B(InEdges[107]), .S(n142), .Z(n873)
         );
    VMW_MUX2I U260 ( .A(\temp684[10] ), .B(InEdges[106]), .S(n142), .Z(n874)
         );
    VMW_MUX2I U261 ( .A(\temp684[0] ), .B(InEdges[96]), .S(n142), .Z(n884) );
    VMW_INV U262 ( .A(n94), .Z(n896) );
    VMW_INV U263 ( .A(n102), .Z(n894) );
    VMW_INV U264 ( .A(n898), .Z(n911) );
    VMW_INV U265 ( .A(n899), .Z(n913) );
    VMW_BUFIZ U266 ( .A(\path[3] ), .E(n909), .Z(\PathData[3] ) );
    VMW_BUFIZ U267 ( .A(\path[1] ), .E(n909), .Z(\PathData[1] ) );
    VMW_BUFIZ U268 ( .A(\path[0] ), .E(n909), .Z(\PathData[0] ) );
    VMW_BUFIZ U269 ( .A(\path[2] ), .E(n909), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n910), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n911), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n912), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n913), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge156[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge156[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge156[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge156[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge156[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge156[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge156[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge156[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge156[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge156[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge156[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge156[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge156[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge156[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge156[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge156[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 lte_55_5 ( .A({\temp594[15] , 
        \temp594[14] , \temp594[13] , \temp594[12] , \temp594[11] , 
        \temp594[10] , \temp594[9] , \temp594[8] , \temp594[7] , \temp594[6] , 
        \temp594[5] , \temp594[4] , \temp594[3] , \temp594[2] , \temp594[1] , 
        \temp594[0] }), .B(InEdges[95:80]), .LEQ(n920), .TC(n920), .GE_GT(n134
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 lte_55_3 ( .A({\temp414[15] , 
        \temp414[14] , \temp414[13] , \temp414[12] , \temp414[11] , 
        \temp414[10] , \temp414[9] , \temp414[8] , \temp414[7] , \temp414[6] , 
        \temp414[5] , \temp414[4] , \temp414[3] , \temp414[2] , \temp414[1] , 
        \temp414[0] }), .B(InEdges[63:48]), .LEQ(n919), .TC(n919), .GE_GT(n118
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 lte_55_4 ( .A({\temp504[15] , 
        \temp504[14] , \temp504[13] , \temp504[12] , \temp504[11] , 
        \temp504[10] , \temp504[9] , \temp504[8] , \temp504[7] , \temp504[6] , 
        \temp504[5] , \temp504[4] , \temp504[3] , \temp504[2] , \temp504[1] , 
        \temp504[0] }), .B(InEdges[79:64]), .LEQ(n918), .TC(n918), .GE_GT(n126
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n917), .TC(n917), .GE_GT(n94) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 lte_55_6 ( .A({\temp684[15] , 
        \temp684[14] , \temp684[13] , \temp684[12] , \temp684[11] , 
        \temp684[10] , \temp684[9] , \temp684[8] , \temp684[7] , \temp684[6] , 
        \temp684[5] , \temp684[4] , \temp684[3] , \temp684[2] , \temp684[1] , 
        \temp684[0] }), .B(InEdges[111:96]), .LEQ(n916), .TC(n916), .GE_GT(
        n142) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp324[15] , 
        \temp324[14] , \temp324[13] , \temp324[12] , \temp324[11] , 
        \temp324[10] , \temp324[9] , \temp324[8] , \temp324[7] , \temp324[6] , 
        \temp324[5] , \temp324[4] , \temp324[3] , \temp324[2] , \temp324[1] , 
        \temp324[0] }), .B(InEdges[47:32]), .LEQ(n915), .TC(n915), .GE_GT(n110
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp230[15] , 
        \temp230[14] , \temp230[13] , \temp230[12] , \temp230[11] , 
        \temp230[10] , \temp230[9] , \temp230[8] , \temp230[7] , \temp230[6] , 
        \temp230[5] , \temp230[4] , \temp230[3] , \temp230[2] , \temp230[1] , 
        \temp230[0] }), .B(InEdges[31:16]), .LEQ(n914), .TC(n914), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_7 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, 
        n107, n108, n109, n110, n111, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n95), .B(B[10]), .Z(n94) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n95), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n102), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n94), .Z(n103) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n102), .C(n106), .D(n103), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n101), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n110), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n102) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n95) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n121, n122, n123, n124, n125, n126, n127, 
        n129, n130, n131, n132, n133, n134, n135, n137, n138, n139, n140, n141, 
        n142, n143, n145, n146, n147, n148, n149, n150, n151, n153, n154, n155, 
        n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
        n168, n169;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n118), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n126), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n134), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n154), .C(n148), .D(n142), .Z(n153) );
    VMW_NAND2 U22 ( .A(n154), .B(A[9]), .Z(n155) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n155), .D(n153), .Z(n156) );
    VMW_NAND2 U24 ( .A(n158), .B(B[12]), .Z(n157) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n160), .C(n156), .D(n150), .Z(n159) );
    VMW_NAND2 U26 ( .A(n160), .B(A[11]), .Z(n161) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n158), .C(n161), .D(n159), .Z(n162) );
    VMW_NAND2 U28 ( .A(n164), .B(B[14]), .Z(n163) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n166), .C(n162), .D(n157), .Z(n165) );
    VMW_NAND2 U30 ( .A(n166), .B(A[13]), .Z(n167) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n164), .C(n167), .D(n165), .Z(n168) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n169), .C(n168), .D(n163), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n158) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n154) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n164) );
    VMW_INV U43 ( .A(B[11]), .Z(n160) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n169) );
    VMW_INV U48 ( .A(B[13]), .Z(n166) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
        n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
        n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
        n217, n218;
    VMW_OAI21 U3 ( .A(B[15]), .B(n170), .C(n171), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n173), .B(B[2]), .Z(n172) );
    VMW_AO22 U5 ( .A(n175), .B(B[0]), .C(n176), .D(B[1]), .Z(n174) );
    VMW_OR2 U6 ( .A(B[2]), .B(n173), .Z(n177) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n176), .C(n177), .D(n174), .Z(n178) );
    VMW_NAND2 U8 ( .A(n180), .B(B[4]), .Z(n179) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n182), .C(n178), .D(n172), .Z(n181) );
    VMW_OR2 U10 ( .A(B[4]), .B(n180), .Z(n183) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n185), .C(n183), .D(n181), .Z(n184) );
    VMW_NAND2 U12 ( .A(n187), .B(B[6]), .Z(n186) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n189), .C(n184), .D(n179), .Z(n188) );
    VMW_OR2 U14 ( .A(B[6]), .B(n187), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n192), .C(n190), .D(n188), .Z(n191) );
    VMW_NAND2 U16 ( .A(n194), .B(B[8]), .Z(n193) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n196), .C(n191), .D(n186), .Z(n195) );
    VMW_OR2 U18 ( .A(B[8]), .B(n194), .Z(n197) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_NAND2 U20 ( .A(n201), .B(B[10]), .Z(n200) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_NAND2 U22 ( .A(n203), .B(A[9]), .Z(n204) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n201), .C(n204), .D(n202), .Z(n205) );
    VMW_NAND2 U24 ( .A(n207), .B(B[12]), .Z(n206) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n209), .C(n205), .D(n200), .Z(n208) );
    VMW_NAND2 U26 ( .A(n209), .B(A[11]), .Z(n210) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n207), .C(n210), .D(n208), .Z(n211) );
    VMW_NAND2 U28 ( .A(n213), .B(B[14]), .Z(n212) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n215), .C(n211), .D(n206), .Z(n214) );
    VMW_NAND2 U30 ( .A(n215), .B(A[13]), .Z(n216) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n213), .C(n216), .D(n214), .Z(n217) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n218), .C(n217), .D(n212), .Z(n171) );
    VMW_INV U33 ( .A(A[12]), .Z(n207) );
    VMW_INV U34 ( .A(B[7]), .Z(n196) );
    VMW_INV U35 ( .A(A[7]), .Z(n199) );
    VMW_INV U36 ( .A(A[3]), .Z(n185) );
    VMW_INV U37 ( .A(B[3]), .Z(n182) );
    VMW_INV U38 ( .A(A[10]), .Z(n201) );
    VMW_INV U39 ( .A(B[9]), .Z(n203) );
    VMW_INV U40 ( .A(A[4]), .Z(n180) );
    VMW_INV U41 ( .A(A[8]), .Z(n194) );
    VMW_INV U42 ( .A(A[14]), .Z(n213) );
    VMW_INV U43 ( .A(B[11]), .Z(n209) );
    VMW_INV U44 ( .A(A[5]), .Z(n192) );
    VMW_INV U45 ( .A(B[5]), .Z(n189) );
    VMW_INV U46 ( .A(A[1]), .Z(n176) );
    VMW_INV U47 ( .A(B[15]), .Z(n218) );
    VMW_INV U48 ( .A(B[13]), .Z(n215) );
    VMW_INV U49 ( .A(A[6]), .Z(n187) );
    VMW_INV U50 ( .A(A[2]), .Z(n173) );
    VMW_INV U51 ( .A(A[0]), .Z(n175) );
    VMW_INV U52 ( .A(A[15]), .Z(n170) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267;
    VMW_OAI21 U3 ( .A(B[15]), .B(n219), .C(n220), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n222), .B(B[2]), .Z(n221) );
    VMW_AO22 U5 ( .A(n224), .B(B[0]), .C(n225), .D(B[1]), .Z(n223) );
    VMW_OR2 U6 ( .A(B[2]), .B(n222), .Z(n226) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n225), .C(n226), .D(n223), .Z(n227) );
    VMW_NAND2 U8 ( .A(n229), .B(B[4]), .Z(n228) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n231), .C(n227), .D(n221), .Z(n230) );
    VMW_OR2 U10 ( .A(B[4]), .B(n229), .Z(n232) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n234), .C(n232), .D(n230), .Z(n233) );
    VMW_NAND2 U12 ( .A(n236), .B(B[6]), .Z(n235) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n238), .C(n233), .D(n228), .Z(n237) );
    VMW_OR2 U14 ( .A(B[6]), .B(n236), .Z(n239) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n241), .C(n239), .D(n237), .Z(n240) );
    VMW_NAND2 U16 ( .A(n243), .B(B[8]), .Z(n242) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n245), .C(n240), .D(n235), .Z(n244) );
    VMW_OR2 U18 ( .A(B[8]), .B(n243), .Z(n246) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n248), .C(n246), .D(n244), .Z(n247) );
    VMW_NAND2 U20 ( .A(n250), .B(B[10]), .Z(n249) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n252), .C(n247), .D(n242), .Z(n251) );
    VMW_NAND2 U22 ( .A(n252), .B(A[9]), .Z(n253) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n250), .C(n253), .D(n251), .Z(n254) );
    VMW_NAND2 U24 ( .A(n256), .B(B[12]), .Z(n255) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n258), .C(n254), .D(n249), .Z(n257) );
    VMW_NAND2 U26 ( .A(n258), .B(A[11]), .Z(n259) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n256), .C(n259), .D(n257), .Z(n260) );
    VMW_NAND2 U28 ( .A(n262), .B(B[14]), .Z(n261) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n264), .C(n260), .D(n255), .Z(n263) );
    VMW_NAND2 U30 ( .A(n264), .B(A[13]), .Z(n265) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n262), .C(n265), .D(n263), .Z(n266) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n267), .C(n266), .D(n261), .Z(n220) );
    VMW_INV U33 ( .A(A[12]), .Z(n256) );
    VMW_INV U34 ( .A(B[7]), .Z(n245) );
    VMW_INV U35 ( .A(A[7]), .Z(n248) );
    VMW_INV U36 ( .A(A[3]), .Z(n234) );
    VMW_INV U37 ( .A(B[3]), .Z(n231) );
    VMW_INV U38 ( .A(A[10]), .Z(n250) );
    VMW_INV U39 ( .A(B[9]), .Z(n252) );
    VMW_INV U40 ( .A(A[4]), .Z(n229) );
    VMW_INV U41 ( .A(A[8]), .Z(n243) );
    VMW_INV U42 ( .A(A[14]), .Z(n262) );
    VMW_INV U43 ( .A(B[11]), .Z(n258) );
    VMW_INV U44 ( .A(A[5]), .Z(n241) );
    VMW_INV U45 ( .A(B[5]), .Z(n238) );
    VMW_INV U46 ( .A(A[1]), .Z(n225) );
    VMW_INV U47 ( .A(B[15]), .Z(n267) );
    VMW_INV U48 ( .A(B[13]), .Z(n264) );
    VMW_INV U49 ( .A(A[6]), .Z(n236) );
    VMW_INV U50 ( .A(A[2]), .Z(n222) );
    VMW_INV U51 ( .A(A[0]), .Z(n224) );
    VMW_INV U52 ( .A(A[15]), .Z(n219) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
        n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316;
    VMW_OAI21 U3 ( .A(B[15]), .B(n268), .C(n269), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n271), .B(B[2]), .Z(n270) );
    VMW_AO22 U5 ( .A(n273), .B(B[0]), .C(n274), .D(B[1]), .Z(n272) );
    VMW_OR2 U6 ( .A(B[2]), .B(n271), .Z(n275) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n274), .C(n275), .D(n272), .Z(n276) );
    VMW_NAND2 U8 ( .A(n278), .B(B[4]), .Z(n277) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n280), .C(n276), .D(n270), .Z(n279) );
    VMW_OR2 U10 ( .A(B[4]), .B(n278), .Z(n281) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n283), .C(n281), .D(n279), .Z(n282) );
    VMW_NAND2 U12 ( .A(n285), .B(B[6]), .Z(n284) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n287), .C(n282), .D(n277), .Z(n286) );
    VMW_OR2 U14 ( .A(B[6]), .B(n285), .Z(n288) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n290), .C(n288), .D(n286), .Z(n289) );
    VMW_NAND2 U16 ( .A(n292), .B(B[8]), .Z(n291) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n294), .C(n289), .D(n284), .Z(n293) );
    VMW_OR2 U18 ( .A(B[8]), .B(n292), .Z(n295) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n297), .C(n295), .D(n293), .Z(n296) );
    VMW_NAND2 U20 ( .A(n299), .B(B[10]), .Z(n298) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n301), .C(n296), .D(n291), .Z(n300) );
    VMW_NAND2 U22 ( .A(n301), .B(A[9]), .Z(n302) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n299), .C(n302), .D(n300), .Z(n303) );
    VMW_NAND2 U24 ( .A(n305), .B(B[12]), .Z(n304) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n307), .C(n303), .D(n298), .Z(n306) );
    VMW_NAND2 U26 ( .A(n307), .B(A[11]), .Z(n308) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n305), .C(n308), .D(n306), .Z(n309) );
    VMW_NAND2 U28 ( .A(n311), .B(B[14]), .Z(n310) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n313), .C(n309), .D(n304), .Z(n312) );
    VMW_NAND2 U30 ( .A(n313), .B(A[13]), .Z(n314) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n311), .C(n314), .D(n312), .Z(n315) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n316), .C(n315), .D(n310), .Z(n269) );
    VMW_INV U33 ( .A(A[12]), .Z(n305) );
    VMW_INV U34 ( .A(B[7]), .Z(n294) );
    VMW_INV U35 ( .A(A[7]), .Z(n297) );
    VMW_INV U36 ( .A(A[3]), .Z(n283) );
    VMW_INV U37 ( .A(B[3]), .Z(n280) );
    VMW_INV U38 ( .A(A[10]), .Z(n299) );
    VMW_INV U39 ( .A(B[9]), .Z(n301) );
    VMW_INV U40 ( .A(A[4]), .Z(n278) );
    VMW_INV U41 ( .A(A[8]), .Z(n292) );
    VMW_INV U42 ( .A(A[14]), .Z(n311) );
    VMW_INV U43 ( .A(B[11]), .Z(n307) );
    VMW_INV U44 ( .A(A[5]), .Z(n290) );
    VMW_INV U45 ( .A(B[5]), .Z(n287) );
    VMW_INV U46 ( .A(A[1]), .Z(n274) );
    VMW_INV U47 ( .A(B[15]), .Z(n316) );
    VMW_INV U48 ( .A(B[13]), .Z(n313) );
    VMW_INV U49 ( .A(A[6]), .Z(n285) );
    VMW_INV U50 ( .A(A[2]), .Z(n271) );
    VMW_INV U51 ( .A(A[0]), .Z(n273) );
    VMW_INV U52 ( .A(A[15]), .Z(n268) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
        n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
        n364, n365;
    VMW_OAI21 U3 ( .A(B[15]), .B(n317), .C(n318), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n320), .B(B[2]), .Z(n319) );
    VMW_AO22 U5 ( .A(n322), .B(B[0]), .C(n323), .D(B[1]), .Z(n321) );
    VMW_OR2 U6 ( .A(B[2]), .B(n320), .Z(n324) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n323), .C(n324), .D(n321), .Z(n325) );
    VMW_NAND2 U8 ( .A(n327), .B(B[4]), .Z(n326) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n329), .C(n325), .D(n319), .Z(n328) );
    VMW_OR2 U10 ( .A(B[4]), .B(n327), .Z(n330) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n332), .C(n330), .D(n328), .Z(n331) );
    VMW_NAND2 U12 ( .A(n334), .B(B[6]), .Z(n333) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n336), .C(n331), .D(n326), .Z(n335) );
    VMW_OR2 U14 ( .A(B[6]), .B(n334), .Z(n337) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n339), .C(n337), .D(n335), .Z(n338) );
    VMW_NAND2 U16 ( .A(n341), .B(B[8]), .Z(n340) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n343), .C(n338), .D(n333), .Z(n342) );
    VMW_OR2 U18 ( .A(B[8]), .B(n341), .Z(n344) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n346), .C(n344), .D(n342), .Z(n345) );
    VMW_NAND2 U20 ( .A(n348), .B(B[10]), .Z(n347) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n350), .C(n345), .D(n340), .Z(n349) );
    VMW_NAND2 U22 ( .A(n350), .B(A[9]), .Z(n351) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n348), .C(n351), .D(n349), .Z(n352) );
    VMW_NAND2 U24 ( .A(n354), .B(B[12]), .Z(n353) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n356), .C(n352), .D(n347), .Z(n355) );
    VMW_NAND2 U26 ( .A(n356), .B(A[11]), .Z(n357) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n354), .C(n357), .D(n355), .Z(n358) );
    VMW_NAND2 U28 ( .A(n360), .B(B[14]), .Z(n359) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n362), .C(n358), .D(n353), .Z(n361) );
    VMW_NAND2 U30 ( .A(n362), .B(A[13]), .Z(n363) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n360), .C(n363), .D(n361), .Z(n364) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n365), .C(n364), .D(n359), .Z(n318) );
    VMW_INV U33 ( .A(A[12]), .Z(n354) );
    VMW_INV U34 ( .A(B[7]), .Z(n343) );
    VMW_INV U35 ( .A(A[7]), .Z(n346) );
    VMW_INV U36 ( .A(A[3]), .Z(n332) );
    VMW_INV U37 ( .A(B[3]), .Z(n329) );
    VMW_INV U38 ( .A(A[10]), .Z(n348) );
    VMW_INV U39 ( .A(B[9]), .Z(n350) );
    VMW_INV U40 ( .A(A[4]), .Z(n327) );
    VMW_INV U41 ( .A(A[8]), .Z(n341) );
    VMW_INV U42 ( .A(A[14]), .Z(n360) );
    VMW_INV U43 ( .A(B[11]), .Z(n356) );
    VMW_INV U44 ( .A(A[5]), .Z(n339) );
    VMW_INV U45 ( .A(B[5]), .Z(n336) );
    VMW_INV U46 ( .A(A[1]), .Z(n323) );
    VMW_INV U47 ( .A(B[15]), .Z(n365) );
    VMW_INV U48 ( .A(B[13]), .Z(n362) );
    VMW_INV U49 ( .A(A[6]), .Z(n334) );
    VMW_INV U50 ( .A(A[2]), .Z(n320) );
    VMW_INV U51 ( .A(A[0]), .Z(n322) );
    VMW_INV U52 ( .A(A[15]), .Z(n317) );
endmodule


module NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
        n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
        n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
        n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
        n413, n414;
    VMW_OAI21 U3 ( .A(B[15]), .B(n366), .C(n367), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n369), .B(B[2]), .Z(n368) );
    VMW_AO22 U5 ( .A(n371), .B(B[0]), .C(n372), .D(B[1]), .Z(n370) );
    VMW_OR2 U6 ( .A(B[2]), .B(n369), .Z(n373) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n372), .C(n373), .D(n370), .Z(n374) );
    VMW_NAND2 U8 ( .A(n376), .B(B[4]), .Z(n375) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n378), .C(n374), .D(n368), .Z(n377) );
    VMW_OR2 U10 ( .A(B[4]), .B(n376), .Z(n379) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n381), .C(n379), .D(n377), .Z(n380) );
    VMW_NAND2 U12 ( .A(n383), .B(B[6]), .Z(n382) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n385), .C(n380), .D(n375), .Z(n384) );
    VMW_OR2 U14 ( .A(B[6]), .B(n383), .Z(n386) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n388), .C(n386), .D(n384), .Z(n387) );
    VMW_NAND2 U16 ( .A(n390), .B(B[8]), .Z(n389) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n392), .C(n387), .D(n382), .Z(n391) );
    VMW_OR2 U18 ( .A(B[8]), .B(n390), .Z(n393) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n395), .C(n393), .D(n391), .Z(n394) );
    VMW_NAND2 U20 ( .A(n397), .B(B[10]), .Z(n396) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n399), .C(n394), .D(n389), .Z(n398) );
    VMW_NAND2 U22 ( .A(n399), .B(A[9]), .Z(n400) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n397), .C(n400), .D(n398), .Z(n401) );
    VMW_NAND2 U24 ( .A(n403), .B(B[12]), .Z(n402) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n405), .C(n401), .D(n396), .Z(n404) );
    VMW_NAND2 U26 ( .A(n405), .B(A[11]), .Z(n406) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n403), .C(n406), .D(n404), .Z(n407) );
    VMW_NAND2 U28 ( .A(n409), .B(B[14]), .Z(n408) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n411), .C(n407), .D(n402), .Z(n410) );
    VMW_NAND2 U30 ( .A(n411), .B(A[13]), .Z(n412) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n409), .C(n412), .D(n410), .Z(n413) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n414), .C(n413), .D(n408), .Z(n367) );
    VMW_INV U33 ( .A(A[12]), .Z(n403) );
    VMW_INV U34 ( .A(B[7]), .Z(n392) );
    VMW_INV U35 ( .A(A[7]), .Z(n395) );
    VMW_INV U36 ( .A(A[3]), .Z(n381) );
    VMW_INV U37 ( .A(B[3]), .Z(n378) );
    VMW_INV U38 ( .A(A[10]), .Z(n397) );
    VMW_INV U39 ( .A(B[9]), .Z(n399) );
    VMW_INV U40 ( .A(A[4]), .Z(n376) );
    VMW_INV U41 ( .A(A[8]), .Z(n390) );
    VMW_INV U42 ( .A(A[14]), .Z(n409) );
    VMW_INV U43 ( .A(B[11]), .Z(n405) );
    VMW_INV U44 ( .A(A[5]), .Z(n388) );
    VMW_INV U45 ( .A(B[5]), .Z(n385) );
    VMW_INV U46 ( .A(A[1]), .Z(n372) );
    VMW_INV U47 ( .A(B[15]), .Z(n414) );
    VMW_INV U48 ( .A(B[13]), .Z(n411) );
    VMW_INV U49 ( .A(A[6]), .Z(n383) );
    VMW_INV U50 ( .A(A[2]), .Z(n369) );
    VMW_INV U51 ( .A(A[0]), .Z(n371) );
    VMW_INV U52 ( .A(A[15]), .Z(n366) );
endmodule


module NodeAux_INDEGREE8_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [5:0] Nid;
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire \temp240[2] , \temp334[3] , \temp424[2] , \temp604[10] , 
        \temp424[14] , n152, \temp694[10] , \temp604[3] , \temp784[12] , n112, 
        \temp424[10] , \temp604[14] , \temp424[6] , \temp240[6] , \temp334[7] , 
        \path[2] , \temp604[7] , \temp694[14] , \path[0] , \temp604[5] , 
        \temp784[14] , \temp424[4] , \temp240[4] , \temp334[5] , \temp424[12] , 
        \temp334[8] , n120, \temp784[10] , \temp240[9] , \temp424[9] , 
        \temp694[12] , \temp604[1] , \temp604[8] , \temp604[12] , \temp334[1] , 
        \temp424[0] , \temp240[0] , \temp240[14] , \temp514[3] , \temp334[10] , 
        \temp694[2] , \temp784[7] , \temp514[13] , \OutEdge166[13] , 
        \OutEdge166[3] , n128, \temp694[6] , \temp784[3] , \temp334[14] , 
        \temp514[7] , \OutEdge166[7] , \temp240[10] , \temp784[8] , 
        \temp514[15] , \OutEdge166[15] , \OutEdge166[5] , n96, \temp514[5] , 
        \temp240[12] , \temp784[1] , \temp694[4] , \temp514[8] , 
        \OutEdge166[11] , \OutEdge166[1] , \temp694[9] , \temp514[11] , 
        \temp334[12] , \temp694[0] , \temp784[5] , \temp514[1] , 
        \OutEdge166[8] , \temp514[9] , \OutEdge166[10] , \OutEdge166[0] , 
        \temp694[8] , \temp514[10] , \temp694[1] , \temp334[13] , \temp514[0] , 
        \temp784[4] , \OutEdge166[9] , \temp514[14] , \temp784[9] , n136, 
        \OutEdge166[14] , \OutEdge166[4] , \temp240[13] , \temp514[4] , 
        \temp784[0] , \temp694[5] , \temp784[2] , \temp334[15] , \temp694[7] , 
        \temp240[11] , \temp514[6] , n144, \OutEdge166[6] , \temp514[2] , n104, 
        \temp240[15] , \temp694[3] , \temp334[11] , \temp784[6] , 
        \temp514[12] , \OutEdge166[12] , \OutEdge166[2] , \temp334[9] , 
        \temp240[8] , \temp424[8] , \temp784[11] , \temp694[13] , \temp604[0] , 
        \temp604[13] , \temp604[9] , \temp334[0] , \temp240[1] , \temp424[1] , 
        \path[1] , \temp604[4] , \temp784[15] , \temp424[5] , \temp240[5] , 
        \temp334[4] , \temp424[13] , \temp424[11] , \temp604[15] , 
        \temp424[7] , \temp240[7] , \temp334[6] , \path[3] , \temp694[15] , 
        \temp604[6] , \temp334[2] , \temp424[3] , \temp240[3] , \temp604[11] , 
        \temp424[15] , \temp604[2] , \temp694[11] , \temp784[13] , n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
        n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
        n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
        n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
        n1024;
    tri \PathData[1] , \PathData[3] , \PathData[2] , \PathData[0] ;
    assign PathData[3] = \PathData[3] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U109 ( .Z(n1019) );
    VMW_PULLDOWN U110 ( .Z(n1018) );
    VMW_PULLDOWN U111 ( .Z(n1021) );
    VMW_PULLDOWN U112 ( .Z(n1022) );
    VMW_PULLDOWN U113 ( .Z(n1017) );
    VMW_PULLDOWN U114 ( .Z(n1024) );
    VMW_PULLDOWN U115 ( .Z(n1020) );
    VMW_PULLDOWN U116 ( .Z(n1023) );
    VMW_NOR2 U117 ( .A(Start), .B(n967), .Z(\OutEdge166[15] ) );
    VMW_NAND2 U118 ( .A(n968), .B(n969), .Z(\OutEdge166[14] ) );
    VMW_NAND2 U119 ( .A(n970), .B(n969), .Z(\OutEdge166[13] ) );
    VMW_NAND2 U120 ( .A(n971), .B(n969), .Z(\OutEdge166[12] ) );
    VMW_NAND2 U121 ( .A(n972), .B(n969), .Z(\OutEdge166[11] ) );
    VMW_NAND2 U122 ( .A(n973), .B(n969), .Z(\OutEdge166[10] ) );
    VMW_NAND2 U123 ( .A(n974), .B(n969), .Z(\OutEdge166[9] ) );
    VMW_NAND2 U124 ( .A(n975), .B(n969), .Z(\OutEdge166[8] ) );
    VMW_NAND2 U125 ( .A(n976), .B(n969), .Z(\OutEdge166[7] ) );
    VMW_NAND2 U126 ( .A(n977), .B(n969), .Z(\OutEdge166[6] ) );
    VMW_NAND2 U127 ( .A(n978), .B(n969), .Z(\OutEdge166[5] ) );
    VMW_NAND2 U128 ( .A(n979), .B(n969), .Z(\OutEdge166[4] ) );
    VMW_NAND2 U129 ( .A(n980), .B(n969), .Z(\OutEdge166[3] ) );
    VMW_NAND2 U130 ( .A(n981), .B(n969), .Z(\OutEdge166[2] ) );
    VMW_NAND2 U131 ( .A(n982), .B(n969), .Z(\OutEdge166[1] ) );
    VMW_NAND2 U132 ( .A(n983), .B(n969), .Z(\OutEdge166[0] ) );
    VMW_AO21 U133 ( .A(n984), .B(n985), .C(n986), .Z(n1016) );
    VMW_AO22 U134 ( .A(\path[3] ), .B(Start), .C(n987), .D(n988), .Z(n1015) );
    VMW_OR4 U135 ( .A(n136), .B(n128), .C(n987), .D(n990), .Z(n989) );
    VMW_OR2 U136 ( .A(n152), .B(n992), .Z(n991) );
    VMW_AO22 U137 ( .A(\temp694[15] ), .B(n993), .C(InEdges[111]), .D(n144), 
        .Z(\temp784[15] ) );
    VMW_OR2 U138 ( .A(n152), .B(n144), .Z(n990) );
    VMW_AND3 U139 ( .A(n969), .B(n994), .C(n995), .Z(n984) );
    VMW_AND4 U140 ( .A(n996), .B(n997), .C(n998), .D(n999), .Z(n987) );
    VMW_INV U141 ( .A(Start), .Z(n969) );
    VMW_OAI22 U142 ( .A(n989), .B(Start), .C(\path[2] ), .D(n969), .Z(n1000)
         );
    VMW_AO22 U143 ( .A(\path[1] ), .B(Start), .C(n990), .D(n969), .Z(n986) );
    VMW_OAI22 U144 ( .A(n991), .B(Start), .C(\path[0] ), .D(n969), .Z(n1001)
         );
    VMW_MUX2I U145 ( .A(\temp784[15] ), .B(InEdges[127]), .S(n152), .Z(n967)
         );
    VMW_NOR2 U146 ( .A(n990), .B(n1002), .Z(n988) );
    VMW_AND3 U147 ( .A(n1004), .B(n1005), .C(n1006), .Z(n1003) );
    VMW_INV U148 ( .A(n120), .Z(n999) );
    VMW_INV U149 ( .A(n136), .Z(n994) );
    VMW_INV U150 ( .A(n112), .Z(n997) );
    VMW_OAI211 U151 ( .A(n96), .B(n104), .C(n997), .D(n999), .Z(n985) );
    VMW_AO21 U152 ( .A(n996), .B(n96), .C(n112), .Z(n1007) );
    VMW_AO21 U153 ( .A(n999), .B(n1007), .C(n128), .Z(n1008) );
    VMW_AOI21 U154 ( .A(n994), .B(n1008), .C(n144), .Z(n992) );
    VMW_AND4 U155 ( .A(n1009), .B(n1010), .C(n1011), .D(n1003), .Z(n1012) );
    VMW_XNOR2 U156 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n1005) );
    VMW_XNOR2 U157 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n1004) );
    VMW_XNOR2 U158 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n1006) );
    VMW_XNOR2 U159 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n1010) );
    VMW_XNOR2 U160 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n1009) );
    VMW_XNOR2 U161 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n1011) );
    VMW_AO22 U162 ( .A(InEdges[9]), .B(n96), .C(OutEdge[9]), .D(n998), .Z(
        \temp240[9] ) );
    VMW_AO22 U163 ( .A(\temp240[9] ), .B(n996), .C(InEdges[25]), .D(n104), .Z(
        \temp334[9] ) );
    VMW_AO22 U164 ( .A(InEdges[41]), .B(n112), .C(\temp334[9] ), .D(n997), .Z(
        \temp424[9] ) );
    VMW_AO22 U165 ( .A(InEdges[57]), .B(n120), .C(\temp424[9] ), .D(n999), .Z(
        \temp514[9] ) );
    VMW_AO22 U166 ( .A(\temp514[9] ), .B(n995), .C(InEdges[73]), .D(n128), .Z(
        \temp604[9] ) );
    VMW_AO22 U167 ( .A(InEdges[89]), .B(n136), .C(\temp604[9] ), .D(n994), .Z(
        \temp694[9] ) );
    VMW_AO22 U168 ( .A(\temp694[9] ), .B(n993), .C(InEdges[105]), .D(n144), 
        .Z(\temp784[9] ) );
    VMW_AO22 U169 ( .A(InEdges[8]), .B(n96), .C(OutEdge[8]), .D(n998), .Z(
        \temp240[8] ) );
    VMW_AO22 U170 ( .A(\temp240[8] ), .B(n996), .C(InEdges[24]), .D(n104), .Z(
        \temp334[8] ) );
    VMW_AO22 U171 ( .A(InEdges[40]), .B(n112), .C(\temp334[8] ), .D(n997), .Z(
        \temp424[8] ) );
    VMW_AO22 U172 ( .A(InEdges[56]), .B(n120), .C(\temp424[8] ), .D(n999), .Z(
        \temp514[8] ) );
    VMW_AO22 U173 ( .A(\temp514[8] ), .B(n995), .C(InEdges[72]), .D(n128), .Z(
        \temp604[8] ) );
    VMW_AO22 U174 ( .A(InEdges[88]), .B(n136), .C(\temp604[8] ), .D(n994), .Z(
        \temp694[8] ) );
    VMW_AO22 U175 ( .A(\temp694[8] ), .B(n993), .C(InEdges[104]), .D(n144), 
        .Z(\temp784[8] ) );
    VMW_AO22 U176 ( .A(InEdges[7]), .B(n96), .C(OutEdge[7]), .D(n998), .Z(
        \temp240[7] ) );
    VMW_AO22 U177 ( .A(\temp240[7] ), .B(n996), .C(InEdges[23]), .D(n104), .Z(
        \temp334[7] ) );
    VMW_AO22 U178 ( .A(InEdges[39]), .B(n112), .C(\temp334[7] ), .D(n997), .Z(
        \temp424[7] ) );
    VMW_AO22 U179 ( .A(InEdges[55]), .B(n120), .C(\temp424[7] ), .D(n999), .Z(
        \temp514[7] ) );
    VMW_AO22 U180 ( .A(\temp514[7] ), .B(n995), .C(InEdges[71]), .D(n128), .Z(
        \temp604[7] ) );
    VMW_AO22 U181 ( .A(InEdges[87]), .B(n136), .C(\temp604[7] ), .D(n994), .Z(
        \temp694[7] ) );
    VMW_AO22 U182 ( .A(\temp694[7] ), .B(n993), .C(InEdges[103]), .D(n144), 
        .Z(\temp784[7] ) );
    VMW_AO22 U183 ( .A(InEdges[6]), .B(n96), .C(OutEdge[6]), .D(n998), .Z(
        \temp240[6] ) );
    VMW_AO22 U184 ( .A(\temp240[6] ), .B(n996), .C(InEdges[22]), .D(n104), .Z(
        \temp334[6] ) );
    VMW_AO22 U185 ( .A(InEdges[38]), .B(n112), .C(\temp334[6] ), .D(n997), .Z(
        \temp424[6] ) );
    VMW_AO22 U186 ( .A(InEdges[54]), .B(n120), .C(\temp424[6] ), .D(n999), .Z(
        \temp514[6] ) );
    VMW_AO22 U187 ( .A(\temp514[6] ), .B(n995), .C(InEdges[70]), .D(n128), .Z(
        \temp604[6] ) );
    VMW_AO22 U188 ( .A(InEdges[86]), .B(n136), .C(\temp604[6] ), .D(n994), .Z(
        \temp694[6] ) );
    VMW_AO22 U189 ( .A(\temp694[6] ), .B(n993), .C(InEdges[102]), .D(n144), 
        .Z(\temp784[6] ) );
    VMW_AO22 U190 ( .A(InEdges[5]), .B(n96), .C(OutEdge[5]), .D(n998), .Z(
        \temp240[5] ) );
    VMW_AO22 U191 ( .A(\temp240[5] ), .B(n996), .C(InEdges[21]), .D(n104), .Z(
        \temp334[5] ) );
    VMW_AO22 U192 ( .A(InEdges[37]), .B(n112), .C(\temp334[5] ), .D(n997), .Z(
        \temp424[5] ) );
    VMW_AO22 U193 ( .A(InEdges[53]), .B(n120), .C(\temp424[5] ), .D(n999), .Z(
        \temp514[5] ) );
    VMW_AO22 U194 ( .A(\temp514[5] ), .B(n995), .C(InEdges[69]), .D(n128), .Z(
        \temp604[5] ) );
    VMW_AO22 U195 ( .A(InEdges[85]), .B(n136), .C(\temp604[5] ), .D(n994), .Z(
        \temp694[5] ) );
    VMW_AO22 U196 ( .A(\temp694[5] ), .B(n993), .C(InEdges[101]), .D(n144), 
        .Z(\temp784[5] ) );
    VMW_AO22 U197 ( .A(InEdges[4]), .B(n96), .C(OutEdge[4]), .D(n998), .Z(
        \temp240[4] ) );
    VMW_AO22 U198 ( .A(\temp240[4] ), .B(n996), .C(InEdges[20]), .D(n104), .Z(
        \temp334[4] ) );
    VMW_AO22 U199 ( .A(InEdges[36]), .B(n112), .C(\temp334[4] ), .D(n997), .Z(
        \temp424[4] ) );
    VMW_AO22 U200 ( .A(InEdges[52]), .B(n120), .C(\temp424[4] ), .D(n999), .Z(
        \temp514[4] ) );
    VMW_AO22 U201 ( .A(\temp514[4] ), .B(n995), .C(InEdges[68]), .D(n128), .Z(
        \temp604[4] ) );
    VMW_AO22 U202 ( .A(InEdges[84]), .B(n136), .C(\temp604[4] ), .D(n994), .Z(
        \temp694[4] ) );
    VMW_AO22 U203 ( .A(\temp694[4] ), .B(n993), .C(InEdges[100]), .D(n144), 
        .Z(\temp784[4] ) );
    VMW_AO22 U204 ( .A(InEdges[3]), .B(n96), .C(OutEdge[3]), .D(n998), .Z(
        \temp240[3] ) );
    VMW_AO22 U205 ( .A(\temp240[3] ), .B(n996), .C(InEdges[19]), .D(n104), .Z(
        \temp334[3] ) );
    VMW_AO22 U206 ( .A(InEdges[35]), .B(n112), .C(\temp334[3] ), .D(n997), .Z(
        \temp424[3] ) );
    VMW_AO22 U207 ( .A(InEdges[51]), .B(n120), .C(\temp424[3] ), .D(n999), .Z(
        \temp514[3] ) );
    VMW_AO22 U208 ( .A(\temp514[3] ), .B(n995), .C(InEdges[67]), .D(n128), .Z(
        \temp604[3] ) );
    VMW_AO22 U209 ( .A(InEdges[83]), .B(n136), .C(\temp604[3] ), .D(n994), .Z(
        \temp694[3] ) );
    VMW_AO22 U210 ( .A(\temp694[3] ), .B(n993), .C(InEdges[99]), .D(n144), .Z(
        \temp784[3] ) );
    VMW_AO22 U211 ( .A(InEdges[2]), .B(n96), .C(OutEdge[2]), .D(n998), .Z(
        \temp240[2] ) );
    VMW_AO22 U212 ( .A(\temp240[2] ), .B(n996), .C(InEdges[18]), .D(n104), .Z(
        \temp334[2] ) );
    VMW_AO22 U213 ( .A(InEdges[34]), .B(n112), .C(\temp334[2] ), .D(n997), .Z(
        \temp424[2] ) );
    VMW_AO22 U214 ( .A(InEdges[50]), .B(n120), .C(\temp424[2] ), .D(n999), .Z(
        \temp514[2] ) );
    VMW_AO22 U215 ( .A(\temp514[2] ), .B(n995), .C(InEdges[66]), .D(n128), .Z(
        \temp604[2] ) );
    VMW_AO22 U216 ( .A(InEdges[82]), .B(n136), .C(\temp604[2] ), .D(n994), .Z(
        \temp694[2] ) );
    VMW_AO22 U217 ( .A(\temp694[2] ), .B(n993), .C(InEdges[98]), .D(n144), .Z(
        \temp784[2] ) );
    VMW_AO22 U218 ( .A(InEdges[1]), .B(n96), .C(OutEdge[1]), .D(n998), .Z(
        \temp240[1] ) );
    VMW_AO22 U219 ( .A(\temp240[1] ), .B(n996), .C(InEdges[17]), .D(n104), .Z(
        \temp334[1] ) );
    VMW_AO22 U220 ( .A(InEdges[33]), .B(n112), .C(\temp334[1] ), .D(n997), .Z(
        \temp424[1] ) );
    VMW_AO22 U221 ( .A(InEdges[49]), .B(n120), .C(\temp424[1] ), .D(n999), .Z(
        \temp514[1] ) );
    VMW_AO22 U222 ( .A(\temp514[1] ), .B(n995), .C(InEdges[65]), .D(n128), .Z(
        \temp604[1] ) );
    VMW_AO22 U223 ( .A(InEdges[81]), .B(n136), .C(\temp604[1] ), .D(n994), .Z(
        \temp694[1] ) );
    VMW_AO22 U224 ( .A(\temp694[1] ), .B(n993), .C(InEdges[97]), .D(n144), .Z(
        \temp784[1] ) );
    VMW_AO22 U225 ( .A(InEdges[15]), .B(n96), .C(OutEdge[15]), .D(n998), .Z(
        \temp240[15] ) );
    VMW_AO22 U226 ( .A(\temp240[15] ), .B(n996), .C(InEdges[31]), .D(n104), 
        .Z(\temp334[15] ) );
    VMW_AO22 U227 ( .A(InEdges[47]), .B(n112), .C(\temp334[15] ), .D(n997), 
        .Z(\temp424[15] ) );
    VMW_AO22 U228 ( .A(InEdges[63]), .B(n120), .C(\temp424[15] ), .D(n999), 
        .Z(\temp514[15] ) );
    VMW_AO22 U229 ( .A(\temp514[15] ), .B(n995), .C(InEdges[79]), .D(n128), 
        .Z(\temp604[15] ) );
    VMW_AO22 U230 ( .A(InEdges[95]), .B(n136), .C(\temp604[15] ), .D(n994), 
        .Z(\temp694[15] ) );
    VMW_AO22 U231 ( .A(InEdges[14]), .B(n96), .C(OutEdge[14]), .D(n998), .Z(
        \temp240[14] ) );
    VMW_AO22 U232 ( .A(\temp240[14] ), .B(n996), .C(InEdges[30]), .D(n104), 
        .Z(\temp334[14] ) );
    VMW_AO22 U233 ( .A(InEdges[46]), .B(n112), .C(\temp334[14] ), .D(n997), 
        .Z(\temp424[14] ) );
    VMW_AO22 U234 ( .A(InEdges[62]), .B(n120), .C(\temp424[14] ), .D(n999), 
        .Z(\temp514[14] ) );
    VMW_AO22 U235 ( .A(\temp514[14] ), .B(n995), .C(InEdges[78]), .D(n128), 
        .Z(\temp604[14] ) );
    VMW_AO22 U236 ( .A(InEdges[94]), .B(n136), .C(\temp604[14] ), .D(n994), 
        .Z(\temp694[14] ) );
    VMW_AO22 U237 ( .A(\temp694[14] ), .B(n993), .C(InEdges[110]), .D(n144), 
        .Z(\temp784[14] ) );
    VMW_AO22 U238 ( .A(InEdges[13]), .B(n96), .C(OutEdge[13]), .D(n998), .Z(
        \temp240[13] ) );
    VMW_AO22 U239 ( .A(\temp240[13] ), .B(n996), .C(InEdges[29]), .D(n104), 
        .Z(\temp334[13] ) );
    VMW_AO22 U240 ( .A(InEdges[45]), .B(n112), .C(\temp334[13] ), .D(n997), 
        .Z(\temp424[13] ) );
    VMW_AO22 U241 ( .A(InEdges[61]), .B(n120), .C(\temp424[13] ), .D(n999), 
        .Z(\temp514[13] ) );
    VMW_AO22 U242 ( .A(\temp514[13] ), .B(n995), .C(InEdges[77]), .D(n128), 
        .Z(\temp604[13] ) );
    VMW_AO22 U243 ( .A(InEdges[93]), .B(n136), .C(\temp604[13] ), .D(n994), 
        .Z(\temp694[13] ) );
    VMW_AO22 U244 ( .A(\temp694[13] ), .B(n993), .C(InEdges[109]), .D(n144), 
        .Z(\temp784[13] ) );
    VMW_AO22 U245 ( .A(InEdges[12]), .B(n96), .C(OutEdge[12]), .D(n998), .Z(
        \temp240[12] ) );
    VMW_AO22 U246 ( .A(\temp240[12] ), .B(n996), .C(InEdges[28]), .D(n104), 
        .Z(\temp334[12] ) );
    VMW_AO22 U247 ( .A(InEdges[44]), .B(n112), .C(\temp334[12] ), .D(n997), 
        .Z(\temp424[12] ) );
    VMW_AO22 U248 ( .A(InEdges[60]), .B(n120), .C(\temp424[12] ), .D(n999), 
        .Z(\temp514[12] ) );
    VMW_AO22 U249 ( .A(\temp514[12] ), .B(n995), .C(InEdges[76]), .D(n128), 
        .Z(\temp604[12] ) );
    VMW_AO22 U250 ( .A(InEdges[92]), .B(n136), .C(\temp604[12] ), .D(n994), 
        .Z(\temp694[12] ) );
    VMW_AO22 U251 ( .A(\temp694[12] ), .B(n993), .C(InEdges[108]), .D(n144), 
        .Z(\temp784[12] ) );
    VMW_AO22 U252 ( .A(InEdges[11]), .B(n96), .C(OutEdge[11]), .D(n998), .Z(
        \temp240[11] ) );
    VMW_AO22 U253 ( .A(\temp240[11] ), .B(n996), .C(InEdges[27]), .D(n104), 
        .Z(\temp334[11] ) );
    VMW_AO22 U254 ( .A(InEdges[43]), .B(n112), .C(\temp334[11] ), .D(n997), 
        .Z(\temp424[11] ) );
    VMW_AO22 U255 ( .A(InEdges[59]), .B(n120), .C(\temp424[11] ), .D(n999), 
        .Z(\temp514[11] ) );
    VMW_AO22 U256 ( .A(\temp514[11] ), .B(n995), .C(InEdges[75]), .D(n128), 
        .Z(\temp604[11] ) );
    VMW_AO22 U257 ( .A(InEdges[91]), .B(n136), .C(\temp604[11] ), .D(n994), 
        .Z(\temp694[11] ) );
    VMW_AO22 U258 ( .A(\temp694[11] ), .B(n993), .C(InEdges[107]), .D(n144), 
        .Z(\temp784[11] ) );
    VMW_AO22 U259 ( .A(InEdges[10]), .B(n96), .C(OutEdge[10]), .D(n998), .Z(
        \temp240[10] ) );
    VMW_AO22 U260 ( .A(\temp240[10] ), .B(n996), .C(InEdges[26]), .D(n104), 
        .Z(\temp334[10] ) );
    VMW_AO22 U261 ( .A(InEdges[42]), .B(n112), .C(\temp334[10] ), .D(n997), 
        .Z(\temp424[10] ) );
    VMW_AO22 U262 ( .A(InEdges[58]), .B(n120), .C(\temp424[10] ), .D(n999), 
        .Z(\temp514[10] ) );
    VMW_AO22 U263 ( .A(\temp514[10] ), .B(n995), .C(InEdges[74]), .D(n128), 
        .Z(\temp604[10] ) );
    VMW_AO22 U264 ( .A(InEdges[90]), .B(n136), .C(\temp604[10] ), .D(n994), 
        .Z(\temp694[10] ) );
    VMW_AO22 U265 ( .A(\temp694[10] ), .B(n993), .C(InEdges[106]), .D(n144), 
        .Z(\temp784[10] ) );
    VMW_AO22 U266 ( .A(InEdges[0]), .B(n96), .C(OutEdge[0]), .D(n998), .Z(
        \temp240[0] ) );
    VMW_AO22 U267 ( .A(\temp240[0] ), .B(n996), .C(InEdges[16]), .D(n104), .Z(
        \temp334[0] ) );
    VMW_AO22 U268 ( .A(InEdges[32]), .B(n112), .C(\temp334[0] ), .D(n997), .Z(
        \temp424[0] ) );
    VMW_AO22 U269 ( .A(InEdges[48]), .B(n120), .C(\temp424[0] ), .D(n999), .Z(
        \temp514[0] ) );
    VMW_AO22 U270 ( .A(\temp514[0] ), .B(n995), .C(InEdges[64]), .D(n128), .Z(
        \temp604[0] ) );
    VMW_AO22 U271 ( .A(InEdges[80]), .B(n136), .C(\temp604[0] ), .D(n994), .Z(
        \temp694[0] ) );
    VMW_AO22 U272 ( .A(\temp694[0] ), .B(n993), .C(InEdges[96]), .D(n144), .Z(
        \temp784[0] ) );
    VMW_MUX2I U273 ( .A(\temp784[9] ), .B(InEdges[121]), .S(n152), .Z(n974) );
    VMW_MUX2I U274 ( .A(\temp784[8] ), .B(InEdges[120]), .S(n152), .Z(n975) );
    VMW_MUX2I U275 ( .A(\temp784[7] ), .B(InEdges[119]), .S(n152), .Z(n976) );
    VMW_MUX2I U276 ( .A(\temp784[6] ), .B(InEdges[118]), .S(n152), .Z(n977) );
    VMW_MUX2I U277 ( .A(\temp784[5] ), .B(InEdges[117]), .S(n152), .Z(n978) );
    VMW_MUX2I U278 ( .A(\temp784[4] ), .B(InEdges[116]), .S(n152), .Z(n979) );
    VMW_MUX2I U279 ( .A(\temp784[3] ), .B(InEdges[115]), .S(n152), .Z(n980) );
    VMW_MUX2I U280 ( .A(\temp784[2] ), .B(InEdges[114]), .S(n152), .Z(n981) );
    VMW_MUX2I U281 ( .A(\temp784[1] ), .B(InEdges[113]), .S(n152), .Z(n982) );
    VMW_MUX2I U282 ( .A(\temp784[14] ), .B(InEdges[126]), .S(n152), .Z(n968)
         );
    VMW_MUX2I U283 ( .A(\temp784[13] ), .B(InEdges[125]), .S(n152), .Z(n970)
         );
    VMW_MUX2I U284 ( .A(\temp784[12] ), .B(InEdges[124]), .S(n152), .Z(n971)
         );
    VMW_MUX2I U285 ( .A(\temp784[11] ), .B(InEdges[123]), .S(n152), .Z(n972)
         );
    VMW_MUX2I U286 ( .A(\temp784[10] ), .B(InEdges[122]), .S(n152), .Z(n973)
         );
    VMW_MUX2I U287 ( .A(\temp784[0] ), .B(InEdges[112]), .S(n152), .Z(n983) );
    VMW_INV U288 ( .A(n96), .Z(n998) );
    VMW_INV U289 ( .A(n104), .Z(n996) );
    VMW_INV U290 ( .A(n128), .Z(n995) );
    VMW_INV U291 ( .A(n144), .Z(n993) );
    VMW_INV U292 ( .A(n984), .Z(n1002) );
    VMW_INV U293 ( .A(n1000), .Z(n1014) );
    VMW_INV U294 ( .A(n1001), .Z(n1013) );
    VMW_BUFIZ U295 ( .A(\path[3] ), .E(n1012), .Z(\PathData[3] ) );
    VMW_BUFIZ U296 ( .A(\path[1] ), .E(n1012), .Z(\PathData[1] ) );
    VMW_BUFIZ U297 ( .A(\path[0] ), .E(n1012), .Z(\PathData[0] ) );
    VMW_BUFIZ U298 ( .A(\path[2] ), .E(n1012), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n1013), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n1014), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[3]  ( .D(n1015), .CP(Clk), .Q(\path[3] ) );
    VMW_FD \path_reg[1]  ( .D(n1016), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge166[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge166[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge166[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge166[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge166[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge166[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge166[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge166[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge166[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge166[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge166[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge166[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge166[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge166[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge166[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge166[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_7 lte_55_2 ( .A({\temp334[15] , 
        \temp334[14] , \temp334[13] , \temp334[12] , \temp334[11] , 
        \temp334[10] , \temp334[9] , \temp334[8] , \temp334[7] , \temp334[6] , 
        \temp334[5] , \temp334[4] , \temp334[3] , \temp334[2] , \temp334[1] , 
        \temp334[0] }), .B(InEdges[47:32]), .LEQ(n1024), .TC(n1024), .GE_GT(
        n112) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_6 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n1023), .TC(n1023), .GE_GT(n96) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_5 lte_55_4 ( .A({\temp514[15] , 
        \temp514[14] , \temp514[13] , \temp514[12] , \temp514[11] , 
        \temp514[10] , \temp514[9] , \temp514[8] , \temp514[7] , \temp514[6] , 
        \temp514[5] , \temp514[4] , \temp514[3] , \temp514[2] , \temp514[1] , 
        \temp514[0] }), .B(InEdges[79:64]), .LEQ(n1022), .TC(n1022), .GE_GT(
        n128) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp604[15] , 
        \temp604[14] , \temp604[13] , \temp604[12] , \temp604[11] , 
        \temp604[10] , \temp604[9] , \temp604[8] , \temp604[7] , \temp604[6] , 
        \temp604[5] , \temp604[4] , \temp604[3] , \temp604[2] , \temp604[1] , 
        \temp604[0] }), .B(InEdges[95:80]), .LEQ(n1021), .TC(n1021), .GE_GT(
        n136) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_3 lte_55_1 ( .A({\temp240[15] , 
        \temp240[14] , \temp240[13] , \temp240[12] , \temp240[11] , 
        \temp240[10] , \temp240[9] , \temp240[8] , \temp240[7] , \temp240[6] , 
        \temp240[5] , \temp240[4] , \temp240[3] , \temp240[2] , \temp240[1] , 
        \temp240[0] }), .B(InEdges[31:16]), .LEQ(n1020), .TC(n1020), .GE_GT(
        n104) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_2 lte_55_7 ( .A({\temp784[15] , 
        \temp784[14] , \temp784[13] , \temp784[12] , \temp784[11] , 
        \temp784[10] , \temp784[9] , \temp784[8] , \temp784[7] , \temp784[6] , 
        \temp784[5] , \temp784[4] , \temp784[3] , \temp784[2] , \temp784[1] , 
        \temp784[0] }), .B(InEdges[127:112]), .LEQ(n1019), .TC(n1019), .GE_GT(
        n152) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_1 lte_55_6 ( .A({\temp694[15] , 
        \temp694[14] , \temp694[13] , \temp694[12] , \temp694[11] , 
        \temp694[10] , \temp694[9] , \temp694[8] , \temp694[7] , \temp694[6] , 
        \temp694[5] , \temp694[4] , \temp694[3] , \temp694[2] , \temp694[1] , 
        \temp694[0] }), .B(InEdges[111:96]), .LEQ(n1018), .TC(n1018), .GE_GT(
        n144) );
    NodeAux_INDEGREE8_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp424[15] , 
        \temp424[14] , \temp424[13] , \temp424[12] , \temp424[11] , 
        \temp424[10] , \temp424[9] , \temp424[8] , \temp424[7] , \temp424[6] , 
        \temp424[5] , \temp424[4] , \temp424[3] , \temp424[2] , \temp424[1] , 
        \temp424[0] }), .B(InEdges[63:48]), .LEQ(n1017), .TC(n1017), .GE_GT(
        n120) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
input  [7:0] WeightAddr;
input  [7:0] Eid;
output [3:0] PathData;
input  [15:0] WeightData;
input  [5:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[15:0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE0_SOURCE0 n_0_0 ( .Nid(Nid), .InEdges(InEdges[1:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE0 n_1_0 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges[63:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE5_SOURCE0 n_5_0 ( .Nid(Nid), .InEdges(InEdges[79:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE0 n_6_0 ( .Nid(Nid), .InEdges(InEdges[95:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE7_SOURCE0 n_7_0 ( .Nid(Nid), .InEdges(InEdges[111:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE8_SOURCE0 n_8_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[47:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE1 n_6_1 ( .Nid(Nid), .InEdges(InEdges[95:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID64 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID65 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID66 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID67 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID68 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID69 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID70 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID71 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID72 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID73 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID74 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID75 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID16_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID76 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID77 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID78 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID79 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID80 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID81 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID17_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID82 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID18_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID83 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID84 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID85 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID86 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID87 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID88 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID89 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID19_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID90 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID91 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID20_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID92 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID93 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID94 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID21_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID95 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID96 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID97 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID98 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID99 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID22_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID23_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID24_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID25_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID26_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID27_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID28_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID29_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID30_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID31_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID32_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID33_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID34_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID35_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID36_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID37_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID38_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID39_INDEGREE0 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [-1:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE0_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule


module Node_NID40_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID41_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID42_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID43_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID44_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID45_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID46_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID47_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID48_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID49_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID50_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID51_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID52_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID53_INDEGREE8 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [127:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE8_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID224 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID225 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID54_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID226 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID227 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID55_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID228 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID229 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID230 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID56_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID231 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID232 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID57_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID233 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID234 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID235 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID236 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID58_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID237 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID238 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID239 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID59_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID240 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID241 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID242 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID243 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID60_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID244 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID245 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID246 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID61_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID247 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID248 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID62_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID249 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID250 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID251 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID252 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID253 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID63_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [5:0] PathAddr;
output [3:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID254 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID255 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [7:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [7:0] WeightAddr;
input  [15:0] WeightData;
input  [5:0] PathAddr;
output [3:0] PathData;
input  Start, Clk;
    wire [95:0] In0;
    wire [15:0] Out0;
    wire [79:0] In1;
    wire [15:0] Out1;
    wire [79:0] In2;
    wire [15:0] Out2;
    wire [15:0] In3;
    wire [15:0] Out3;
    wire [95:0] In4;
    wire [15:0] Out4;
    wire [127:0] In5;
    wire [15:0] Out5;
    wire [79:0] In6;
    wire [15:0] Out6;
    wire [47:0] In7;
    wire [15:0] Out7;
    wire [31:0] In8;
    wire [15:0] Out8;
    wire [63:0] In9;
    wire [15:0] Out9;
    wire [95:0] In10;
    wire [15:0] Out10;
    wire [47:0] In11;
    wire [15:0] Out11;
    wire [79:0] In12;
    wire [15:0] Out12;
    wire [79:0] In13;
    wire [15:0] Out13;
    wire [127:0] In14;
    wire [15:0] Out14;
    wire [63:0] In15;
    wire [15:0] Out15;
    wire [95:0] In16;
    wire [15:0] Out16;
    wire [15:0] In17;
    wire [15:0] Out17;
    wire [111:0] In18;
    wire [15:0] Out18;
    wire [31:0] In19;
    wire [15:0] Out19;
    wire [47:0] In20;
    wire [15:0] Out20;
    wire [79:0] In21;
    wire [15:0] Out21;
    wire [47:0] In22;
    wire [15:0] Out22;
    wire [47:0] In23;
    wire [15:0] Out23;
    wire [111:0] In24;
    wire [15:0] Out24;
    wire [15:0] In25;
    wire [15:0] Out25;
    wire [31:0] In26;
    wire [15:0] Out26;
    wire [111:0] In27;
    wire [15:0] Out27;
    wire [47:0] In28;
    wire [15:0] Out28;
    wire [31:0] In29;
    wire [15:0] Out29;
    wire [95:0] In30;
    wire [15:0] Out30;
    wire [127:0] In31;
    wire [15:0] Out31;
    wire [47:0] In32;
    wire [15:0] Out32;
    wire [15:0] In33;
    wire [15:0] Out33;
    wire [47:0] In34;
    wire [15:0] Out34;
    wire [95:0] In35;
    wire [15:0] Out35;
    wire [47:0] In36;
    wire [15:0] Out36;
    wire [31:0] In37;
    wire [15:0] Out37;
    wire [79:0] In38;
    wire [15:0] Out38;
    wire [-1:0] In39;
    wire [15:0] Out39;
    wire [63:0] In40;
    wire [15:0] Out40;
    wire [47:0] In41;
    wire [15:0] Out41;
    wire [79:0] In42;
    wire [15:0] Out42;
    wire [63:0] In43;
    wire [15:0] Out43;
    wire [79:0] In44;
    wire [15:0] Out44;
    wire [31:0] In45;
    wire [15:0] Out45;
    wire [79:0] In46;
    wire [15:0] Out46;
    wire [79:0] In47;
    wire [15:0] Out47;
    wire [15:0] In48;
    wire [15:0] Out48;
    wire [79:0] In49;
    wire [15:0] Out49;
    wire [63:0] In50;
    wire [15:0] Out50;
    wire [79:0] In51;
    wire [15:0] Out51;
    wire [79:0] In52;
    wire [15:0] Out52;
    wire [127:0] In53;
    wire [15:0] Out53;
    wire [31:0] In54;
    wire [15:0] Out54;
    wire [47:0] In55;
    wire [15:0] Out55;
    wire [31:0] In56;
    wire [15:0] Out56;
    wire [63:0] In57;
    wire [15:0] Out57;
    wire [47:0] In58;
    wire [15:0] Out58;
    wire [63:0] In59;
    wire [15:0] Out59;
    wire [47:0] In60;
    wire [15:0] Out60;
    wire [31:0] In61;
    wire [15:0] Out61;
    wire [79:0] In62;
    wire [15:0] Out62;
    wire [31:0] In63;
    wire [15:0] Out63;

    Node_NID0_INDEGREE6 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out59), .OutEdge(In0[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out48), .OutEdge(In0[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out43), .OutEdge(In0[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out15), .OutEdge(In0[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out12), .OutEdge(In0[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out5), .OutEdge(In0[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE5 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out52), .OutEdge(In1[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out38), .OutEdge(In1[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out28), .OutEdge(In1[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out20), .OutEdge(In1[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out3), .OutEdge(In1[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE5 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out58), .OutEdge(In2[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out36), .OutEdge(In2[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out29), .OutEdge(In2[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out23), .OutEdge(In2[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out3), .OutEdge(In2[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE1 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out8), .OutEdge(In3[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE6 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out44), .OutEdge(In4[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out39), .OutEdge(In4[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out34), .OutEdge(In4[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out30), .OutEdge(In4[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out23), .OutEdge(In4[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out8), .OutEdge(In4[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE8 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out60), .OutEdge(In5[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out58), .OutEdge(In5[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out50), .OutEdge(In5[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out49), .OutEdge(In5[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out41), .OutEdge(In5[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out36), .OutEdge(In5[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out18), .OutEdge(In5[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out9), .OutEdge(In5[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE5 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out45), .OutEdge(In6[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out38), .OutEdge(In6[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out34), .OutEdge(In6[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out29), .OutEdge(In6[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out21), .OutEdge(In6[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE3 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out52), .OutEdge(In7[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out29), .OutEdge(In7[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out14), .OutEdge(In7[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE2 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out50), .OutEdge(In8[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out23), .OutEdge(In8[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE4 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out54), .OutEdge(In9[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out47), .OutEdge(In9[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out40), .OutEdge(In9[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out36), .OutEdge(In9[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE6 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out38), .OutEdge(In10[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out24), .OutEdge(In10[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out22), .OutEdge(In10[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out20), .OutEdge(In10[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out18), .OutEdge(In10[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out7), .OutEdge(In10[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE3 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out36), .OutEdge(In11[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out20), .OutEdge(In11[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out19), .OutEdge(In11[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE5 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out59), .OutEdge(In12[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out58), .OutEdge(In12[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out28), .OutEdge(In12[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out24), .OutEdge(In12[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out7), .OutEdge(In12[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE5 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out60), .OutEdge(In13[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out39), .OutEdge(In13[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out14), .OutEdge(In13[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out8), .OutEdge(In13[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out3), .OutEdge(In13[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE8 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID64 e64 ( .InEdge(Out52), .OutEdge(In14[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID65 e65 ( .InEdge(Out51), .OutEdge(In14[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID66 e66 ( .InEdge(Out49), .OutEdge(In14[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID67 e67 ( .InEdge(Out47), .OutEdge(In14[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID68 e68 ( .InEdge(Out42), .OutEdge(In14[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID69 e69 ( .InEdge(Out39), .OutEdge(In14[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID70 e70 ( .InEdge(Out36), .OutEdge(In14[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID71 e71 ( .InEdge(Out29), .OutEdge(In14[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE4 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID72 e72 ( .InEdge(Out54), .OutEdge(In15[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID73 e73 ( .InEdge(Out48), .OutEdge(In15[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID74 e74 ( .InEdge(Out46), .OutEdge(In15[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID75 e75 ( .InEdge(Out11), .OutEdge(In15[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID16_INDEGREE6 n16 ( .InEdges(In16), .OutEdge(Out16),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID76 e76 ( .InEdge(Out60), .OutEdge(In16[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID77 e77 ( .InEdge(Out54), .OutEdge(In16[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID78 e78 ( .InEdge(Out52), .OutEdge(In16[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID79 e79 ( .InEdge(Out34), .OutEdge(In16[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID80 e80 ( .InEdge(Out19), .OutEdge(In16[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID81 e81 ( .InEdge(Out18), .OutEdge(In16[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID17_INDEGREE1 n17 ( .InEdges(In17), .OutEdge(Out17),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID82 e82 ( .InEdge(Out41), .OutEdge(In17[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID18_INDEGREE7 n18 ( .InEdges(In18), .OutEdge(Out18),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID83 e83 ( .InEdge(Out52), .OutEdge(In18[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID84 e84 ( .InEdge(Out50), .OutEdge(In18[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID85 e85 ( .InEdge(Out44), .OutEdge(In18[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID86 e86 ( .InEdge(Out32), .OutEdge(In18[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID87 e87 ( .InEdge(Out29), .OutEdge(In18[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID88 e88 ( .InEdge(Out20), .OutEdge(In18[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID89 e89 ( .InEdge(Out11), .OutEdge(In18[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID19_INDEGREE2 n19 ( .InEdges(In19), .OutEdge(Out19),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID90 e90 ( .InEdge(Out47), .OutEdge(In19[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID91 e91 ( .InEdge(Out13), .OutEdge(In19[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID20_INDEGREE3 n20 ( .InEdges(In20), .OutEdge(Out20),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID92 e92 ( .InEdge(Out44), .OutEdge(In20[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID93 e93 ( .InEdge(Out28), .OutEdge(In20[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID94 e94 ( .InEdge(Out5), .OutEdge(In20[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID21_INDEGREE5 n21 ( .InEdges(In21), .OutEdge(Out21),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID95 e95 ( .InEdge(Out46), .OutEdge(In21[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID96 e96 ( .InEdge(Out44), .OutEdge(In21[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID97 e97 ( .InEdge(Out32), .OutEdge(In21[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID98 e98 ( .InEdge(Out31), .OutEdge(In21[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID99 e99 ( .InEdge(Out22), .OutEdge(In21[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID22_INDEGREE3 n22 ( .InEdges(In22), .OutEdge(Out22),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID100 e100 ( .InEdge(Out55), .OutEdge(In22[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID101 e101 ( .InEdge(Out49), .OutEdge(In22[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID102 e102 ( .InEdge(Out5), .OutEdge(In22[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID23_INDEGREE3 n23 ( .InEdges(In23), .OutEdge(Out23),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID103 e103 ( .InEdge(Out61), .OutEdge(In23[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID104 e104 ( .InEdge(Out55), .OutEdge(In23[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID105 e105 ( .InEdge(Out18), .OutEdge(In23[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID24_INDEGREE7 n24 ( .InEdges(In24), .OutEdge(Out24),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID106 e106 ( .InEdge(Out63), .OutEdge(In24[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID107 e107 ( .InEdge(Out42), .OutEdge(In24[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID108 e108 ( .InEdge(Out35), .OutEdge(In24[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID109 e109 ( .InEdge(Out31), .OutEdge(In24[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID110 e110 ( .InEdge(Out14), .OutEdge(In24[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID111 e111 ( .InEdge(Out8), .OutEdge(In24[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID112 e112 ( .InEdge(Out0), .OutEdge(In24[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID25_INDEGREE1 n25 ( .InEdges(In25), .OutEdge(Out25),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID113 e113 ( .InEdge(Out28), .OutEdge(In25[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID26_INDEGREE2 n26 ( .InEdges(In26), .OutEdge(Out26),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID114 e114 ( .InEdge(Out39), .OutEdge(In26[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID115 e115 ( .InEdge(Out0), .OutEdge(In26[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID27_INDEGREE7 n27 ( .InEdges(In27), .OutEdge(Out27),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID116 e116 ( .InEdge(Out59), .OutEdge(In27[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID117 e117 ( .InEdge(Out52), .OutEdge(In27[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID118 e118 ( .InEdge(Out34), .OutEdge(In27[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID119 e119 ( .InEdge(Out33), .OutEdge(In27[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID120 e120 ( .InEdge(Out18), .OutEdge(In27[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID121 e121 ( .InEdge(Out17), .OutEdge(In27[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID122 e122 ( .InEdge(Out13), .OutEdge(In27[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID28_INDEGREE3 n28 ( .InEdges(In28), .OutEdge(Out28),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID123 e123 ( .InEdge(Out49), .OutEdge(In28[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID124 e124 ( .InEdge(Out42), .OutEdge(In28[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID125 e125 ( .InEdge(Out21), .OutEdge(In28[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID29_INDEGREE2 n29 ( .InEdges(In29), .OutEdge(Out29),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID126 e126 ( .InEdge(Out38), .OutEdge(In29[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID127 e127 ( .InEdge(Out33), .OutEdge(In29[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID30_INDEGREE6 n30 ( .InEdges(In30), .OutEdge(Out30),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID128 e128 ( .InEdge(Out63), .OutEdge(In30[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID129 e129 ( .InEdge(Out38), .OutEdge(In30[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID130 e130 ( .InEdge(Out37), .OutEdge(In30[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID131 e131 ( .InEdge(Out22), .OutEdge(In30[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID132 e132 ( .InEdge(Out2), .OutEdge(In30[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID133 e133 ( .InEdge(Out0), .OutEdge(In30[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID31_INDEGREE8 n31 ( .InEdges(In31), .OutEdge(Out31),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID134 e134 ( .InEdge(Out56), .OutEdge(In31[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID135 e135 ( .InEdge(Out48), .OutEdge(In31[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID136 e136 ( .InEdge(Out46), .OutEdge(In31[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID137 e137 ( .InEdge(Out44), .OutEdge(In31[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID138 e138 ( .InEdge(Out43), .OutEdge(In31[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID139 e139 ( .InEdge(Out29), .OutEdge(In31[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID140 e140 ( .InEdge(Out18), .OutEdge(In31[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID141 e141 ( .InEdge(Out14), .OutEdge(In31[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID32_INDEGREE3 n32 ( .InEdges(In32), .OutEdge(Out32),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID142 e142 ( .InEdge(Out58), .OutEdge(In32[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID143 e143 ( .InEdge(Out39), .OutEdge(In32[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID144 e144 ( .InEdge(Out12), .OutEdge(In32[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID33_INDEGREE1 n33 ( .InEdges(In33), .OutEdge(Out33),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID145 e145 ( .InEdge(Out57), .OutEdge(In33[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID34_INDEGREE3 n34 ( .InEdges(In34), .OutEdge(Out34),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID146 e146 ( .InEdge(Out42), .OutEdge(In34[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID147 e147 ( .InEdge(Out37), .OutEdge(In34[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID148 e148 ( .InEdge(Out12), .OutEdge(In34[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID35_INDEGREE6 n35 ( .InEdges(In35), .OutEdge(Out35),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID149 e149 ( .InEdge(Out58), .OutEdge(In35[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID150 e150 ( .InEdge(Out54), .OutEdge(In35[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID151 e151 ( .InEdge(Out51), .OutEdge(In35[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID152 e152 ( .InEdge(Out20), .OutEdge(In35[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID153 e153 ( .InEdge(Out5), .OutEdge(In35[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID154 e154 ( .InEdge(Out0), .OutEdge(In35[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID36_INDEGREE3 n36 ( .InEdges(In36), .OutEdge(Out36),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID155 e155 ( .InEdge(Out63), .OutEdge(In36[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID156 e156 ( .InEdge(Out37), .OutEdge(In36[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID157 e157 ( .InEdge(Out3), .OutEdge(In36[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID37_INDEGREE2 n37 ( .InEdges(In37), .OutEdge(Out37),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID158 e158 ( .InEdge(Out44), .OutEdge(In37[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID159 e159 ( .InEdge(Out24), .OutEdge(In37[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID38_INDEGREE5 n38 ( .InEdges(In38), .OutEdge(Out38),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID160 e160 ( .InEdge(Out43), .OutEdge(In38[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID161 e161 ( .InEdge(Out24), .OutEdge(In38[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID162 e162 ( .InEdge(Out13), .OutEdge(In38[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID163 e163 ( .InEdge(Out10), .OutEdge(In38[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID164 e164 ( .InEdge(Out2), .OutEdge(In38[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID39_INDEGREE0 n39 ( .InEdges(In39), .OutEdge(Out39),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );

    Node_NID40_INDEGREE4 n40 ( .InEdges(In40), .OutEdge(Out40),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID165 e165 ( .InEdge(Out51), .OutEdge(In40[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID166 e166 ( .InEdge(Out27), .OutEdge(In40[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID167 e167 ( .InEdge(Out17), .OutEdge(In40[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID168 e168 ( .InEdge(Out12), .OutEdge(In40[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID41_INDEGREE3 n41 ( .InEdges(In41), .OutEdge(Out41),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID169 e169 ( .InEdge(Out32), .OutEdge(In41[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID170 e170 ( .InEdge(Out16), .OutEdge(In41[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID171 e171 ( .InEdge(Out5), .OutEdge(In41[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID42_INDEGREE5 n42 ( .InEdges(In42), .OutEdge(Out42),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID172 e172 ( .InEdge(Out50), .OutEdge(In42[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID173 e173 ( .InEdge(Out46), .OutEdge(In42[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID174 e174 ( .InEdge(Out32), .OutEdge(In42[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID175 e175 ( .InEdge(Out22), .OutEdge(In42[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID176 e176 ( .InEdge(Out13), .OutEdge(In42[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID43_INDEGREE4 n43 ( .InEdges(In43), .OutEdge(Out43),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID177 e177 ( .InEdge(Out51), .OutEdge(In43[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID178 e178 ( .InEdge(Out46), .OutEdge(In43[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID179 e179 ( .InEdge(Out24), .OutEdge(In43[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID180 e180 ( .InEdge(Out0), .OutEdge(In43[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID44_INDEGREE5 n44 ( .InEdges(In44), .OutEdge(Out44),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID181 e181 ( .InEdge(Out49), .OutEdge(In44[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID182 e182 ( .InEdge(Out33), .OutEdge(In44[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID183 e183 ( .InEdge(Out31), .OutEdge(In44[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID184 e184 ( .InEdge(Out27), .OutEdge(In44[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID185 e185 ( .InEdge(Out22), .OutEdge(In44[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID45_INDEGREE2 n45 ( .InEdges(In45), .OutEdge(Out45),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID186 e186 ( .InEdge(Out39), .OutEdge(In45[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID187 e187 ( .InEdge(Out12), .OutEdge(In45[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID46_INDEGREE5 n46 ( .InEdges(In46), .OutEdge(Out46),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID188 e188 ( .InEdge(Out50), .OutEdge(In46[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID189 e189 ( .InEdge(Out42), .OutEdge(In46[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID190 e190 ( .InEdge(Out31), .OutEdge(In46[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID191 e191 ( .InEdge(Out28), .OutEdge(In46[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID192 e192 ( .InEdge(Out16), .OutEdge(In46[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID47_INDEGREE5 n47 ( .InEdges(In47), .OutEdge(Out47),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID193 e193 ( .InEdge(Out59), .OutEdge(In47[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID194 e194 ( .InEdge(Out42), .OutEdge(In47[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID195 e195 ( .InEdge(Out39), .OutEdge(In47[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID196 e196 ( .InEdge(Out36), .OutEdge(In47[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID197 e197 ( .InEdge(Out13), .OutEdge(In47[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID48_INDEGREE1 n48 ( .InEdges(In48), .OutEdge(Out48),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID198 e198 ( .InEdge(Out47), .OutEdge(In48[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID49_INDEGREE5 n49 ( .InEdges(In49), .OutEdge(Out49),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID199 e199 ( .InEdge(Out59), .OutEdge(In49[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID200 e200 ( .InEdge(Out55), .OutEdge(In49[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID201 e201 ( .InEdge(Out43), .OutEdge(In49[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID202 e202 ( .InEdge(Out42), .OutEdge(In49[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID203 e203 ( .InEdge(Out21), .OutEdge(In49[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID50_INDEGREE4 n50 ( .InEdges(In50), .OutEdge(Out50),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID204 e204 ( .InEdge(Out51), .OutEdge(In50[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID205 e205 ( .InEdge(Out49), .OutEdge(In50[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID206 e206 ( .InEdge(Out37), .OutEdge(In50[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID207 e207 ( .InEdge(Out8), .OutEdge(In50[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID51_INDEGREE5 n51 ( .InEdges(In51), .OutEdge(Out51),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID208 e208 ( .InEdge(Out55), .OutEdge(In51[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID209 e209 ( .InEdge(Out48), .OutEdge(In51[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID210 e210 ( .InEdge(Out44), .OutEdge(In51[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID211 e211 ( .InEdge(Out38), .OutEdge(In51[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID212 e212 ( .InEdge(Out14), .OutEdge(In51[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID52_INDEGREE5 n52 ( .InEdges(In52), .OutEdge(Out52),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID213 e213 ( .InEdge(Out49), .OutEdge(In52[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID214 e214 ( .InEdge(Out43), .OutEdge(In52[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID215 e215 ( .InEdge(Out34), .OutEdge(In52[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID216 e216 ( .InEdge(Out32), .OutEdge(In52[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID217 e217 ( .InEdge(Out21), .OutEdge(In52[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID53_INDEGREE8 n53 ( .InEdges(In53), .OutEdge(Out53),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID218 e218 ( .InEdge(Out60), .OutEdge(In53[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID219 e219 ( .InEdge(Out41), .OutEdge(In53[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID220 e220 ( .InEdge(Out34), .OutEdge(In53[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID221 e221 ( .InEdge(Out33), .OutEdge(In53[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID222 e222 ( .InEdge(Out32), .OutEdge(In53[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID223 e223 ( .InEdge(Out23), .OutEdge(In53[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID224 e224 ( .InEdge(Out21), .OutEdge(In53[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID225 e225 ( .InEdge(Out0), .OutEdge(In53[127:112]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID54_INDEGREE2 n54 ( .InEdges(In54), .OutEdge(Out54),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID226 e226 ( .InEdge(Out41), .OutEdge(In54[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID227 e227 ( .InEdge(Out31), .OutEdge(In54[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID55_INDEGREE3 n55 ( .InEdges(In55), .OutEdge(Out55),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID228 e228 ( .InEdge(Out57), .OutEdge(In55[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID229 e229 ( .InEdge(Out28), .OutEdge(In55[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID230 e230 ( .InEdge(Out14), .OutEdge(In55[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID56_INDEGREE2 n56 ( .InEdges(In56), .OutEdge(Out56),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID231 e231 ( .InEdge(Out43), .OutEdge(In56[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID232 e232 ( .InEdge(Out14), .OutEdge(In56[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID57_INDEGREE4 n57 ( .InEdges(In57), .OutEdge(Out57),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID233 e233 ( .InEdge(Out47), .OutEdge(In57[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID234 e234 ( .InEdge(Out38), .OutEdge(In57[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID235 e235 ( .InEdge(Out32), .OutEdge(In57[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID236 e236 ( .InEdge(Out31), .OutEdge(In57[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID58_INDEGREE3 n58 ( .InEdges(In58), .OutEdge(Out58),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID237 e237 ( .InEdge(Out60), .OutEdge(In58[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID238 e238 ( .InEdge(Out46), .OutEdge(In58[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID239 e239 ( .InEdge(Out19), .OutEdge(In58[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID59_INDEGREE4 n59 ( .InEdges(In59), .OutEdge(Out59),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID240 e240 ( .InEdge(Out60), .OutEdge(In59[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID241 e241 ( .InEdge(Out54), .OutEdge(In59[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID242 e242 ( .InEdge(Out20), .OutEdge(In59[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID243 e243 ( .InEdge(Out5), .OutEdge(In59[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID60_INDEGREE3 n60 ( .InEdges(In60), .OutEdge(Out60),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID244 e244 ( .InEdge(Out41), .OutEdge(In60[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID245 e245 ( .InEdge(Out26), .OutEdge(In60[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID246 e246 ( .InEdge(Out8), .OutEdge(In60[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID61_INDEGREE2 n61 ( .InEdges(In61), .OutEdge(Out61),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID247 e247 ( .InEdge(Out28), .OutEdge(In61[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID248 e248 ( .InEdge(Out15), .OutEdge(In61[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID62_INDEGREE5 n62 ( .InEdges(In62), .OutEdge(Out62),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID249 e249 ( .InEdge(Out61), .OutEdge(In62[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID250 e250 ( .InEdge(Out60), .OutEdge(In62[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID251 e251 ( .InEdge(Out55), .OutEdge(In62[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID252 e252 ( .InEdge(Out33), .OutEdge(In62[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID253 e253 ( .InEdge(Out0), .OutEdge(In62[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID63_INDEGREE2 n63 ( .InEdges(In63), .OutEdge(Out63),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID254 e254 ( .InEdge(Out46), .OutEdge(In63[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID255 e255 ( .InEdge(Out34), .OutEdge(In63[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
