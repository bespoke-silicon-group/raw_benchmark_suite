
module Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Load, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  Clk, Reset, RD, WR, ScanEnable, Load;
    wire \Out[31] , \Out[5] , n175, n190, n217, n182, n222, n167, n205, n199, 
        n185, n160, n219, n169, n210, n202, n224, n172, n203, n197, \Out[24] , 
        \Out[17] , n161, n184, \Out[30] , n196, n218, \Out[29] , \Out[22] , 
        \Out[20] , \Out[13] , \Out[8] , \Out[1] , n173, n168, n211, \Out[11] , 
        n216, \Out[2] , n183, \Out[18] , \Out[3] , n174, n191, \Out[26] , 
        \Out[15] , n166, n223, \Out[7] , n204, n198, n193, \Out[27] , 
        \Out[14] , n214, n176, \Out[23] , \Out[10] , \Out[6] , n188, n206, 
        n221, \Out[28] , \Out[19] , n164, n181, \Out[0] , n186, \Out[21] , 
        \Out[12] , \Out[9] , n163, n178, n213, n201, \Out[25] , \Out[16] , 
        \Out[4] , n171, n208, n194, n179, n200, n162, n187, n209, n195, n170, 
        n212, n215, n192, n189, n177, n180, n165, n220, n207;
    assign ScanOut[31] = \Out[31] ;
    assign ScanOut[30] = \Out[30] ;
    assign ScanOut[29] = \Out[29] ;
    assign ScanOut[28] = \Out[28] ;
    assign ScanOut[27] = \Out[27] ;
    assign ScanOut[26] = \Out[26] ;
    assign ScanOut[25] = \Out[25] ;
    assign ScanOut[24] = \Out[24] ;
    assign ScanOut[23] = \Out[23] ;
    assign ScanOut[22] = \Out[22] ;
    assign ScanOut[21] = \Out[21] ;
    assign ScanOut[20] = \Out[20] ;
    assign ScanOut[19] = \Out[19] ;
    assign ScanOut[18] = \Out[18] ;
    assign ScanOut[17] = \Out[17] ;
    assign ScanOut[16] = \Out[16] ;
    assign ScanOut[15] = \Out[15] ;
    assign ScanOut[14] = \Out[14] ;
    assign ScanOut[13] = \Out[13] ;
    assign ScanOut[12] = \Out[12] ;
    assign ScanOut[11] = \Out[11] ;
    assign ScanOut[10] = \Out[10] ;
    assign ScanOut[9] = \Out[9] ;
    assign ScanOut[8] = \Out[8] ;
    assign ScanOut[7] = \Out[7] ;
    assign ScanOut[6] = \Out[6] ;
    assign ScanOut[5] = \Out[5] ;
    assign ScanOut[4] = \Out[4] ;
    assign ScanOut[3] = \Out[3] ;
    assign ScanOut[2] = \Out[2] ;
    assign ScanOut[1] = \Out[1] ;
    assign ScanOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AO21 U54 ( .A(\Out[27] ), .B(n160), .C(n188), .Z(n197) );
    VMW_AO21 U73 ( .A(ScanIn[26]), .B(ScanEnable), .C(Reset), .Z(n187) );
    VMW_AO21 U68 ( .A(ScanIn[30]), .B(ScanEnable), .C(Reset), .Z(n191) );
    VMW_AO21 U28 ( .A(\Out[1] ), .B(n160), .C(n162), .Z(n223) );
    VMW_AO21 U33 ( .A(\Out[6] ), .B(n160), .C(n167), .Z(n218) );
    VMW_AO21 U34 ( .A(\Out[7] ), .B(n160), .C(n168), .Z(n217) );
    VMW_AO21 U41 ( .A(\Out[14] ), .B(n160), .C(n175), .Z(n210) );
    VMW_AO21 U46 ( .A(\Out[19] ), .B(n160), .C(n180), .Z(n205) );
    VMW_AO21 U61 ( .A(ScanIn[8]), .B(ScanEnable), .C(Reset), .Z(n169) );
    VMW_AO21 U84 ( .A(ScanIn[16]), .B(ScanEnable), .C(Reset), .Z(n177) );
    VMW_AO21 U66 ( .A(ScanIn[3]), .B(ScanEnable), .C(Reset), .Z(n164) );
    VMW_AO21 U83 ( .A(ScanIn[17]), .B(ScanEnable), .C(Reset), .Z(n178) );
    VMW_AO21 U35 ( .A(\Out[8] ), .B(n160), .C(n169), .Z(n216) );
    VMW_AO21 U48 ( .A(\Out[21] ), .B(n160), .C(n182), .Z(n203) );
    VMW_AO21 U53 ( .A(\Out[26] ), .B(n160), .C(n187), .Z(n198) );
    VMW_AO21 U91 ( .A(ScanIn[0]), .B(ScanEnable), .C(Reset), .Z(n161) );
    VMW_AO21 U74 ( .A(ScanIn[25]), .B(ScanEnable), .C(Reset), .Z(n186) );
    VMW_FD \Out_reg[25]  ( .D(n199), .CP(Clk), .Q(\Out[25] ) );
    VMW_FD \Out_reg[16]  ( .D(n208), .CP(Clk), .Q(\Out[16] ) );
    VMW_AO21 U27 ( .A(\Out[0] ), .B(n160), .C(n161), .Z(n224) );
    VMW_AO21 U40 ( .A(\Out[13] ), .B(n160), .C(n174), .Z(n211) );
    VMW_AO21 U82 ( .A(ScanIn[18]), .B(ScanEnable), .C(Reset), .Z(n179) );
    VMW_FD \Out_reg[5]  ( .D(n219), .CP(Clk), .Q(\Out[5] ) );
    VMW_AO21 U52 ( .A(\Out[25] ), .B(n160), .C(n186), .Z(n199) );
    VMW_AO21 U67 ( .A(ScanIn[31]), .B(ScanEnable), .C(Reset), .Z(n192) );
    VMW_AO21 U75 ( .A(ScanIn[24]), .B(ScanEnable), .C(Reset), .Z(n185) );
    VMW_FD \Out_reg[12]  ( .D(n212), .CP(Clk), .Q(\Out[12] ) );
    VMW_AO21 U90 ( .A(ScanIn[10]), .B(ScanEnable), .C(Reset), .Z(n171) );
    VMW_FD \Out_reg[21]  ( .D(n203), .CP(Clk), .Q(\Out[21] ) );
    VMW_FD \Out_reg[8]  ( .D(n216), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO21 U29 ( .A(\Out[2] ), .B(n160), .C(n163), .Z(n222) );
    VMW_AO21 U47 ( .A(\Out[20] ), .B(n160), .C(n181), .Z(n204) );
    VMW_AO21 U49 ( .A(\Out[22] ), .B(n160), .C(n183), .Z(n202) );
    VMW_FD \Out_reg[31]  ( .D(n193), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n196), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n223), .CP(Clk), .Q(\Out[1] ) );
    VMW_AO21 U55 ( .A(\Out[28] ), .B(n160), .C(n189), .Z(n196) );
    VMW_AO21 U69 ( .A(ScanIn[2]), .B(ScanEnable), .C(Reset), .Z(n163) );
    VMW_FD \Out_reg[19]  ( .D(n205), .CP(Clk), .Q(\Out[19] ) );
    VMW_AO21 U72 ( .A(ScanIn[27]), .B(ScanEnable), .C(Reset), .Z(n188) );
    VMW_FD \Out_reg[3]  ( .D(n221), .CP(Clk), .Q(\Out[3] ) );
    VMW_FD \Out_reg[23]  ( .D(n201), .CP(Clk), .Q(\Out[23] ) );
    VMW_FD \Out_reg[10]  ( .D(n214), .CP(Clk), .Q(\Out[10] ) );
    VMW_AO21 U60 ( .A(ScanIn[9]), .B(ScanEnable), .C(Reset), .Z(n170) );
    VMW_FD \Out_reg[7]  ( .D(n217), .CP(Clk), .Q(\Out[7] ) );
    VMW_AO21 U32 ( .A(\Out[5] ), .B(n160), .C(n166), .Z(n219) );
    VMW_AO21 U85 ( .A(ScanIn[15]), .B(ScanEnable), .C(Reset), .Z(n176) );
    VMW_FD \Out_reg[27]  ( .D(n197), .CP(Clk), .Q(\Out[27] ) );
    VMW_FD \Out_reg[14]  ( .D(n210), .CP(Clk), .Q(\Out[14] ) );
    VMW_AO21 U30 ( .A(\Out[3] ), .B(n160), .C(n164), .Z(n221) );
    VMW_AO21 U39 ( .A(\Out[12] ), .B(n160), .C(n173), .Z(n212) );
    VMW_AO21 U57 ( .A(\Out[30] ), .B(n160), .C(n191), .Z(n194) );
    VMW_FD \Out_reg[6]  ( .D(n218), .CP(Clk), .Q(\Out[6] ) );
    VMW_AO21 U70 ( .A(ScanIn[29]), .B(ScanEnable), .C(Reset), .Z(n190) );
    VMW_AO21 U79 ( .A(ScanIn[20]), .B(ScanEnable), .C(Reset), .Z(n181) );
    VMW_FD \Out_reg[26]  ( .D(n198), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n209), .CP(Clk), .Q(\Out[15] ) );
    VMW_FD \Out_reg[18]  ( .D(n206), .CP(Clk), .Q(\Out[18] ) );
    VMW_AO21 U31 ( .A(\Out[4] ), .B(n160), .C(n165), .Z(n220) );
    VMW_AO21 U36 ( .A(\Out[9] ), .B(n160), .C(n170), .Z(n215) );
    VMW_AO21 U37 ( .A(\Out[10] ), .B(n160), .C(n171), .Z(n214) );
    VMW_AO21 U42 ( .A(\Out[15] ), .B(n160), .C(n176), .Z(n209) );
    VMW_AO21 U45 ( .A(\Out[18] ), .B(n160), .C(n179), .Z(n206) );
    VMW_AO21 U87 ( .A(ScanIn[13]), .B(ScanEnable), .C(Reset), .Z(n174) );
    VMW_FD \Out_reg[2]  ( .D(n222), .CP(Clk), .Q(\Out[2] ) );
    VMW_FD \Out_reg[11]  ( .D(n213), .CP(Clk), .Q(\Out[11] ) );
    VMW_AO21 U62 ( .A(ScanIn[7]), .B(ScanEnable), .C(Reset), .Z(n168) );
    VMW_FD \Out_reg[22]  ( .D(n202), .CP(Clk), .Q(\Out[22] ) );
    VMW_AO21 U65 ( .A(ScanIn[4]), .B(ScanEnable), .C(Reset), .Z(n165) );
    VMW_FD \Out_reg[20]  ( .D(n204), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n211), .CP(Clk), .Q(\Out[13] ) );
    VMW_AO21 U80 ( .A(ScanIn[1]), .B(ScanEnable), .C(Reset), .Z(n162) );
    VMW_FD \Out_reg[9]  ( .D(n215), .CP(Clk), .Q(\Out[9] ) );
    VMW_AO21 U50 ( .A(\Out[23] ), .B(n160), .C(n184), .Z(n201) );
    VMW_NOR2 U59 ( .A(ScanEnable), .B(Load), .Z(n160) );
    VMW_FD \Out_reg[30]  ( .D(n194), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n224), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n195), .CP(Clk), .Q(\Out[29] ) );
    VMW_AO21 U77 ( .A(ScanIn[22]), .B(ScanEnable), .C(Reset), .Z(n183) );
    VMW_AO21 U89 ( .A(ScanIn[11]), .B(ScanEnable), .C(Reset), .Z(n172) );
    VMW_FD \Out_reg[24]  ( .D(n200), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n207), .CP(Clk), .Q(\Out[17] ) );
    VMW_FD \Out_reg[4]  ( .D(n220), .CP(Clk), .Q(\Out[4] ) );
    VMW_AO21 U58 ( .A(\Out[31] ), .B(n160), .C(n192), .Z(n193) );
    VMW_AO21 U38 ( .A(\Out[11] ), .B(n160), .C(n172), .Z(n213) );
    VMW_AO21 U43 ( .A(\Out[16] ), .B(n160), .C(n177), .Z(n208) );
    VMW_AO21 U64 ( .A(ScanIn[5]), .B(ScanEnable), .C(Reset), .Z(n166) );
    VMW_AO21 U81 ( .A(ScanIn[19]), .B(ScanEnable), .C(Reset), .Z(n180) );
    VMW_AO21 U51 ( .A(\Out[24] ), .B(n160), .C(n185), .Z(n200) );
    VMW_AO21 U76 ( .A(ScanIn[23]), .B(ScanEnable), .C(Reset), .Z(n184) );
    VMW_AO21 U88 ( .A(ScanIn[12]), .B(ScanEnable), .C(Reset), .Z(n173) );
    VMW_AO21 U44 ( .A(\Out[17] ), .B(n160), .C(n178), .Z(n207) );
    VMW_AO21 U56 ( .A(\Out[29] ), .B(n160), .C(n190), .Z(n195) );
    VMW_AO21 U71 ( .A(ScanIn[28]), .B(ScanEnable), .C(Reset), .Z(n189) );
    VMW_AO21 U63 ( .A(ScanIn[6]), .B(ScanEnable), .C(Reset), .Z(n167) );
    VMW_AO21 U86 ( .A(ScanIn[14]), .B(ScanEnable), .C(Reset), .Z(n175) );
    VMW_AO21 U78 ( .A(ScanIn[21]), .B(ScanEnable), .C(Reset), .Z(n182) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n55, n72, n97, n20, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n115, n107, n90, n52, n75, 
        n98, n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, 
        n101, n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, 
        n113, n94, n23, n103, n16, n111, n31, n36, n44, n63, n86, n43, n64, 
        n81, n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, 
        n19, n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n62, 
        n87, n17, n30, n79, n110;
    VMW_AO21 U3 ( .A(n15), .B(A[31]), .C(n16), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(n115), .Z(n16) );
    VMW_INV U68 ( .A(A[30]), .Z(n110) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n74), .D(n68), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(A[6]), .Z(n30) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(B[13]), .Z(n58) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(A[28]), .Z(n103) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n77), .B(B[20]), .Z(n76) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n98) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n72) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n62) );
    VMW_NAND2 U60 ( .A(n110), .B(B[30]), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n90) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n75), .C(n73), .D(n71), .Z(n74) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n75) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n86) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n76), .Z(n85) );
    VMW_NAND2 U62 ( .A(n112), .B(A[29]), .Z(n113) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U102 ( .A(B[2]), .Z(n21) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n72), .C(n66), .D(n61), .Z(n71) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[20]), .Z(n77) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n112) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n77), .C(n81), .D(n79), .Z(n82) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n15), .C(n114), .D(n109), .Z(n115) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(A[25]), .Z(n101) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n73) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n80) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, n182, 
        n129, n185, n147, n160, n120, n132, n202, n169, n210, n155, n172, n197, 
        n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, n211, 
        n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, n193, 
        n198, n151, n176, n124, n188, n206, n136, n143, n158, n144, n163, n164, 
        n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, n138, 
        n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, n170, 
        n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, n165, 
        n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n116), .C(n117), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n119), .C(B[0]), .Z(n120) );
    VMW_AO22 U6 ( .A(A[2]), .B(n122), .C(n120), .D(A[0]), .Z(n121) );
    VMW_OR2 U14 ( .A(B[6]), .B(n131), .Z(n134) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n147), .C(n142), .D(n137), .Z(n146) );
    VMW_OR2 U54 ( .A(B[26]), .B(n195), .Z(n198) );
    VMW_INV U73 ( .A(B[27]), .Z(n204) );
    VMW_INV U96 ( .A(A[16]), .Z(n163) );
    VMW_INV U68 ( .A(A[30]), .Z(n212) );
    VMW_NAND2 U28 ( .A(n157), .B(B[14]), .Z(n156) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_OAI22 U7 ( .A(n118), .B(n121), .C(A[2]), .D(n122), .Z(n123) );
    VMW_NAND2 U8 ( .A(n125), .B(B[4]), .Z(n124) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n133), .C(n129), .D(n124), .Z(n132) );
    VMW_OR2 U34 ( .A(B[16]), .B(n163), .Z(n166) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n179), .C(n174), .D(n169), .Z(n178) );
    VMW_NAND2 U46 ( .A(n185), .B(A[21]), .Z(n186) );
    VMW_NAND2 U61 ( .A(n209), .B(A[29]), .Z(n210) );
    VMW_INV U84 ( .A(A[4]), .Z(n125) );
    VMW_INV U101 ( .A(B[2]), .Z(n122) );
    VMW_INV U66 ( .A(B[7]), .Z(n140) );
    VMW_INV U83 ( .A(B[15]), .Z(n165) );
    VMW_INV U98 ( .A(A[26]), .Z(n195) );
    VMW_NAND2 U26 ( .A(n153), .B(A[11]), .Z(n154) );
    VMW_NAND2 U48 ( .A(n189), .B(B[24]), .Z(n188) );
    VMW_AO21 U9 ( .A(B[3]), .B(n127), .C(n123), .Z(n126) );
    VMW_NAND2 U12 ( .A(n131), .B(B[6]), .Z(n130) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n168), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n197), .C(n193), .D(n188), .Z(n196) );
    VMW_INV U91 ( .A(A[28]), .Z(n202) );
    VMW_INV U74 ( .A(A[3]), .Z(n127) );
    VMW_INV U99 ( .A(B[23]), .Z(n191) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U40 ( .A(n177), .B(B[20]), .Z(n176) );
    VMW_INV U82 ( .A(A[15]), .Z(n168) );
    VMW_NAND2 U52 ( .A(n195), .B(B[26]), .Z(n194) );
    VMW_INV U67 ( .A(A[7]), .Z(n143) );
    VMW_INV U75 ( .A(B[25]), .Z(n197) );
    VMW_INV U90 ( .A(B[11]), .Z(n153) );
    VMW_NAND2 U20 ( .A(n145), .B(B[10]), .Z(n144) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n191), .C(n187), .D(n182), .Z(n190) );
    VMW_INV U69 ( .A(B[17]), .Z(n172) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n183), .C(n186), .D(n184), .Z(n187) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n200), .C(n198), .D(n196), .Z(n199) );
    VMW_INV U72 ( .A(A[27]), .Z(n207) );
    VMW_INV U97 ( .A(B[13]), .Z(n159) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n209), .C(n206), .D(n201), .Z(n208) );
    VMW_INV U100 ( .A(A[6]), .Z(n131) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n136), .C(n134), .D(n132), .Z(n135) );
    VMW_INV U85 ( .A(A[24]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n140), .C(n135), .D(n130), .Z(n139) );
    VMW_NAND2 U22 ( .A(n147), .B(A[9]), .Z(n148) );
    VMW_NAND2 U32 ( .A(n163), .B(B[16]), .Z(n162) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n175), .C(n173), .D(n171), .Z(n174) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n204), .C(n199), .D(n194), .Z(n203) );
    VMW_INV U70 ( .A(A[17]), .Z(n175) );
    VMW_INV U95 ( .A(B[31]), .Z(n116) );
    VMW_NAND2 U30 ( .A(n159), .B(A[13]), .Z(n160) );
    VMW_INV U79 ( .A(A[10]), .Z(n145) );
    VMW_INV U87 ( .A(B[21]), .Z(n185) );
    VMW_OR2 U10 ( .A(B[4]), .B(n125), .Z(n128) );
    VMW_NAND2 U42 ( .A(n179), .B(A[19]), .Z(n180) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n185), .C(n181), .D(n176), .Z(n184) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n151) );
    VMW_INV U80 ( .A(B[9]), .Z(n147) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n127), .C(n128), .D(n126), .Z(n129) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n143), .C(n141), .D(n139), .Z(n142) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n153), .C(n149), .D(n144), .Z(n152) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n172), .C(n167), .D(n162), .Z(n171) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n207), .C(n205), .D(n203), .Z(n206) );
    VMW_INV U89 ( .A(A[14]), .Z(n157) );
    VMW_NAND2 U50 ( .A(n191), .B(A[23]), .Z(n192) );
    VMW_INV U77 ( .A(A[20]), .Z(n177) );
    VMW_INV U92 ( .A(A[5]), .Z(n136) );
    VMW_OR2 U58 ( .A(B[28]), .B(n202), .Z(n205) );
    VMW_NAND2 U36 ( .A(n170), .B(B[18]), .Z(n169) );
    VMW_INV U81 ( .A(B[29]), .Z(n209) );
    VMW_NOR2 U4 ( .A(n119), .B(B[1]), .Z(n118) );
    VMW_OR2 U18 ( .A(B[8]), .B(n138), .Z(n141) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n177), .C(n180), .D(n178), .Z(n181) );
    VMW_AO22 U64 ( .A(n211), .B(n213), .C(A[31]), .D(n116), .Z(n117) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n189), .C(n192), .D(n190), .Z(n193) );
    VMW_INV U76 ( .A(A[25]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n145), .C(n148), .D(n146), .Z(n149) );
    VMW_NAND2 U24 ( .A(n151), .B(B[12]), .Z(n150) );
    VMW_INV U88 ( .A(A[18]), .Z(n170) );
    VMW_INV U93 ( .A(B[5]), .Z(n133) );
    VMW_OR2 U38 ( .A(B[18]), .B(n170), .Z(n173) );
    VMW_NAND2 U44 ( .A(n183), .B(B[22]), .Z(n182) );
    VMW_NAND2 U56 ( .A(n202), .B(B[28]), .Z(n201) );
    VMW_INV U94 ( .A(A[1]), .Z(n119) );
    VMW_INV U71 ( .A(A[22]), .Z(n183) );
    VMW_NAND2 U63 ( .A(n212), .B(B[30]), .Z(n213) );
    VMW_INV U86 ( .A(A[8]), .Z(n138) );
    VMW_NAND2 U16 ( .A(n138), .B(B[8]), .Z(n137) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_INV U78 ( .A(B[19]), .Z(n179) );
endmodule


module Merge_Node_DWIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Load, 
    Out, In1, In2, Read1, Read2 );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [31:0] In1;
output [31:0] Out;
input  [31:0] In2;
input  Clk, Reset, RD, WR, Load;
output Read1, Read2;
    wire n337, n339, n217, n287, n330, n317, n245, n262, n279, n230, n222, 
        n219, n257, n270, n239, n295, n305, n322, n292, n325, n302, n250, n277, 
        n225, n289, n319, n237, n259, n265, n242, n336, n218, n224, n280, n310, 
        n251, n276, n288, n318, n293, n303, n324, n338, n216, n231, n236, n243, 
        n264, n281, n311, n258, n278, n223, n238, n244, n263, n286, n316, n294, 
        n331, n304, n323, n256, n271, n70, n215, n214, n228, n284, n333, n314, 
        n246, n261, n221, n233, n328, n226, n248, n254, n268, n78, n273, n253, 
        n291, n296, n321, n301, n306, n326, n274, n227, n234, n241, n298, n308, 
        n266, n283, n313, n334, n249, n252, n275, n282, n290, n300, n327, n312, 
        n335, n235, n240, n267, n299, n309, n232, n329, n247, n260, n332, n229, 
        n285, n315, n297, n307, n320, n255, n272, n220, n269;
    VMW_PULLDOWN U36 ( .Z(n337) );
    VMW_PULLUP U37 ( .Z(n336) );
    VMW_PULLUP U39 ( .Z(n338) );
    VMW_OAI21 U40 ( .A(n70), .B(n215), .C(Load), .Z(n214) );
    VMW_AO21 U41 ( .A(n215), .B(n217), .C(Reset), .Z(n216) );
    VMW_AOI211 U46 ( .A(n219), .B(In2[5]), .C(n228), .D(n216), .Z(n227) );
    VMW_AOI211 U54 ( .A(n219), .B(In2[27]), .C(n244), .D(n216), .Z(n243) );
    VMW_AOI211 U73 ( .A(n219), .B(In2[0]), .C(n282), .D(n216), .Z(n281) );
    VMW_AO22 U113 ( .A(Out[22]), .B(n293), .C(n294), .D(In1[22]), .Z(n254) );
    VMW_INV U134 ( .A(n225), .Z(n329) );
    VMW_AOI211 U61 ( .A(n219), .B(In2[20]), .C(n258), .D(n216), .Z(n257) );
    VMW_AOI211 U68 ( .A(n219), .B(In2[14]), .C(n272), .D(n216), .Z(n271) );
    VMW_AO22 U96 ( .A(Out[9]), .B(n293), .C(n294), .D(In1[9]), .Z(n220) );
    VMW_AO22 U108 ( .A(Out[27]), .B(n293), .C(n294), .D(In1[27]), .Z(n244) );
    VMW_INV U141 ( .A(n239), .Z(n306) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_1 r140 ( .A(In1), .B(In2), .LEQ(n338), 
        .TC(n339), .GE_GT(n70) );
    VMW_AND4 U84 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(n285
        ) );
    VMW_INV U148 ( .A(n253), .Z(n313) );
    VMW_INV U153 ( .A(n263), .Z(n317) );
    VMW_AO22 U101 ( .A(Out[4]), .B(n293), .C(n294), .D(In1[4]), .Z(n230) );
    VMW_AO22 U126 ( .A(Out[10]), .B(n293), .C(n294), .D(In1[10]), .Z(n280) );
    VMW_AOI211 U48 ( .A(n219), .B(In2[3]), .C(n232), .D(n216), .Z(n231) );
    VMW_AOI211 U66 ( .A(n219), .B(In2[16]), .C(n268), .D(n216), .Z(n267) );
    VMW_AO22 U106 ( .A(Out[29]), .B(n293), .C(n294), .D(In1[29]), .Z(n240) );
    VMW_AO22 U121 ( .A(Out[15]), .B(n293), .C(n294), .D(In1[15]), .Z(n270) );
    VMW_AND4 U83 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(n286
        ) );
    VMW_AO22 U98 ( .A(Out[7]), .B(n293), .C(n294), .D(In1[7]), .Z(n224) );
    VMW_OAI21 U128 ( .A(n78), .B(n217), .C(Load), .Z(n303) );
    VMW_INV U154 ( .A(n265), .Z(n318) );
    VMW_AOI211 U53 ( .A(n219), .B(In2[28]), .C(n242), .D(n216), .Z(n241) );
    VMW_AND4 U91 ( .A(n302), .B(n301), .C(n300), .D(n299), .Z(n292) );
    VMW_INV U146 ( .A(n249), .Z(n311) );
    VMW_INV U161 ( .A(n279), .Z(n325) );
    VMW_AND5 U74 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(n287), .Z(n217)
         );
    VMW_AO22 U114 ( .A(Out[21]), .B(n293), .C(n294), .D(In1[21]), .Z(n256) );
    VMW_INV U133 ( .A(n223), .Z(n328) );
    VMW_AND4 U82 ( .A(n298), .B(n297), .C(n296), .D(n295), .Z(n287) );
    VMW_AO22 U99 ( .A(Out[6]), .B(n293), .C(n294), .D(In1[6]), .Z(n226) );
    VMW_INV U155 ( .A(n267), .Z(n319) );
    VMW_FD \Out_reg[16]  ( .D(n319), .CP(Clk), .Q(Out[16]) );
    VMW_FD \Out_reg[25]  ( .D(n310), .CP(Clk), .Q(Out[25]) );
    VMW_FD \Out_reg[5]  ( .D(n330), .CP(Clk), .Q(Out[5]) );
    VMW_AOI211 U47 ( .A(n219), .B(In2[4]), .C(n230), .D(n216), .Z(n229) );
    VMW_AOI211 U49 ( .A(n219), .B(In2[31]), .C(n234), .D(n216), .Z(n233) );
    VMW_AOI211 U52 ( .A(n219), .B(In2[29]), .C(n240), .D(n216), .Z(n239) );
    VMW_AOI211 U67 ( .A(n219), .B(In2[15]), .C(n270), .D(n216), .Z(n269) );
    VMW_AO22 U107 ( .A(Out[28]), .B(n293), .C(n294), .D(In1[28]), .Z(n242) );
    VMW_AO22 U120 ( .A(Out[16]), .B(n293), .C(n294), .D(In1[16]), .Z(n268) );
    VMW_AND5 U75 ( .A(n288), .B(n289), .C(n290), .D(n291), .E(n292), .Z(n215)
         );
    VMW_AO22 U115 ( .A(Out[20]), .B(n293), .C(n294), .D(In1[20]), .Z(n258) );
    VMW_INV U132 ( .A(n221), .Z(n327) );
    VMW_FD \Out_reg[12]  ( .D(n323), .CP(Clk), .Q(Out[12]) );
    VMW_AND4 U90 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(n302
        ) );
    VMW_FD \Out_reg[21]  ( .D(n314), .CP(Clk), .Q(Out[21]) );
    VMW_INV U129 ( .A(n214), .Z(Read1) );
    VMW_INV U147 ( .A(n251), .Z(n312) );
    VMW_FD \Out_reg[8]  ( .D(n327), .CP(Clk), .Q(Out[8]) );
    VMW_INV U160 ( .A(n277), .Z(n324) );
    VMW_FD \Out_reg[31]  ( .D(n304), .CP(Clk), .Q(Out[31]) );
    VMW_FD \Out_reg[28]  ( .D(n307), .CP(Clk), .Q(Out[28]) );
    VMW_FD \Out_reg[1]  ( .D(n334), .CP(Clk), .Q(Out[1]) );
    VMW_AOI211 U55 ( .A(n219), .B(In2[26]), .C(n246), .D(n216), .Z(n245) );
    VMW_AOI211 U69 ( .A(n219), .B(In2[13]), .C(n274), .D(n216), .Z(n273) );
    VMW_AO22 U109 ( .A(Out[26]), .B(n293), .C(n294), .D(In1[26]), .Z(n246) );
    VMW_FD \Out_reg[19]  ( .D(n316), .CP(Clk), .Q(Out[19]) );
    VMW_AOI211 U72 ( .A(n219), .B(In2[10]), .C(n280), .D(n216), .Z(n279) );
    VMW_AO22 U97 ( .A(Out[8]), .B(n293), .C(n294), .D(In1[8]), .Z(n222) );
    VMW_INV U140 ( .A(n237), .Z(n333) );
    VMW_FD \Out_reg[3]  ( .D(n332), .CP(Clk), .Q(Out[3]) );
    VMW_AO22 U112 ( .A(Out[23]), .B(n293), .C(n294), .D(In1[23]), .Z(n252) );
    VMW_INV U135 ( .A(n227), .Z(n330) );
    VMW_FD \Out_reg[10]  ( .D(n325), .CP(Clk), .Q(Out[10]) );
    VMW_FD \Out_reg[23]  ( .D(n312), .CP(Clk), .Q(Out[23]) );
    VMW_AOI211 U60 ( .A(n219), .B(In2[21]), .C(n256), .D(n216), .Z(n255) );
    VMW_FD \Out_reg[7]  ( .D(n328), .CP(Clk), .Q(Out[7]) );
    VMW_AO22 U100 ( .A(Out[5]), .B(n293), .C(n294), .D(In1[5]), .Z(n228) );
    VMW_AO22 U127 ( .A(Out[0]), .B(n293), .C(n294), .D(In1[0]), .Z(n282) );
    VMW_AOI211 U57 ( .A(n219), .B(In2[24]), .C(n250), .D(n216), .Z(n249) );
    VMW_AND4 U85 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(n284
        ) );
    VMW_INV U149 ( .A(n255), .Z(n314) );
    VMW_INV U137 ( .A(n231), .Z(n332) );
    VMW_INV U152 ( .A(n261), .Z(n316) );
    VMW_FD \Out_reg[27]  ( .D(n308), .CP(Clk), .Q(Out[27]) );
    VMW_FD \Out_reg[14]  ( .D(n321), .CP(Clk), .Q(Out[14]) );
    VMW_FD \Out_reg[6]  ( .D(n329), .CP(Clk), .Q(Out[6]) );
    VMW_AOI211 U70 ( .A(n219), .B(In2[12]), .C(n276), .D(n216), .Z(n275) );
    VMW_AO22 U110 ( .A(Out[25]), .B(n293), .C(n294), .D(In1[25]), .Z(n248) );
    VMW_INV U159 ( .A(n275), .Z(n323) );
    VMW_AOI211 U42 ( .A(n219), .B(In2[9]), .C(n220), .D(n216), .Z(n218) );
    VMW_AOI211 U45 ( .A(n219), .B(In2[6]), .C(n226), .D(n216), .Z(n225) );
    VMW_AND4 U79 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n296) );
    VMW_AND4 U95 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(n288
        ) );
    VMW_AO22 U119 ( .A(Out[17]), .B(n293), .C(n294), .D(In1[17]), .Z(n266) );
    VMW_INV U142 ( .A(n241), .Z(n307) );
    VMW_FD \Out_reg[26]  ( .D(n309), .CP(Clk), .Q(Out[26]) );
    VMW_FD \Out_reg[15]  ( .D(n320), .CP(Clk), .Q(Out[15]) );
    VMW_FD \Out_reg[18]  ( .D(n317), .CP(Clk), .Q(Out[18]) );
    VMW_AND4 U87 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n299) );
    VMW_INV U150 ( .A(n257), .Z(n315) );
    VMW_FD \Out_reg[2]  ( .D(n333), .CP(Clk), .Q(Out[2]) );
    VMW_AO22 U125 ( .A(Out[11]), .B(n293), .C(n294), .D(In1[11]), .Z(n278) );
    VMW_FD \Out_reg[11]  ( .D(n324), .CP(Clk), .Q(Out[11]) );
    VMW_AOI211 U62 ( .A(n219), .B(In2[1]), .C(n260), .D(n216), .Z(n259) );
    VMW_FD \Out_reg[22]  ( .D(n313), .CP(Clk), .Q(Out[22]) );
    VMW_AOI211 U65 ( .A(n219), .B(In2[17]), .C(n266), .D(n216), .Z(n265) );
    VMW_AO22 U102 ( .A(Out[3]), .B(n293), .C(n294), .D(In1[3]), .Z(n232) );
    VMW_AO22 U105 ( .A(Out[2]), .B(n293), .C(n294), .D(In1[2]), .Z(n238) );
    VMW_FD \Out_reg[20]  ( .D(n315), .CP(Clk), .Q(Out[20]) );
    VMW_FD \Out_reg[13]  ( .D(n322), .CP(Clk), .Q(Out[13]) );
    VMW_AND4 U80 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n297)
         );
    VMW_AO22 U122 ( .A(Out[14]), .B(n293), .C(n294), .D(In1[14]), .Z(n272) );
    VMW_INV U157 ( .A(n271), .Z(n321) );
    VMW_FD \Out_reg[9]  ( .D(n326), .CP(Clk), .Q(Out[9]) );
    VMW_AOI211 U50 ( .A(n219), .B(In2[30]), .C(n236), .D(n216), .Z(n235) );
    VMW_AOI211 U59 ( .A(n219), .B(In2[22]), .C(n254), .D(n216), .Z(n253) );
    VMW_INV U139 ( .A(n235), .Z(n305) );
    VMW_FD \Out_reg[30]  ( .D(n305), .CP(Clk), .Q(Out[30]) );
    VMW_FD \Out_reg[0]  ( .D(n335), .CP(Clk), .Q(Out[0]) );
    VMW_FD \Out_reg[29]  ( .D(n306), .CP(Clk), .Q(Out[29]) );
    VMW_AND2 U77 ( .A(n70), .B(Load), .Z(n294) );
    VMW_AND4 U89 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n301)
         );
    VMW_AND4 U92 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(n291
        ) );
    VMW_INV U145 ( .A(n247), .Z(n310) );
    VMW_INV U162 ( .A(n281), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n311), .CP(Clk), .Q(Out[24]) );
    VMW_FD \Out_reg[17]  ( .D(n318), .CP(Clk), .Q(Out[17]) );
    VMW_AO22 U117 ( .A(Out[19]), .B(n293), .C(n294), .D(In1[19]), .Z(n262) );
    VMW_FD \Out_reg[4]  ( .D(n331), .CP(Clk), .Q(Out[4]) );
    VMW_AOI211 U58 ( .A(n219), .B(In2[23]), .C(n252), .D(n216), .Z(n251) );
    VMW_INV U130 ( .A(Load), .Z(n293) );
    VMW_INV U138 ( .A(n233), .Z(n304) );
    VMW_INV U156 ( .A(n269), .Z(n320) );
    VMW_PULLDOWN U38 ( .Z(n339) );
    VMW_AOI211 U43 ( .A(n219), .B(In2[8]), .C(n222), .D(n216), .Z(n221) );
    VMW_AOI211 U64 ( .A(n219), .B(In2[18]), .C(n264), .D(n216), .Z(n263) );
    VMW_AND4 U81 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(n298
        ) );
    VMW_AO22 U104 ( .A(Out[30]), .B(n293), .C(n294), .D(In1[30]), .Z(n236) );
    VMW_AOI211 U51 ( .A(n219), .B(In2[2]), .C(n238), .D(n216), .Z(n237) );
    VMW_NOR2 U76 ( .A(n293), .B(n70), .Z(n219) );
    VMW_AO22 U116 ( .A(Out[1]), .B(n293), .C(n294), .D(In1[1]), .Z(n260) );
    VMW_AO22 U123 ( .A(Out[13]), .B(n293), .C(n294), .D(In1[13]), .Z(n274) );
    VMW_AND4 U88 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n300) );
    VMW_AND4 U93 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(n290
        ) );
    VMW_INV U131 ( .A(n218), .Z(n326) );
    VMW_INV U143 ( .A(n243), .Z(n308) );
    VMW_INV U144 ( .A(n245), .Z(n309) );
    VMW_INV U163 ( .A(n303), .Z(Read2) );
    VMW_INV U158 ( .A(n273), .Z(n322) );
    VMW_AOI211 U44 ( .A(n219), .B(In2[7]), .C(n224), .D(n216), .Z(n223) );
    VMW_AOI211 U56 ( .A(n219), .B(In2[25]), .C(n248), .D(n216), .Z(n247) );
    VMW_AND4 U94 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(n289
        ) );
    VMW_INV U136 ( .A(n229), .Z(n331) );
    VMW_AOI211 U71 ( .A(n219), .B(In2[11]), .C(n278), .D(n216), .Z(n277) );
    VMW_AO22 U111 ( .A(Out[24]), .B(n293), .C(n294), .D(In1[24]), .Z(n250) );
    VMW_AO22 U124 ( .A(Out[12]), .B(n293), .C(n294), .D(In1[12]), .Z(n276) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_0 lte_86 ( .A(In1), .B(In2), .LEQ(n336), 
        .TC(n337), .LT_LE(n78) );
    VMW_AOI211 U63 ( .A(n219), .B(In2[19]), .C(n262), .D(n216), .Z(n261) );
    VMW_AND4 U78 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n295) );
    VMW_AND4 U86 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(n283
        ) );
    VMW_AO22 U103 ( .A(Out[31]), .B(n293), .C(n294), .D(In1[31]), .Z(n234) );
    VMW_AO22 U118 ( .A(Out[18]), .B(n293), .C(n294), .D(In1[18]), .Z(n264) );
    VMW_INV U151 ( .A(n259), .Z(n334) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n28, n84, n33, n38, n56, n71, n113, n94, n23, n103, n16, 
        n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, n104, n18, n24, 
        n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, n50, n77, n89, n92, 
        n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, n87, n17, n30, n79, 
        n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n94), .Z(n97) );
    VMW_INV U73 ( .A(B[27]), .Z(n104) );
    VMW_INV U96 ( .A(A[16]), .Z(n62) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n78), .C(n73), .D(n68), .Z(n77) );
    VMW_NAND2 U46 ( .A(n84), .B(A[21]), .Z(n85) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(B[2]), .Z(n21) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(A[26]), .Z(n94) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n88), .B(B[24]), .Z(n87) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n96), .C(n92), .D(n87), .Z(n95) );
    VMW_INV U91 ( .A(A[28]), .Z(n102) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(B[23]), .Z(n90) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n76), .B(B[20]), .Z(n75) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n94), .B(B[26]), .Z(n93) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n96) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n90), .C(n86), .D(n81), .Z(n89) );
    VMW_INV U69 ( .A(B[17]), .Z(n71) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n82), .C(n85), .D(n83), .Z(n86) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n99), .C(n97), .D(n95), .Z(n98) );
    VMW_INV U72 ( .A(A[27]), .Z(n107) );
    VMW_INV U97 ( .A(B[13]), .Z(n58) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n106), .D(n101), .Z(n109) );
    VMW_INV U100 ( .A(A[6]), .Z(n30) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n74), .C(n72), .D(n70), .Z(n73) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n104), .C(n98), .D(n93), .Z(n103) );
    VMW_INV U70 ( .A(A[17]), .Z(n74) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n84) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n78), .B(A[19]), .Z(n79) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n84), .C(n80), .D(n75), .Z(n83) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n71), .C(n66), .D(n61), .Z(n70) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n107), .C(n105), .D(n103), .Z(n106) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n90), .B(A[23]), .Z(n91) );
    VMW_INV U77 ( .A(A[20]), .Z(n76) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n102), .Z(n105) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n110) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n76), .C(n79), .D(n77), .Z(n80) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n88), .C(n91), .D(n89), .Z(n92) );
    VMW_INV U76 ( .A(A[25]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n72) );
    VMW_NAND2 U44 ( .A(n82), .B(B[22]), .Z(n81) );
    VMW_NAND2 U56 ( .A(n102), .B(B[28]), .Z(n101) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n82) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n78) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n115, n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, 
        n182, n129, n185, n147, n160, n132, n202, n120, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, 
        n211, n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, 
        n193, n198, n151, n176, n124, n188, n206, n136, n144, n143, n158, n164, 
        n163, n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, 
        n138, n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, 
        n170, n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, 
        n165, n159, n137, n207;
    VMW_AO21 U3 ( .A(n115), .B(A[31]), .C(n116), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n118), .C(B[0]), .Z(n119) );
    VMW_AO22 U6 ( .A(A[2]), .B(n121), .C(n119), .D(A[0]), .Z(n120) );
    VMW_OR2 U14 ( .A(B[6]), .B(n130), .Z(n133) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n146), .C(n141), .D(n136), .Z(n145) );
    VMW_OR2 U54 ( .A(B[26]), .B(n194), .Z(n197) );
    VMW_INV U73 ( .A(B[27]), .Z(n203) );
    VMW_INV U96 ( .A(n213), .Z(n116) );
    VMW_INV U68 ( .A(A[30]), .Z(n208) );
    VMW_NAND2 U28 ( .A(n156), .B(B[14]), .Z(n155) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI22 U7 ( .A(n117), .B(n120), .C(A[2]), .D(n121), .Z(n122) );
    VMW_NAND2 U8 ( .A(n124), .B(B[4]), .Z(n123) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n132), .C(n128), .D(n123), .Z(n131) );
    VMW_OR2 U34 ( .A(B[16]), .B(n162), .Z(n165) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n178), .C(n173), .D(n168), .Z(n177) );
    VMW_NAND2 U46 ( .A(n184), .B(A[21]), .Z(n185) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n210), .C(n205), .D(n200), .Z(n209) );
    VMW_INV U84 ( .A(A[4]), .Z(n124) );
    VMW_INV U101 ( .A(A[6]), .Z(n130) );
    VMW_INV U66 ( .A(B[7]), .Z(n139) );
    VMW_INV U83 ( .A(B[15]), .Z(n164) );
    VMW_INV U98 ( .A(B[13]), .Z(n158) );
    VMW_NAND2 U26 ( .A(n152), .B(A[11]), .Z(n153) );
    VMW_NAND2 U48 ( .A(n188), .B(B[24]), .Z(n187) );
    VMW_AO21 U9 ( .A(B[3]), .B(n126), .C(n122), .Z(n125) );
    VMW_NAND2 U12 ( .A(n130), .B(B[6]), .Z(n129) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n167), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U91 ( .A(A[28]), .Z(n201) );
    VMW_INV U74 ( .A(A[3]), .Z(n126) );
    VMW_INV U99 ( .A(A[26]), .Z(n194) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U40 ( .A(n176), .B(B[20]), .Z(n175) );
    VMW_INV U82 ( .A(A[15]), .Z(n167) );
    VMW_NAND2 U52 ( .A(n194), .B(B[26]), .Z(n193) );
    VMW_INV U67 ( .A(A[7]), .Z(n142) );
    VMW_INV U75 ( .A(B[25]), .Z(n196) );
    VMW_INV U90 ( .A(B[11]), .Z(n152) );
    VMW_NAND2 U20 ( .A(n144), .B(B[10]), .Z(n143) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_INV U69 ( .A(B[17]), .Z(n171) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U72 ( .A(A[27]), .Z(n206) );
    VMW_INV U97 ( .A(A[16]), .Z(n162) );
    VMW_NAND2 U60 ( .A(n208), .B(B[30]), .Z(n207) );
    VMW_INV U100 ( .A(B[23]), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n135), .C(n133), .D(n131), .Z(n134) );
    VMW_INV U85 ( .A(A[24]), .Z(n188) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n139), .C(n134), .D(n129), .Z(n138) );
    VMW_NAND2 U22 ( .A(n146), .B(A[9]), .Z(n147) );
    VMW_NAND2 U32 ( .A(n162), .B(B[16]), .Z(n161) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n174), .C(n172), .D(n170), .Z(n173) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_INV U70 ( .A(A[17]), .Z(n174) );
    VMW_INV U95 ( .A(B[31]), .Z(n115) );
    VMW_NAND2 U30 ( .A(n158), .B(A[13]), .Z(n159) );
    VMW_INV U79 ( .A(A[10]), .Z(n144) );
    VMW_INV U87 ( .A(B[21]), .Z(n184) );
    VMW_OR2 U10 ( .A(B[4]), .B(n124), .Z(n127) );
    VMW_NAND2 U42 ( .A(n178), .B(A[19]), .Z(n179) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n184), .C(n180), .D(n175), .Z(n183) );
    VMW_NAND2 U62 ( .A(n210), .B(A[29]), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n150) );
    VMW_INV U102 ( .A(B[2]), .Z(n121) );
    VMW_INV U80 ( .A(B[9]), .Z(n146) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n126), .C(n127), .D(n125), .Z(n128) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n142), .C(n140), .D(n138), .Z(n141) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n152), .C(n148), .D(n143), .Z(n151) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n171), .C(n166), .D(n161), .Z(n170) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n206), .C(n204), .D(n202), .Z(n205) );
    VMW_INV U89 ( .A(A[14]), .Z(n156) );
    VMW_NAND2 U50 ( .A(n190), .B(A[23]), .Z(n191) );
    VMW_INV U77 ( .A(A[20]), .Z(n176) );
    VMW_INV U92 ( .A(A[5]), .Z(n135) );
    VMW_OR2 U58 ( .A(B[28]), .B(n201), .Z(n204) );
    VMW_NAND2 U36 ( .A(n169), .B(B[18]), .Z(n168) );
    VMW_INV U81 ( .A(B[29]), .Z(n210) );
    VMW_NOR2 U4 ( .A(n118), .B(B[1]), .Z(n117) );
    VMW_OR2 U18 ( .A(B[8]), .B(n137), .Z(n140) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n176), .C(n179), .D(n177), .Z(n180) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n115), .C(n212), .D(n207), .Z(n213) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_INV U76 ( .A(A[25]), .Z(n199) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n144), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U24 ( .A(n150), .B(B[12]), .Z(n149) );
    VMW_INV U88 ( .A(A[18]), .Z(n169) );
    VMW_INV U93 ( .A(B[5]), .Z(n132) );
    VMW_OR2 U38 ( .A(B[18]), .B(n169), .Z(n172) );
    VMW_NAND2 U44 ( .A(n182), .B(B[22]), .Z(n181) );
    VMW_NAND2 U56 ( .A(n201), .B(B[28]), .Z(n200) );
    VMW_INV U94 ( .A(A[1]), .Z(n118) );
    VMW_INV U71 ( .A(A[22]), .Z(n182) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n208), .C(n211), .D(n209), .Z(n212) );
    VMW_INV U86 ( .A(A[8]), .Z(n137) );
    VMW_NAND2 U16 ( .A(n137), .B(B[8]), .Z(n136) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_INV U78 ( .A(B[19]), .Z(n178) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, In1, In2, Read1, 
    Read2, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Read1, Read2;
    wire \Out[31] , n100, n245, n287, n317, n330, n262, n279, n362, n345, n357, 
        n339, n270, n257, n295, n305, n322, n292, n325, n302, n250, n277, n350, 
        n289, n319, n259, n342, n365, n265, n359, n356, \Out[5] , n280, n310, 
        n337, n288, n318, n351, \Out[24] , \Out[17] , n276, n251, \Out[30] , 
        n293, n303, n324, n281, n336, n311, \Out[29] , \Out[8] , \Out[1] , 
        n358, n243, n264, n258, n343, n364, \Out[20] , \Out[13] , \Out[26] , 
        \Out[22] , \Out[11] , \Out[18] , \Out[3] , n344, n278, n363, n244, 
        n263, n286, n316, n331, \Out[15] , n294, n304, n323, n256, n108, n271, 
        \Out[27] , \Out[14] , \Out[7] , n338, n284, n314, n333, n246, n261, 
        n361, n346, \Out[6] , n328, \Out[28] , \Out[23] , \Out[10] , \Out[19] , 
        \Out[2] , n268, n354, n368, n254, n273, n321, n306, n296, \Out[9] , 
        \Out[0] , n291, n301, n326, n348, n274, n253, n248, n353, \Out[25] , 
        \Out[21] , \Out[12] , \Out[16] , \Out[4] , n366, n298, n308, n341, 
        n266, n283, n313, n334, n249, n352, n349, n252, n275, n282, n290, n300, 
        n312, n327, n335, n267, n315, n367, n340, n299, n309, n329, n360, n347, 
        n247, n260, n332, n285, n269, n255, n297, n307, n320, n272, n355;
    assign ScanEnable = WR;
    assign DataOut[31] = \Out[31] ;
    assign DataOut[30] = \Out[30] ;
    assign DataOut[29] = \Out[29] ;
    assign DataOut[28] = \Out[28] ;
    assign DataOut[27] = \Out[27] ;
    assign DataOut[26] = \Out[26] ;
    assign DataOut[25] = \Out[25] ;
    assign DataOut[24] = \Out[24] ;
    assign DataOut[23] = \Out[23] ;
    assign DataOut[22] = \Out[22] ;
    assign DataOut[21] = \Out[21] ;
    assign DataOut[20] = \Out[20] ;
    assign DataOut[19] = \Out[19] ;
    assign DataOut[18] = \Out[18] ;
    assign DataOut[17] = \Out[17] ;
    assign DataOut[16] = \Out[16] ;
    assign DataOut[15] = \Out[15] ;
    assign DataOut[14] = \Out[14] ;
    assign DataOut[13] = \Out[13] ;
    assign DataOut[12] = \Out[12] ;
    assign DataOut[11] = \Out[11] ;
    assign DataOut[10] = \Out[10] ;
    assign DataOut[9] = \Out[9] ;
    assign DataOut[8] = \Out[8] ;
    assign DataOut[7] = \Out[7] ;
    assign DataOut[6] = \Out[6] ;
    assign DataOut[5] = \Out[5] ;
    assign DataOut[4] = \Out[4] ;
    assign DataOut[3] = \Out[3] ;
    assign DataOut[2] = \Out[2] ;
    assign DataOut[1] = \Out[1] ;
    assign DataOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AND2 U54 ( .A(DataIn[24]), .B(ScanEnable), .Z(ScanOut[24]) );
    VMW_AND2 U73 ( .A(DataIn[5]), .B(ScanEnable), .Z(ScanOut[5]) );
    VMW_AND5 U113 ( .A(n317), .B(n318), .C(n319), .D(n320), .E(n321), .Z(n246)
         );
    VMW_AO22 U134 ( .A(\Out[9] ), .B(n322), .C(n323), .D(In1[9]), .Z(n249) );
    VMW_AND2 U68 ( .A(DataIn[10]), .B(ScanEnable), .Z(ScanOut[10]) );
    VMW_AOI211 U96 ( .A(n248), .B(In2[23]), .C(n281), .D(n245), .Z(n280) );
    VMW_INV U198 ( .A(n306), .Z(n353) );
    VMW_AOI211 U108 ( .A(n248), .B(In2[12]), .C(n305), .D(n245), .Z(n304) );
    VMW_AO22 U141 ( .A(\Out[31] ), .B(n322), .C(n323), .D(In1[31]), .Z(n263)
         );
    VMW_OAI21 U166 ( .A(n108), .B(n246), .C(RD), .Z(n332) );
    VMW_INV U183 ( .A(n276), .Z(n339) );
    VMW_OAI21 U46 ( .A(n100), .B(n244), .C(RD), .Z(n243) );
    VMW_AND2 U61 ( .A(DataIn[17]), .B(ScanEnable), .Z(ScanOut[17]) );
    VMW_AOI211 U84 ( .A(n248), .B(In2[5]), .C(n257), .D(n245), .Z(n256) );
    VMW_AO22 U148 ( .A(\Out[25] ), .B(n322), .C(n323), .D(In1[25]), .Z(n277)
         );
    VMW_AO22 U153 ( .A(\Out[20] ), .B(n322), .C(n323), .D(In1[20]), .Z(n287)
         );
    VMW_INV U174 ( .A(n258), .Z(n360) );
    VMW_INV U191 ( .A(n292), .Z(n346) );
    VMW_AOI211 U101 ( .A(n248), .B(In2[19]), .C(n291), .D(n245), .Z(n290) );
    VMW_AND4 U126 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n329)
         );
    VMW_AND2 U48 ( .A(DataIn[30]), .B(ScanEnable), .Z(ScanOut[30]) );
    VMW_AND2 U66 ( .A(DataIn[12]), .B(ScanEnable), .Z(ScanOut[12]) );
    VMW_AOI211 U106 ( .A(n248), .B(In2[14]), .C(n301), .D(n245), .Z(n300) );
    VMW_AND4 U121 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(
        n320) );
    VMW_AOI211 U83 ( .A(n248), .B(In2[6]), .C(n255), .D(n245), .Z(n254) );
    VMW_INV U168 ( .A(RD), .Z(n322) );
    VMW_AOI211 U98 ( .A(n248), .B(In2[21]), .C(n285), .D(n245), .Z(n284) );
    VMW_AND4 U128 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(
        n331) );
    VMW_AO22 U154 ( .A(\Out[1] ), .B(n322), .C(n323), .D(In1[1]), .Z(n289) );
    VMW_INV U173 ( .A(n256), .Z(n359) );
    VMW_INV U184 ( .A(n278), .Z(n340) );
    VMW_INV U196 ( .A(n302), .Z(n351) );
    VMW_AND2 U53 ( .A(DataIn[25]), .B(ScanEnable), .Z(ScanOut[25]) );
    VMW_AOI211 U91 ( .A(n248), .B(In2[28]), .C(n271), .D(n245), .Z(n270) );
    VMW_AO22 U146 ( .A(\Out[27] ), .B(n322), .C(n323), .D(In1[27]), .Z(n273)
         );
    VMW_AO22 U161 ( .A(\Out[13] ), .B(n322), .C(n323), .D(In1[13]), .Z(n303)
         );
    VMW_AND2 U74 ( .A(DataIn[4]), .B(ScanEnable), .Z(ScanOut[4]) );
    VMW_NOR2 U114 ( .A(n322), .B(n100), .Z(n248) );
    VMW_AND4 U133 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(
        n312) );
    VMW_AOI211 U99 ( .A(n248), .B(In2[20]), .C(n287), .D(n245), .Z(n286) );
    VMW_INV U197 ( .A(n304), .Z(n352) );
    VMW_AO22 U155 ( .A(\Out[19] ), .B(n322), .C(n323), .D(In1[19]), .Z(n291)
         );
    VMW_FD \Out_reg[16]  ( .D(n348), .CP(Clk), .Q(\Out[16] ) );
    VMW_INV U172 ( .A(n254), .Z(n358) );
    VMW_FD \Out_reg[25]  ( .D(n339), .CP(Clk), .Q(\Out[25] ) );
    VMW_AND2 U47 ( .A(DataIn[31]), .B(ScanEnable), .Z(ScanOut[31]) );
    VMW_AND2 U49 ( .A(DataIn[29]), .B(ScanEnable), .Z(ScanOut[29]) );
    VMW_AND2 U52 ( .A(DataIn[26]), .B(ScanEnable), .Z(ScanOut[26]) );
    VMW_AND2 U67 ( .A(DataIn[11]), .B(ScanEnable), .Z(ScanOut[11]) );
    VMW_AOI211 U82 ( .A(n248), .B(In2[7]), .C(n253), .D(n245), .Z(n252) );
    VMW_INV U169 ( .A(n247), .Z(n355) );
    VMW_AOI211 U107 ( .A(n248), .B(In2[13]), .C(n303), .D(n245), .Z(n302) );
    VMW_AND4 U120 ( .A(n327), .B(n326), .C(n325), .D(n324), .Z(n321) );
    VMW_FD \Out_reg[5]  ( .D(n359), .CP(Clk), .Q(\Out[5] ) );
    VMW_AND2 U75 ( .A(DataIn[3]), .B(ScanEnable), .Z(ScanOut[3]) );
    VMW_AND2 U115 ( .A(n100), .B(RD), .Z(n323) );
    VMW_AND4 U132 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(
        n313) );
    VMW_FD \Out_reg[12]  ( .D(n352), .CP(Clk), .Q(\Out[12] ) );
    VMW_AOI211 U90 ( .A(n248), .B(In2[29]), .C(n269), .D(n245), .Z(n268) );
    VMW_FD \Out_reg[21]  ( .D(n343), .CP(Clk), .Q(\Out[21] ) );
    VMW_AND4 U129 ( .A(n331), .B(n330), .C(n329), .D(n328), .Z(n316) );
    VMW_AO22 U147 ( .A(\Out[26] ), .B(n322), .C(n323), .D(In1[26]), .Z(n275)
         );
    VMW_FD \Out_reg[8]  ( .D(n356), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO22 U160 ( .A(\Out[14] ), .B(n322), .C(n323), .D(In1[14]), .Z(n301)
         );
    VMW_INV U185 ( .A(n280), .Z(n341) );
    VMW_FD \Out_reg[31]  ( .D(n333), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n336), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n363), .CP(Clk), .Q(\Out[1] ) );
    VMW_AND2 U55 ( .A(DataIn[23]), .B(ScanEnable), .Z(ScanOut[23]) );
    VMW_AND2 U69 ( .A(ScanEnable), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AOI211 U109 ( .A(n248), .B(In2[11]), .C(n307), .D(n245), .Z(n306) );
    VMW_INV U182 ( .A(n274), .Z(n338) );
    VMW_FD \Out_reg[19]  ( .D(n345), .CP(Clk), .Q(\Out[19] ) );
    VMW_AND2 U72 ( .A(DataIn[6]), .B(ScanEnable), .Z(ScanOut[6]) );
    VMW_AOI211 U97 ( .A(n248), .B(In2[22]), .C(n283), .D(n245), .Z(n282) );
    VMW_AO22 U140 ( .A(\Out[3] ), .B(n322), .C(n323), .D(In1[3]), .Z(n261) );
    VMW_INV U167 ( .A(n243), .Z(Read1) );
    VMW_FD \Out_reg[3]  ( .D(n361), .CP(Clk), .Q(\Out[3] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 r141 ( .A(In1), .B(
        In2), .LEQ(n365), .TC(n366), .GE_GT(n100) );
    VMW_AND5 U112 ( .A(n312), .B(n313), .C(n314), .D(n315), .E(n316), .Z(n244)
         );
    VMW_AO22 U135 ( .A(\Out[8] ), .B(n322), .C(n323), .D(In1[8]), .Z(n251) );
    VMW_FD \Out_reg[10]  ( .D(n354), .CP(Clk), .Q(\Out[10] ) );
    VMW_FD \Out_reg[23]  ( .D(n341), .CP(Clk), .Q(\Out[23] ) );
    VMW_AND2 U60 ( .A(DataIn[18]), .B(ScanEnable), .Z(ScanOut[18]) );
    VMW_INV U199 ( .A(n308), .Z(n354) );
    VMW_FD \Out_reg[7]  ( .D(n357), .CP(Clk), .Q(\Out[7] ) );
    VMW_AOI211 U100 ( .A(n248), .B(In2[1]), .C(n289), .D(n245), .Z(n288) );
    VMW_AND4 U127 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n330)
         );
    VMW_AOI211 U85 ( .A(n248), .B(In2[4]), .C(n259), .D(n245), .Z(n258) );
    VMW_AO22 U149 ( .A(\Out[24] ), .B(n322), .C(n323), .D(In1[24]), .Z(n279)
         );
    VMW_AO22 U152 ( .A(\Out[21] ), .B(n322), .C(n323), .D(In1[21]), .Z(n285)
         );
    VMW_INV U175 ( .A(n260), .Z(n361) );
    VMW_FD \Out_reg[14]  ( .D(n350), .CP(Clk), .Q(\Out[14] ) );
    VMW_FD \Out_reg[27]  ( .D(n337), .CP(Clk), .Q(\Out[27] ) );
    VMW_PULLDOWN U42 ( .Z(n366) );
    VMW_PULLUP U45 ( .Z(n367) );
    VMW_AND2 U57 ( .A(DataIn[21]), .B(ScanEnable), .Z(ScanOut[21]) );
    VMW_AO22 U137 ( .A(\Out[6] ), .B(n322), .C(n323), .D(In1[6]), .Z(n255) );
    VMW_INV U190 ( .A(n290), .Z(n345) );
    VMW_FD \Out_reg[6]  ( .D(n358), .CP(Clk), .Q(\Out[6] ) );
    VMW_AND2 U70 ( .A(DataIn[8]), .B(ScanEnable), .Z(ScanOut[8]) );
    VMW_AO21 U79 ( .A(n246), .B(n244), .C(Reset), .Z(n245) );
    VMW_AOI211 U95 ( .A(n248), .B(In2[24]), .C(n279), .D(n245), .Z(n278) );
    VMW_AOI211 U110 ( .A(n248), .B(In2[10]), .C(n309), .D(n245), .Z(n308) );
    VMW_AO22 U159 ( .A(\Out[15] ), .B(n322), .C(n323), .D(In1[15]), .Z(n299)
         );
    VMW_AND4 U119 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(
        n327) );
    VMW_AO22 U142 ( .A(\Out[30] ), .B(n322), .C(n323), .D(In1[30]), .Z(n265)
         );
    VMW_AO22 U165 ( .A(\Out[0] ), .B(n322), .C(n323), .D(In1[0]), .Z(n311) );
    VMW_INV U180 ( .A(n270), .Z(n336) );
    VMW_FD \Out_reg[26]  ( .D(n338), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n349), .CP(Clk), .Q(\Out[15] ) );
    VMW_INV U192 ( .A(n294), .Z(n347) );
    VMW_FD \Out_reg[18]  ( .D(n346), .CP(Clk), .Q(\Out[18] ) );
    VMW_AOI211 U87 ( .A(n248), .B(In2[31]), .C(n263), .D(n245), .Z(n262) );
    VMW_AO22 U150 ( .A(\Out[23] ), .B(n322), .C(n323), .D(In1[23]), .Z(n281)
         );
    VMW_INV U177 ( .A(n264), .Z(n334) );
    VMW_FD \Out_reg[2]  ( .D(n362), .CP(Clk), .Q(\Out[2] ) );
    VMW_AND4 U125 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n328)
         );
    VMW_FD \Out_reg[11]  ( .D(n353), .CP(Clk), .Q(\Out[11] ) );
    VMW_AND2 U62 ( .A(DataIn[16]), .B(ScanEnable), .Z(ScanOut[16]) );
    VMW_FD \Out_reg[22]  ( .D(n342), .CP(Clk), .Q(\Out[22] ) );
    VMW_AND2 U65 ( .A(DataIn[13]), .B(ScanEnable), .Z(ScanOut[13]) );
    VMW_AOI211 U102 ( .A(n248), .B(In2[18]), .C(n293), .D(n245), .Z(n292) );
    VMW_AOI211 U105 ( .A(n248), .B(In2[15]), .C(n299), .D(n245), .Z(n298) );
    VMW_INV U189 ( .A(n288), .Z(n363) );
    VMW_FD \Out_reg[20]  ( .D(n344), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n351), .CP(Clk), .Q(\Out[13] ) );
    VMW_PULLUP U43 ( .Z(n365) );
    VMW_AND2 U50 ( .A(DataIn[28]), .B(ScanEnable), .Z(ScanOut[28]) );
    VMW_AND2 U59 ( .A(DataIn[19]), .B(ScanEnable), .Z(ScanOut[19]) );
    VMW_AOI211 U80 ( .A(n248), .B(In2[9]), .C(n249), .D(n245), .Z(n247) );
    VMW_AND4 U122 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(
        n319) );
    VMW_AO22 U139 ( .A(\Out[4] ), .B(n322), .C(n323), .D(In1[4]), .Z(n259) );
    VMW_AO22 U157 ( .A(\Out[17] ), .B(n322), .C(n323), .D(In1[17]), .Z(n295)
         );
    VMW_INV U170 ( .A(n250), .Z(n356) );
    VMW_FD \Out_reg[9]  ( .D(n355), .CP(Clk), .Q(\Out[9] ) );
    VMW_INV U195 ( .A(n300), .Z(n350) );
    VMW_FD \Out_reg[30]  ( .D(n334), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n364), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n335), .CP(Clk), .Q(\Out[29] ) );
    VMW_AND2 U77 ( .A(DataIn[1]), .B(ScanEnable), .Z(ScanOut[1]) );
    VMW_AOI211 U89 ( .A(n248), .B(In2[2]), .C(n267), .D(n245), .Z(n266) );
    VMW_INV U187 ( .A(n284), .Z(n343) );
    VMW_AOI211 U92 ( .A(n248), .B(In2[27]), .C(n273), .D(n245), .Z(n272) );
    VMW_AO22 U145 ( .A(\Out[28] ), .B(n322), .C(n323), .D(In1[28]), .Z(n271)
         );
    VMW_AO22 U162 ( .A(\Out[12] ), .B(n322), .C(n323), .D(In1[12]), .Z(n305)
         );
    VMW_INV U179 ( .A(n268), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n340), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n347), .CP(Clk), .Q(\Out[17] ) );
    VMW_AND4 U117 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n325)
         );
    VMW_FD \Out_reg[4]  ( .D(n360), .CP(Clk), .Q(\Out[4] ) );
    VMW_INV U200 ( .A(n310), .Z(n364) );
    VMW_AND2 U58 ( .A(DataIn[20]), .B(ScanEnable), .Z(ScanOut[20]) );
    VMW_AND4 U130 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(
        n315) );
    VMW_AO22 U138 ( .A(\Out[5] ), .B(n322), .C(n323), .D(In1[5]), .Z(n257) );
    VMW_INV U194 ( .A(n298), .Z(n349) );
    VMW_AND2 U64 ( .A(DataIn[14]), .B(ScanEnable), .Z(ScanOut[14]) );
    VMW_AOI211 U81 ( .A(n248), .B(In2[8]), .C(n251), .D(n245), .Z(n250) );
    VMW_AO22 U156 ( .A(\Out[18] ), .B(n322), .C(n323), .D(In1[18]), .Z(n293)
         );
    VMW_INV U171 ( .A(n252), .Z(n357) );
    VMW_AOI211 U104 ( .A(n248), .B(In2[16]), .C(n297), .D(n245), .Z(n296) );
    VMW_PULLDOWN U44 ( .Z(n368) );
    VMW_AND2 U51 ( .A(DataIn[27]), .B(ScanEnable), .Z(ScanOut[27]) );
    VMW_AND2 U76 ( .A(DataIn[2]), .B(ScanEnable), .Z(ScanOut[2]) );
    VMW_AND4 U116 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n324)
         );
    VMW_AND4 U123 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(
        n318) );
    VMW_AND2 U56 ( .A(DataIn[22]), .B(ScanEnable), .Z(ScanOut[22]) );
    VMW_AOI211 U88 ( .A(n248), .B(In2[30]), .C(n265), .D(n245), .Z(n264) );
    VMW_AOI211 U93 ( .A(n248), .B(In2[26]), .C(n275), .D(n245), .Z(n274) );
    VMW_AND4 U131 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(
        n314) );
    VMW_INV U201 ( .A(n332), .Z(Read2) );
    VMW_INV U178 ( .A(n266), .Z(n362) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 lte_43 ( .A(In1), 
        .B(In2), .LEQ(n367), .TC(n368), .LT_LE(n108) );
    VMW_AOI211 U94 ( .A(n248), .B(In2[25]), .C(n277), .D(n245), .Z(n276) );
    VMW_AO22 U143 ( .A(\Out[2] ), .B(n322), .C(n323), .D(In1[2]), .Z(n267) );
    VMW_AO22 U144 ( .A(\Out[29] ), .B(n322), .C(n323), .D(In1[29]), .Z(n269)
         );
    VMW_AO22 U163 ( .A(\Out[11] ), .B(n322), .C(n323), .D(In1[11]), .Z(n307)
         );
    VMW_INV U181 ( .A(n272), .Z(n337) );
    VMW_INV U186 ( .A(n282), .Z(n342) );
    VMW_AO22 U158 ( .A(\Out[16] ), .B(n322), .C(n323), .D(In1[16]), .Z(n297)
         );
    VMW_AO22 U164 ( .A(\Out[10] ), .B(n322), .C(n323), .D(In1[10]), .Z(n309)
         );
    VMW_AO22 U136 ( .A(\Out[7] ), .B(n322), .C(n323), .D(In1[7]), .Z(n253) );
    VMW_AND2 U71 ( .A(DataIn[7]), .B(ScanEnable), .Z(ScanOut[7]) );
    VMW_AOI211 U111 ( .A(n248), .B(In2[0]), .C(n311), .D(n245), .Z(n310) );
    VMW_AND4 U124 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(
        n317) );
    VMW_AND2 U63 ( .A(DataIn[15]), .B(ScanEnable), .Z(ScanOut[15]) );
    VMW_AND2 U78 ( .A(DataIn[0]), .B(ScanEnable), .Z(ScanOut[0]) );
    VMW_AOI211 U86 ( .A(n248), .B(In2[3]), .C(n261), .D(n245), .Z(n260) );
    VMW_AOI211 U103 ( .A(n248), .B(In2[17]), .C(n295), .D(n245), .Z(n294) );
    VMW_INV U188 ( .A(n286), .Z(n344) );
    VMW_AND4 U118 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n326)
         );
    VMW_AO22 U151 ( .A(\Out[22] ), .B(n322), .C(n323), .D(In1[22]), .Z(n283)
         );
    VMW_INV U176 ( .A(n262), .Z(n333) );
    VMW_INV U193 ( .A(n296), .Z(n348) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \Level1Out10[15] , \Level1Out33[24] , \Level1Out46[14] , 
        \Level1Out209[18] , \Level2Out246[28] , \Level4Out116[1] , 
        \Level1Out65[25] , \ScanLink213[0] , \Level2Out210[30] , 
        \Level2Out246[31] , \Level2Out8[24] , \Level2Out210[29] , 
        \Level1Out53[20] , \Level1Out70[11] , \ScanLink173[5] , 
        \ScanLink0[13] , \Level1Out11[2] , \ScanLink24[18] , \Level1Out26[10] , 
        \ScanLink50[8] , \ScanLink51[31] , \ScanLink72[19] , \ScanLink51[28] , 
        \ScanLink89[18] , \Level1Load154[0] , \ScanLink219[19] , 
        \Level1Out233[8] , \Level2Out78[2] , \Level2Out122[2] , 
        \Level4Out0[18] , \Level1Out182[8] , \ScanLink210[3] , 
        \Level2Out242[7] , \Level8Out248[7] , \Level1Out12[1] , 
        \Level64Out128[25] , \Level1Out26[23] , \ScanLink29[3] , 
        \Level1Out68[9] , \Level1Out137[9] , \ScanLink170[6] , 
        \Level8Out128[2] , \Level1Out70[22] , \Level4Out172[5] , 
        \ScanLink0[20] , \Level1Out10[26] , \Level1Out33[17] , 
        \Level1Out53[13] , \Level1Out46[27] , \Level1Out75[6] , 
        \Level4Out212[0] , \Level1Out65[16] , \Level2Out8[17] , 
        \Level1Load86[0] , \ScanLink117[1] , \Level1Out129[5] , 
        \Level1Out142[19] , \Level1Out161[31] , \Level64Out128[16] , 
        \Level1Out137[29] , \Level2Out178[19] , \Level2Out194[0] , 
        \ScanLink114[2] , \Level1Out114[18] , \Level1Out137[30] , 
        \Level1Out161[28] , \Level1Out249[0] , \ScanLink1[19] , 
        \Level1Out1[7] , \Level1Out2[23] , \ScanLink19[22] , \Level1Load28[0] , 
        \Level1Out76[5] , \ScanLink104[19] , \ScanLink127[31] , 
        \ScanLink127[28] , \ScanLink152[18] , \ScanLink171[30] , 
        \Level2Out146[6] , \Level8Out8[6] , \ScanLink171[29] , 
        \Level2Out226[3] , \ScanLink84[0] , \ScanLink212[26] , 
        \Level2Out52[15] , \ScanLink79[26] , \ScanLink181[24] , 
        \Level1Out187[5] , \ScanLink244[27] , \ScanLink194[10] , 
        \ScanLink231[17] , \ScanLink251[13] , \Level2Out64[10] , 
        \ScanLink224[23] , \ScanLink207[12] , \Level1Out228[9] , 
        \Level2Out32[11] , \Level1Out2[10] , \ScanLink9[6] , \ScanLink55[5] , 
        \ScanLink56[6] , \Level1Out241[12] , \Level1Out149[15] , 
        \Level1Out155[3] , \Level1Out191[25] , \Level1Out234[22] , 
        \Level2Out188[14] , \Level16Out144[15] , \Level32Out192[5] , 
        \Level16Out112[14] , \ScanLink168[4] , \Level1Out202[27] , 
        \ScanLink208[1] , \Level1Out217[13] , \Level2Out238[27] , 
        \Level1Out254[26] , \Level1Out184[11] , \Level1Out221[16] , 
        \Level1Out235[6] , \Level2Out106[25] , \Level4Out48[1] , 
        \Level1Out156[0] , \Level1Out199[9] , \Level32Out64[28] , 
        \Level2Load44[0] , \Level2Out150[24] , \Level32Out32[30] , 
        \Level32Out64[31] , \Level32Out32[29] , \ScanLink97[13] , 
        \Level1Out129[11] , \Level1Out236[5] , \Level2Out130[20] , 
        \Level2Out166[21] , \Level2Out244[9] , \ScanLink32[2] , 
        \Level1Out38[31] , \Level1Out38[28] , \ScanLink82[27] , 
        \ScanLink87[3] , \Level1Out184[6] , \ScanLink139[10] , 
        \ScanLink159[14] , \ScanLink176[8] , \Level2Out60[0] , 
        \Level1Out202[14] , \Level1Out131[7] , \Level2Out238[14] , 
        \Level1Out184[22] , \Level1Out221[25] , \Level1Out254[15] , 
        \Level1Out191[16] , \Level16Out144[26] , \Level1Out234[11] , 
        \Level1Out251[2] , \Level1Out6[21] , \ScanLink15[7] , \ScanLink19[11] , 
        \ScanLink79[15] , \ScanLink181[17] , \Level1Out217[20] , 
        \Level1Out241[21] , \Level2Out188[27] , \Level16Out112[27] , 
        \ScanLink224[10] , \Level4Out32[9] , \ScanLink194[23] , 
        \ScanLink207[21] , \ScanLink251[20] , \Level2Out64[23] , 
        \ScanLink212[15] , \Level2Out32[22] , \ScanLink231[24] , 
        \Level2Out52[26] , \ScanLink31[1] , \Level1Out73[8] , \ScanLink82[14] , 
        \ScanLink159[27] , \ScanLink244[14] , \Level8Out16[31] , 
        \Level8Out16[28] , \Level8Out40[29] , \Level1Out95[28] , 
        \ScanLink97[20] , \Level8Out40[30] , \ScanLink139[23] , 
        \Level2Out140[8] , \Level1Out49[2] , \ScanLink86[25] , 
        \Level1Out95[31] , \Level1Out129[22] , \Level2Out130[13] , 
        \Level2Out166[12] , \ScanLink128[26] , \Level1Out132[4] , 
        \Level1Out149[26] , \Level16Out48[19] , \Level128Out0[30] , 
        \Level1Out252[1] , \Level2Out106[16] , \Level2Out150[17] , 
        \Level128Out0[29] , \Level2Out20[2] , \Level1Out91[19] , 
        \ScanLink93[11] , \ScanLink148[22] , \Level2Out134[22] , 
        \Level1Out158[23] , \Level2Out0[0] , \Level2Out162[23] , 
        \Level1Out116[2] , \Level1Out138[27] , \Level2Out102[27] , 
        \Level2Out154[26] , \Level1Out49[30] , \Level1Out49[29] , 
        \Level1Out206[25] , \Level1Out85[8] , \Level16Out176[12] , 
        \ScanLink128[6] , \Level1Out250[24] , \Level4Out188[14] , 
        \Level1Out180[13] , \Level1Out225[14] , \Level1Out245[10] , 
        \Level8Load136[0] , \ScanLink16[4] , \Level1Out30[9] , 
        \ScanLink68[10] , \Level1Out98[7] , \Level1Out115[1] , 
        \Level1Out195[27] , \Level8Out184[31] , \Level1Out230[20] , 
        \ScanLink185[26] , \Level1Out213[11] , \ScanLink248[3] , 
        \Level8Out184[28] , \ScanLink255[11] , \Level2Out60[12] , 
        \ScanLink220[21] , \ScanLink135[9] , \ScanLink203[10] , 
        \Level2Out36[13] , \ScanLink216[24] , \Level2Out56[17] , 
        \ScanLink240[25] , \ScanLink71[3] , \Level1Out138[14] , 
        \ScanLink190[12] , \ScanLink235[15] , \Level2Out96[0] , 
        \ScanLink180[8] , \Level2Out102[14] , \Level2Out154[15] , 
        \Level1Out212[3] , \Level1Out158[10] , \Level1Out172[6] , 
        \Level2Out134[11] , \Level2Out162[10] , \Level2Out44[6] , 
        \ScanLink93[22] , \Level1Out2[4] , \ScanLink86[16] , \ScanLink128[15] , 
        \ScanLink148[11] , \ScanLink4[22] , \ScanLink4[11] , \Level1Out6[12] , 
        \ScanLink68[23] , \ScanLink216[17] , \Level2Out56[24] , 
        \ScanLink185[15] , \ScanLink190[21] , \ScanLink235[26] , 
        \ScanLink240[16] , \Level1Out195[14] , \ScanLink203[23] , 
        \ScanLink220[12] , \ScanLink231[8] , \Level2Out60[21] , 
        \ScanLink255[22] , \Level2Out36[20] , \Level1Out211[0] , 
        \Level1Out230[13] , \Level1Out245[23] , \Level1Load7[0] , 
        \ScanLink72[0] , \Level1Out171[5] , \Level1Out206[16] , 
        \Level1Out213[22] , \Level16Out176[21] , \Level1Out180[20] , 
        \Level1Out225[27] , \Level1Out250[17] , \Level4Out188[27] , 
        \Level1Out52[3] , \Level1Out110[30] , \Level1Out133[18] , 
        \Level1Out146[28] , \Level1Out110[29] , \ScanLink130[4] , 
        \Level1Out146[31] , \Level1Out165[19] , \Level8Out168[0] , 
        \ScanLink250[1] , \Level16Out32[27] , \Level16Out64[26] , 
        \Level128Out0[5] , \Level8Out208[5] , \Level1Out7[9] , \ScanLink13[9] , 
        \Level1Load70[0] , \Level1Out80[5] , \Level2Out202[5] , 
        \ScanLink100[31] , \ScanLink123[19] , \ScanLink156[29] , 
        \Level2Out162[0] , \Level1Out14[17] , \Level1Out22[12] , 
        \Level1Out51[0] , \Level1Out57[22] , \Level1Out74[13] , 
        \Level1Out83[6] , \ScanLink100[28] , \ScanLink156[30] , 
        \ScanLink175[18] , \Level2Out28[18] , \Level2Out38[0] , 
        \Level8Load16[0] , \Level4Out184[5] , \Level4Out236[6] , 
        \Level8Out216[9] , \ScanLink133[7] , \Level4Out4[6] , 
        \Level1Out37[26] , \Level1Out42[16] , \Level4Out156[3] , 
        \Level1Out61[27] , \ScanLink253[2] , \Level1Out174[8] , 
        \ScanLink186[6] , \Level4Out4[30] , \Level4Out4[29] , 
        \Level1Load213[0] , \Level2Out106[4] , \Level16Out64[15] , 
        \ScanLink154[0] , \Level8Out80[3] , \Level1Out209[2] , 
        \Level2Out42[8] , \ScanLink5[31] , \ScanLink5[28] , \Level1Out7[18] , 
        \Level1Out14[24] , \Level1Out35[4] , \Level1Out36[7] , 
        \Level1Out37[15] , \Level1Out169[7] , \Level16Out32[14] , 
        \ScanLink234[5] , \Level1Out42[25] , \Level2Load202[0] , 
        \Level2Out242[19] , \ScanLink20[30] , \Level1Out22[21] , 
        \Level1Out61[14] , \Level2Out214[18] , \Level4Out252[2] , 
        \ScanLink69[1] , \ScanLink157[3] , \Level2Out118[8] , 
        \Level1Out74[20] , \Level4Out132[7] , \Level1Out57[11] , 
        \ScanLink237[6] , \ScanLink20[29] , \ScanLink76[28] , 
        \Level1Out28[14] , \ScanLink55[19] , \ScanLink185[5] , 
        \ScanLink76[31] , \Level1Out212[28] , \Level8Load64[0] , 
        \Level8Out112[8] , \ScanLink193[1] , \Level1Out212[31] , 
        \Level1Out231[19] , \Level1Out244[30] , \Level2Out228[28] , 
        \Level16Out80[15] , \Level2Out228[31] , \ScanLink17[26] , 
        \ScanLink18[2] , \Level1Out20[3] , \Level1Out23[0] , \Level1Out48[10] , 
        \Level1Out244[29] , \Level2Out6[20] , \Level8Out216[13] , 
        \ScanLink69[29] , \Level2Out98[6] , \Level8Out240[12] , 
        \Level8Out88[25] , \ScanLink69[30] , \ScanLink92[31] , 
        \ScanLink141[7] , \Level4Out244[6] , \Level128Out128[13] , 
        \ScanLink202[30] , \ScanLink202[29] , \ScanLink221[18] , 
        \ScanLink254[31] , \ScanLink221[2] , \ScanLink254[28] , 
        \Level4Out124[3] , \ScanLink92[28] , \ScanLink142[4] , 
        \Level8Out96[7] , \Level1Out28[27] , \Level1Out47[4] , \ScanLink61[9] , 
        \Level1Out85[14] , \Level1Out202[9] , \ScanLink222[1] , 
        \Level4Out144[30] , \Level8Out128[11] , \Level1Out90[20] , 
        \ScanLink190[2] , \Level4Out112[28] , \Level2Out110[0] , 
        \Level4Out112[31] , \Level4Out144[29] , \ScanLink125[3] , 
        \Level2Out42[29] , \Level4Out220[2] , \Level2Out14[31] , 
        \Level2Out42[30] , \Level1Out48[23] , \Level1Out118[4] , 
        \Level2Out14[28] , \Level4Out140[7] , \Level8Out88[16] , 
        \Level1Out181[19] , \ScanLink191[18] , \ScanLink245[6] , 
        \Level2Out6[13] , \Level128Out128[20] , \Level2Out198[31] , 
        \Level2Out198[28] , \Level8Out160[8] , \Level8Out216[20] , 
        \Level8Out240[21] , \Level1Out95[2] , \Level4Out192[1] , 
        \Level1Out44[7] , \Level1Out59[8] , \Level1Out96[1] , 
        \Level1Out159[29] , \Level2Out116[19] , \Level16Out80[26] , 
        \Level2Out214[1] , \Level4Out52[29] , \Level1Out85[27] , 
        \Level1Out90[13] , \Level1Out159[30] , \Level2Out140[18] , 
        \Level2Out174[4] , \Level4Out52[30] , \Level1Out106[8] , 
        \Level8Out128[22] , \Level2Out30[8] , \ScanLink126[0] , 
        \ScanLink149[28] , \ScanLink21[23] , \ScanLink149[31] , 
        \ScanLink246[5] , \Level1Out38[1] , \ScanLink54[13] , 
        \Level1Out207[4] , \ScanLink209[16] , \Level8Load144[0] , 
        \ScanLink77[22] , \ScanLink34[17] , \ScanLink62[16] , 
        \Level1Out167[1] , \ScanLink41[27] , \ScanLink64[4] , \ScanLink147[9] , 
        \ScanLink188[0] , \Level4Out252[25] , \Level1Out152[25] , 
        \Level1Out219[17] , \Level2Out186[10] , \Level2Out236[23] , 
        \Level4Out204[24] , \Level2Out52[2] , \Level2Out108[2] , 
        \Level2Out200[26] , \Level4Out232[21] , \Level8Out208[18] , 
        \Level1Out127[15] , \Level1Out171[14] , \Level2Out168[25] , 
        \Level32Out192[14] , \Level1Out8[25] , \ScanLink17[15] , 
        \Level1Out23[18] , \Level1Out56[28] , \ScanLink67[7] , 
        \ScanLink101[11] , \Level1Out104[24] , \Level1Out111[10] , 
        \Level1Out164[20] , \Level1Out219[8] , \Level1Out132[21] , 
        \Level1Out147[11] , \Level2Out108[21] , \Level16Out192[21] , 
        \ScanLink174[21] , \Level2Out80[4] , \ScanLink122[20] , 
        \ScanLink157[10] , \ScanLink159[5] , \ScanLink142[24] , 
        \Level1Out204[7] , \ScanLink99[17] , \ScanLink137[14] , 
        \ScanLink114[25] , \ScanLink161[15] , \Level1Out164[2] , 
        \Level1Out219[24] , \ScanLink239[0] , \Level2Out84[21] , 
        \Level1Out56[31] , \Level1Out75[19] , \Level2Out186[23] , 
        \ScanLink62[25] , \ScanLink243[8] , \Level2Out8[8] , 
        \Level2Out200[15] , \Level2Out236[10] , \Level4Out232[12] , 
        \Level4Out252[16] , \Level4Out204[17] , \ScanLink21[10] , 
        \ScanLink34[24] , \ScanLink41[14] , \ScanLink54[20] , 
        \ScanLink209[25] , \ScanLink27[5] , \Level1Out42[9] , \ScanLink77[11] , 
        \ScanLink99[24] , \Level1Out103[5] , \ScanLink114[16] , 
        \ScanLink137[27] , \ScanLink142[17] , \Level2Out84[12] , 
        \Level1Out100[6] , \ScanLink101[22] , \ScanLink161[26] , 
        \ScanLink174[12] , \Level1Out111[23] , \ScanLink122[13] , 
        \ScanLink157[23] , \Level4Load228[0] , \Level1Out132[12] , 
        \Level1Out164[13] , \Level2Out36[6] , \Level2Out108[12] , 
        \Level16Out192[12] , \Level1Out104[17] , \Level1Out127[26] , 
        \Level1Out147[22] , \Level2Out168[16] , \Level1Out152[16] , 
        \Level8Out136[30] , \Level8Out160[28] , \ScanLink146[26] , 
        \Level1Out171[27] , \Level8Out136[29] , \Level32Out192[27] , 
        \Level8Out160[31] , \Level1Out27[29] , \ScanLink88[21] , 
        \ScanLink110[27] , \Level1Out124[0] , \ScanLink133[16] , 
        \ScanLink165[17] , \Level2Load36[0] , \Level2Out80[23] , 
        \ScanLink170[23] , \Level2Out236[9] , \Level1Out100[26] , 
        \ScanLink104[8] , \ScanLink105[13] , \Level1Out115[12] , 
        \ScanLink119[7] , \ScanLink126[22] , \ScanLink153[12] , 
        \Level1Out160[22] , \Level1Out244[5] , \Level1Out123[17] , 
        \Level1Out136[23] , \Level1Out143[13] , \Level4Out168[25] , 
        \Level4Out48[13] , \Level1Out156[27] , \Level2Out12[0] , 
        \Level4Out28[17] , \Level1Out175[16] , \Level4Out108[21] , 
        \Level2Out182[12] , \Level1Out52[19] , \Level1Out71[31] , 
        \Level2Out148[0] , \Level2Out252[25] , \ScanLink13[24] , 
        \Level1Out27[30] , \Level2Out204[24] , \Level4Out236[23] , 
        \ScanLink39[9] , \Level1Out71[28] , \Level1Out208[21] , 
        \Level2Out228[5] , \Level2Out232[21] , \Level4Out200[26] , 
        \ScanLink24[6] , \ScanLink30[15] , \ScanLink66[14] , \Level1Out127[3] , 
        \ScanLink45[25] , \Level2Out58[13] , \ScanLink25[21] , 
        \ScanLink218[20] , \ScanLink50[11] , \Level1Out247[6] , 
        \Level2Out38[17] , \ScanLink73[20] , \Level8Out8[10] , 
        \Level1Out78[3] , \Level1Out123[24] , \Level1Out156[14] , 
        \Level4Out28[24] , \Level1Out192[2] , \ScanLink200[9] , 
        \Level1Out8[16] , \ScanLink13[17] , \ScanLink25[12] , \ScanLink40[2] , 
        \ScanLink43[1] , \ScanLink88[12] , \ScanLink91[7] , \Level1Out100[15] , 
        \Level1Out175[25] , \ScanLink105[20] , \Level1Out115[21] , 
        \Level4Out108[12] , \Level1Out136[10] , \Level1Out160[11] , 
        \Level4Out168[16] , \Level4Out48[20] , \Level1Out143[20] , 
        \Level2Out76[4] , \Level1Out140[4] , \ScanLink170[10] , 
        \ScanLink126[11] , \ScanLink153[21] , \Level2Out132[8] , 
        \ScanLink50[22] , \ScanLink110[14] , \ScanLink133[25] , 
        \ScanLink146[15] , \Level1Out220[1] , \Level1Load188[0] , 
        \Level2Out80[10] , \ScanLink165[24] , \Level2Load228[0] , 
        \Level2Out38[24] , \ScanLink66[27] , \ScanLink73[13] , 
        \Level8Out8[23] , \Level1Out143[7] , \Level2Out68[8] , 
        \ScanLink30[26] , \ScanLink45[16] , \ScanLink218[13] , 
        \Level16Out0[6] , \ScanLink92[4] , \Level1Out223[2] , 
        \Level1Load239[0] , \Level2Out58[20] , \Level1Out191[1] , 
        \Level1Out208[12] , \Level2Out232[12] , \Level4Out40[9] , 
        \Level4Out200[15] , \Level2Out182[21] , \Level2Out252[16] , 
        \Level2Out204[17] , \ScanLink22[8] , \Level1Out60[1] , 
        \Level1Out81[16] , \Level1Out94[22] , \Level1Out128[31] , 
        \Level1Out128[28] , \Level4Out236[10] , \Level2Out112[28] , 
        \Level2Out144[30] , \Level4Out56[18] , \Level2Out144[29] , 
        \Level2Out150[2] , \Level2Out112[31] , \ScanLink102[6] , 
        \ScanLink138[29] , \Level2Out182[4] , \Level2Out230[7] , 
        \ScanLink138[30] , \Level1Out63[2] , \ScanLink195[29] , 
        \Level2Out10[19] , \Level2Out46[18] , \Level4Out164[1] , 
        \ScanLink101[5] , \ScanLink195[30] , \Level4Out204[4] , 
        \Level1Out185[28] , \Level2Out2[22] , \Level4Out228[28] , 
        \Level1Out39[22] , \Level1Out185[31] , \Level4Out228[31] , 
        \ScanLink58[0] , \Level1Out59[26] , \Level8Out224[14] , 
        \ScanLink97[9] , \Level1Load126[0] , \Level1Out241[8] , 
        \Level1Out81[25] , \ScanLink96[19] , \ScanLink166[2] , 
        \ScanLink206[7] , \Level2Out134[6] , \Level4Out116[19] , 
        \ScanLink0[30] , \ScanLink1[23] , \ScanLink1[10] , \Level1Out3[30] , 
        \ScanLink4[3] , \ScanLink7[0] , \Level1Out94[11] , \Level1Out189[3] , 
        \Level2Out254[3] , \Level4Out140[18] , \Level32Out0[31] , 
        \Level32Out0[28] , \Level64Out128[7] , \Level1Out3[29] , 
        \Level1Out59[15] , \Level1Out145[9] , \Level8Out224[27] , 
        \Level1Out216[19] , \Level1Out235[31] , \Level2Load98[0] , 
        \Level1Out240[18] , \Level1Out3[20] , \ScanLink5[21] , \ScanLink5[12] , 
        \Level1Out15[14] , \ScanLink18[31] , \ScanLink18[28] , 
        \Level1Out39[11] , \ScanLink89[5] , \Level1Out235[28] , 
        \Level2Out2[11] , \Level1Out158[6] , \Level4Out100[5] , 
        \ScanLink205[4] , \Level1Out60[24] , \ScanLink165[1] , 
        \ScanLink206[18] , \ScanLink225[30] , \ScanLink225[29] , 
        \Level1Out238[3] , \ScanLink250[19] , \ScanLink21[19] , 
        \Level1Out23[11] , \Level1Out36[25] , \Level1Out43[15] , 
        \Level1Out41[3] , \Level1Out56[21] , \ScanLink243[1] , 
        \Level2Out236[19] , \ScanLink54[29] , \Level1Load63[0] , 
        \Level1Out75[10] , \Level4Load156[0] , \Level8Out208[22] , 
        \ScanLink123[4] , \Level2Out8[1] , \ScanLink54[30] , \ScanLink77[18] , 
        \Level8Out96[14] , \Level1Out90[6] , \Level1Out93[5] , 
        \Level2Out28[3] , \Level2Out172[3] , \Level2Out212[6] , 
        \ScanLink240[2] , \Level1Out9[6] , \Level1Out42[0] , \ScanLink120[7] , 
        \Level8Out136[20] , \Level8Out160[21] , \Level1Out167[8] , 
        \Level1Load200[0] , \Level1Out15[27] , \Level1Out23[22] , 
        \Level1Out38[8] , \ScanLink195[6] , \Level8Out96[27] , 
        \Level1Out56[12] , \ScanLink227[5] , \Level2Out186[19] , 
        \Level4Out64[6] , \Level4Out232[31] , \Level1Out75[23] , 
        \ScanLink79[2] , \Level4Out232[28] , \Level8Out208[11] , 
        \Level1Out25[7] , \Level1Out36[16] , \Level1Out60[17] , 
        \ScanLink188[9] , \ScanLink147[0] , \Level1Out43[26] , 
        \Level1Out111[19] , \Level1Out132[31] , \Level1Out164[29] , 
        \Level2Out108[31] , \Level16Out192[31] , \Level1Out132[28] , 
        \Level1Out147[18] , \Level1Out164[30] , \Level2Out108[28] , 
        \Level16Out192[28] , \Level1Out179[4] , \ScanLink224[6] , 
        \Level8Out160[12] , \ScanLink7[9] , \Level1Out7[22] , \Level1Out26[4] , 
        \ScanLink69[13] , \ScanLink101[18] , \ScanLink122[30] , 
        \ScanLink144[3] , \ScanLink174[28] , \Level1Out219[1] , 
        \Level8Out136[13] , \ScanLink239[9] , \Level2Out84[31] , 
        \Level2Out116[7] , \Level2Out84[28] , \ScanLink122[29] , 
        \ScanLink157[19] , \ScanLink174[31] , \ScanLink196[5] , 
        \ScanLink241[26] , \Level2Out74[25] , \Level128Out128[30] , 
        \Level1Out88[4] , \ScanLink184[25] , \ScanLink191[11] , 
        \ScanLink202[13] , \ScanLink217[27] , \ScanLink234[16] , 
        \Level2Out22[24] , \Level128Out128[29] , \Level2Out42[20] , 
        \ScanLink221[22] , \ScanLink254[12] , \Level2Out14[21] , 
        \Level1Out105[2] , \Level2Out228[12] , \Level4Out192[8] , 
        \Level1Out212[12] , \Level8Out200[4] , \Level1Out244[13] , 
        \Level1Out7[11] , \Level1Out48[19] , \Level1Out59[1] , 
        \Level1Out96[8] , \Level1Out106[1] , \ScanLink138[5] , 
        \Level1Out194[24] , \Level1Out231[23] , \Level1Out251[27] , 
        \Level8Out240[31] , \Level1Out139[24] , \Level1Out181[10] , 
        \Level1Out207[26] , \Level1Out224[17] , \Level2Out198[21] , 
        \Level8Out160[1] , \Level8Out216[29] , \Level8Out240[28] , 
        \Level2Out120[15] , \Level2Out248[16] , \Level4Out112[12] , 
        \Level8Out216[30] , \Level4Out32[24] , \Level4Out64[25] , 
        \Level4Out144[13] , \Level1Out159[20] , \Level2Out176[14] , 
        \Level4Out124[17] , \Level2Out116[10] , \Level2Out214[8] , 
        \Level4Out52[20] , \ScanLink62[3] , \ScanLink87[26] , \ScanLink92[12] , 
        \ScanLink149[21] , \Level2Out140[11] , \Level4Out172[16] , 
        \ScanLink126[9] , \ScanLink129[25] , \Level2Out30[1] , 
        \Level1Out181[23] , \Level1Out224[24] , \Level1Out251[14] , 
        \Level2Out6[29] , \Level1Out207[15] , \Level2Out248[25] , 
        \Level4Load96[0] , \Level1Out161[6] , \Level2Out6[30] , 
        \Level2Out198[12] , \ScanLink193[8] , \Level1Out194[17] , 
        \Level1Out212[21] , \Level1Out231[10] , \Level2Out228[21] , 
        \Level16Out80[7] , \Level1Out201[3] , \Level1Out244[20] , 
        \Level8Out104[5] , \Level1Out19[3] , \Level1Out23[9] , 
        \ScanLink69[20] , \ScanLink184[16] , \ScanLink202[20] , 
        \Level8Out88[2] , \ScanLink221[11] , \Level2Out42[13] , 
        \ScanLink254[21] , \Level2Out14[12] , \ScanLink191[22] , 
        \ScanLink234[25] , \ScanLink58[9] , \ScanLink61[0] , \ScanLink87[15] , 
        \ScanLink217[14] , \ScanLink241[15] , \Level2Out74[16] , 
        \Level2Out22[17] , \ScanLink222[8] , \Level1Out90[30] , 
        \ScanLink92[21] , \ScanLink129[16] , \ScanLink149[12] , 
        \Level2Out54[5] , \Level4Out52[13] , \Level1Out159[13] , 
        \Level1Out162[5] , \Level2Out116[23] , \Level4Out124[24] , 
        \Level2Out110[9] , \Level2Out140[22] , \Level4Out172[25] , 
        \ScanLink83[24] , \Level1Out90[29] , \Level1Out139[17] , 
        \Level1Out202[0] , \Level2Out120[26] , \Level4Out64[16] , 
        \Level8Out128[18] , \Level4Out112[21] , \Level2Out86[3] , 
        \Level2Out176[27] , \Level4Out144[20] , \Level4Out32[17] , 
        \ScanLink97[0] , \ScanLink158[17] , \Level2Out70[3] , \ScanLink96[10] , 
        \ScanLink138[13] , \Level1Out128[12] , \Level1Out194[5] , 
        \Level2Out112[12] , \Level4Out120[15] , \Level4Out56[22] , 
        \Level1Out39[18] , \ScanLink45[6] , \Level1Out94[18] , 
        \Level1Out226[6] , \Level4Out176[14] , \Level32Out0[21] , 
        \Level2Out124[17] , \Level2Out144[13] , \Level4Out116[10] , 
        \Level4Out60[27] , \Level1Out146[3] , \Level1Out148[16] , 
        \Level4Out36[26] , \ScanLink178[7] , \Level1Out255[25] , 
        \Level2Out172[16] , \Level4Out140[11] , \Level4Out228[12] , 
        \Level2Out2[18] , \Level1Out185[12] , \Level1Out220[15] , 
        \Level1Out225[5] , \Level8Out120[3] , \Level1Out203[24] , 
        \Level1Out145[0] , \Level1Out216[10] , \ScanLink218[2] , 
        \Level8Out240[6] , \Level1Out3[13] , \ScanLink18[21] , \ScanLink46[5] , 
        \Level1Out240[11] , \ScanLink78[25] , \ScanLink165[8] , 
        \Level1Out190[26] , \Level1Out235[21] , \Level4Out248[16] , 
        \ScanLink206[11] , \Level2Out46[22] , \ScanLink180[27] , 
        \ScanLink225[20] , \ScanLink250[10] , \Level2Out10[23] , 
        \ScanLink18[12] , \ScanLink21[2] , \ScanLink94[3] , \ScanLink195[13] , 
        \Level1Out197[6] , \ScanLink245[24] , \Level2Out70[27] , 
        \ScanLink213[25] , \ScanLink230[14] , \Level2Out26[26] , 
        \Level4Load60[0] , \Level1Out122[7] , \Level1Out128[21] , 
        \Level1Out148[25] , \Level1Out242[2] , \Level2Out124[24] , 
        \Level4Out60[14] , \Level2Out172[25] , \Level4Out116[23] , 
        \Level4Out36[15] , \Level4Out140[22] , \Level4Out56[11] , 
        \Level2Out112[21] , \Level4Out120[26] , \Level2Out144[20] , 
        \Level4Out176[27] , \Level1Out60[8] , \ScanLink138[20] , 
        \Level32Out0[12] , \Level2Out14[7] , \ScanLink83[17] , 
        \ScanLink96[23] , \ScanLink158[24] , \ScanLink195[20] , 
        \ScanLink230[27] , \ScanLink78[16] , \ScanLink180[14] , 
        \ScanLink206[22] , \ScanLink213[16] , \ScanLink245[17] , 
        \Level2Out70[14] , \Level2Out26[15] , \ScanLink225[13] , 
        \Level2Out10[10] , \Level2Out46[11] , \Level1Out190[15] , 
        \Level1Out216[23] , \ScanLink250[23] , \Level4Out164[8] , 
        \Level1Out235[12] , \Level4Out248[25] , \Level8Out0[7] , 
        \Level1Out241[1] , \ScanLink22[1] , \Level1Out185[21] , 
        \Level1Out240[22] , \Level8Out144[7] , \Level1Out220[26] , 
        \Level1Out255[16] , \Level4Out228[21] , \Level1Out115[31] , 
        \Level1Out115[28] , \Level1Out121[4] , \Level1Out203[17] , 
        \Level8Out224[2] , \Level1Out143[30] , \ScanLink160[5] , 
        \Level4Out48[30] , \Level8Out152[26] , \Level1Out160[18] , 
        \Level8Out104[27] , \Level1Out136[19] , \Level1Out143[29] , 
        \Level4Out48[29] , \ScanLink200[0] , \ScanLink1[7] , \ScanLink2[4] , 
        \ScanLink105[29] , \Level1Load147[0] , \Level1Out220[8] , 
        \Level2Out80[19] , \Level2Out252[4] , \ScanLink43[8] , 
        \ScanLink105[30] , \ScanLink153[31] , \ScanLink170[19] , 
        \ScanLink126[18] , \Level2Out132[1] , \ScanLink153[28] , 
        \Level2Out58[30] , \Level2Out68[1] , \Level2Out58[29] , 
        \Level1Out11[16] , \Level1Out27[13] , \Level1Out52[23] , 
        \Level4Out92[6] , \Level2Out182[28] , \Level1Out64[26] , 
        \Level1Out71[12] , \ScanLink163[6] , \Level2Out182[31] , 
        \Level4Out236[19] , \Level2Load156[0] , \Level1Out32[27] , 
        \Level1Out47[17] , \Level4Out40[0] , \ScanLink88[31] , 
        \ScanLink88[28] , \Level1Out191[8] , \ScanLink203[3] , 
        \Level32Out32[3] , \Level2Out236[0] , \Level1Out124[9] , 
        \Level2Out156[5] , \Level2Out12[9] , \Level4Out108[31] , 
        \Level1Out2[19] , \Level1Out11[25] , \Level1Out66[6] , 
        \ScanLink104[1] , \Level4Out108[28] , \Level1Out139[6] , 
        \Level2Out184[3] , \Level8Out104[14] , \Level8Out152[15] , 
        \ScanLink25[31] , \ScanLink25[28] , \Level1Out27[20] , 
        \Level1Out32[14] , \Level1Out64[15] , \Level1Out208[31] , 
        \Level2Out232[31] , \ScanLink107[2] , \Level2Out232[28] , 
        \Level1Out47[24] , \Level1Out208[28] , \Level1Out65[5] , 
        \ScanLink39[0] , \Level1Out52[10] , \Level4Out24[4] , 
        \Level1Out71[21] , \Level1Load95[0] , \Level2Out148[9] , 
        \ScanLink50[18] , \ScanLink73[30] , \ScanLink73[29] , 
        \Level1Out217[30] , \ScanLink218[30] , \Level8Out8[19] , 
        \ScanLink218[29] , \Level1Out234[18] , \Level1Out241[28] , 
        \Level1Out9[26] , \ScanLink12[27] , \Level1Out14[6] , \Level1Out17[5] , 
        \ScanLink19[18] , \Level1Out38[21] , \Level1Out58[25] , 
        \Level1Out217[29] , \Level1Out241[31] , \ScanLink111[6] , 
        \ScanLink31[8] , \Level1Out70[2] , \Level1Out73[1] , \ScanLink97[29] , 
        \ScanLink207[31] , \ScanLink224[19] , \ScanLink207[28] , 
        \ScanLink251[29] , \Level4Out32[0] , \ScanLink251[30] , 
        \Level2Load124[0] , \Level1Out80[15] , \ScanLink97[30] , 
        \ScanLink112[5] , \Level1Load135[0] , \Level2Out192[7] , 
        \Level2Out220[4] , \Level8Out16[21] , \Level8Out40[20] , 
        \Level32Out32[13] , \Level32Out64[12] , \Level128Out0[20] , 
        \Level1Out252[8] , \Level2Out140[1] , \Level1Out95[21] , 
        \Level2Out64[19] , \Level16Out48[10] , \Level1Out38[12] , 
        \ScanLink84[9] , \ScanLink175[2] , \Level1Out228[0] , 
        \Level2Out32[18] , \Level1Out148[5] , \Level4Out56[4] , 
        \ScanLink194[19] , \ScanLink215[7] , \Level1Out58[16] , 
        \ScanLink99[6] , \Level1Out184[18] , \Level4Out84[2] , 
        \Level1Out80[26] , \Level1Out95[12] , \ScanLink208[8] , 
        \Level1Out129[18] , \Level2Out130[30] , \Level2Out130[29] , 
        \Level2Out166[31] , \Level2Out244[0] , \Level16Out48[23] , 
        \Level1Out156[9] , \Level1Out199[0] , \Level2Out166[28] , 
        \Level4Out48[8] , \Level32Out64[21] , \Level2Out124[5] , 
        \ScanLink176[1] , \Level8Out40[13] , \Level32Out32[20] , 
        \Level128Out0[13] , \Level2Out60[9] , \ScanLink24[22] , 
        \ScanLink48[3] , \ScanLink139[19] , \ScanLink216[4] , 
        \Level8Out16[12] , \Level1Out68[0] , \ScanLink72[23] , 
        \ScanLink31[16] , \ScanLink51[12] , \Level8Out152[3] , \ScanLink34[5] , 
        \ScanLink44[26] , \ScanLink219[23] , \ScanLink67[17] , 
        \Level8Out232[6] , \ScanLink117[8] , \Level1Out137[0] , 
        \Level1Out209[22] , \Level2Out196[25] , \Level2Out238[6] , 
        \Level2Out246[12] , \Level2Out210[13] , \Level4Out84[14] , 
        \Level4Out212[9] , \Level2Out158[3] , \Level1Out174[15] , 
        \Level2Out226[16] , \Level4Load12[0] , \Level4Out192[27] , 
        \ScanLink0[29] , \Level1Out101[25] , \Level1Out157[24] , 
        \Level1Out249[9] , \Level2Out118[14] , \ScanLink4[18] , 
        \Level1Out4[3] , \Level1Out7[0] , \Level1Out9[15] , \ScanLink37[6] , 
        \Level1Load49[0] , \Level1Out122[14] , \Level1Out137[20] , 
        \Level1Out142[10] , \Level2Out178[10] , \Level2Out194[9] , 
        \ScanLink89[22] , \ScanLink109[4] , \Level1Out114[11] , 
        \Level1Out161[21] , \ScanLink127[21] , \ScanLink152[11] , 
        \ScanLink171[20] , \Level1Out254[6] , \Level4Out0[22] , 
        \ScanLink104[10] , \Level2Out94[14] , \ScanLink111[24] , 
        \Level1Out134[3] , \ScanLink164[14] , \ScanLink147[25] , 
        \Level1Out53[30] , \Level1Out70[18] , \ScanLink132[15] , 
        \ScanLink12[14] , \Level1Out26[19] , \Level1Out53[29] , 
        \Level4Out192[14] , \ScanLink31[25] , \ScanLink44[15] , 
        \ScanLink82[7] , \Level1Out181[2] , \Level1Out209[11] , 
        \Level2Out226[25] , \Level4Out116[8] , \Level2Out196[16] , 
        \Level2Out246[21] , \ScanLink213[9] , \Level2Out210[20] , 
        \Level4Out84[27] , \ScanLink219[10] , \ScanLink67[24] , 
        \Level1Out233[1] , \Level8Out136[7] , \Level1Out12[8] , 
        \ScanLink24[11] , \ScanLink50[1] , \ScanLink51[21] , \ScanLink72[10] , 
        \Level1Out153[4] , \ScanLink53[2] , \ScanLink111[17] , 
        \ScanLink127[12] , \ScanLink132[26] , \ScanLink164[27] , 
        \ScanLink147[16] , \Level1Out230[2] , \ScanLink152[22] , 
        \Level4Out0[11] , \ScanLink89[11] , \ScanLink104[23] , 
        \Level2Out94[27] , \Level1Out150[7] , \ScanLink171[13] , 
        \Level4Out108[4] , \Level1Out137[13] , \Level1Out142[23] , 
        \Level2Out66[7] , \Level2Out178[23] , \ScanLink77[4] , \ScanLink81[4] , 
        \Level1Out101[16] , \Level1Out114[22] , \Level1Out161[12] , 
        \Level1Out174[26] , \ScanLink98[14] , \Level1Out122[27] , 
        \Level1Out157[17] , \Level1Out182[1] , \Level2Out118[27] , 
        \ScanLink115[26] , \ScanLink160[16] , \Level1Out174[1] , 
        \ScanLink143[27] , \ScanLink229[3] , \ScanLink100[12] , 
        \ScanLink123[23] , \ScanLink136[17] , \ScanLink149[6] , 
        \ScanLink156[13] , \ScanLink175[22] , \Level1Out214[4] , 
        \Level4Out4[20] , \Level2Out90[7] , \Level1Out110[13] , 
        \Level1Out133[22] , \Level1Out146[12] , \Level2Out90[16] , 
        \Level1Out165[23] , \Level1Out170[17] , \Level1Out22[31] , 
        \Level1Out105[27] , \ScanLink154[9] , \Level1Out126[16] , 
        \Level1Out153[26] , \Level2Out42[1] , \Level2Out118[1] , 
        \Level4Out196[25] , \Level1Out22[28] , \ScanLink69[8] , 
        \Level1Out74[29] , \Level2Out222[14] , \Level1Out57[18] , 
        \Level1Out218[14] , \Level1Out74[30] , \Level2Out192[27] , 
        \Level2Out214[11] , \Level2Out242[10] , \Level4Out80[16] , 
        \ScanLink16[25] , \ScanLink35[14] , \ScanLink198[3] , \ScanLink40[24] , 
        \ScanLink74[7] , \Level2Out28[22] , \ScanLink20[20] , \Level1Out28[2] , 
        \ScanLink63[15] , \ScanLink76[21] , \Level1Out177[2] , 
        \Level2Out48[26] , \ScanLink55[10] , \ScanLink208[15] , 
        \Level16Out96[3] , \Level1Out217[7] , \Level8Out112[1] , 
        \Level1Out105[14] , \Level1Out126[25] , \Level1Out170[24] , 
        \Level1Out153[15] , \ScanLink250[8] , \Level1Out110[20] , 
        \Level1Out133[11] , \Level1Out146[21] , \Level2Out26[5] , 
        \ScanLink123[10] , \Level1Out165[10] , \Level2Out162[9] , 
        \Level8Out168[9] , \ScanLink156[20] , \Level4Out4[13] , 
        \Level1Out6[31] , \Level1Out6[28] , \ScanLink10[3] , \ScanLink13[0] , 
        \ScanLink55[23] , \ScanLink76[12] , \ScanLink98[27] , 
        \ScanLink100[21] , \Level1Out110[5] , \ScanLink175[11] , 
        \Level2Out90[25] , \Level4Out148[6] , \ScanLink115[15] , 
        \ScanLink136[24] , \ScanLink160[25] , \Level4Out228[3] , 
        \ScanLink143[14] , \Level2Out6[7] , \Level1Out113[6] , 
        \ScanLink208[26] , \Level8Out216[0] , \Level2Out48[15] , 
        \Level1Load11[0] , \ScanLink16[16] , \ScanLink20[13] , 
        \ScanLink35[27] , \ScanLink40[17] , \Level2Out28[11] , 
        \ScanLink63[26] , \Level8Out176[5] , \Level2Out38[9] , 
        \Level1Out30[0] , \Level1Out51[9] , \Level1Out218[27] , 
        \Level2Out192[14] , \Level2Out242[23] , \Level16Out192[2] , 
        \Level2Out214[22] , \Level4Out80[25] , \Level4Out196[16] , 
        \Level1Out84[17] , \Level1Out91[23] , \Level2Out100[3] , 
        \Level2Out222[27] , \Level2Out134[18] , \Level1Out158[19] , 
        \Level2Out162[19] , \Level2Out96[9] , \ScanLink180[1] , 
        \ScanLink232[2] , \Level1Out33[3] , \ScanLink148[18] , 
        \ScanLink152[7] , \Level8Out24[26] , \Level8Out72[27] , 
        \ScanLink151[4] , \ScanLink190[31] , \ScanLink231[1] , 
        \Level2Out36[30] , \Level4Out72[2] , \Level2Out36[29] , 
        \Level2Out60[28] , \Level2Out60[31] , \ScanLink190[28] , 
        \Level2Out88[5] , \Level4Load124[0] , \Level1Out49[13] , 
        \Level1Out180[30] , \Level1Out180[29] , \Level16Out176[28] , 
        \Level16Out176[31] , \Level1Out29[17] , \ScanLink72[9] , 
        \ScanLink183[2] , \Level1Out211[9] , \Level8Out184[12] , 
        \Level1Out54[4] , \ScanLink93[18] , \Level8Out72[14] , 
        \ScanLink136[3] , \ScanLink256[6] , \Level8Out24[15] , 
        \Level8Load248[0] , \Level1Out84[24] , \Level2Out164[7] , 
        \Level1Out86[2] , \Level1Out91[10] , \Level2Out0[9] , 
        \Level2Out204[2] , \Level1Out230[29] , \Level1Out245[19] , 
        \ScanLink7[4] , \Level1Out29[24] , \Level1Out39[26] , 
        \Level1Out49[20] , \Level1Out115[8] , \Level8Out184[21] , 
        \Level1Out213[18] , \Level1Out230[30] , \Level1Out57[7] , 
        \ScanLink68[19] , \Level1Out85[1] , \Level1Out108[7] , 
        \Level4Out16[6] , \ScanLink255[18] , \ScanLink255[5] , 
        \Level32Out64[5] , \Level1Out59[22] , \ScanLink135[0] , 
        \ScanLink203[19] , \ScanLink220[28] , \Level1Out190[18] , 
        \ScanLink220[31] , \Level4Out248[31] , \Level4Out248[28] , 
        \Level8Out224[10] , \Level1Out39[15] , \Level1Out60[5] , 
        \Level1Out63[6] , \ScanLink101[1] , \Level1Out121[9] , 
        \Level2Out2[26] , \Level2Out26[18] , \Level4Out204[0] , 
        \Level2Out70[19] , \ScanLink180[19] , \Level4Out164[5] , 
        \ScanLink78[31] , \ScanLink78[28] , \Level1Out81[12] , 
        \Level1Load90[0] , \ScanLink102[2] , \Level2Out182[0] , 
        \Level1Out148[28] , \ScanLink158[30] , \ScanLink158[29] , 
        \Level2Out172[28] , \Level2Out230[3] , \Level2Out124[30] , 
        \Level4Out36[18] , \Level2Out172[31] , \Level4Out60[19] , 
        \Level1Out94[26] , \Level1Out148[31] , \Level2Out124[29] , 
        \Level2Out150[6] , \ScanLink165[5] , \Level1Out238[7] , 
        \Level1Out158[2] , \ScanLink213[28] , \ScanLink245[30] , 
        \ScanLink245[29] , \Level4Out100[1] , \ScanLink205[0] , 
        \ScanLink213[31] , \ScanLink230[19] , \ScanLink46[8] , 
        \Level1Load142[0] , \Level1Out203[30] , \Level1Out203[29] , 
        \Level1Out255[31] , \Level1Out220[18] , \Level1Out255[28] , 
        \Level2Out2[15] , \Level1Out225[8] , \ScanLink89[1] , 
        \Level64Out128[3] , \Level1Out59[11] , \Level8Out224[23] , 
        \Level1Out94[15] , \Level2Out254[7] , \Level4Out120[18] , 
        \Level4Out176[19] , \Level16Load192[0] , \ScanLink4[7] , 
        \ScanLink58[4] , \Level1Out81[21] , \Level1Out189[7] , 
        \Level2Out134[2] , \ScanLink83[30] , \ScanLink83[29] , 
        \ScanLink166[6] , \Level1Out194[8] , \ScanLink206[3] , \ScanLink0[17] , 
        \ScanEnable[0] , \ScanLink2[9] , \Level1Out8[21] , \Level1Out11[31] , 
        \ScanLink13[20] , \ScanLink24[2] , \ScanLink25[25] , \ScanLink73[24] , 
        \Level1Out78[7] , \Level8Out8[14] , \ScanLink30[11] , \ScanLink50[15] , 
        \Level1Out247[2] , \Level2Out38[13] , \ScanLink45[21] , 
        \Level2Out58[17] , \ScanLink218[24] , \Level1Out32[19] , 
        \ScanLink66[10] , \Level1Out127[7] , \Level2Out232[25] , 
        \Level4Out200[22] , \Level1Out11[28] , \Level1Out47[29] , 
        \Level1Out208[25] , \Level2Out228[1] , \Level1Out65[8] , 
        \Level1Out47[30] , \Level1Out64[18] , \Level2Out148[4] , 
        \Level4Out236[27] , \Level1Out8[12] , \ScanLink27[1] , 
        \ScanLink88[25] , \Level1Out100[22] , \Level1Out175[12] , 
        \Level2Out182[16] , \Level2Out204[20] , \Level4Out24[9] , 
        \Level2Out252[21] , \Level4Out108[25] , \Level1Out115[16] , 
        \Level1Out123[13] , \Level1Out156[23] , \Level2Out12[4] , 
        \Level4Out28[13] , \Level1Out136[27] , \Level1Out143[17] , 
        \Level4Out48[17] , \Level8Out104[19] , \Level1Out160[26] , 
        \Level8Out152[18] , \ScanLink119[3] , \ScanLink153[16] , 
        \Level4Out168[21] , \ScanLink126[26] , \ScanLink170[27] , 
        \Level1Out244[1] , \ScanLink105[17] , \ScanLink110[23] , 
        \Level1Out124[4] , \ScanLink165[13] , \ScanLink146[22] , 
        \Level2Out80[27] , \Level2Out156[8] , \ScanLink133[12] , 
        \Level2Out204[13] , \Level4Out236[14] , \ScanLink13[13] , 
        \ScanLink30[22] , \ScanLink45[12] , \ScanLink92[0] , \Level1Out191[5] , 
        \Level1Out208[16] , \Level2Out182[25] , \Level2Out252[12] , 
        \Level2Out232[16] , \Level4Out200[11] , \ScanLink218[17] , 
        \ScanLink66[23] , \Level1Out223[6] , \Level16Out0[2] , 
        \Level2Out58[24] , \ScanLink25[16] , \ScanLink40[6] , \ScanLink50[26] , 
        \ScanLink73[17] , \Level1Out143[3] , \Level8Out8[27] , 
        \Level2Out38[20] , \ScanLink43[5] , \ScanLink110[10] , 
        \ScanLink126[15] , \ScanLink133[21] , \ScanLink165[20] , 
        \Level2Out80[14] , \Level2Out252[9] , \ScanLink146[11] , 
        \Level1Out220[5] , \ScanLink153[25] , \ScanLink105[24] , 
        \ScanLink4[26] , \ScanLink4[15] , \Level1Out14[13] , \Level1Out15[19] , 
        \ScanLink17[22] , \Level1Out26[9] , \ScanLink67[3] , \ScanLink88[16] , 
        \Level1Out140[0] , \ScanLink170[14] , \Level2Load52[0] , 
        \ScanLink91[3] , \Level1Out100[11] , \Level1Out115[25] , 
        \Level1Out136[14] , \Level4Out48[24] , \Level1Out143[24] , 
        \Level2Out76[0] , \ScanLink160[8] , \Level1Out160[15] , 
        \Level4Out168[12] , \Level1Out175[21] , \Level4Out108[16] , 
        \ScanLink99[13] , \Level1Out123[20] , \Level1Out156[10] , 
        \Level1Out192[6] , \Level4Out28[20] , \ScanLink114[21] , 
        \ScanLink161[11] , \Level1Out164[6] , \ScanLink239[4] , 
        \Level2Out84[25] , \ScanLink142[20] , \ScanLink101[15] , 
        \ScanLink122[24] , \ScanLink137[10] , \ScanLink157[14] , 
        \ScanLink159[1] , \ScanLink174[25] , \ScanLink196[8] , 
        \Level1Out204[3] , \Level2Out80[0] , \Level1Out104[20] , 
        \Level1Out111[14] , \Level1Out132[25] , \Level1Out147[15] , 
        \Level1Out179[9] , \Level2Out108[25] , \Level16Out192[25] , 
        \Level1Out164[24] , \Level1Out171[10] , \Level32Out192[10] , 
        \Level1Out152[21] , \Level2Out52[6] , \ScanLink34[13] , 
        \Level1Out127[11] , \ScanLink188[4] , \Level1Out219[13] , 
        \ScanLink227[8] , \Level2Out108[6] , \Level2Out168[21] , 
        \Level2Out186[14] , \Level2Out200[22] , \Level4Out232[25] , 
        \Level2Out236[27] , \Level4Out204[20] , \Level4Out252[21] , 
        \ScanLink41[23] , \ScanLink64[0] , \ScanLink17[11] , \ScanLink21[27] , 
        \Level1Out38[5] , \ScanLink62[12] , \ScanLink77[26] , 
        \Level1Out167[5] , \ScanLink21[14] , \ScanLink54[24] , 
        \ScanLink54[17] , \Level1Out207[0] , \ScanLink209[12] , 
        \ScanLink77[15] , \ScanLink99[20] , \Level1Out100[2] , 
        \ScanLink101[26] , \Level1Out104[13] , \Level1Out111[27] , 
        \Level1Out127[22] , \Level1Out171[23] , \Level32Out192[23] , 
        \Level2Out168[12] , \Level1Out132[16] , \Level1Out152[12] , 
        \Level1Out147[26] , \Level2Out36[2] , \Level2Out108[16] , 
        \Level16Out192[16] , \ScanLink122[17] , \Level1Out164[17] , 
        \ScanLink157[27] , \ScanLink174[16] , \ScanLink114[12] , 
        \Level2Out84[16] , \ScanLink137[23] , \ScanLink161[22] , 
        \ScanLink142[13] , \Level8Out96[19] , \Level1Out103[1] , 
        \ScanLink209[21] , \ScanLink34[20] , \ScanLink41[10] , 
        \ScanLink62[21] , \Level8Load120[0] , \Level1Out36[28] , 
        \Level1Out43[18] , \Level1Out93[8] , \Level1Out60[30] , 
        \Level2Out236[14] , \Level4Out204[13] , \Level1Out60[29] , 
        \Level4Out252[12] , \ScanLink18[6] , \Level1Out20[7] , 
        \Level1Out36[31] , \Level1Out85[10] , \Level1Out90[24] , 
        \ScanLink123[9] , \Level1Load205[0] , \Level1Out219[20] , 
        \Level2Out200[11] , \Level4Out232[16] , \Level2Out110[4] , 
        \Level2Out186[27] , \Level4Out172[28] , \Level4Out124[30] , 
        \Level1Out162[8] , \Level4Out172[31] , \Level4Out124[29] , 
        \Level8Out128[15] , \ScanLink87[18] , \ScanLink190[6] , 
        \ScanLink222[5] , \Level2Out54[8] , \Level1Out23[4] , \ScanLink141[3] , 
        \ScanLink142[0] , \ScanLink217[19] , \ScanLink221[6] , 
        \Level4Out124[7] , \Level8Out96[3] , \Level4Out244[2] , 
        \ScanLink234[31] , \Level128Out128[17] , \ScanLink234[28] , 
        \Level2Out98[2] , \Level8Out88[21] , \ScanLink241[18] , 
        \Level2Load214[0] , \Level1Out28[10] , \Level1Out48[14] , 
        \Level1Out207[18] , \ScanLink193[5] , \Level1Out224[30] , 
        \Level2Out248[28] , \Level1Out224[29] , \Level2Out248[31] , 
        \Level8Out240[16] , \Level1Out251[19] , \Level8Out216[17] , 
        \Level2Out6[24] , \Level16Out80[11] , \Level8Out104[8] , 
        \ScanLink246[1] , \Level1Out28[23] , \Level1Out44[3] , 
        \ScanLink126[4] , \ScanLink129[28] , \ScanLink129[31] , 
        \Level1Load66[0] , \Level1Out139[29] , \Level2Out176[19] , 
        \Level4Out32[29] , \Level4Out64[31] , \Level1Out85[23] , 
        \Level2Out120[18] , \Level2Out174[0] , \Level4Out32[30] , 
        \Level1Out90[17] , \Level1Out139[30] , \Level4Out64[28] , 
        \Level8Out128[26] , \Level1Out96[5] , \Level2Out214[5] , 
        \Level1Out194[29] , \Level16Out80[22] , \Level1Out47[0] , 
        \Level1Out48[27] , \Level1Out194[30] , \Level4Out192[5] , 
        \Level8Out200[9] , \Level8Out240[25] , \Level1Out95[6] , 
        \Level1Out118[0] , \ScanLink138[8] , \Level2Out6[17] , 
        \Level2Out22[29] , \Level2Out74[31] , \Level8Out216[24] , 
        \Level128Out128[24] , \Level2Out74[28] , \Level4Out140[3] , 
        \ScanLink245[2] , \Level8Out88[12] , \Level2Out22[30] , 
        \Level1Out61[23] , \Level1Out88[9] , \ScanLink184[28] , 
        \ScanLink125[7] , \Level4Out220[6] , \ScanLink184[31] , 
        \Level4Out80[28] , \Level1Out22[16] , \Level1Out37[22] , 
        \Level1Out42[12] , \Level4Out156[7] , \Level1Out51[4] , 
        \Level1Out57[26] , \ScanLink253[6] , \Level2Out192[19] , 
        \Level4Out80[31] , \Level4Out4[2] , \Level1Out74[17] , 
        \Level1Out80[1] , \Level1Out83[2] , \ScanLink133[3] , 
        \Level4Out236[2] , \Level2Out38[4] , \Level2Out48[18] , 
        \Level4Out184[1] , \Level1Out110[8] , \Level2Out90[28] , 
        \Level8Out176[8] , \ScanLink115[18] , \ScanLink136[30] , 
        \ScanLink136[29] , \Level2Out90[31] , \Level2Out162[4] , 
        \ScanLink143[19] , \ScanLink160[31] , \Level2Out202[1] , 
        \Level1Out126[28] , \ScanLink160[28] , \Level1Out153[18] , 
        \Level1Out170[30] , \Level16Out32[23] , \ScanLink250[5] , 
        \Level8Out208[1] , \Level1Out14[20] , \ScanLink16[31] , 
        \ScanLink16[28] , \Level1Out52[7] , \Level1Out105[19] , 
        \Level1Out126[31] , \ScanLink130[0] , \Level1Out170[29] , 
        \Level16Out64[22] , \Level128Out0[1] , \Level2Out26[8] , 
        \Level8Out168[4] , \ScanLink35[19] , \ScanLink40[30] , 
        \ScanLink63[18] , \Level1Out22[25] , \ScanLink40[29] , 
        \ScanLink185[1] , \ScanLink208[18] , \Level8Load72[0] , 
        \Level1Out57[15] , \Level1Out218[19] , \ScanLink237[2] , 
        \Level2Out222[19] , \Level4Out132[3] , \Level4Out196[31] , 
        \Level2Load78[0] , \ScanLink69[5] , \Level1Out74[24] , 
        \Level4Out196[28] , \Level4Out252[6] , \Level1Out35[0] , 
        \Level1Out37[11] , \Level1Out61[10] , \ScanLink157[7] , 
        \Level1Out42[21] , \Level1Out169[3] , \ScanLink234[1] , 
        \Level1Out6[25] , \Level1Load14[0] , \Level1Out36[3] , 
        \ScanLink154[4] , \Level16Out32[10] , \Level16Out64[11] , 
        \Level1Out209[6] , \Level8Out80[7] , \Level2Out106[0] , 
        \Level1Out29[30] , \Level1Out29[29] , \ScanLink68[14] , 
        \ScanLink77[9] , \ScanLink98[19] , \ScanLink186[2] , \Level1Out214[9] , 
        \ScanLink240[21] , \Level1Out98[3] , \ScanLink185[22] , 
        \ScanLink190[16] , \ScanLink235[11] , \ScanLink255[8] , 
        \Level32Out64[8] , \ScanLink203[14] , \ScanLink216[20] , 
        \Level2Out56[13] , \ScanLink255[15] , \Level2Out36[17] , 
        \Level2Out60[16] , \ScanLink220[25] , \Level1Out115[5] , 
        \Level1Out213[15] , \ScanLink248[7] , \ScanLink15[3] , \ScanLink16[0] , 
        \Level1Out245[14] , \Level1Out84[29] , \ScanLink128[2] , 
        \Level1Out195[23] , \Level1Out230[24] , \Level1Out250[20] , 
        \Level4Out188[10] , \Level1Out180[17] , \Level1Out225[10] , 
        \Level1Out206[21] , \Level16Out176[16] , \Level2Out154[22] , 
        \Level1Out49[6] , \Level1Out84[30] , \Level1Out116[6] , 
        \Level2Out102[23] , \Level1Out138[23] , \Level1Out158[27] , 
        \Level2Out162[27] , \Level2Out134[26] , \Level1Out1[3] , 
        \Level1Out2[0] , \Level1Out6[16] , \Level1Out54[9] , \ScanLink86[21] , 
        \ScanLink93[15] , \ScanLink148[26] , \Level2Out0[4] , 
        \Level8Out24[18] , \Level8Out72[19] , \Level2Out20[6] , 
        \ScanLink72[4] , \ScanLink128[22] , \Level1Out180[24] , 
        \Level1Out225[23] , \Level1Out250[13] , \Level4Out188[23] , 
        \Level1Out171[1] , \Level1Out206[12] , \Level16Out176[25] , 
        \Level1Out195[10] , \Level1Out213[26] , \Level1Out211[4] , 
        \Level1Out230[17] , \Level8Load152[0] , \ScanLink68[27] , 
        \ScanLink185[11] , \ScanLink203[27] , \Level1Out245[27] , 
        \Level2Out36[24] , \ScanLink220[16] , \ScanLink255[26] , 
        \Level2Out60[25] , \Level2Out88[8] , \ScanLink190[25] , 
        \ScanLink235[22] , \ScanLink240[12] , \ScanLink86[12] , 
        \ScanLink151[9] , \ScanLink216[13] , \Level2Out56[20] , 
        \ScanLink128[11] , \Level1Out2[27] , \ScanLink9[2] , \ScanLink71[7] , 
        \ScanLink93[26] , \ScanLink148[15] , \Level1Load168[0] , 
        \Level2Out44[2] , \Level1Out158[14] , \Level2Out162[14] , 
        \Level1Out172[2] , \ScanLink82[23] , \Level1Out138[10] , 
        \Level1Out212[7] , \Level2Out134[15] , \Level2Out154[11] , 
        \Level2Out96[4] , \Level2Out102[10] , \ScanLink87[7] , 
        \ScanLink159[10] , \Level2Out60[4] , \ScanLink97[17] , 
        \ScanLink139[14] , \ScanLink55[1] , \Level1Out129[15] , 
        \Level1Out184[2] , \ScanLink216[9] , \Level2Out166[25] , 
        \Level1Out236[1] , \Level2Out130[24] , \Level2Out124[8] , 
        \Level2Out150[20] , \Level1Out149[11] , \Level2Out106[21] , 
        \Level4Out48[5] , \Level1Out155[7] , \Level1Out156[4] , 
        \ScanLink168[0] , \Level1Out254[22] , \Level1Out184[15] , 
        \Level1Out221[12] , \Level1Out202[23] , \Level1Out235[2] , 
        \Level2Out238[23] , \Level2Out188[10] , \Level16Out112[10] , 
        \ScanLink208[5] , \Level1Out217[17] , \Level1Out241[16] , 
        \Level1Out2[14] , \Level1Out17[8] , \ScanLink56[2] , \ScanLink181[20] , 
        \Level1Out191[21] , \Level32Out192[1] , \ScanLink207[16] , 
        \Level1Out234[26] , \Level2Out32[15] , \Level16Out144[11] , 
        \ScanLink251[17] , \Level2Out64[14] , \ScanLink224[27] , 
        \ScanLink19[26] , \ScanLink79[22] , \Level4Out56[9] , \ScanLink19[15] , 
        \ScanLink31[5] , \Level1Out80[18] , \ScanLink84[4] , \Level1Out148[8] , 
        \ScanLink244[23] , \Level1Out187[1] , \ScanLink194[14] , 
        \ScanLink231[13] , \ScanLink212[22] , \Level2Out52[11] , 
        \Level1Out252[5] , \Level2Out150[13] , \Level1Out129[26] , 
        \Level1Out149[22] , \Level2Out220[9] , \Level2Out106[12] , 
        \Level1Out132[0] , \Level2Load20[0] , \Level2Out166[16] , 
        \ScanLink82[10] , \ScanLink97[24] , \ScanLink112[8] , 
        \ScanLink139[27] , \Level2Out130[17] , \ScanLink159[23] , 
        \ScanLink194[27] , \ScanLink231[20] , \Level1Out58[31] , 
        \Level1Out58[28] , \ScanLink79[11] , \ScanLink181[13] , 
        \ScanLink207[25] , \ScanLink212[11] , \ScanLink244[10] , 
        \Level2Out32[26] , \Level2Out52[22] , \ScanLink224[14] , 
        \Level1Out217[24] , \ScanLink251[24] , \Level2Out64[27] , 
        \Level2Out188[23] , \Level16Out112[23] , \Level16Out144[22] , 
        \Level1Out191[12] , \Level1Out234[15] , \Level1Out241[25] , 
        \Level1Out251[6] , \Level1Out12[5] , \ScanLink32[6] , 
        \Level1Out184[26] , \Level1Out221[21] , \Level1Out254[11] , 
        \Level1Out131[3] , \Level1Out202[10] , \Level2Out238[10] , 
        \ScanLink170[2] , \Level8Out128[6] , \Level64Out128[21] , 
        \ScanLink210[7] , \Level8Out248[3] , \ScanLink12[19] , 
        \ScanLink67[29] , \ScanLink81[9] , \Level2Out78[6] , \Level2Out122[6] , 
        \Level2Out242[3] , \Level4Out108[9] , \ScanLink31[31] , 
        \ScanLink31[28] , \ScanLink44[18] , \ScanLink67[30] , 
        \Level1Out53[24] , \Level1Out153[9] , \ScanLink0[24] , 
        \Level1Out9[18] , \Level1Out11[6] , \Level1Out26[14] , 
        \Level2Out226[28] , \Level1Out70[15] , \ScanLink173[1] , 
        \Level1Out10[11] , \Level1Out65[21] , \Level2Out226[31] , 
        \Level4Out192[19] , \Level2Out8[20] , \Level1Out33[20] , 
        \Level1Out46[10] , \Level4Out116[5] , \ScanLink109[9] , 
        \ScanLink213[4] , \Level2Out94[19] , \Level2Out226[7] , 
        \ScanLink111[30] , \ScanLink147[28] , \Level2Out146[2] , 
        \ScanLink111[29] , \ScanLink132[18] , \ScanLink147[31] , 
        \ScanLink164[19] , \Level1Out157[29] , \Level2Out118[19] , 
        \Level1Out10[22] , \Level1Out76[1] , \Level1Out101[31] , 
        \Level1Out101[28] , \Level1Out122[19] , \Level1Out157[30] , 
        \Level8Out8[2] , \Level1Out174[18] , \ScanLink114[6] , 
        \Level1Out129[1] , \Level1Out249[4] , \Level2Out194[4] , 
        \Level64Out128[12] , \Level1Out26[27] , \Level1Out33[13] , 
        \Level1Out65[12] , \Level2Out8[13] , \Level2Out196[31] , 
        \Level4Out84[19] , \Level4Out212[4] , \ScanLink117[5] , 
        \Level2Out196[28] , \Level1Out46[23] , \Level1Out75[2] , 
        \Level4Out172[1] , \Level1Load2[0] , \Level1Out2[9] , \ScanLink29[7] , 
        \Level1Out53[17] , \Level1Out29[13] , \ScanLink34[8] , 
        \Level1Out70[26] , \Level1Load130[0] , \Level8Out184[16] , 
        \Level1Out33[7] , \Level1Out49[17] , \ScanLink183[6] , 
        \Level1Out195[19] , \Level1Load216[0] , \Level1Out171[8] , 
        \Level2Out88[1] , \Level2Out56[30] , \Level1Out30[4] , 
        \ScanLink151[0] , \Level2Out56[29] , \ScanLink152[3] , 
        \ScanLink185[18] , \ScanLink231[5] , \Level4Out72[6] , 
        \Level8Out24[22] , \Level8Out72[23] , \Level1Out84[13] , 
        \ScanLink128[18] , \ScanLink232[6] , \Level2Out154[18] , 
        \Level1Out91[27] , \Level1Out138[19] , \ScanLink180[5] , 
        \Level2Out100[7] , \Level2Out102[19] , \ScanLink135[4] , 
        \Level1Out4[7] , \Level1Out14[29] , \ScanLink16[21] , \ScanLink16[9] , 
        \Level1Out29[20] , \Level1Out49[24] , \Level1Out57[3] , 
        \Level1Out108[3] , \ScanLink240[28] , \Level4Out16[2] , 
        \Level4Load140[0] , \Level1Out206[31] , \ScanLink216[30] , 
        \ScanLink235[18] , \ScanLink255[1] , \Level32Out64[1] , 
        \ScanLink216[29] , \ScanLink240[31] , \Level1Out225[19] , 
        \Level1Out250[29] , \Level4Out188[19] , \Level1Out206[28] , 
        \Level1Out250[30] , \Level1Out85[5] , \Level1Load75[0] , 
        \Level8Out184[25] , \ScanLink20[24] , \Level1Out54[0] , 
        \Level1Out84[20] , \Level1Out86[6] , \Level2Out204[6] , 
        \Level1Out91[14] , \Level2Out164[3] , \ScanLink86[28] , 
        \ScanLink86[31] , \ScanLink136[7] , \ScanLink256[2] , 
        \Level8Out24[11] , \Level8Out72[10] , \Level2Out48[22] , 
        \Level1Out28[6] , \ScanLink55[14] , \ScanLink185[8] , 
        \ScanLink208[11] , \Level16Out96[7] , \Level1Out217[3] , 
        \Level8Out112[5] , \ScanLink76[25] , \ScanLink35[10] , 
        \ScanLink63[11] , \Level1Out177[6] , \ScanLink40[20] , \ScanLink74[3] , 
        \Level2Out28[26] , \Level4Load80[0] , \Level2Out214[15] , 
        \Level1Out7[4] , \Level1Out14[30] , \Level1Out37[18] , 
        \Level1Out42[31] , \Level1Out61[19] , \Level4Out80[12] , 
        \ScanLink198[7] , \Level1Out35[9] , \Level1Out42[28] , 
        \Level2Out192[23] , \Level2Out242[14] , \Level1Out126[12] , 
        \Level1Out153[22] , \Level1Out218[10] , \Level2Out222[10] , 
        \Level2Out42[5] , \Level2Out118[5] , \Level4Out196[21] , 
        \Level1Out170[13] , \Level16Out32[19] , \Level16Out64[18] , 
        \ScanLink10[7] , \ScanLink16[12] , \ScanLink63[22] , \ScanLink77[0] , 
        \ScanLink100[16] , \Level1Out105[23] , \Level1Out110[17] , 
        \Level1Out165[27] , \Level1Out133[26] , \Level1Out146[16] , 
        \ScanLink234[8] , \ScanLink175[26] , \Level2Out90[12] , 
        \Level2Out90[3] , \ScanLink123[27] , \ScanLink156[17] , 
        \ScanLink143[23] , \ScanLink149[2] , \Level1Out214[0] , 
        \Level4Out4[24] , \Level2Out106[9] , \ScanLink98[10] , 
        \ScanLink136[13] , \Level1Load109[0] , \ScanLink115[22] , 
        \ScanLink160[12] , \Level1Out174[5] , \ScanLink229[7] , 
        \Level1Out218[23] , \Level2Out192[10] , \Level2Out214[26] , 
        \Level2Out222[23] , \Level4Out80[21] , \Level4Out196[12] , 
        \Level2Out242[27] , \Level16Out192[6] , \ScanLink35[23] , 
        \ScanLink40[13] , \Level2Out28[15] , \ScanLink55[27] , 
        \ScanLink208[22] , \Level8Out176[1] , \Level2Out48[11] , 
        \ScanLink13[4] , \ScanLink20[17] , \ScanLink76[16] , \Level4Out184[8] , 
        \Level1Out80[8] , \ScanLink98[23] , \Level1Out113[2] , 
        \ScanLink115[11] , \ScanLink136[20] , \Level4Out228[7] , 
        \Level8Out216[4] , \ScanLink143[10] , \Level2Out6[3] , 
        \Level2Out202[8] , \ScanLink100[25] , \ScanLink160[21] , 
        \Level2Out90[21] , \Level1Out110[1] , \ScanLink175[15] , 
        \Level4Out148[2] , \ScanLink123[14] , \ScanLink156[24] , 
        \Level4Out4[17] , \Level2Load118[0] , \ScanLink37[2] , 
        \Level1Out105[10] , \Level1Out110[24] , \Level1Out126[21] , 
        \ScanLink130[9] , \Level1Out165[14] , \Level1Out133[15] , 
        \Level1Out146[25] , \Level2Out26[1] , \Level1Out153[11] , 
        \Level8Out208[8] , \ScanLink147[21] , \Level1Out170[20] , 
        \Level128Out0[8] , \Level1Out76[8] , \ScanLink89[26] , 
        \ScanLink111[20] , \ScanLink132[11] , \Level1Out134[7] , 
        \ScanLink164[10] , \ScanLink171[24] , \ScanLink104[14] , 
        \ScanLink109[0] , \ScanLink152[15] , \Level2Out94[10] , 
        \Level1Out114[15] , \ScanLink127[25] , \Level1Out161[25] , 
        \Level1Out254[2] , \Level4Out0[26] , \Level1Out122[10] , 
        \Level1Out129[8] , \Level1Out142[14] , \Level1Out137[24] , 
        \Level2Out178[14] , \Level1Out157[20] , \Level2Out118[10] , 
        \Level1Out101[21] , \Level1Out174[11] , \Level2Out226[12] , 
        \Level4Out172[8] , \ScanLink1[27] , \ScanLink1[14] , \ScanLink1[3] , 
        \Level1Out9[22] , \Level2Out158[7] , \Level4Out192[23] , 
        \Level1Out9[11] , \Level1Out10[18] , \ScanLink12[23] , 
        \Level1Out209[26] , \Level2Out196[21] , \Level2Out210[17] , 
        \Level4Out84[10] , \Level2Out238[2] , \Level2Out246[16] , 
        \ScanLink12[10] , \ScanLink24[26] , \ScanLink31[12] , \ScanLink67[13] , 
        \Level8Out232[2] , \Level1Out137[4] , \ScanLink34[1] , 
        \ScanLink44[22] , \ScanLink219[27] , \ScanLink24[15] , \ScanLink50[5] , 
        \ScanLink51[25] , \ScanLink51[16] , \Level8Out152[7] , \ScanLink53[6] , 
        \Level1Out68[4] , \ScanLink72[27] , \ScanLink81[0] , 
        \Level1Out101[12] , \Level1Out122[23] , \Level1Out157[13] , 
        \Level1Out182[5] , \Level2Out118[23] , \Level1Out174[22] , 
        \ScanLink89[15] , \ScanLink104[27] , \Level1Out114[26] , 
        \Level1Out137[17] , \Level1Out161[16] , \Level64Out128[31] , 
        \Level1Out142[27] , \Level2Out66[3] , \Level2Out178[27] , 
        \Level64Out128[28] , \Level1Out150[3] , \ScanLink171[17] , 
        \Level2Out94[23] , \Level4Out108[0] , \ScanLink127[16] , 
        \ScanLink152[26] , \Level4Out0[15] , \ScanLink111[13] , 
        \ScanLink132[22] , \ScanLink147[12] , \Level1Out230[6] , 
        \ScanLink164[23] , \ScanLink67[20] , \ScanLink72[14] , 
        \Level1Out153[0] , \ScanLink31[21] , \ScanLink44[11] , 
        \ScanLink219[14] , \Level1Out65[28] , \Level1Out233[5] , 
        \Level8Out136[3] , \Level4Out84[23] , \Level1Out33[30] , 
        \Level2Out210[24] , \Level1Out33[29] , \Level1Out46[19] , 
        \ScanLink82[3] , \Level2Out8[29] , \Level4Load76[0] , 
        \Level1Out209[15] , \Level1Out65[31] , \Level2Out196[12] , 
        \Level2Out246[25] , \ScanLink173[8] , \Level1Out181[6] , 
        \Level2Out8[30] , \Level2Out226[21] , \Level4Out192[10] , 
        \Level1Out11[12] , \Level1Out14[2] , \Level1Out38[25] , 
        \Level1Out70[6] , \Level1Out80[11] , \Level1Out95[25] , 
        \Level1Out132[9] , \Level2Out140[5] , \Level16Out48[14] , 
        \Level32Out32[17] , \Level128Out0[24] , \ScanLink82[19] , 
        \Level2Out220[0] , \Level8Out16[25] , \Level32Out64[16] , 
        \ScanLink112[1] , \Level2Out192[3] , \Level8Out40[24] , 
        \Level1Out73[5] , \ScanLink79[18] , \Level1Load83[0] , 
        \ScanLink231[29] , \Level4Out32[4] , \ScanLink244[19] , 
        \ScanLink111[2] , \ScanLink212[18] , \ScanLink231[30] , 
        \Level1Out202[19] , \Level1Out221[28] , \Level1Out254[18] , 
        \Level1Out221[31] , \Level2Out238[19] , \Level32Load96[0] , 
        \ScanLink48[7] , \Level1Out58[21] , \ScanLink216[0] , \Level4Load0[0] , 
        \Level8Out16[16] , \Level1Out17[1] , \Level1Out38[16] , 
        \ScanLink55[8] , \Level1Out80[22] , \ScanLink159[19] , 
        \ScanLink176[5] , \Level8Out40[17] , \Level2Out124[1] , 
        \Level2Out106[31] , \Level128Out0[17] , \Level1Out58[12] , 
        \Level1Out95[16] , \Level1Out149[18] , \Level2Out150[29] , 
        \Level32Out32[24] , \Level32Out64[25] , \Level1Load151[0] , 
        \Level1Out199[4] , \Level2Out106[28] , \Level2Out150[30] , 
        \Level2Out244[4] , \Level16Out48[27] , \Level1Out236[8] , 
        \Level2Out188[19] , \Level4Out84[6] , \Level16Out112[19] , 
        \ScanLink99[2] , \Level1Out191[31] , \Level1Out191[28] , 
        \Level16Out144[18] , \Level32Out192[8] , \ScanLink168[9] , 
        \Level1Out148[1] , \Level4Out56[0] , \ScanLink175[6] , 
        \Level1Out187[8] , \ScanLink215[3] , \Level2Out52[18] , 
        \Level2Load140[0] , \ScanLink181[30] , \Level1Out228[4] , 
        \Level1Out32[23] , \Level1Out47[13] , \ScanLink181[29] , 
        \Level4Out40[4] , \Level4Out200[18] , \Level1Out64[22] , 
        \ScanLink203[7] , \Level32Out32[7] , \Level1Out27[17] , 
        \Level1Out52[27] , \Level1Out71[16] , \ScanLink92[9] , 
        \ScanLink163[2] , \Level2Out38[30] , \ScanLink2[0] , \Level2Out38[29] , 
        \Level4Out92[2] , \Level2Out68[5] , \Level2Out132[5] , 
        \Level1Out100[18] , \ScanLink110[19] , \ScanLink133[31] , 
        \Level1Out140[9] , \Level2Out252[0] , \Level1Out123[30] , 
        \ScanLink133[28] , \ScanLink165[29] , \ScanLink146[18] , 
        \ScanLink165[30] , \Level1Out123[29] , \Level1Out175[28] , 
        \Level4Out28[30] , \Level1Out156[19] , \Level1Out175[31] , 
        \ScanLink200[4] , \Level4Out28[29] , \Level1Out8[31] , 
        \Level1Out8[28] , \ScanLink13[30] , \ScanLink30[18] , \ScanLink160[1] , 
        \Level2Out76[9] , \Level8Out104[23] , \Level8Out152[22] , 
        \ScanLink13[29] , \ScanLink45[28] , \ScanLink45[31] , \ScanLink66[19] , 
        \Level2Out204[29] , \Level1Out27[24] , \ScanLink39[4] , 
        \Level1Out71[25] , \Level2Out252[31] , \Level2Load132[0] , 
        \Level2Out204[30] , \Level1Out11[21] , \Level1Out32[10] , 
        \Level1Out52[14] , \Level2Out252[28] , \Level4Out24[0] , 
        \Level1Out47[20] , \Level2Out228[8] , \Level1Out65[1] , 
        \Level1Out64[11] , \ScanLink104[5] , \ScanLink107[6] , 
        \Level1Out139[2] , \Level8Out104[10] , \Level2Out184[7] , 
        \Level4Out168[31] , \Level8Out152[11] , \Level4Out168[28] , 
        \Level1Out3[24] , \ScanLink18[25] , \ScanLink27[8] , \Level1Out66[2] , 
        \Level2Out156[1] , \ScanLink94[7] , \Level1Load123[0] , 
        \Level1Out244[8] , \Level2Out236[4] , \ScanLink213[21] , 
        \Level2Out26[22] , \Level4Out100[8] , \ScanLink78[21] , 
        \ScanLink180[23] , \ScanLink195[17] , \Level1Out197[2] , 
        \ScanLink245[20] , \Level2Out70[23] , \ScanLink205[9] , 
        \ScanLink230[10] , \ScanLink225[24] , \ScanLink250[14] , 
        \Level2Out10[27] , \ScanLink206[15] , \Level2Out46[26] , 
        \Level1Out240[15] , \ScanLink46[1] , \Level1Out59[18] , 
        \ScanLink89[8] , \Level1Out145[4] , \Level1Out190[22] , 
        \Level1Out235[25] , \Level4Out248[12] , \Level1Out216[14] , 
        \ScanLink218[6] , \Level8Out240[2] , \ScanLink178[3] , 
        \Level1Out203[20] , \Level1Out255[21] , \Level4Out228[16] , 
        \Level1Out185[16] , \Level8Out120[7] , \Level1Out220[11] , 
        \Level1Out225[1] , \ScanLink1[25] , \ScanLink1[16] , \Level1Out3[17] , 
        \Level1Out19[7] , \ScanLink45[2] , \Level1Out81[31] , 
        \Level1Out81[28] , \Level1Out146[7] , \Level1Out148[12] , 
        \Level4Out36[22] , \Level4Out140[15] , \Level2Out172[12] , 
        \Level4Out116[14] , \Level2Out124[13] , \Level4Out60[23] , 
        \Level1Out128[16] , \Level1Out226[2] , \Level32Out0[25] , 
        \Level2Out112[16] , \Level2Out144[17] , \Level4Out176[10] , 
        \Level4Out120[11] , \Level4Out56[26] , \ScanLink22[5] , 
        \ScanLink83[20] , \ScanLink96[14] , \ScanLink97[4] , \Level1Out194[1] , 
        \ScanLink138[17] , \ScanLink158[13] , \Level2Out70[7] , 
        \Level1Out121[0] , \Level1Out203[13] , \Level8Out224[6] , 
        \Level1Out185[25] , \Level1Out220[22] , \Level1Out255[12] , 
        \Level4Out228[25] , \Level1Out190[11] , \Level1Out235[16] , 
        \Level4Out248[21] , \Level1Out240[26] , \Level1Out241[5] , 
        \Level8Out144[3] , \ScanLink5[25] , \ScanLink5[16] , \Level1Out7[26] , 
        \ScanLink18[16] , \ScanLink78[12] , \ScanLink180[10] , 
        \Level1Out216[27] , \Level8Out224[19] , \ScanLink225[17] , 
        \Level8Out0[3] , \Level2Out10[14] , \ScanLink101[8] , 
        \ScanLink206[26] , \ScanLink250[27] , \ScanLink213[12] , 
        \Level2Out26[11] , \Level2Out46[15] , \Level4Out204[9] , 
        \ScanLink195[24] , \ScanLink230[23] , \ScanLink21[6] , 
        \ScanLink83[13] , \ScanLink158[20] , \ScanLink245[13] , 
        \Level2Out70[10] , \Level2Out182[9] , \ScanLink96[27] , 
        \Level2Out14[3] , \ScanLink138[24] , \Level2Out144[24] , 
        \Level4Out176[23] , \Level1Out59[5] , \ScanLink87[22] , 
        \Level1Out122[3] , \Level1Out128[25] , \Level4Out56[15] , 
        \Level32Out0[16] , \Level2Out112[25] , \ScanLink129[21] , 
        \Level1Out148[21] , \Level2Out172[21] , \Level4Out120[22] , 
        \Level4Out36[11] , \Level4Out140[26] , \Level1Out242[6] , 
        \Level2Out124[20] , \Level4Out60[10] , \Level4Out116[27] , 
        \Level2Out30[5] , \ScanLink92[16] , \ScanLink149[25] , 
        \ScanLink246[8] , \Level1Out159[24] , \Level2Out140[15] , 
        \Level4Out172[12] , \Level4Out124[13] , \Level2Out116[14] , 
        \Level4Out52[24] , \Level1Out106[5] , \Level4Out32[20] , 
        \ScanLink138[1] , \Level1Out139[20] , \Level4Out144[17] , 
        \Level1Out207[22] , \Level2Out120[11] , \Level2Out174[9] , 
        \Level2Out176[10] , \Level4Out112[16] , \Level2Out198[25] , 
        \Level4Out64[21] , \Level1Out251[23] , \Level2Out248[12] , 
        \Level1Out181[14] , \Level8Out160[5] , \Level1Out224[13] , 
        \Level1Out7[15] , \Level1Out47[9] , \Level1Out105[6] , 
        \Level1Out194[20] , \Level1Out231[27] , \Level1Out244[17] , 
        \Level2Out228[16] , \ScanLink184[21] , \Level1Out212[16] , 
        \ScanLink221[26] , \ScanLink254[16] , \Level8Out200[0] , 
        \Level2Out14[25] , \ScanLink61[4] , \ScanLink69[17] , \Level1Out88[0] , 
        \ScanLink202[17] , \Level2Out42[24] , \ScanLink217[23] , 
        \ScanLink241[22] , \Level2Out22[20] , \Level2Out74[21] , 
        \Level1Out85[19] , \Level1Out118[9] , \Level1Out139[13] , 
        \ScanLink191[15] , \ScanLink234[12] , \Level2Out86[7] , 
        \Level2Out176[23] , \Level4Out144[24] , \Level2Out120[22] , 
        \Level4Out32[13] , \Level4Out64[12] , \Level1Out202[4] , 
        \Level2Out140[26] , \Level4Out112[25] , \Level4Out172[21] , 
        \ScanLink69[24] , \ScanLink87[11] , \ScanLink92[25] , 
        \Level1Out159[17] , \Level2Out116[27] , \Level4Out52[17] , 
        \Level4Out124[20] , \Level1Out162[1] , \Level2Out54[1] , 
        \ScanLink129[12] , \ScanLink142[9] , \ScanLink149[16] , 
        \ScanLink217[10] , \Level8Out88[31] , \Level2Out22[13] , 
        \Level8Out88[28] , \ScanLink184[12] , \ScanLink191[26] , 
        \ScanLink221[15] , \ScanLink234[21] , \ScanLink241[11] , 
        \Level2Out14[16] , \Level2Out74[12] , \Level1Out194[13] , 
        \ScanLink202[24] , \ScanLink254[25] , \Level1Out231[14] , 
        \Level2Out42[17] , \Level16Out80[18] , \Level1Out201[7] , 
        \Level16Out80[3] , \Level1Out28[19] , \Level1Out212[25] , 
        \Level1Out244[24] , \Level8Out104[1] , \Level8Out88[6] , 
        \Level2Out228[25] , \Level1Out42[4] , \ScanLink62[7] , 
        \Level1Out161[2] , \Level1Out207[11] , \Level2Out248[21] , 
        \Level2Out198[16] , \Level1Out181[27] , \Level1Out224[20] , 
        \Level1Out251[10] , \ScanLink120[3] , \ScanLink240[6] , 
        \Level8Out136[24] , \Level1Out15[10] , \ScanLink17[18] , 
        \ScanLink34[29] , \ScanLink41[19] , \Level1Out90[2] , 
        \Level2Out212[2] , \Level8Out160[25] , \ScanLink99[30] , 
        \ScanLink99[29] , \Level2Out172[7] , \ScanLink62[31] , 
        \ScanLink62[28] , \Level2Out28[7] , \Level1Out23[15] , 
        \ScanLink34[30] , \Level1Out41[7] , \Level1Out56[25] , 
        \Level1Out75[14] , \Level1Out93[1] , \Level1Out103[8] , 
        \ScanLink209[31] , \Level8Out96[10] , \ScanLink209[28] , 
        \Level1Out219[30] , \Level8Out208[26] , \ScanLink123[0] , 
        \Level1Out219[29] , \Level2Out8[5] , \Level2Out200[18] , 
        \Level1Out36[21] , \Level1Out43[11] , \Level1Out60[20] , 
        \ScanLink243[5] , \Level1Out104[29] , \ScanLink114[31] , 
        \ScanLink114[28] , \ScanLink142[30] , \ScanLink159[8] , 
        \ScanLink196[1] , \Level2Out80[9] , \ScanLink161[18] , 
        \ScanLink142[29] , \Level2Out116[3] , \ScanLink137[19] , 
        \Level1Out152[31] , \Level1Out171[19] , \Level2Out168[31] , 
        \Level32Out192[19] , \ScanLink144[7] , \Level1Out152[28] , 
        \Level1Out219[5] , \Level8Out136[17] , \Level8Out160[16] , 
        \Level1Out9[2] , \Level1Out15[23] , \Level1Out25[3] , \Level1Out26[0] , 
        \Level1Out104[30] , \Level2Out168[28] , \Level1Out127[18] , 
        \Level1Out36[12] , \Level1Out179[0] , \ScanLink224[2] , 
        \Level1Out43[22] , \Level4Load132[0] , \Level4Out204[29] , 
        \Level4Out252[31] , \Level1Out23[26] , \Level1Out60[13] , 
        \Level4Out204[30] , \Level1Out75[27] , \ScanLink147[4] , 
        \Level4Out252[28] , \Level8Out208[15] , \ScanLink79[6] , 
        \Level1Out56[16] , \ScanLink227[1] , \Level4Out64[2] , 
        \Level8Out96[23] , \ScanLink64[9] , \ScanLink195[2] , 
        \Level1Out207[9] , \ScanLink91[8] , \ScanLink160[3] , 
        \Level1Load195[0] , \Level8Out104[21] , \Level8Out152[20] , 
        \Level4Out168[19] , \ScanLink200[6] , \ScanLink1[1] , \ScanLink2[2] , 
        \Level2Out132[7] , \Level2Out252[2] , \ScanLink13[18] , 
        \ScanLink30[30] , \ScanLink30[29] , \ScanLink45[19] , \ScanLink66[31] , 
        \Level16Out0[9] , \ScanLink66[28] , \Level2Out68[7] , 
        \Level1Out143[8] , \Level1Out8[19] , \ScanLink163[0] , 
        \Level1Load224[0] , \Level2Load184[0] , \Level4Out92[0] , 
        \Level2Out204[18] , \Level1Out11[10] , \Level1Out27[15] , 
        \Level1Out71[14] , \Level1Out32[21] , \Level1Out52[25] , 
        \Level2Out252[19] , \Level1Out47[11] , \ScanLink203[5] , 
        \Level32Out32[5] , \Level4Out40[6] , \Level1Out64[20] , 
        \Level1Out66[0] , \Level1Out100[29] , \ScanLink104[7] , 
        \ScanLink110[31] , \ScanLink110[28] , \ScanLink119[8] , 
        \Level2Out236[6] , \ScanLink133[19] , \ScanLink146[30] , 
        \ScanLink165[18] , \ScanLink146[29] , \Level2Out156[3] , 
        \Level1Out123[18] , \Level1Out156[31] , \Level1Out175[19] , 
        \Level1Out100[30] , \Level1Out156[28] , \Level4Out28[18] , 
        \Level1Out1[8] , \Level1Out3[26] , \Level1Out11[23] , 
        \Level1Out32[12] , \Level1Out47[22] , \Level1Out139[0] , 
        \Level2Out184[5] , \Level8Out104[12] , \Level4Load172[0] , 
        \Level8Out152[13] , \Level1Out65[3] , \Level1Out64[13] , 
        \Level4Out200[29] , \ScanLink107[4] , \Level4Out200[30] , 
        \Level1Out19[5] , \ScanLink24[9] , \Level1Out27[26] , \ScanLink39[6] , 
        \Level1Out71[27] , \Level1Out52[16] , \Level4Out24[2] , 
        \Level1Out247[9] , \Level2Out38[18] , \Level1Load47[0] , 
        \ScanLink83[22] , \ScanLink158[11] , \ScanLink96[16] , 
        \Level1Out194[3] , \ScanLink206[8] , \Level2Out70[5] , \ScanLink97[6] , 
        \Level1Out128[14] , \ScanLink138[15] , \Level1Out226[0] , 
        \Level2Out144[15] , \Level4Out176[12] , \Level32Out0[27] , 
        \Level4Out56[24] , \ScanLink45[0] , \Level1Out146[5] , 
        \Level2Out112[14] , \Level2Out172[10] , \Level4Out120[13] , 
        \Level1Out148[10] , \Level4Out140[17] , \Level4Out36[20] , 
        \ScanLink46[3] , \ScanLink178[1] , \Level1Out185[14] , 
        \Level1Out203[22] , \Level2Out124[11] , \Level2Out134[9] , 
        \Level4Out60[21] , \Level4Out116[16] , \Level1Out220[13] , 
        \Level8Out120[5] , \Level1Out225[3] , \Level1Out255[23] , 
        \Level4Out228[14] , \Level8Out224[31] , \Level1Out190[20] , 
        \Level1Out235[27] , \Level4Out248[10] , \Level1Out3[15] , 
        \ScanLink18[27] , \ScanLink78[23] , \Level1Out145[6] , 
        \Level1Out240[17] , \Level8Out224[28] , \ScanLink180[21] , 
        \Level1Out216[16] , \Level8Out240[0] , \ScanLink218[4] , 
        \Level2Out10[25] , \Level64Out128[8] , \ScanLink225[26] , 
        \ScanLink94[5] , \ScanLink206[17] , \ScanLink250[16] , 
        \Level2Out46[24] , \Level1Out158[9] , \ScanLink213[23] , 
        \Level2Out26[20] , \ScanLink195[15] , \ScanLink230[12] , 
        \Level1Out197[0] , \ScanLink18[14] , \ScanLink21[4] , 
        \Level1Out81[19] , \Level1Out148[23] , \ScanLink245[22] , 
        \Level2Out70[21] , \Level1Out242[4] , \Level2Out172[23] , 
        \Level2Out230[8] , \Level4Out36[13] , \Level4Out140[24] , 
        \Level2Out124[22] , \Level4Out116[25] , \Level4Out60[12] , 
        \ScanLink83[11] , \ScanLink96[25] , \Level1Out122[1] , 
        \Level2Out144[26] , \Level4Out176[21] , \Level32Out0[14] , 
        \Level4Out120[20] , \Level1Out128[27] , \Level2Out112[27] , 
        \Level4Out56[17] , \ScanLink102[9] , \Level2Out14[1] , 
        \ScanLink138[26] , \ScanLink158[22] , \ScanLink213[10] , 
        \Level2Out26[13] , \ScanLink78[10] , \ScanLink180[12] , 
        \ScanLink195[26] , \ScanLink230[21] , \ScanLink245[11] , 
        \Level2Out70[12] , \ScanLink250[25] , \Level2Out10[16] , 
        \ScanLink225[15] , \ScanLink206[24] , \Level2Out46[17] , 
        \Level1Out241[7] , \ScanLink5[27] , \ScanLink5[14] , \Level1Out7[24] , 
        \ScanLink22[7] , \Level1Out59[30] , \Level1Out190[13] , 
        \Level1Out240[24] , \Level8Out144[1] , \Level1Out235[14] , 
        \Level4Out248[23] , \Level1Out59[29] , \Level8Out0[1] , 
        \Level1Out121[2] , \Level1Out216[25] , \Level8Out224[4] , 
        \Level1Out203[11] , \Level1Out255[10] , \Level4Out228[27] , 
        \ScanLink69[15] , \Level1Out185[27] , \Level1Out220[20] , 
        \ScanLink217[21] , \Level2Out22[22] , \Level8Out88[19] , 
        \Level1Out88[2] , \ScanLink184[23] , \ScanLink191[17] , 
        \ScanLink234[10] , \ScanLink241[20] , \ScanLink245[9] , 
        \Level2Out74[23] , \Level4Out140[8] , \ScanLink221[24] , 
        \Level2Out14[27] , \Level1Out194[22] , \ScanLink202[15] , 
        \ScanLink254[14] , \Level2Out42[26] , \Level16Out80[29] , 
        \Level1Out231[25] , \Level1Out244[15] , \Level1Out7[17] , 
        \Level1Out28[31] , \Level1Out28[28] , \Level1Out105[4] , 
        \Level16Out80[30] , \Level1Out212[14] , \Level8Out200[2] , 
        \Level2Out228[14] , \Level1Out44[8] , \Level1Out59[7] , 
        \Level1Out85[31] , \Level1Out106[7] , \ScanLink138[3] , 
        \Level1Out181[16] , \Level1Out207[20] , \Level2Out248[10] , 
        \Level1Out224[11] , \Level2Out198[27] , \Level8Out160[7] , 
        \Level1Out139[22] , \Level1Out251[21] , \Level2Out176[12] , 
        \Level4Out144[15] , \Level4Out32[22] , \Level1Out85[28] , 
        \Level2Out120[13] , \Level4Out64[23] , \Level4Out112[14] , 
        \Level2Out140[17] , \Level4Out52[26] , \Level4Out172[10] , 
        \ScanLink92[14] , \Level1Out159[26] , \Level2Out116[16] , 
        \Level4Out124[11] , \ScanLink129[23] , \ScanLink149[27] , 
        \ScanLink62[5] , \ScanLink87[20] , \Level1Out161[0] , \Level2Out30[7] , 
        \Level2Out198[14] , \Level1Out207[13] , \Level1Out251[12] , 
        \Level2Out248[23] , \Level1Out181[25] , \Level1Out224[22] , 
        \Level1Out201[5] , \Level1Out244[26] , \Level8Out88[4] , 
        \Level8Out104[3] , \Level1Out15[12] , \Level1Out36[23] , 
        \ScanLink61[6] , \ScanLink69[26] , \ScanLink141[8] , \ScanLink184[10] , 
        \Level1Out194[11] , \Level16Out80[1] , \Level1Out212[27] , 
        \Level1Out231[16] , \Level2Out228[27] , \ScanLink254[27] , 
        \ScanLink202[26] , \ScanLink221[17] , \Level2Out14[14] , 
        \Level2Out42[15] , \Level4Load44[0] , \ScanLink217[12] , 
        \Level2Out22[11] , \Level4Out244[9] , \ScanLink241[13] , 
        \Level2Out74[10] , \Level2Out98[9] , \ScanLink87[13] , 
        \ScanLink129[10] , \ScanLink191[24] , \ScanLink234[23] , 
        \ScanLink92[27] , \ScanLink149[14] , \Level2Out54[3] , 
        \Level8Out96[8] , \Level1Out139[11] , \Level1Out159[15] , 
        \Level1Out162[3] , \Level2Out140[24] , \Level4Out172[23] , 
        \Level2Out116[25] , \Level4Out124[22] , \Level4Out32[11] , 
        \Level4Out52[15] , \Level1Out202[6] , \Level2Out86[5] , 
        \Level2Out176[21] , \Level4Out144[26] , \Level4Out112[27] , 
        \Level2Out120[20] , \Level4Out64[10] , \Level4Out204[18] , 
        \Level1Out43[13] , \ScanLink243[7] , \Level1Out23[17] , 
        \Level1Out41[5] , \Level1Out60[22] , \Level4Out252[19] , 
        \Level1Out75[16] , \ScanLink123[2] , \Level2Out8[7] , 
        \Level8Out208[24] , \Level1Out56[27] , \Level1Out90[0] , 
        \Level1Out93[3] , \Level4Load184[0] , \Level8Out96[12] , 
        \Level1Out100[9] , \Level2Out28[5] , \Level2Out172[5] , 
        \Level1Out104[18] , \ScanLink114[19] , \ScanLink161[29] , 
        \Level2Out212[0] , \ScanLink137[31] , \ScanLink137[28] , 
        \ScanLink142[18] , \ScanLink161[30] , \Level1Out171[28] , 
        \Level32Out192[28] , \Level1Out127[30] , \Level1Out152[19] , 
        \Level8Out136[26] , \Level1Out171[31] , \ScanLink240[4] , 
        \Level32Out192[31] , \Level8Out160[27] , \Level1Out9[0] , 
        \ScanLink17[30] , \ScanLink41[28] , \Level1Out42[6] , 
        \Level1Out127[29] , \Level2Out168[19] , \ScanLink120[1] , 
        \Level2Out36[9] , \ScanLink17[29] , \ScanLink34[18] , \ScanLink41[31] , 
        \ScanLink62[19] , \ScanLink195[0] , \ScanLink209[19] , 
        \Level8Out96[21] , \Level1Out15[21] , \Level1Out23[24] , 
        \Level1Out56[14] , \Level1Out75[25] , \ScanLink79[4] , 
        \Level2Load172[0] , \Level8Out208[17] , \ScanLink227[3] , 
        \Level2Out200[29] , \Level1Out219[18] , \Level2Out200[30] , 
        \Level4Out64[0] , \Level1Out25[1] , \Level1Out43[20] , 
        \Level1Out36[10] , \Level1Out60[11] , \ScanLink147[6] , 
        \Level1Out26[2] , \ScanLink144[5] , \Level1Out179[2] , 
        \ScanLink224[0] , \Level1Out219[7] , \Level8Out136[15] , 
        \ScanLink67[8] , \ScanLink99[18] , \Level8Out160[14] , 
        \Level1Out84[11] , \Level1Out91[25] , \Level1Load163[0] , 
        \ScanLink196[3] , \Level2Out116[1] , \Level1Out204[8] , 
        \Level1Out172[9] , \ScanLink180[7] , \Level2Out100[5] , 
        \ScanLink86[19] , \ScanLink152[1] , \ScanLink232[4] , 
        \Level8Out24[20] , \Level1Out4[5] , \Level1Out7[6] , \ScanLink15[8] , 
        \Level1Out29[11] , \Level1Out30[6] , \Level1Out33[5] , 
        \ScanLink231[7] , \Level2Out44[9] , \Level8Out72[21] , 
        \Level4Out72[4] , \Level1Out49[15] , \ScanLink151[2] , 
        \ScanLink235[29] , \ScanLink240[19] , \Level2Out88[3] , 
        \ScanLink216[18] , \ScanLink235[30] , \Level1Out225[31] , 
        \Level1Out225[28] , \Level1Out250[18] , \Level4Out188[28] , 
        \Level4Out188[31] , \Level1Out206[19] , \Level1Out54[2] , 
        \ScanLink128[30] , \ScanLink183[4] , \Level8Out184[14] , 
        \ScanLink256[0] , \Level8Out24[13] , \Level8Out72[12] , 
        \ScanLink128[29] , \ScanLink136[5] , \Level1Out138[31] , 
        \Level2Out154[29] , \Level1Out29[22] , \Level1Out84[22] , 
        \Level2Out102[31] , \Level2Out164[1] , \Level1Out86[4] , 
        \Level1Out138[28] , \Level2Out154[30] , \Level2Out102[28] , 
        \Level1Out91[16] , \Level1Load111[0] , \Level2Out204[4] , 
        \Level1Out195[31] , \Level8Out184[27] , \Level1Out36[8] , 
        \Level1Out49[26] , \ScanLink128[9] , \Level1Out195[28] , 
        \Level1Out57[1] , \Level1Out85[7] , \Level1Out108[1] , 
        \ScanLink135[6] , \ScanLink185[30] , \ScanLink255[3] , 
        \Level32Out64[3] , \Level2Out56[18] , \Level2Load100[0] , 
        \Level4Out16[0] , \ScanLink185[29] , \ScanLink77[2] , \Level1Out98[8] , 
        \ScanLink98[12] , \ScanLink115[20] , \ScanLink136[11] , 
        \ScanLink143[21] , \Level1Out174[7] , \ScanLink229[5] , 
        \ScanLink100[14] , \ScanLink160[10] , \Level1Out110[15] , 
        \ScanLink123[25] , \ScanLink149[0] , \ScanLink175[24] , 
        \Level2Out90[10] , \Level2Out90[1] , \ScanLink156[15] , 
        \ScanLink186[9] , \Level1Out214[2] , \Level4Out4[26] , 
        \Level1Out126[10] , \Level1Out133[24] , \Level1Out165[25] , 
        \Level1Out169[8] , \Level1Out146[14] , \Level1Out105[21] , 
        \Level1Out153[20] , \Level2Out42[7] , \Level1Out170[11] , 
        \ScanLink198[5] , \Level1Out218[12] , \ScanLink237[9] , 
        \Level2Out118[7] , \Level2Out222[12] , \Level4Out132[8] , 
        \Level4Out196[23] , \Level4Out80[10] , \Level1Out9[20] , 
        \ScanLink10[5] , \ScanLink13[6] , \ScanLink16[23] , \ScanLink63[13] , 
        \Level2Out192[21] , \Level2Out214[17] , \Level2Out242[16] , 
        \Level1Out177[4] , \ScanLink20[26] , \ScanLink35[12] , 
        \ScanLink40[22] , \ScanLink74[1] , \Level2Out28[24] , \ScanLink55[16] , 
        \ScanLink208[13] , \Level1Out217[1] , \Level2Out48[20] , 
        \Level8Out112[7] , \Level16Out96[5] , \Level1Out28[4] , 
        \ScanLink76[27] , \ScanLink100[27] , \Level1Out105[12] , 
        \Level1Out126[23] , \Level1Out153[13] , \Level16Out64[30] , 
        \Level1Out170[22] , \Level16Out32[28] , \Level16Out64[29] , 
        \Level1Out110[26] , \Level1Out165[16] , \Level16Out32[31] , 
        \Level1Out110[3] , \Level1Out133[17] , \Level1Out146[27] , 
        \Level2Out26[3] , \ScanLink175[17] , \ScanLink156[26] , 
        \Level2Out90[23] , \Level4Out148[0] , \ScanLink98[21] , 
        \ScanLink123[16] , \ScanLink136[22] , \ScanLink143[12] , 
        \Level4Out4[15] , \Level2Out6[1] , \Level4Out228[5] , 
        \ScanLink115[13] , \ScanLink160[23] , \Level1Out10[30] , 
        \Level1Out10[29] , \ScanLink12[21] , \Level1Out14[18] , 
        \ScanLink16[10] , \ScanLink20[15] , \Level2Out48[13] , 
        \ScanLink55[25] , \ScanLink208[20] , \ScanLink76[14] , 
        \Level1Out113[0] , \Level8Out216[6] , \ScanLink35[21] , 
        \ScanLink63[20] , \Level1Out83[9] , \Level8Out176[3] , 
        \Level1Out37[30] , \ScanLink40[11] , \Level2Out28[17] , 
        \Level2Out214[24] , \Level4Out80[23] , \ScanLink24[24] , 
        \Level1Out37[29] , \Level1Out61[28] , \Level4Load36[0] , 
        \Level1Out42[19] , \Level1Out61[31] , \Level2Out192[12] , 
        \Level2Out242[25] , \ScanLink51[14] , \ScanLink133[8] , 
        \Level1Out218[21] , \Level2Out222[21] , \Level16Out192[4] , 
        \Level4Out4[9] , \Level4Out196[10] , \Level4Out236[9] , 
        \Level8Out152[5] , \ScanLink67[11] , \Level1Out68[6] , 
        \ScanLink72[25] , \Level1Out137[6] , \Level8Out232[0] , 
        \ScanLink31[10] , \ScanLink34[3] , \ScanLink44[20] , \ScanLink219[25] , 
        \Level1Out46[31] , \Level1Out65[19] , \Level1Out46[28] , 
        \Level2Out8[18] , \Level4Out84[12] , \Level2Out210[15] , 
        \Level1Out75[9] , \Level1Out209[24] , \Level2Out246[14] , 
        \Level2Out196[23] , \Level1Out33[18] , \Level2Out158[5] , 
        \Level2Out226[10] , \Level2Out238[0] , \ScanLink37[0] , 
        \ScanLink89[24] , \Level1Out101[23] , \Level1Out122[12] , 
        \Level4Out192[21] , \Level1Out157[22] , \Level8Out8[9] , 
        \Level2Out118[12] , \ScanLink104[16] , \Level1Out114[17] , 
        \Level1Out174[13] , \Level1Out137[26] , \Level1Out161[27] , 
        \Level1Out142[16] , \Level2Out178[16] , \Level64Out128[19] , 
        \Level2Out94[12] , \ScanLink171[26] , \ScanLink109[2] , 
        \ScanLink127[27] , \ScanLink152[17] , \Level1Out254[0] , 
        \Level4Out0[24] , \ScanLink111[22] , \ScanLink132[13] , 
        \Level1Out134[5] , \ScanLink147[23] , \Level2Out146[9] , 
        \Level1Load149[0] , \ScanLink164[12] , \Level2Out226[23] , 
        \Level1Out9[13] , \Level4Out192[12] , \Level1Out1[1] , \ScanLink4[24] , 
        \ScanLink4[17] , \ScanLink9[9] , \ScanLink12[12] , \ScanLink82[1] , 
        \Level2Out210[26] , \Level4Out84[21] , \Level1Out181[4] , 
        \Level2Out196[10] , \Level1Out209[17] , \Level2Out246[27] , 
        \Level1Out14[0] , \Level1Out17[3] , \ScanLink24[17] , \ScanLink31[23] , 
        \ScanLink67[22] , \Level8Out136[1] , \ScanLink44[13] , 
        \Level1Out233[7] , \ScanLink50[7] , \ScanLink219[16] , 
        \Level1Out38[27] , \ScanLink51[27] , \ScanLink53[4] , \ScanLink72[16] , 
        \Level1Out153[2] , \ScanLink89[17] , \ScanLink111[11] , 
        \ScanLink132[20] , \ScanLink147[10] , \Level1Out230[4] , 
        \ScanLink164[21] , \Level2Out242[8] , \ScanLink171[15] , 
        \ScanLink104[25] , \Level1Out150[1] , \Level2Out94[21] , 
        \ScanLink152[24] , \Level4Out108[2] , \Level1Out58[23] , 
        \ScanLink81[2] , \Level1Out114[24] , \ScanLink127[14] , 
        \Level2Load158[0] , \Level1Out161[14] , \ScanLink170[9] , 
        \Level4Out0[17] , \Level1Out122[21] , \Level1Out137[15] , 
        \Level1Out142[25] , \Level2Out66[1] , \Level2Out178[25] , 
        \Level1Out157[11] , \Level2Out118[21] , \Level8Out248[8] , 
        \Level1Out182[7] , \Level128Load0[0] , \Level1Out101[10] , 
        \Level1Out174[20] , \Level2Out188[28] , \Level16Out112[28] , 
        \Level16Out144[30] , \Level1Out191[19] , \Level2Out188[31] , 
        \Level16Out112[31] , \Level16Out144[29] , \Level1Out70[4] , 
        \Level1Out73[7] , \Level1Out131[8] , \ScanLink111[0] , 
        \Level2Out52[30] , \ScanLink112[3] , \ScanLink181[18] , 
        \Level2Out52[29] , \Level4Out32[6] , \ScanLink79[30] , 
        \Level1Out80[13] , \Level1Out149[30] , \ScanLink159[31] , 
        \ScanLink159[28] , \Level8Out16[27] , \Level2Out192[1] , 
        \Level8Out40[26] , \Level1Out95[27] , \Level1Out149[29] , 
        \Level2Out150[18] , \Level32Out32[15] , \Level128Out0[26] , 
        \Level2Out106[19] , \Level32Out64[14] , \Level2Out220[2] , 
        \Level16Out48[16] , \ScanLink175[4] , \Level2Out140[7] , 
        \Level1Out228[6] , \Level1Load35[0] , \Level1Out38[14] , 
        \ScanLink79[29] , \Level4Load100[0] , \Level1Out148[3] , 
        \Level1Out202[31] , \ScanLink212[30] , \ScanLink212[29] , 
        \ScanLink215[1] , \ScanLink231[18] , \ScanLink244[28] , 
        \Level4Out56[2] , \ScanLink244[31] , \Level1Out202[28] , 
        \Level1Out221[19] , \Level1Out235[9] , \Level1Out254[29] , 
        \Level2Out238[31] , \Level1Out254[30] , \Level2Out238[28] , 
        \ScanLink56[9] , \Level1Out58[10] , \Level4Out84[4] , \ScanLink99[0] , 
        \Level1Out80[20] , \Level1Out95[14] , \Level2Out244[6] , 
        \Level16Out48[25] , \Level2Out124[3] , \Level32Out32[26] , 
        \Level128Out0[15] , \Level1Out199[6] , \Level32Out64[27] , 
        \ScanLink48[5] , \ScanLink82[31] , \ScanLink82[28] , \Level8Out16[14] , 
        \ScanLink176[7] , \Level8Out40[15] , \Level1Out184[9] , 
        \ScanLink216[2] , \Level1Out52[5] , \ScanLink130[2] , 
        \Level8Out168[6] , \ScanLink250[7] , \Level8Out208[3] , 
        \Level1Out14[11] , \ScanLink16[19] , \ScanLink35[31] , 
        \Level1Out80[3] , \ScanLink98[31] , \Level16Out32[21] , 
        \Level16Out64[20] , \Level128Out0[3] , \ScanLink98[28] , 
        \Level2Out6[8] , \Level2Out162[6] , \Level2Out202[3] , 
        \Level4Out148[9] , \Level1Out22[14] , \ScanLink35[28] , 
        \ScanLink63[29] , \Level1Out83[0] , \Level2Out38[6] , \ScanLink40[18] , 
        \ScanLink63[30] , \Level1Out51[6] , \Level1Out113[9] , 
        \ScanLink208[29] , \ScanLink208[30] , \Level4Out184[3] , 
        \Level1Out57[24] , \Level2Out222[28] , \Level1Out74[15] , 
        \ScanLink133[1] , \Level1Out218[28] , \Level4Out4[0] , 
        \Level2Out222[31] , \Level4Out196[19] , \Level4Out236[0] , 
        \Level1Out218[31] , \Level1Out36[1] , \Level1Out37[20] , 
        \Level1Out61[21] , \Level1Out42[10] , \ScanLink253[4] , 
        \ScanLink115[30] , \ScanLink136[18] , \ScanLink149[9] , 
        \Level2Out90[19] , \Level4Out156[5] , \Level2Out90[8] , 
        \ScanLink186[0] , \ScanLink115[29] , \ScanLink143[28] , 
        \Level2Out106[2] , \ScanLink143[31] , \ScanLink160[19] , 
        \Level1Out105[31] , \Level1Out126[19] , \Level1Out153[29] , 
        \Level16Out32[12] , \Level1Out6[27] , \Level1Out14[22] , 
        \Level1Out61[12] , \Level1Out105[28] , \ScanLink154[6] , 
        \Level8Out80[5] , \Level1Out153[30] , \Level1Out170[18] , 
        \Level1Out209[4] , \Level1Out169[1] , \Level16Out64[13] , 
        \ScanLink234[3] , \ScanLink157[5] , \Level2Out192[31] , 
        \ScanLink15[1] , \Level1Out22[27] , \Level1Out35[2] , 
        \Level1Out42[23] , \Level4Out80[19] , \Level4Out252[4] , 
        \Level1Out37[13] , \Level1Out57[17] , \ScanLink237[0] , 
        \Level2Out192[28] , \Level4Out132[1] , \Level1Out49[4] , 
        \ScanLink69[7] , \ScanLink74[8] , \Level1Out74[26] , 
        \Level1Load170[0] , \ScanLink185[3] , \Level1Out217[8] , 
        \Level2Out48[30] , \Level2Out48[29] , \ScanLink86[23] , 
        \Level2Out20[4] , \ScanLink93[17] , \ScanLink128[20] , 
        \ScanLink148[24] , \ScanLink256[9] , \Level2Out162[25] , 
        \Level1Out158[25] , \Level2Out0[6] , \Level2Out134[24] , 
        \ScanLink16[2] , \Level1Out115[7] , \Level1Out116[4] , 
        \Level1Out138[21] , \Level2Out154[20] , \Level2Out164[8] , 
        \ScanLink128[0] , \Level1Out180[15] , \Level2Out102[21] , 
        \Level1Out225[12] , \Level1Out206[23] , \Level1Out250[22] , 
        \Level4Out188[12] , \Level16Out176[14] , \Level1Out213[17] , 
        \ScanLink248[5] , \Level1Out195[21] , \Level1Out230[26] , 
        \Level1Out245[16] , \Level1Out57[8] , \ScanLink203[16] , 
        \Level2Out36[15] , \ScanLink68[16] , \Level1Out98[1] , 
        \ScanLink185[20] , \ScanLink220[27] , \Level1Out108[8] , 
        \ScanLink255[17] , \Level2Out60[14] , \ScanLink71[5] , 
        \Level1Out84[18] , \ScanLink190[14] , \ScanLink216[22] , 
        \ScanLink235[13] , \ScanLink240[23] , \Level4Out16[9] , 
        \Level2Out56[11] , \Level1Out138[12] , \Level1Out212[5] , 
        \Level2Out102[12] , \Level2Out154[13] , \Level1Out158[16] , 
        \Level1Out172[0] , \Level2Out96[6] , \Level2Load60[0] , 
        \Level2Out134[17] , \Level2Out162[16] , \ScanLink148[17] , 
        \ScanLink152[8] , \Level8Out72[31] , \Level8Out24[29] , 
        \Level1Out2[25] , \Level1Out2[2] , \ScanLink68[25] , \ScanLink86[10] , 
        \ScanLink93[24] , \Level2Out44[0] , \Level8Out24[30] , 
        \Level8Out72[28] , \ScanLink128[13] , \ScanLink240[10] , 
        \ScanLink190[27] , \ScanLink235[20] , \Level2Out56[22] , 
        \Level1Out6[14] , \Level1Out29[18] , \ScanLink185[13] , 
        \ScanLink203[25] , \ScanLink216[11] , \Level2Out36[26] , 
        \ScanLink220[14] , \ScanLink255[24] , \Level2Out60[27] , 
        \Level1Out211[6] , \Level1Out213[24] , \Level1Out245[25] , 
        \ScanLink19[24] , \ScanLink72[6] , \Level1Out195[12] , 
        \Level1Out230[15] , \Level1Out250[11] , \Level4Out188[21] , 
        \Level1Out171[3] , \Level1Out180[26] , \Level1Out225[21] , 
        \Level1Out187[3] , \ScanLink194[16] , \Level1Out206[10] , 
        \ScanLink215[8] , \Level16Out176[27] , \ScanLink231[11] , 
        \ScanLink56[0] , \Level1Out58[19] , \ScanLink79[20] , \ScanLink84[6] , 
        \ScanLink244[21] , \ScanLink181[22] , \ScanLink207[14] , 
        \ScanLink212[20] , \Level2Out52[13] , \ScanLink224[25] , 
        \Level2Out32[17] , \Level1Out155[5] , \ScanLink251[15] , 
        \Level2Out64[16] , \ScanLink208[7] , \Level1Out217[15] , 
        \Level2Out188[12] , \Level16Out112[12] , \ScanLink99[9] , 
        \Level1Out191[23] , \Level1Out234[24] , \Level16Out144[13] , 
        \Level32Out192[3] , \Level1Out2[16] , \ScanLink9[0] , \ScanLink55[3] , 
        \ScanLink168[2] , \Level1Out184[17] , \Level1Out241[14] , 
        \Level1Out221[10] , \Level1Out202[21] , \Level1Out235[0] , 
        \Level1Out254[20] , \Level2Out238[21] , \Level1Out80[30] , 
        \Level1Out80[29] , \Level2Out150[22] , \Level1Out149[13] , 
        \Level1Out156[6] , \Level2Out106[23] , \ScanLink87[5] , 
        \Level1Out129[17] , \Level4Out48[7] , \Level1Out236[3] , 
        \Level2Out166[27] , \Level2Out130[26] , \ScanLink97[15] , 
        \ScanLink139[16] , \Level1Out184[0] , \Level2Load96[0] , 
        \Level1Out14[9] , \ScanLink32[4] , \ScanLink82[21] , \Level2Out60[6] , 
        \ScanLink159[12] , \Level1Out254[13] , \Level1Out131[1] , 
        \Level1Out184[24] , \Level1Out221[23] , \Level2Out238[12] , 
        \Level1Out202[12] , \Level1Out217[26] , \Level2Out188[21] , 
        \Level16Out112[21] , \Level1Out251[4] , \Level8Load112[0] , 
        \Level1Out10[13] , \ScanLink19[17] , \ScanLink79[13] , 
        \ScanLink181[11] , \Level1Out191[10] , \Level1Out234[17] , 
        \Level1Out241[27] , \ScanLink207[27] , \Level16Out144[20] , 
        \ScanLink224[16] , \ScanLink251[26] , \Level2Out32[24] , 
        \Level2Out64[25] , \ScanLink31[7] , \ScanLink82[12] , \ScanLink111[9] , 
        \ScanLink194[25] , \ScanLink244[12] , \ScanLink231[22] , 
        \Level2Out52[20] , \ScanLink212[13] , \ScanLink97[26] , 
        \ScanLink139[25] , \ScanLink159[21] , \Level2Out192[8] , 
        \Level1Load128[0] , \Level1Out129[24] , \Level1Out132[2] , 
        \Level2Out166[14] , \Level2Out130[15] , \Level1Out149[20] , 
        \Level1Out252[7] , \Level2Out106[10] , \Level2Out150[11] , 
        \Level4Out84[28] , \Level1Out11[4] , \Level1Out33[22] , 
        \Level1Out65[23] , \ScanLink82[8] , \Level2Out8[22] , 
        \Level2Out196[19] , \Level4Out84[31] , \Level1Out46[12] , 
        \ScanLink213[6] , \Level4Out116[7] , \Level1Out26[16] , 
        \Level2Load226[0] , \ScanLink0[15] , \Level1Out53[26] , 
        \Level1Out70[17] , \ScanLink173[3] , \Level1Load186[0] , 
        \ScanLink111[18] , \ScanLink132[29] , \ScanLink147[19] , 
        \Level1Out150[8] , \Level2Out78[4] , \Level8Out136[8] , 
        \Level1Load237[0] , \Level2Out94[28] , \Level2Out122[4] , 
        \Level2Out94[31] , \ScanLink164[31] , \ScanLink164[28] , 
        \ScanLink132[30] , \Level2Out242[1] , \Level1Out157[18] , 
        \Level1Out174[30] , \Level8Out248[1] , \ScanLink210[5] , 
        \Level2Out118[28] , \ScanLink12[31] , \ScanLink12[28] , 
        \Level1Out12[7] , \Level1Out101[19] , \Level1Out122[28] , 
        \Level1Out174[29] , \Level2Out118[31] , \Level1Out122[31] , 
        \ScanLink170[0] , \Level8Out128[4] , \Level64Out128[23] , 
        \ScanLink44[30] , \Level2Out66[8] , \ScanLink67[18] , 
        \Level8Out232[9] , \ScanLink44[29] , \ScanLink31[19] , 
        \Level1Out53[15] , \Level8Load32[0] , \ScanLink0[26] , 
        \Level1Out9[30] , \Level2Load38[0] , \Level4Out192[31] , 
        \Level1Out9[29] , \Level1Out26[25] , \Level2Out226[19] , 
        \ScanLink29[5] , \Level1Out70[24] , \Level4Out172[3] , 
        \Level4Out192[28] , \Level1Out10[20] , \Level1Out65[10] , 
        \ScanLink117[7] , \Level2Out8[11] , \Level4Out212[6] , 
        \Level1Out33[11] , \Level1Out46[21] , \Level1Out75[0] , 
        \Level1Out76[3] , \Level1Out129[3] , \Level2Out194[6] , 
        \Level2Out238[9] , \Level64Out128[10] , \Level8Out8[0] , 
        \ScanLink37[9] , \ScanLink114[4] , \Level1Out249[6] , 
        \Level1Out39[24] , \Level1Load54[0] , \Level1Out60[7] , 
        \Level1Out81[10] , \Level1Out94[24] , \Level1Out254[9] , 
        \Level2Out146[0] , \Level2Out226[5] , \Level1Out122[8] , 
        \Level1Load245[0] , \Level4Out120[30] , \Level4Out176[28] , 
        \Level2Out150[4] , \Level2Out230[1] , \Level4Out120[29] , 
        \Level4Out176[31] , \ScanLink83[18] , \Level2Out182[2] , 
        \Level1Out63[4] , \ScanLink78[19] , \ScanLink102[0] , \Level2Out14[8] , 
        \ScanLink101[3] , \Level4Out164[7] , \ScanLink213[19] , 
        \ScanLink230[31] , \Level4Out204[2] , \Level2Load254[0] , 
        \ScanLink230[28] , \ScanLink245[18] , \ScanLink58[6] , 
        \Level1Out59[20] , \Level1Out203[18] , \Level1Out220[30] , 
        \Level1Out220[29] , \Level1Out255[19] , \Level2Out2[24] , 
        \Level8Out0[8] , \Level8Out144[8] , \Level8Out224[12] , 
        \ScanLink206[1] , \ScanLink158[18] , \ScanLink166[4] , 
        \Level1Out189[5] , \Level2Out172[19] , \Level4Out60[31] , 
        \ScanLink0[18] , \ScanLink1[8] , \ScanLink4[5] , \ScanLink7[6] , 
        \Level1Load26[0] , \ScanLink45[9] , \Level1Out148[19] , 
        \Level4Out36[29] , \Level4Out60[28] , \Level2Out134[0] , 
        \Level1Out59[13] , \Level1Out81[23] , \ScanLink89[3] , 
        \Level1Out94[17] , \Level1Out226[9] , \Level2Out124[18] , 
        \Level4Out36[30] , \Level2Out254[5] , \Level1Out190[30] , 
        \Level1Out190[29] , \Level4Out248[19] , \Level8Out224[21] , 
        \Level8Out240[9] , \Level1Out8[23] , \ScanLink27[3] , 
        \Level1Out39[17] , \Level64Out128[1] , \ScanLink110[21] , 
        \Level1Out124[6] , \Level1Out158[0] , \ScanLink178[8] , 
        \Level8Load40[0] , \Level2Out2[17] , \Level2Out26[29] , 
        \Level2Out70[31] , \ScanLink165[7] , \ScanLink180[31] , 
        \ScanLink180[28] , \Level1Out197[9] , \Level2Out26[30] , 
        \ScanLink205[2] , \Level2Out70[28] , \Level4Out100[3] , 
        \Level1Out238[5] , \Level2Out80[25] , \ScanLink165[11] , 
        \Level1Out66[9] , \ScanLink88[27] , \ScanLink105[15] , 
        \ScanLink119[1] , \ScanLink126[24] , \ScanLink133[10] , 
        \ScanLink146[20] , \ScanLink153[14] , \Level1Out244[3] , 
        \ScanLink170[25] , \Level1Out100[20] , \Level1Out115[14] , 
        \Level1Out136[25] , \Level1Out139[9] , \Level1Out143[15] , 
        \Level4Out48[15] , \Level4Out168[23] , \Level1Out160[24] , 
        \Level1Out175[10] , \Level4Out108[27] , \Level1Out123[11] , 
        \Level1Out156[21] , \Level2Out12[6] , \Level4Out28[11] , 
        \Level2Out148[6] , \Level2Out204[22] , \ScanLink13[22] , 
        \ScanLink24[0] , \ScanLink45[23] , \Level1Out208[27] , 
        \Level2Out182[14] , \Level2Out252[23] , \Level4Out236[25] , 
        \Level2Out228[3] , \Level2Out232[27] , \Level4Out200[20] , 
        \ScanLink218[26] , \ScanLink30[13] , \ScanLink66[12] , 
        \Level1Load88[0] , \Level2Out58[15] , \Level1Out127[5] , 
        \ScanLink25[27] , \ScanLink50[17] , \ScanLink73[26] , \Level1Out78[5] , 
        \Level8Out8[16] , \Level1Out247[0] , \Level2Out38[11] , 
        \ScanLink43[7] , \ScanLink91[1] , \Level1Out100[13] , 
        \Level1Out175[23] , \Level4Out108[14] , \Level1Out115[27] , 
        \Level1Out123[22] , \Level1Out156[12] , \Level1Out192[4] , 
        \Level4Out28[22] , \Level1Out136[16] , \Level1Out143[26] , 
        \Level8Out152[30] , \Level2Out76[2] , \Level8Out104[28] , 
        \Level1Out160[17] , \Level4Out48[26] , \Level8Out152[29] , 
        \Level4Out168[10] , \Level8Out104[31] , \ScanLink153[27] , 
        \ScanLink88[14] , \ScanLink126[17] , \ScanLink170[16] , 
        \ScanLink105[26] , \Level1Out140[2] , \ScanLink110[12] , 
        \ScanLink165[22] , \Level2Out80[16] , \ScanLink133[23] , 
        \ScanLink146[13] , \Level1Out220[7] , \Level1Out143[1] , 
        \Level1Out2[31] , \Level1Out2[28] , \Level1Out8[10] , 
        \Level1Out11[19] , \ScanLink13[11] , \ScanLink25[14] , \ScanLink40[4] , 
        \ScanLink73[15] , \Level4Out92[9] , \Level8Out8[25] , \ScanLink30[20] , 
        \ScanLink50[24] , \Level2Out38[22] , \Level16Out0[0] , 
        \ScanLink45[10] , \Level1Out223[4] , \Level2Out58[26] , 
        \Level8Load160[0] , \ScanLink218[15] , \Level1Out32[31] , 
        \Level1Out32[28] , \ScanLink66[21] , \Level4Out200[13] , 
        \Level1Out47[18] , \Level1Out64[30] , \Level1Out191[7] , 
        \Level2Out232[14] , \Level1Out208[14] , \Level1Out64[29] , 
        \ScanLink92[2] , \ScanLink163[9] , \Level1Load9[0] , \Level1Out9[9] , 
        \Level1Out38[7] , \Level2Out182[27] , \Level2Out204[11] , 
        \Level4Out236[16] , \Level2Out252[10] , \ScanLink54[15] , 
        \ScanLink77[24] , \Level8Out96[28] , \ScanLink195[9] , 
        \Level1Out207[2] , \ScanLink209[10] , \Level8Out96[31] , 
        \Level1Out15[31] , \ScanLink17[20] , \ScanLink21[25] , 
        \ScanLink34[11] , \ScanLink41[21] , \ScanLink64[2] , \ScanLink62[10] , 
        \Level1Out167[7] , \Level1Out25[8] , \Level1Out43[29] , 
        \Level1Out15[28] , \Level1Out36[19] , \Level2Out236[25] , 
        \Level1Out43[30] , \ScanLink188[6] , \Level4Out204[22] , 
        \Level1Out60[18] , \Level4Out252[23] , \ScanLink17[13] , 
        \ScanLink34[22] , \ScanLink67[1] , \ScanLink99[11] , \ScanLink101[17] , 
        \Level1Out104[22] , \Level1Out219[11] , \Level2Out108[4] , 
        \Level2Out200[20] , \Level4Out232[27] , \Level2Out186[16] , 
        \Level4Out64[9] , \Level1Out111[16] , \Level1Out127[13] , 
        \Level1Out171[12] , \Level2Out168[23] , \Level32Out192[12] , 
        \Level1Out132[27] , \Level1Out152[23] , \Level2Out52[4] , 
        \Level1Out147[17] , \ScanLink224[9] , \Level2Out108[27] , 
        \Level16Out192[27] , \ScanLink122[26] , \ScanLink159[3] , 
        \Level1Out164[26] , \ScanLink157[16] , \Level1Out204[1] , 
        \ScanLink114[23] , \Level1Out164[4] , \ScanLink174[27] , 
        \Level2Out80[2] , \ScanLink239[6] , \Level2Out84[27] , 
        \ScanLink161[13] , \ScanLink137[12] , \ScanLink142[22] , 
        \Level1Out219[22] , \Level2Out116[8] , \Level2Out186[25] , 
        \Level2Out200[13] , \Level4Out232[14] , \Level2Out236[16] , 
        \Level4Out204[11] , \Level4Out252[10] , \ScanLink41[12] , 
        \ScanLink62[23] , \Level1Out14[4] , \ScanLink18[4] , \Level1Out20[5] , 
        \ScanLink21[16] , \ScanLink77[17] , \Level1Out103[3] , 
        \Level1Out23[6] , \Level1Out28[12] , \ScanLink54[26] , 
        \ScanLink209[23] , \Level1Out90[9] , \ScanLink99[22] , 
        \Level1Out100[0] , \ScanLink114[10] , \ScanLink161[20] , 
        \ScanLink122[15] , \ScanLink137[21] , \ScanLink142[11] , 
        \Level2Out84[14] , \Level2Out212[9] , \ScanLink157[25] , 
        \ScanLink174[14] , \Level2Load12[0] , \ScanLink101[24] , 
        \Level1Out104[11] , \Level1Out111[25] , \ScanLink120[8] , 
        \Level1Out132[14] , \Level1Out147[24] , \Level2Out36[0] , 
        \Level2Out108[14] , \Level16Out192[14] , \Level1Out164[15] , 
        \Level1Out171[21] , \Level32Out192[21] , \Level1Out127[20] , 
        \Level1Out152[10] , \ScanLink193[7] , \Level2Out168[10] , 
        \Level1Out194[18] , \Level16Out80[13] , \Level16Out80[8] , 
        \Level1Out48[16] , \Level1Out161[9] , \Level8Out240[14] , 
        \ScanLink141[1] , \Level2Out6[26] , \Level8Out216[15] , 
        \Level128Out128[15] , \Level2Out22[18] , \Level4Out244[0] , 
        \ScanLink184[19] , \ScanLink221[4] , \Level2Out74[19] , 
        \Level2Out98[0] , \Level8Out88[23] , \Level4Out124[5] , 
        \Level1Out28[21] , \Level1Out47[2] , \Level1Out85[12] , 
        \ScanLink129[19] , \ScanLink142[2] , \Level8Out96[1] , 
        \Level1Out139[18] , \ScanLink222[7] , \Level2Out120[30] , 
        \Level4Out32[18] , \Level2Out176[28] , \ScanLink190[4] , 
        \Level2Out120[29] , \Level1Out90[26] , \Level2Out176[31] , 
        \Level4Out64[19] , \Level8Out128[17] , \Level2Out110[6] , 
        \Level1Out48[25] , \Level1Out118[2] , \ScanLink125[5] , 
        \ScanLink217[28] , \Level4Out220[4] , \ScanLink241[30] , 
        \Level128Out128[26] , \Level8Out88[10] , \ScanLink217[31] , 
        \ScanLink234[19] , \ScanLink245[0] , \ScanLink241[29] , 
        \Level4Out140[1] , \Level1Out95[4] , \Level1Out207[29] , 
        \Level2Out248[19] , \Level1Load102[0] , \Level1Out251[31] , 
        \Level1Out207[30] , \Level8Out240[27] , \Level1Out224[18] , 
        \Level1Out251[28] , \Level8Out216[26] , \Level2Out6[15] , 
        \Level4Out192[7] , \Level16Out80[20] , \Level1Out44[1] , 
        \Level1Out85[21] , \Level1Out90[15] , \Level4Out172[19] , 
        \Level1Out96[7] , \Level2Out174[2] , \Level2Out214[7] , 
        \Level4Out124[18] , \Level8Out128[24] , \ScanLink87[30] , 
        \ScanLink126[6] , \ScanLink87[29] , \ScanLink246[3] , \ScanLink32[9] , 
        \Level1Out38[23] , \Level1Out70[0] , \Level1Out80[17] , 
        \Level1Out95[23] , \Level1Out129[30] , \Level2Out130[18] , 
        \Level1Out129[29] , \Level2Out140[3] , \Level16Out48[12] , 
        \Level2Out166[19] , \Level2Out220[6] , \Level32Out64[10] , 
        \Level2Out192[5] , \Level8Out40[22] , \Level32Out32[11] , 
        \Level128Out0[22] , \Level8Out16[23] , \Level1Out73[3] , 
        \ScanLink111[4] , \ScanLink112[7] , \ScanLink139[31] , 
        \ScanLink139[28] , \Level2Out32[30] , \Level2Out64[28] , 
        \Level2Out32[29] , \Level2Out64[31] , \Level4Out32[2] , 
        \ScanLink194[31] , \Level4Load164[0] , \ScanLink194[28] , 
        \Level1Out184[30] , \ScanLink48[1] , \Level1Load51[0] , 
        \Level1Out184[29] , \Level1Out58[27] , \Level1Out251[9] , 
        \ScanLink87[8] , \ScanLink97[18] , \ScanLink216[6] , 
        \Level8Load208[0] , \ScanLink176[3] , \Level8Out16[10] , 
        \Level8Out40[11] , \Level1Out80[24] , \Level1Load183[0] , 
        \Level1Out199[2] , \Level2Out124[7] , \Level32Out32[22] , 
        \Level32Out64[23] , \Level128Out0[11] , \Level1Out95[10] , 
        \ScanLink99[4] , \Level2Out244[2] , \Level16Out48[21] , 
        \Level1Out234[29] , \Level2Load192[0] , \Level1Out58[14] , 
        \Level1Out155[8] , \Level1Load232[0] , \Level1Out241[19] , 
        \Level1Out234[30] , \Level1Out217[18] , \Level1Out9[24] , 
        \Level1Out17[7] , \ScanLink19[30] , \Level1Out38[10] , 
        \Level4Out84[0] , \ScanLink19[29] , \Level1Out148[7] , 
        \ScanLink215[5] , \Level4Out56[6] , \ScanLink224[28] , 
        \Level1Out26[31] , \ScanLink29[8] , \ScanLink37[4] , \ScanLink111[26] , 
        \Level1Out134[1] , \ScanLink175[0] , \ScanLink207[19] , 
        \ScanLink224[31] , \ScanLink251[18] , \Level1Out228[2] , 
        \ScanLink164[16] , \Level1Out70[29] , \ScanLink89[20] , 
        \ScanLink104[12] , \ScanLink109[6] , \ScanLink132[17] , 
        \ScanLink147[27] , \ScanLink127[23] , \ScanLink152[13] , 
        \Level1Out254[4] , \Level4Out0[20] , \ScanLink171[22] , 
        \Level2Out94[16] , \Level2Out226[8] , \Level1Out101[27] , 
        \Level1Out114[13] , \Level1Out137[22] , \Level1Out142[12] , 
        \Level2Out178[12] , \Level1Out161[23] , \ScanLink114[9] , 
        \Level1Out122[16] , \Level1Out174[17] , \Level1Out157[26] , 
        \Level2Out118[16] , \Level2Out158[1] , \Level4Out192[25] , 
        \ScanLink12[25] , \Level1Out26[28] , \Level1Out53[18] , 
        \Level1Out70[30] , \ScanLink31[14] , \ScanLink34[7] , \ScanLink44[24] , 
        \Level1Out209[20] , \Level2Out226[14] , \Level2Out196[27] , 
        \Level2Out246[10] , \Level2Out210[11] , \Level2Out238[4] , 
        \Level4Out84[16] , \ScanLink219[21] , \ScanLink67[15] , 
        \Level1Out137[2] , \Level8Out232[4] , \ScanLink24[20] , 
        \ScanLink51[10] , \Level1Out68[2] , \ScanLink72[21] , 
        \Level8Out152[1] , \ScanLink81[6] , \Level1Out101[14] , 
        \Level1Out174[24] , \Level1Out157[15] , \Level1Out182[3] , 
        \ScanLink210[8] , \Level2Out118[25] , \ScanLink4[30] , \Level1Out4[1] , 
        \Level1Out9[17] , \ScanLink12[16] , \ScanLink24[13] , \ScanLink50[3] , 
        \ScanLink53[0] , \Level1Out114[20] , \Level1Out122[25] , 
        \Level1Out137[11] , \Level1Out142[21] , \Level2Out66[5] , 
        \Level2Out178[21] , \Level1Out161[10] , \Level8Out128[9] , 
        \ScanLink152[20] , \ScanLink72[12] , \ScanLink89[13] , 
        \ScanLink127[10] , \Level2Out122[9] , \ScanLink171[11] , 
        \Level4Out0[13] , \ScanLink104[21] , \Level1Out150[5] , 
        \ScanLink111[15] , \ScanLink164[25] , \Level2Out94[25] , 
        \Level4Out108[6] , \ScanLink132[24] , \ScanLink147[14] , 
        \Level1Out230[0] , \Level1Out153[6] , \ScanLink31[27] , 
        \ScanLink51[23] , \Level8Out136[5] , \ScanLink44[17] , 
        \Level1Out233[3] , \ScanLink219[12] , \ScanLink67[26] , 
        \Level2Out78[9] , \ScanLink82[5] , \Level1Out181[0] , 
        \Level2Out196[14] , \Level1Out209[13] , \Level2Out246[23] , 
        \Level2Out210[22] , \Level4Out84[25] , \Level4Out192[16] , 
        \Level1Out11[9] , \ScanLink16[27] , \ScanLink20[22] , \Level1Out28[0] , 
        \Level2Out226[27] , \ScanLink55[12] , \ScanLink76[23] , 
        \ScanLink208[17] , \Level1Out217[5] , \Level2Out48[24] , 
        \Level8Out112[3] , \Level16Out96[1] , \ScanLink35[16] , 
        \ScanLink40[26] , \ScanLink74[5] , \Level2Out28[20] , \ScanLink63[17] , 
        \Level1Out177[0] , \ScanLink157[8] , \ScanLink198[1] , 
        \Level2Out192[25] , \Level2Out242[12] , \Level1Out7[2] , 
        \Level1Out105[25] , \Level1Out218[16] , \Level2Out118[3] , 
        \Level2Out214[13] , \Level4Out80[14] , \Level4Out252[9] , 
        \Level4Load52[0] , \Level4Out196[27] , \Level2Out222[16] , 
        \Level1Out170[15] , \Level1Out209[9] , \Level8Out80[8] , 
        \ScanLink4[29] , \Level1Out126[14] , \Level1Out153[24] , 
        \Level2Out42[3] , \ScanLink10[1] , \ScanLink16[14] , \Level1Out22[19] , 
        \Level1Out57[30] , \ScanLink77[6] , \ScanLink98[16] , 
        \ScanLink100[10] , \Level1Out110[11] , \Level1Out133[20] , 
        \Level1Out146[10] , \ScanLink123[21] , \Level1Out165[21] , 
        \ScanLink149[4] , \ScanLink156[11] , \Level1Out214[6] , 
        \Level4Out4[22] , \Level2Out90[14] , \ScanLink115[24] , 
        \Level1Out174[3] , \ScanLink175[20] , \Level2Out90[5] , 
        \ScanLink229[1] , \ScanLink160[14] , \ScanLink136[15] , 
        \ScanLink143[25] , \Level4Out196[14] , \Level1Out74[18] , 
        \Level2Out222[25] , \ScanLink35[25] , \Level1Out57[29] , 
        \Level1Out218[25] , \ScanLink253[9] , \Level2Out192[16] , 
        \Level2Out214[20] , \Level2Out242[21] , \Level4Out156[8] , 
        \Level16Out192[0] , \Level4Out80[27] , \Level8Out176[7] , 
        \ScanLink40[15] , \Level2Out28[13] , \ScanLink63[24] , 
        \ScanLink76[10] , \Level1Out113[4] , \Level8Out216[2] , 
        \ScanLink13[2] , \ScanLink20[11] , \Level2Out48[17] , \ScanLink55[21] , 
        \ScanLink208[24] , \ScanLink98[25] , \ScanLink115[17] , 
        \ScanLink160[27] , \ScanLink136[26] , \ScanLink143[16] , 
        \Level2Out6[5] , \Level4Out228[1] , \ScanLink156[22] , \ScanLink1[31] , 
        \ScanLink1[28] , \ScanLink1[21] , \ScanLink1[12] , \ScanLink1[5] , 
        \Level1Out3[22] , \ScanLink5[23] , \ScanLink5[10] , \Level1Out6[19] , 
        \Level1Out52[8] , \ScanLink100[23] , \Level1Out110[7] , 
        \ScanLink123[12] , \ScanLink175[13] , \Level4Out4[11] , 
        \Level2Out90[27] , \Level1Out146[23] , \Level4Out148[4] , 
        \Level1Out105[16] , \Level1Out110[22] , \Level1Out133[13] , 
        \Level2Out26[7] , \Level1Out165[12] , \Level1Out170[26] , 
        \Level1Out126[27] , \Level1Out153[17] , \ScanLink183[0] , 
        \Level1Out245[28] , \Level1Out29[26] , \Level1Out29[15] , 
        \Level1Out213[30] , \Level1Out230[18] , \Level1Out245[31] , 
        \Level1Out30[2] , \Level1Out33[1] , \Level1Out49[11] , 
        \Level1Out213[29] , \Level8Out184[10] , \ScanLink68[31] , 
        \ScanLink151[6] , \ScanLink68[28] , \Level2Out88[7] , 
        \ScanLink203[31] , \ScanLink231[3] , \ScanLink255[29] , 
        \ScanLink203[28] , \ScanLink220[19] , \ScanLink255[30] , 
        \Level4Out72[0] , \Level2Load164[0] , \Level8Out72[25] , 
        \Level1Out49[22] , \Level1Out57[5] , \ScanLink71[8] , 
        \Level1Out84[15] , \ScanLink93[30] , \ScanLink93[29] , 
        \ScanLink152[5] , \Level1Load175[0] , \ScanLink232[0] , 
        \Level8Out24[24] , \ScanLink180[3] , \Level1Out212[8] , 
        \Level1Out91[21] , \Level2Out100[1] , \Level1Out108[5] , 
        \ScanLink135[2] , \Level2Out60[19] , \Level2Out36[18] , 
        \ScanLink190[19] , \ScanLink255[7] , \Level32Out64[7] , 
        \Level4Out16[4] , \Level4Load192[0] , \Level1Out85[3] , 
        \Level16Out176[19] , \Level1Out180[18] , \ScanLink248[8] , 
        \Level8Out184[23] , \Level1Out42[2] , \Level1Out49[9] , 
        \Level1Out86[0] , \Level1Out91[12] , \Level1Out158[31] , 
        \Level2Out134[29] , \Level2Out162[31] , \Level2Out162[28] , 
        \Level1Out54[6] , \Level1Out84[26] , \Level1Out116[9] , 
        \Level1Out158[28] , \Level2Out134[30] , \Level2Out204[0] , 
        \Level2Out164[5] , \ScanLink136[1] , \Level1Out111[28] , 
        \ScanLink120[5] , \ScanLink148[30] , \ScanLink256[4] , 
        \Level2Out20[9] , \Level8Out72[16] , \ScanLink148[29] , 
        \Level8Out24[17] , \Level1Out164[18] , \Level1Out147[30] , 
        \Level2Out108[19] , \Level16Out192[19] , \Level1Out111[31] , 
        \Level1Out132[19] , \Level1Out147[29] , \ScanLink240[0] , 
        \Level8Out160[23] , \Level1Out15[16] , \Level1Out23[13] , 
        \Level1Out41[1] , \Level1Out90[4] , \Level8Out136[22] , 
        \Level1Out93[7] , \ScanLink101[30] , \ScanLink101[29] , 
        \Level1Load107[0] , \Level2Out84[19] , \Level2Out212[4] , 
        \ScanLink157[31] , \ScanLink174[19] , \ScanLink122[18] , 
        \ScanLink157[28] , \Level2Out172[1] , \Level2Out28[1] , 
        \Level8Out96[16] , \Level1Out56[23] , \Level2Out186[28] , 
        \Level1Out75[12] , \ScanLink123[6] , \Level2Out8[3] , 
        \Level2Out186[31] , \Level4Out232[19] , \Level8Out208[20] , 
        \Level1Out26[6] , \Level1Out36[27] , \Level1Out60[26] , 
        \Level2Load116[0] , \Level1Out43[17] , \ScanLink243[3] , 
        \Level1Out164[9] , \ScanLink196[7] , \Level2Out116[5] , 
        \Level2Out52[9] , \Level1Out7[20] , \Level1Out9[4] , \Level1Out15[25] , 
        \Level1Out60[15] , \ScanLink144[1] , \Level8Out160[10] , 
        \Level1Out179[6] , \Level1Out219[3] , \Level8Out136[11] , 
        \ScanLink224[4] , \ScanLink147[2] , \Level2Out236[31] , 
        \Level1Out23[20] , \Level1Out25[5] , \Level1Out43[24] , 
        \Level1Out36[14] , \Level1Out56[10] , \ScanLink227[7] , 
        \Level2Out236[28] , \Level4Out64[4] , \ScanLink54[18] , 
        \Level1Out75[21] , \Level8Out208[13] , \ScanLink77[30] , 
        \ScanLink79[0] , \ScanLink195[4] , \Level2Out108[9] , \ScanLink18[9] , 
        \ScanLink21[31] , \ScanLink21[28] , \ScanLink77[29] , 
        \Level8Out96[25] , \ScanLink87[24] , \Level2Out30[3] , 
        \ScanLink129[27] , \Level1Out48[31] , \Level1Out59[3] , 
        \ScanLink92[10] , \ScanLink149[23] , \Level4Out52[22] , 
        \Level1Out90[18] , \Level1Out159[22] , \Level2Out116[12] , 
        \Level2Out140[13] , \Level4Out124[15] , \Level4Out172[14] , 
        \Level1Out106[3] , \Level2Out120[17] , \Level4Out64[27] , 
        \Level8Out128[29] , \Level2Out176[16] , \Level4Out112[10] , 
        \Level8Out128[30] , \Level1Out139[26] , \Level1Out181[12] , 
        \Level1Out224[15] , \Level4Out32[26] , \Level4Out144[11] , 
        \Level8Out160[3] , \Level1Out48[28] , \ScanLink138[7] , 
        \Level1Out251[25] , \Level2Out6[18] , \Level2Out248[14] , 
        \Level1Out95[9] , \Level1Out207[24] , \Level1Out105[0] , 
        \Level2Out198[23] , \Level1Out194[26] , \Level1Out212[10] , 
        \Level2Out228[10] , \Level8Out200[6] , \Level1Out231[21] , 
        \Level1Out7[13] , \Level1Out20[8] , \ScanLink61[2] , \ScanLink69[11] , 
        \Level1Out88[6] , \ScanLink125[8] , \ScanLink202[11] , 
        \Level1Out244[11] , \ScanLink184[27] , \Level2Out14[23] , 
        \Level2Out42[22] , \Level4Out220[9] , \ScanLink221[20] , 
        \ScanLink254[10] , \Level1Out139[15] , \ScanLink190[9] , 
        \ScanLink191[13] , \ScanLink234[14] , \Level1Out202[2] , 
        \ScanLink217[25] , \ScanLink241[24] , \Level2Out74[27] , 
        \Level4Load20[0] , \Level2Out22[26] , \Level4Out112[23] , 
        \Level2Out120[24] , \Level4Out32[15] , \Level4Out64[14] , 
        \Level1Out159[11] , \Level2Out86[1] , \Level4Out144[22] , 
        \Level2Out176[25] , \Level1Out162[7] , \Level4Out124[26] , 
        \Level2Out116[21] , \Level4Out52[11] , \ScanLink92[23] , 
        \ScanLink149[10] , \Level2Out140[20] , \Level4Out172[27] , 
        \ScanLink69[22] , \ScanLink87[17] , \Level2Out54[7] , 
        \ScanLink129[14] , \Level1Load218[0] , \ScanLink241[17] , 
        \Level2Out74[14] , \ScanLink184[14] , \ScanLink191[20] , 
        \ScanLink234[27] , \ScanLink202[22] , \ScanLink217[16] , 
        \Level128Out128[18] , \Level2Out22[15] , \Level2Out42[11] , 
        \ScanLink221[9] , \ScanLink254[23] , \Level2Out14[10] , 
        \Level1Out201[1] , \Level1Out212[23] , \ScanLink221[13] , 
        \Level2Out228[23] , \Level4Out124[8] , \Level8Out88[0] , 
        \ScanLink18[23] , \ScanLink62[1] , \Level1Out194[15] , 
        \Level1Out244[22] , \Level8Out104[7] , \Level1Out231[12] , 
        \Level1Out251[16] , \Level16Out80[5] , \Level1Out161[4] , 
        \Level1Out181[21] , \Level1Out224[26] , \Level2Out198[10] , 
        \Level8Out216[18] , \ScanLink195[11] , \Level1Out207[17] , 
        \Level8Out240[19] , \ScanLink230[16] , \Level2Out248[27] , 
        \Level1Out197[4] , \ScanLink46[7] , \ScanLink78[27] , \ScanLink94[1] , 
        \ScanLink245[26] , \Level2Out70[25] , \ScanLink180[25] , 
        \ScanLink206[13] , \ScanLink213[27] , \Level2Out26[24] , 
        \Level1Out238[8] , \Level2Out46[20] , \ScanLink225[22] , 
        \Level2Out10[21] , \Level1Out145[2] , \ScanLink250[12] , 
        \Level1Out216[12] , \ScanLink218[0] , \Level8Out240[4] , 
        \Level1Out190[24] , \Level1Out235[23] , \Level1Out240[13] , 
        \Level4Out248[14] , \Level1Out3[11] , \ScanLink4[8] , \ScanLink45[4] , 
        \ScanLink178[5] , \Level1Out185[10] , \Level1Out220[17] , 
        \Level8Out120[1] , \Level1Out203[26] , \Level1Out225[7] , 
        \Level1Out255[27] , \Level4Out228[10] , \Level1Out146[1] , 
        \Level1Out189[8] , \Level2Out124[15] , \Level4Out60[25] , 
        \Level4Out116[12] , \Level2Out172[14] , \Level4Out140[13] , 
        \Level1Out148[14] , \Level4Out36[24] , \Level1Out19[1] , 
        \Level1Out128[10] , \Level4Out56[20] , \ScanLink22[3] , 
        \Level1Out39[30] , \ScanLink83[26] , \ScanLink96[12] , \ScanLink97[2] , 
        \Level1Out226[4] , \Level2Out112[10] , \Level2Out144[11] , 
        \Level2Out254[8] , \Level4Out120[17] , \Level4Out176[16] , 
        \Level32Out0[23] , \ScanLink138[11] , \Level1Out194[7] , 
        \Level2Out70[1] , \ScanLink158[15] , \ScanLink166[9] , 
        \Level1Out255[14] , \Level4Out228[23] , \Level2Out2[29] , 
        \Level1Out39[29] , \Level1Out185[23] , \Level1Out220[24] , 
        \Level1Out121[6] , \Level2Out2[30] , \Level8Out224[0] , 
        \Level1Out203[15] , \Level1Out216[21] , \Level8Out0[5] , 
        \Level1Out240[20] , \Level1Out241[3] , \Level8Out144[5] , 
        \Level1Out11[14] , \ScanLink18[10] , \ScanLink78[14] , 
        \ScanLink180[16] , \Level1Out190[17] , \ScanLink206[20] , 
        \Level1Out235[10] , \Level2Out46[13] , \Level4Out248[27] , 
        \ScanLink250[21] , \ScanLink225[11] , \Level2Out10[12] , 
        \ScanLink21[0] , \Level1Out63[9] , \ScanLink245[15] , 
        \Level2Out70[16] , \ScanLink83[15] , \ScanLink195[22] , 
        \ScanLink230[25] , \ScanLink213[14] , \Level2Out26[17] , 
        \Level1Out94[30] , \ScanLink96[21] , \ScanLink138[22] , 
        \ScanLink158[26] , \Level1Out122[5] , \Level2Out14[5] , 
        \Level2Out112[23] , \Level4Out120[24] , \Level1Out128[23] , 
        \Level4Out56[13] , \Level1Out94[29] , \Level1Out148[27] , 
        \Level1Out242[0] , \Level2Out144[22] , \Level4Out176[25] , 
        \Level32Out0[10] , \Level2Out150[9] , \Level4Out116[21] , 
        \Level2Out124[26] , \Level4Out60[16] , \Level2Out172[27] , 
        \Level4Out36[17] , \Level4Out140[20] , \Level1Load23[0] , 
        \ScanLink25[19] , \Level1Out27[11] , \Level1Out32[25] , 
        \Level1Out64[24] , \Level2Out232[19] , \Level1Out47[15] , 
        \ScanLink203[1] , \Level32Out32[1] , \Level1Out208[19] , 
        \Level4Out40[2] , \Level4Load116[0] , \ScanLink40[9] , 
        \Level1Out52[21] , \Level1Out71[10] , \ScanLink163[4] , 
        \ScanLink50[29] , \Level8Out8[31] , \ScanLink2[6] , \ScanLink50[30] , 
        \ScanLink73[18] , \Level8Out8[28] , \ScanLink88[19] , 
        \ScanLink218[18] , \Level1Out223[9] , \Level2Out68[3] , 
        \Level4Out92[4] , \Level64Load128[0] , \Level1Out192[9] , 
        \Level2Out132[3] , \Level2Out252[6] , \ScanLink200[2] , 
        \Level1Out11[27] , \Level1Out27[22] , \Level1Out52[12] , 
        \Level1Out78[8] , \Level1Out127[8] , \ScanLink160[7] , 
        \Level4Out108[19] , \Level8Out152[24] , \Level8Out104[25] , 
        \Level1Load240[0] , \Level2Out58[18] , \Level2Out182[19] , 
        \Level4Out24[6] , \Level4Out236[31] , \ScanLink39[2] , 
        \Level1Out64[17] , \Level1Out71[23] , \Level4Out236[28] , 
        \ScanLink107[0] , \Level1Out32[16] , \Level1Out47[26] , 
        \Level1Out65[7] , \Level1Out66[4] , \Level1Out115[19] , 
        \Level1Out136[31] , \Level1Out136[28] , \Level1Out139[4] , 
        \Level1Out160[29] , \Level2Out184[1] , \Level8Out152[17] , 
        \Level4Out48[18] , \Level8Out104[16] , \Level1Out143[18] , 
        \Level1Out160[30] , \ScanLink5[19] , \Level1Out7[30] , \ScanLink18[0] , 
        \Level1Out20[1] , \Level1Out85[16] , \Level1Out90[22] , 
        \ScanLink104[3] , \ScanLink105[18] , \Level2Out80[31] , 
        \Level2Out80[28] , \Level2Out156[7] , \ScanLink126[30] , 
        \ScanLink126[29] , \ScanLink170[28] , \Level2Out236[2] , 
        \ScanLink153[19] , \Level1Out159[18] , \ScanLink170[31] , 
        \Level2Out116[28] , \Level2Out116[31] , \Level2Out140[30] , 
        \Level4Out52[18] , \ScanLink190[0] , \Level2Out110[2] , 
        \Level2Out140[29] , \ScanLink142[6] , \ScanLink222[3] , 
        \Level2Out86[8] , \Level8Out128[13] , \ScanLink149[19] , 
        \Level8Out96[5] , \Level1Out23[2] , \ScanLink221[0] , 
        \Level2Out42[18] , \Level2Out14[19] , \Level4Out124[1] , 
        \Level1Out28[16] , \Level1Out48[12] , \ScanLink62[8] , 
        \ScanLink141[5] , \ScanLink191[29] , \Level2Out98[4] , 
        \Level8Out88[27] , \Level128Out128[11] , \ScanLink191[30] , 
        \Level4Out244[4] , \Level2Out6[22] , \Level1Out181[31] , 
        \Level1Out181[28] , \Level2Out198[19] , \Level8Out216[11] , 
        \Level8Out240[10] , \Level1Load166[0] , \ScanLink193[3] , 
        \Level1Out201[8] , \Level8Out88[9] , \Level16Out80[17] , 
        \Level1Out28[25] , \Level1Out44[5] , \ScanLink92[19] , 
        \ScanLink246[7] , \Level1Out85[25] , \ScanLink126[2] , 
        \Level2Out174[6] , \Level8Out128[20] , \Level4Out112[19] , 
        \Level1Out90[11] , \Level1Out96[3] , \Level4Out144[18] , 
        \Level2Out214[3] , \Level1Out105[9] , \Level1Out212[19] , 
        \Level1Out231[31] , \Level2Out228[19] , \Level4Out192[3] , 
        \Level1Out7[29] , \Level1Out231[28] , \Level16Out80[24] , 
        \Level1Out244[18] , \ScanLink17[24] , \Level1Out23[30] , 
        \Level1Out23[29] , \Level1Out47[6] , \Level1Out48[21] , 
        \Level2Out6[11] , \Level8Out216[22] , \ScanLink69[18] , 
        \Level1Out95[0] , \Level8Out240[23] , \Level1Out118[6] , 
        \ScanLink125[1] , \ScanLink221[30] , \ScanLink245[4] , 
        \Level8Out88[14] , \Level4Out140[5] , \Level128Out128[22] , 
        \ScanLink202[18] , \ScanLink221[29] , \Level4Out220[0] , 
        \Level1Out56[19] , \ScanLink67[5] , \ScanLink254[19] , 
        \Level1Out75[31] , \ScanLink99[15] , \ScanLink114[27] , 
        \ScanLink137[16] , \ScanLink142[26] , \Level1Out164[0] , 
        \ScanLink239[2] , \Level2Load76[0] , \Level2Out84[23] , 
        \ScanLink101[13] , \ScanLink161[17] , \Level1Out104[26] , 
        \Level1Out111[12] , \ScanLink122[22] , \ScanLink174[23] , 
        \Level2Out80[6] , \ScanLink157[12] , \ScanLink159[7] , 
        \Level1Out204[5] , \Level1Out127[17] , \Level1Out132[23] , 
        \Level1Out164[22] , \Level1Out147[13] , \Level2Out108[23] , 
        \Level16Out192[23] , \Level2Out168[27] , \Level1Out152[27] , 
        \Level2Out52[0] , \Level8Out160[19] , \ScanLink144[8] , 
        \Level1Out171[16] , \Level8Out136[18] , \Level32Out192[16] , 
        \Level1Out219[15] , \Level1Out75[28] , \ScanLink79[9] , 
        \Level2Out186[12] , \Level2Out108[0] , \ScanLink62[14] , 
        \ScanLink188[2] , \Level2Out200[24] , \Level4Out232[23] , 
        \Level2Load4[0] , \Level4Out252[27] , \Level2Out236[21] , 
        \Level4Out204[26] , \Level1Out167[3] , \ScanLink21[21] , 
        \ScanLink34[15] , \ScanLink41[25] , \ScanLink64[6] , \ScanLink54[11] , 
        \Level1Out207[6] , \ScanLink209[14] , \Level1Out38[3] , 
        \ScanLink77[20] , \Level1Out152[14] , \ScanLink240[9] , 
        \Level1Out8[27] , \ScanLink13[26] , \ScanLink17[17] , \ScanLink21[12] , 
        \ScanLink99[26] , \Level1Out100[4] , \Level1Out104[15] , 
        \Level1Out127[24] , \Level1Out171[25] , \Level2Out168[14] , 
        \Level32Out192[25] , \Level1Out111[21] , \Level1Out164[11] , 
        \Level1Out132[10] , \Level1Out147[20] , \Level2Out36[4] , 
        \Level2Out108[10] , \Level16Out192[10] , \ScanLink174[10] , 
        \ScanLink101[20] , \ScanLink122[11] , \ScanLink157[21] , 
        \ScanLink137[25] , \ScanLink142[15] , \Level2Out172[8] , 
        \ScanLink114[14] , \ScanLink161[24] , \Level2Out84[10] , 
        \ScanLink54[22] , \ScanLink209[27] , \ScanLink77[13] , 
        \Level1Out103[7] , \ScanLink25[23] , \ScanLink34[26] , 
        \ScanLink62[27] , \Level2Out28[8] , \ScanLink41[16] , \Level1Out41[8] , 
        \Level2Out236[12] , \Level4Out204[15] , \Level4Out252[14] , 
        \ScanLink50[13] , \Level1Out219[26] , \Level2Out186[21] , 
        \Level8Out208[30] , \Level1Out247[4] , \Level2Out200[17] , 
        \Level4Out232[10] , \Level8Out208[29] , \Level2Out38[15] , 
        \Level8Load104[0] , \ScanLink66[16] , \ScanLink73[22] , 
        \Level1Out78[1] , \Level8Out8[12] , \Level1Out127[1] , \ScanLink24[4] , 
        \ScanLink45[27] , \ScanLink218[22] , \ScanLink30[17] , 
        \ScanLink107[9] , \Level2Out58[11] , \Level1Out208[23] , 
        \Level2Out148[2] , \Level2Out182[10] , \Level2Out228[7] , 
        \Level2Out232[23] , \Level4Out200[24] , \Level2Out252[27] , 
        \Level2Out204[26] , \Level4Out236[21] , \Level1Out123[15] , 
        \Level1Out156[25] , \Level2Out12[2] , \Level4Out28[15] , 
        \Level1Out100[24] , \Level1Out175[14] , \Level4Out108[23] , 
        \Level1Out3[18] , \Level1Out8[14] , \ScanLink27[7] , \ScanLink88[23] , 
        \ScanLink105[11] , \Level1Out115[10] , \Level4Out168[27] , 
        \Level1Out136[21] , \Level1Out160[20] , \Level2Out184[8] , 
        \Level1Out143[11] , \Level4Out48[11] , \ScanLink170[21] , 
        \ScanLink119[5] , \ScanLink126[20] , \ScanLink153[10] , 
        \Level1Out244[7] , \Level1Out27[18] , \ScanLink110[25] , 
        \Level1Out124[2] , \ScanLink133[14] , \ScanLink146[24] , 
        \ScanLink165[15] , \Level2Out80[21] , \Level2Out182[23] , 
        \Level1Out52[28] , \Level2Out252[14] , \Level4Out236[12] , 
        \ScanLink13[15] , \Level1Out52[31] , \Level2Out204[15] , 
        \Level1Out71[19] , \ScanLink92[6] , \Level1Out191[3] , 
        \ScanLink203[8] , \Level2Out232[10] , \Level4Out200[17] , 
        \Level32Out32[8] , \Level1Out208[10] , \ScanLink25[10] , 
        \ScanLink30[24] , \ScanLink66[25] , \ScanLink40[0] , \ScanLink45[14] , 
        \Level1Out223[0] , \Level2Out58[22] , \Level16Out0[4] , 
        \ScanLink218[11] , \ScanLink43[3] , \ScanLink50[20] , 
        \Level2Out38[26] , \ScanLink73[11] , \Level1Out143[5] , 
        \ScanLink88[10] , \ScanLink110[16] , \ScanLink133[27] , 
        \ScanLink146[17] , \Level1Out220[3] , \Level8Out8[21] , 
        \ScanLink165[26] , \ScanLink170[12] , \Level2Out80[12] , 
        \ScanLink105[22] , \Level1Out140[6] , \ScanLink153[23] , 
        \Level1Out59[24] , \ScanLink91[5] , \Level1Out115[23] , 
        \ScanLink126[13] , \Level1Out160[13] , \Level4Out168[14] , 
        \Level1Out123[26] , \Level1Out136[12] , \Level1Out143[22] , 
        \Level2Out76[6] , \Level1Out156[16] , \Level1Out192[0] , 
        \Level2Load80[0] , \Level4Out48[22] , \Level4Out28[26] , 
        \Level4Out108[10] , \Level1Out100[17] , \Level1Out175[27] , 
        \Level1Out240[30] , \Level8Load24[0] , \Level8Out224[16] , 
        \Level1Out216[28] , \ScanLink7[2] , \ScanLink18[19] , 
        \Level1Out39[20] , \Level1Out216[31] , \Level1Out240[29] , 
        \Level1Out235[19] , \Level2Out2[20] , \Level8Out224[9] , 
        \ScanLink21[9] , \Level1Out60[3] , \Level1Out63[0] , \ScanLink96[31] , 
        \ScanLink101[7] , \ScanLink102[4] , \ScanLink206[30] , 
        \ScanLink206[29] , \ScanLink250[31] , \Level4Out204[6] , 
        \ScanLink250[28] , \ScanLink225[18] , \Level4Out164[3] , 
        \Level1Out81[14] , \ScanLink96[28] , \Level2Out182[6] , 
        \Level1Out94[20] , \Level1Out242[9] , \Level2Out230[5] , 
        \Level4Out116[31] , \Level4Out116[28] , \Level4Out140[30] , 
        \Level4Out140[29] , \Level32Load192[0] , \Level1Out39[13] , 
        \Level1Load42[0] , \Level32Out0[19] , \ScanLink94[8] , 
        \Level1Out158[4] , \ScanLink165[3] , \Level2Out10[31] , 
        \Level2Out150[0] , \Level1Load190[0] , \Level1Out238[1] , 
        \Level2Out10[28] , \Level2Out46[29] , \Level2Out46[30] , 
        \Level2Load230[0] , \ScanLink195[18] , \ScanLink205[6] , 
        \Level4Out100[7] , \Level1Out185[19] , \Level8Out120[8] , 
        \Level2Out2[13] , \Level4Out228[19] , \Level1Out59[17] , 
        \ScanLink218[9] , \Level8Out224[25] , \Level64Out128[5] , 
        \Level1Out19[8] , \ScanLink89[7] , \Level1Out128[19] , 
        \Level4Out56[29] , \Level1Out81[27] , \Level1Out94[13] , 
        \Level2Out112[19] , \Level2Out144[18] , \Level2Out254[1] , 
        \Level4Out56[30] , \Level1Load221[0] , \Level2Out134[4] , 
        \Level1Out146[8] , \Level1Out189[1] , \ScanLink0[11] , \ScanLink4[1] , 
        \Level1Out12[3] , \ScanLink58[2] , \ScanLink166[0] , \Level2Out70[8] , 
        \ScanLink138[18] , \Level1Out142[28] , \ScanLink206[5] , 
        \Level64Out128[27] , \Level1Out114[30] , \Level1Out137[18] , 
        \Level1Out114[29] , \Level1Out142[31] , \Level1Out161[19] , 
        \Level2Out178[28] , \Level8Out128[0] , \ScanLink170[4] , 
        \ScanLink210[1] , \Level2Out178[31] , \Level8Out248[5] , 
        \Level1Out11[0] , \Level1Load30[0] , \ScanLink53[9] , 
        \ScanLink152[29] , \Level1Out230[9] , \Level2Out242[5] , 
        \ScanLink104[31] , \ScanLink127[19] , \Level2Out122[0] , 
        \Level1Out70[13] , \ScanLink104[28] , \ScanLink152[30] , 
        \ScanLink171[18] , \ScanLink173[7] , \Level2Out78[0] , 
        \Level8Load56[0] , \Level1Out26[12] , \ScanLink0[22] , 
        \Level1Out10[17] , \Level1Out33[26] , \Level1Out53[22] , 
        \Level1Out46[16] , \Level1Out181[9] , \ScanLink213[2] , 
        \Level4Out116[3] , \Level1Out65[27] , \Level2Out8[26] , 
        \Level1Out76[7] , \ScanLink89[30] , \Level4Out0[29] , \ScanLink89[29] , 
        \Level2Out226[1] , \Level4Out0[30] , \ScanLink114[0] , 
        \Level1Out134[8] , \Level1Load253[0] , \Level2Out146[4] , 
        \Level1Out249[2] , \Level8Out8[4] , \Level1Out10[24] , 
        \Level1Out33[15] , \Level1Out46[25] , \Level1Out129[7] , 
        \Level2Out194[2] , \Level64Out128[14] , \Level2Load242[0] , 
        \Level2Out246[19] , \Level1Out75[4] , \Level1Out209[29] , 
        \Level1Out65[14] , \ScanLink117[3] , \Level1Out209[30] , 
        \Level2Out8[15] , \Level2Out210[18] , \ScanLink29[1] , 
        \Level4Out212[2] , \Level1Out53[11] , \Level1Out70[20] , 
        \Level2Out158[8] , \Level1Out0[27] , \Level1Out0[14] , \Level1Out0[8] , 
        \Level1Out1[5] , \Level1Out2[21] , \ScanLink9[4] , \ScanLink24[30] , 
        \Level1Out26[21] , \Level4Out172[7] , \ScanLink72[28] , 
        \ScanLink24[29] , \ScanLink51[19] , \ScanLink72[31] , 
        \Level8Out152[8] , \ScanLink82[25] , \ScanLink159[16] , 
        \ScanLink219[31] , \ScanLink219[28] , \Level8Out16[19] , 
        \Level8Out40[18] , \ScanLink97[11] , \Level1Out184[4] , 
        \Level2Out60[2] , \Level1Out38[19] , \ScanLink48[8] , \ScanLink87[1] , 
        \ScanLink139[12] , \ScanLink55[7] , \Level1Out95[19] , 
        \Level1Out236[7] , \Level1Out129[13] , \Level2Out130[22] , 
        \Level16Out48[31] , \Level1Out149[17] , \Level1Out156[2] , 
        \Level2Out166[23] , \Level16Out48[28] , \Level2Out106[27] , 
        \Level4Out48[3] , \Level128Out0[18] , \Level1Out202[25] , 
        \Level2Out150[26] , \ScanLink56[4] , \ScanLink168[6] , 
        \Level1Out184[13] , \Level2Out238[25] , \Level1Out221[14] , 
        \Level1Out235[4] , \Level8Load176[0] , \Level1Out254[24] , 
        \Level1Out191[27] , \Level1Out234[20] , \Level16Out144[17] , 
        \Level32Out192[7] , \Level1Out241[10] , \Level1Out2[12] , 
        \ScanLink19[20] , \ScanLink79[24] , \Level1Out155[1] , 
        \ScanLink181[26] , \ScanLink208[3] , \Level1Out217[11] , 
        \ScanLink224[21] , \Level2Out188[16] , \Level4Out84[9] , 
        \Level16Out112[16] , \ScanLink84[2] , \ScanLink175[9] , 
        \ScanLink251[11] , \Level2Out64[12] , \ScanLink207[10] , 
        \Level2Out32[13] , \Level1Out187[7] , \ScanLink194[12] , 
        \ScanLink212[24] , \Level2Out52[17] , \ScanLink231[15] , 
        \ScanLink19[13] , \ScanLink31[3] , \Level1Out149[24] , 
        \ScanLink244[25] , \Level2Out106[14] , \Level32Out64[19] , 
        \Level1Out252[3] , \Level2Out130[11] , \Level2Out150[15] , 
        \Level32Out32[18] , \Level1Out70[9] , \ScanLink97[22] , 
        \Level1Out129[20] , \Level1Out132[6] , \Level2Out166[10] , 
        \ScanLink82[16] , \ScanLink139[21] , \ScanLink159[25] , 
        \ScanLink212[17] , \Level2Out52[24] , \ScanLink79[17] , 
        \ScanLink181[15] , \ScanLink194[21] , \ScanLink244[16] , 
        \ScanLink224[12] , \ScanLink231[26] , \ScanLink251[22] , 
        \Level2Out64[21] , \ScanLink207[23] , \Level2Out32[20] , 
        \Level1Out241[23] , \Level1Out251[0] , \Level1Out2[6] , 
        \Level1Out6[23] , \ScanLink16[6] , \ScanLink32[0] , \Level1Out131[5] , 
        \Level1Out191[14] , \Level1Out234[13] , \Level1Out217[22] , 
        \Level2Out188[25] , \Level16Out112[25] , \Level16Out144[24] , 
        \Level2Out238[16] , \Level1Out202[16] , \Level1Out254[17] , 
        \ScanLink68[12] , \Level1Load68[0] , \Level1Out184[20] , 
        \ScanLink216[26] , \Level1Out221[27] , \Level2Out56[15] , 
        \Level1Out98[5] , \ScanLink185[24] , \ScanLink190[10] , 
        \ScanLink220[23] , \ScanLink235[17] , \ScanLink240[27] , 
        \ScanLink203[12] , \ScanLink255[13] , \Level2Out60[10] , 
        \Level2Out36[11] , \Level1Out195[25] , \Level1Out230[22] , 
        \Level1Out6[10] , \ScanLink15[5] , \Level1Out115[3] , 
        \Level1Out245[12] , \Level1Out116[0] , \ScanLink128[4] , 
        \Level1Out180[11] , \Level1Out206[27] , \Level1Out213[13] , 
        \ScanLink248[1] , \Level16Out176[10] , \Level1Out225[16] , 
        \Level1Out250[26] , \Level4Out188[16] , \Level1Out138[25] , 
        \Level2Out102[25] , \Level1Out49[18] , \Level1Out49[0] , 
        \Level1Out86[9] , \Level2Out0[2] , \Level2Out154[24] , 
        \Level2Out134[20] , \Level2Out162[21] , \ScanLink86[27] , 
        \ScanLink93[13] , \Level1Out158[21] , \Level2Out204[9] , 
        \ScanLink128[24] , \ScanLink148[20] , \ScanLink136[8] , 
        \Level1Out171[7] , \Level2Out20[0] , \ScanLink72[2] , 
        \Level1Out206[14] , \Level1Out250[15] , \Level4Out188[25] , 
        \Level16Out176[23] , \Level1Out180[22] , \ScanLink183[9] , 
        \Level1Out211[2] , \Level1Out225[25] , \ScanLink185[17] , 
        \Level1Out195[16] , \Level1Out230[11] , \Level1Out245[21] , 
        \Level1Out213[20] , \Level8Out184[19] , \ScanLink220[10] , 
        \ScanLink255[20] , \Level2Out60[23] , \ScanLink203[21] , 
        \Level4Out72[9] , \Level2Out36[22] , \Level2Out56[26] , 
        \Level1Out33[8] , \ScanLink216[15] , \ScanLink240[14] , 
        \ScanLink68[21] , \ScanLink86[14] , \ScanLink128[17] , 
        \ScanLink190[23] , \ScanLink235[24] , \ScanLink232[9] , 
        \ScanLink93[20] , \ScanLink148[13] , \Level2Out44[4] , \ScanLink2[24] , 
        \ScanLink4[20] , \ScanLink4[13] , \ScanLink10[8] , \Level1Out14[15] , 
        \Level1Out37[24] , \ScanLink71[1] , \Level1Out91[28] , 
        \Level2Out134[13] , \Level1Out91[31] , \Level1Out158[12] , 
        \Level2Out100[8] , \Level1Out172[4] , \Level1Out138[16] , 
        \Level2Out102[16] , \Level2Out162[12] , \Level1Out212[1] , 
        \Level2Out96[2] , \Level2Out154[17] , \Level2Out214[30] , 
        \Level1Out42[14] , \ScanLink253[0] , \Level4Out156[1] , 
        \Level2Out242[28] , \Level16Out192[9] , \Level1Out22[10] , 
        \Level1Out51[2] , \Level1Out61[25] , \Level2Out214[29] , 
        \Level1Out74[11] , \ScanLink133[5] , \Level2Out242[31] , 
        \Level4Out236[4] , \ScanLink55[31] , \Level1Out57[20] , 
        \Level4Out4[4] , \ScanLink76[19] , \Level4Out184[7] , \ScanLink20[18] , 
        \ScanLink55[28] , \Level1Out80[7] , \Level1Out83[4] , 
        \Level1Load114[0] , \Level2Out38[2] , \Level2Out162[2] , 
        \Level4Out4[18] , \ScanLink250[3] , \Level2Out202[7] , 
        \Level4Out228[8] , \Level8Out208[7] , \Level16Out64[24] , 
        \Level128Out0[7] , \Level1Out4[8] , \Level1Out14[26] , 
        \Level1Out22[23] , \Level1Out28[9] , \Level1Out52[1] , 
        \Level16Out32[25] , \ScanLink130[6] , \Level8Out168[2] , 
        \Level1Out177[9] , \Level2Out28[30] , \Level2Out28[29] , 
        \Level1Out57[13] , \ScanLink69[3] , \Level1Out74[22] , 
        \ScanLink185[7] , \Level16Out96[8] , \ScanLink237[4] , 
        \Level1Out35[6] , \Level1Out42[27] , \Level4Out132[5] , 
        \Level1Out37[17] , \Level1Out61[16] , \ScanLink157[1] , 
        \ScanLink198[8] , \Level4Out252[0] , \Level1Out36[5] , 
        \Level1Out110[18] , \Level1Out133[29] , \Level1Out169[5] , 
        \ScanLink234[7] , \Level1Out146[19] , \Level1Out165[31] , 
        \Level1Out133[30] , \ScanLink154[2] , \Level1Out165[28] , 
        \Level1Out209[0] , \Level8Out80[1] , \Level16Out64[17] , 
        \Level16Out32[16] , \Level1Out56[1] , \Level1Out84[7] , 
        \ScanLink100[19] , \ScanLink123[28] , \ScanLink229[8] , 
        \Level2Out106[6] , \ScanLink156[18] , \ScanLink186[4] , 
        \ScanLink175[30] , \ScanLink113[30] , \ScanLink113[29] , 
        \ScanLink123[31] , \ScanLink175[29] , \ScanLink145[31] , 
        \ScanLink166[19] , \ScanLink129[9] , \ScanLink130[18] , 
        \ScanLink145[28] , \Level2Out166[2] , \Level8Out32[3] , 
        \Level1Out89[27] , \Level1Out109[1] , \ScanLink254[3] , 
        \Level2Out96[19] , \Level2Out206[7] , \Level1Out99[8] , 
        \Level1Out103[28] , \ScanLink134[6] , \Level1Out155[30] , 
        \Level8Out144[26] , \Level1Out176[18] , \Level1Out103[31] , 
        \Level8Out112[27] , \Level1Out120[19] , \ScanLink2[17] , 
        \Level1Out12[22] , \Level1Out24[27] , \Level1Out51[17] , 
        \Level1Out72[26] , \Level1Out155[29] , \Level4Out152[1] , 
        \Level32Out96[21] , \Level1Out31[13] , \Level1Out44[23] , 
        \Level1Out55[2] , \Level2Out194[28] , \Level4Out0[4] , 
        \Level1Out67[12] , \ScanLink137[5] , \Level2Out194[31] , 
        \Level64Out192[26] , \ScanLink14[8] , \Level4Out220[19] , 
        \Level4Out232[4] , \Level1Out87[4] , \Level2Out18[28] , 
        \Level4Out180[7] , \Level1Load110[0] , \Level2Out18[31] , 
        \Level8Out144[15] , \ScanLink10[19] , \Level1Out32[5] , 
        \ScanLink230[7] , \Level8Out112[14] , \ScanLink33[28] , 
        \Level1Out89[14] , \ScanLink150[2] , \Level4Out148[29] , 
        \Level1Out173[9] , \ScanLink182[4] , \Level2Out102[6] , 
        \Level4Out148[30] , \Level4Out128[9] , \Level8Out56[7] , 
        \ScanLink181[7] , \ScanLink46[18] , \ScanLink65[30] , 
        \Level1Out12[11] , \Level1Out31[20] , \ScanLink33[31] , 
        \ScanLink65[29] , \ScanLink233[4] , \Level2Out58[6] , 
        \Level1Out44[10] , \Level4Out136[5] , \Level64Out192[15] , 
        \Level1Out67[21] , \ScanLink153[1] , \Level1Out248[29] , 
        \Level2Out224[31] , \ScanLink11[5] , \Level1Out24[14] , 
        \Level1Out72[15] , \Level1Out248[30] , \Level2Out224[28] , 
        \Level1Out31[6] , \Level1Out51[24] , \Level32Out96[12] , 
        \ScanLink12[6] , \ScanLink38[24] , \ScanLink58[20] , \ScanLink80[10] , 
        \Level1Out82[18] , \Level1Out82[9] , \Level1Out108[17] , 
        \Level2Out132[17] , \Level4Out100[10] , \Level1Out112[0] , 
        \Level4Out76[27] , \Level2Out164[16] , \Level4Out20[26] , 
        \Level4Out156[11] , \Level1Out168[13] , \Level2Out104[12] , 
        \Level4Out136[15] , \Level2Out200[9] , \Level4Out40[22] , 
        \Level4Out16[23] , \Level2Out4[2] , \Level2Out152[13] , 
        \Level4Out160[14] , \ScanLink95[24] , \ScanLink178[12] , 
        \ScanLink118[16] , \ScanLink132[8] , \Level2Out24[0] , 
        \Level2Out88[12] , \ScanLink183[13] , \ScanLink226[14] , 
        \ScanLink253[24] , \Level2Out66[27] , \Level8Out0[21] , 
        \ScanLink205[25] , \Level2Out30[26] , \Level2Out50[22] , 
        \Level1Out111[3] , \ScanLink196[27] , \ScanLink210[11] , 
        \ScanLink246[10] , \ScanLink233[20] , \Level1Out200[10] , 
        \Level4Out208[17] , \Level1Out186[26] , \Level1Out223[21] , 
        \Level1Out243[25] , \Level1Out5[5] , \Level1Out79[19] , 
        \ScanLink95[17] , \ScanLink118[25] , \Level1Out193[12] , 
        \Level1Out236[15] , \Level1Out215[24] , \ScanLink236[9] , 
        \Level2Out88[21] , \ScanLink199[5] , \Level128Out128[3] , 
        \ScanLink9[31] , \ScanLink75[1] , \ScanLink80[23] , \Level2Out40[4] , 
        \Level1Out176[4] , \ScanLink178[21] , \Level4Out40[11] , 
        \Level2Out104[21] , \Level4Out68[5] , \Level2Out152[20] , 
        \Level4Out136[26] , \Level4Out160[27] , \Level1Out108[24] , 
        \Level1Out168[20] , \Level1Out216[1] , \Level2Out104[8] , 
        \Level4Out16[10] , \Level4Out76[14] , \ScanLink9[28] , 
        \Level1Out29[4] , \Level2Out132[24] , \Level4Out100[23] , 
        \Level2Out164[25] , \Level4Out156[22] , \ScanLink76[2] , 
        \Level1Out193[21] , \Level1Out236[26] , \Level2Out92[2] , 
        \Level4Out20[15] , \Level1Out243[16] , \Level1Out4[25] , 
        \Level1Out4[16] , \Level1Out6[6] , \Level1Out37[8] , \ScanLink38[17] , 
        \ScanLink148[0] , \Level1Out175[7] , \Level1Out215[17] , 
        \ScanLink228[5] , \ScanLink187[9] , \Level1Out200[23] , 
        \Level1Out215[2] , \Level4Out208[24] , \Level1Out186[15] , 
        \ScanLink210[22] , \Level1Out223[12] , \Level2Out50[11] , 
        \Level32Out160[7] , \Level1Out168[8] , \ScanLink196[14] , 
        \ScanLink233[13] , \ScanLink183[20] , \ScanLink226[27] , 
        \ScanLink246[23] , \Level4Out76[9] , \Level8Out0[12] , 
        \ScanLink58[13] , \ScanLink253[17] , \Level2Out66[14] , 
        \ScanLink205[16] , \Level2Out30[15] , \Level8Load184[0] , 
        \ScanLink29[21] , \ScanLink29[12] , \ScanLink49[16] , \ScanLink52[4] , 
        \Level1Out151[1] , \Level1Out197[10] , \Level1Out231[4] , 
        \Level1Out247[27] , \Level2Out208[17] , \Level1Out232[17] , 
        \Level1Out211[26] , \Level8Out200[29] , \Level8Out200[30] , 
        \Level1Out204[12] , \Level4Out80[9] , \ScanLink171[9] , 
        \Level1Out182[24] , \Level1Out252[13] , \Level1Out227[23] , 
        \ScanLink214[13] , \Level2Out54[20] , \Level1Out183[7] , 
        \ScanLink192[25] , \ScanLink242[12] , \Level32Out224[4] , 
        \ScanLink237[22] , \Level2Out62[25] , \ScanLink187[11] , 
        \ScanLink222[16] , \ScanLink51[7] , \ScanLink80[2] , \ScanLink83[1] , 
        \ScanLink91[26] , \ScanLink169[24] , \ScanLink201[27] , 
        \Level2Out34[24] , \Level1Load148[0] , \Level2Out64[2] , 
        \Level64Out0[15] , \ScanLink84[12] , \ScanLink109[20] , 
        \Level1Out180[4] , \Level1Out119[21] , \Level1Out232[7] , 
        \Level2Out100[10] , \Level4Out132[17] , \Level4Out44[20] , 
        \Level4Out12[21] , \Level1Out179[25] , \Level2Out156[11] , 
        \Level4Out164[16] , \Level1Out152[2] , \Level2Out136[15] , 
        \Level4Out104[12] , \Level4Out24[24] , \Level4Out72[25] , 
        \ScanLink187[22] , \ScanLink222[25] , \Level2Out160[14] , 
        \Level4Out152[13] , \ScanLink201[14] , \Level2Out62[16] , 
        \Level2Out34[17] , \ScanLink36[0] , \ScanLink49[25] , 
        \ScanLink214[20] , \ScanLink108[2] , \ScanLink192[16] , 
        \Level2Out54[13] , \Level1Out204[21] , \ScanLink237[11] , 
        \ScanLink242[21] , \Level1Out255[0] , \Level1Out182[17] , 
        \Level1Out197[23] , \Level1Out227[10] , \Level1Out232[24] , 
        \Level1Out252[20] , \Level2Out208[24] , \ScanLink6[26] , 
        \ScanLink8[9] , \ScanLink14[31] , \ScanLink35[3] , \Level1Out69[6] , 
        \Level1Out135[5] , \Level1Out211[15] , \Level1Out247[14] , 
        \Level2Out188[0] , \Level1Out179[16] , \Level2Out136[26] , 
        \Level4Out72[16] , \Level4Out104[21] , \Level1Out86[30] , 
        \Level1Out136[6] , \Level2Out160[27] , \Level4Out24[17] , 
        \Level4Out152[20] , \Level8Out168[19] , \Level2Out100[23] , 
        \Level4Out44[13] , \Level1Out119[12] , \Level2Out156[22] , 
        \Level4Out28[7] , \Level4Out132[24] , \ScanLink37[19] , 
        \ScanLink42[29] , \Level1Out74[9] , \Level1Out86[29] , 
        \Level4Out164[25] , \Level4Out12[12] , \ScanLink84[21] , 
        \ScanLink109[13] , \ScanLink91[15] , \ScanLink169[17] , 
        \ScanLink229[30] , \ScanLink229[29] , \Level64Out0[26] , 
        \Level64Out64[11] , \ScanLink14[28] , \ScanLink42[30] , 
        \ScanLink61[18] , \Level1Out198[6] , \Level8Out80[14] , 
        \Level1Out15[0] , \Level1Out16[20] , \Level1Out35[11] , 
        \Level1Out40[21] , \Level8Out248[23] , \Level1Out63[10] , 
        \ScanLink177[7] , \Level16Out64[8] , \Level1Out20[25] , 
        \ScanLink49[5] , \Level1Out76[24] , \Level1Out239[28] , 
        \Level1Out55[15] , \Level1Out239[31] , \Level2Load58[0] , 
        \Level1Out185[9] , \ScanLink217[2] , \Level2Out220[19] , 
        \Level4Out112[3] , \Level1Out16[3] , \Level1Out98[11] , 
        \ScanLink174[4] , \Level1Out229[6] , \Level1Out16[13] , 
        \Level1Out20[16] , \Level1Load34[0] , \ScanLink57[9] , \ScanLink98[0] , 
        \Level1Out149[3] , \ScanLink214[1] , \Level1Out234[9] , 
        \Level8Out120[20] , \Level8Out176[21] , \Level2Out246[5] , 
        \Level8Out72[1] , \Level64Load0[0] , \Level2Out126[0] , 
        \Level1Out76[17] , \ScanLink113[3] , \Level2Load246[0] , 
        \Level4Out216[2] , \Level1Out35[22] , \Level1Out55[26] , 
        \Level1Out71[4] , \Level8Out248[10] , \Level1Out40[12] , 
        \Level1Out189[31] , \Level2Out190[19] , \Level4Out224[31] , 
        \Level4Out176[7] , \Level4Out224[28] , \Level1Out63[23] , 
        \Level1Out189[28] , \ScanLink199[30] , \ScanLink199[29] , 
        \Level2Out18[4] , \Level8Out80[27] , \Level16Out160[9] , 
        \Level64Out64[22] , \ScanLink0[1] , \ScanLink6[15] , \Level1Out72[7] , 
        \ScanLink117[18] , \ScanLink134[30] , \ScanLink162[28] , 
        \Level1Out130[8] , \ScanLink134[29] , \ScanLink141[19] , 
        \ScanLink162[31] , \Level2Out222[1] , \Level8Out16[5] , 
        \Level2Out92[31] , \Level2Out142[4] , \Level2Out92[28] , 
        \Level1Out98[22] , \ScanLink110[0] , \Level8Out176[12] , 
        \Level1Out172[29] , \Level8Out120[13] , \Level1Out107[19] , 
        \Level1Out124[31] , \Level2Out190[2] , \Level2Out148[29] , 
        \ScanLink25[9] , \ScanLink38[6] , \Level1Out64[3] , \Level1Out124[28] , 
        \Level1Out151[18] , \Level1Out172[30] , \Level2Out148[30] , 
        \ScanLink106[4] , \ScanLink108[19] , \Level8Out64[27] , 
        \Level8Out32[26] , \Level16Out208[4] , \Level1Out92[17] , 
        \Level1Out246[9] , \Level2Out186[6] , \Level2Out234[5] , 
        \Level1Load46[0] , \Level1Out87[23] , \Level1Out118[18] , 
        \Level2Out122[18] , \Level1Out67[0] , \Level1Out69[16] , 
        \Level2Out154[0] , \Level2Out174[19] , \ScanLink105[7] , 
        \ScanLink118[8] , \Level1Out196[30] , \Level2Out4[17] , 
        \Level8Out192[12] , \Level16Out160[28] , \Level1Out196[29] , 
        \Level16Out160[31] , \ScanLink186[31] , \Level4Out200[6] , 
        \Level16Out16[8] , \Level1Out87[10] , \Level1Out138[0] , 
        \ScanLink186[28] , \Level2Out20[30] , \Level2Out20[29] , 
        \Level2Out76[28] , \Level4Out160[3] , \Level2Out76[31] , 
        \Level1Out142[8] , \Level2Out250[1] , \Level8Out64[5] , \ScanLink3[2] , 
        \ScanLink28[18] , \ScanLink85[18] , \Level1Out92[24] , 
        \Level16Out208[18] , \ScanLink162[0] , \Level1Load225[0] , 
        \Level2Out130[4] , \ScanLink202[5] , \Level2Out74[8] , 
        \Level16Load144[0] , \Level8Out64[14] , \ScanLink161[3] , 
        \Level1Load194[0] , \ScanLink236[28] , \ScanLink243[18] , 
        \Level8Out32[15] , \Level2Load234[0] , \ScanLink215[19] , 
        \ScanLink236[31] , \Level1Out69[25] , \ScanLink90[8] , 
        \ScanLink201[6] , \Level1Out253[19] , \Level4Out104[7] , 
        \Level2Out4[24] , \Level1Out226[29] , \ScanLink15[11] , 
        \ScanLink23[7] , \Level1Out99[31] , \Level1Out113[27] , 
        \Level1Out166[17] , \Level1Out205[18] , \Level8Out192[21] , 
        \Level16Out112[9] , \Level1Out226[30] , \Level1Out130[16] , 
        \Level1Out145[26] , \Level1Out150[12] , \Level2Out16[2] , 
        \Level16Out240[21] , \Level1Out99[28] , \Level1Out125[22] , 
        \ScanLink103[26] , \Level1Out106[13] , \Level1Out173[23] , 
        \Level2Out180[8] , \ScanLink116[12] , \ScanLink135[23] , 
        \ScanLink140[13] , \Level1Out240[7] , \ScanLink163[22] , 
        \Level2Out86[16] , \Level1Out120[2] , \ScanLink176[16] , 
        \ScanLink120[17] , \ScanLink155[27] , \ScanLink248[14] , 
        \Level1Out17[19] , \ScanLink20[4] , \ScanLink23[14] , \ScanLink36[20] , 
        \ScanLink60[21] , \ScanLink198[23] , \Level1Out243[4] , 
        \ScanLink43[10] , \ScanLink56[24] , \ScanLink75[15] , 
        \Level1Out123[1] , \Level2Out68[23] , \ScanLink103[9] , 
        \ScanLink228[10] , \Level2Out184[27] , \Level32Out128[17] , 
        \Level64Out0[5] , \Level2Out202[11] , \Level2Out254[10] , 
        \Level4Out96[16] , \Level1Out238[11] , \Level1Out34[31] , 
        \Level4Out180[25] , \Level16Out128[22] , \Level1Out34[28] , 
        \Level1Out62[29] , \Level1Out188[22] , \Level2Out234[14] , 
        \Level1Out41[18] , \ScanLink47[3] , \Level1Out62[30] , 
        \ScanLink103[15] , \ScanLink120[24] , \ScanLink176[25] , 
        \Level1Out224[3] , \ScanLink135[10] , \ScanLink155[14] , 
        \ScanLink179[1] , \Level1Out106[20] , \ScanLink116[21] , 
        \ScanLink140[20] , \ScanLink219[4] , \Level2Out86[25] , 
        \Level1Out125[11] , \Level1Out144[6] , \ScanLink163[11] , 
        \Level1Out150[21] , \Level2Out72[6] , \ScanLink15[22] , 
        \Level1Out18[5] , \ScanLink23[27] , \ScanLink56[17] , \ScanLink95[5] , 
        \Level1Out113[14] , \Level1Out173[10] , \ScanLink96[6] , 
        \Level1Out130[25] , \Level1Out166[24] , \Level1Out196[0] , 
        \Level2Load84[0] , \Level16Out240[12] , \Level1Out145[15] , 
        \Level1Out159[9] , \Level1Out188[11] , \Level4Out88[1] , 
        \Level1Out195[3] , \ScanLink207[8] , \Level2Out234[27] , 
        \Level2Out248[3] , \Level4Out180[16] , \Level16Out128[11] , 
        \Level2Out254[23] , \Level1Out238[22] , \Level2Out184[14] , 
        \Level32Out128[24] , \Level2Out128[6] , \Level2Out202[22] , 
        \Level4Out96[25] , \Level1Out227[0] , \ScanLink75[26] , 
        \ScanLink60[12] , \Level1Out147[5] , \ScanLink198[10] , 
        \ScanLink228[23] , \Level2Out68[10] , \ScanLink248[27] , 
        \ScanLink36[13] , \ScanLink43[23] , \ScanLink44[0] , 
        \Level1Out199[14] , \Level1Out229[27] , \Level4Out184[27] , 
        \Level1Out249[23] , \Level2Load0[0] , \Level2Out180[25] , 
        \Level2Out230[16] , \Level2Out206[13] , \Level2Out250[12] , 
        \Level4Out92[14] , \ScanLink11[20] , \ScanLink11[13] , 
        \ScanLink27[16] , \ScanLink52[26] , \ScanLink60[6] , \ScanLink71[17] , 
        \Level1Out163[3] , \ScanLink189[15] , \ScanLink32[22] , 
        \ScanLink64[23] , \ScanLink239[26] , \Level1Out203[6] , 
        \ScanLink47[12] , \ScanLink63[5] , \ScanLink107[24] , 
        \Level1Out160[0] , \ScanLink172[14] , \Level2Load72[0] , 
        \ScanLink64[10] , \Level1Out102[11] , \ScanLink112[10] , 
        \ScanLink124[15] , \ScanLink151[25] , \ScanLink131[21] , 
        \ScanLink144[11] , \Level1Out200[5] , \ScanLink167[20] , 
        \Level1Out121[20] , \Level1Out154[10] , \Level2Out82[14] , 
        \Level2Out84[6] , \Level16Out224[27] , \Level1Out177[21] , 
        \Level2Out138[11] , \Level1Out107[7] , \Level1Out117[25] , 
        \ScanLink140[8] , \Level1Out162[15] , \Level32Out224[12] , 
        \Level2Out158[15] , \Level1Out134[14] , \Level1Out141[24] , 
        \ScanLink239[15] , \Level2Out56[0] , \ScanLink27[25] , 
        \ScanLink32[11] , \ScanLink47[21] , \ScanLink52[15] , \Level1Out58[7] , 
        \ScanLink71[24] , \ScanLink189[26] , \Level1Out199[27] , 
        \Level2Out180[16] , \Level2Out250[21] , \ScanLink0[8] , \ScanLink5[5] , 
        \ScanLink6[6] , \ScanLink8[22] , \Level1Out13[31] , \Level1Out13[28] , 
        \Level1Out45[30] , \Level1Out66[18] , \Level1Out249[10] , 
        \Level4Out92[27] , \Level2Out168[4] , \Level2Out206[20] , 
        \Level1Out229[14] , \Level4Out184[14] , \Level1Out30[19] , 
        \Level1Out45[29] , \Level1Out45[8] , \Level2Out208[1] , 
        \Level1Out18[24] , \Level1Out27[2] , \ScanLink59[19] , 
        \Level1Out89[2] , \Level1Out117[16] , \Level2Out230[25] , 
        \Level1Out134[27] , \Level1Out162[26] , \Level2Out158[26] , 
        \Level32Out224[21] , \ScanLink244[9] , \Level1Out141[17] , 
        \Level16Out16[30] , \Level1Out102[22] , \Level1Out121[13] , 
        \Level1Out154[23] , \Level2Out32[4] , \Level16Out224[14] , 
        \Level16Out16[29] , \Level1Out104[4] , \ScanLink112[23] , 
        \ScanLink131[12] , \Level1Out177[12] , \Level2Out138[22] , 
        \ScanLink144[22] , \Level2Out176[8] , \Level2Out82[27] , 
        \ScanLink107[17] , \ScanLink167[13] , \ScanLink124[26] , 
        \ScanLink139[3] , \ScanLink172[27] , \ScanLink151[16] , 
        \Level8Out48[18] , \Level1Out178[2] , \ScanLink211[31] , 
        \ScanLink225[0] , \ScanLink232[19] , \ScanLink211[28] , 
        \ScanLink247[29] , \Level4Out120[1] , \Level1Out218[7] , 
        \ScanLink247[30] , \ScanLink145[5] , \Level4Out240[4] , 
        \ScanLink66[8] , \Level1Out78[20] , \ScanLink197[3] , 
        \Level1Out201[30] , \Level1Out205[8] , \Level1Out222[18] , 
        \Level2Out0[15] , \Level2Out218[18] , \Level1Out83[21] , 
        \Level1Load162[0] , \Level1Out201[29] , \Level64Out64[2] , 
        \Level2Out114[2] , \ScanLink8[11] , \Level1Out8[0] , \ScanLink194[0] , 
        \Level2Out82[8] , \Level8Out40[3] , \Level16Out48[6] , 
        \Level1Out18[17] , \Level1Out24[1] , \ScanLink78[4] , 
        \Level1Out96[15] , \ScanLink226[3] , \Level8Out56[20] , 
        \Level4Out8[30] , \Level16Out128[3] , \ScanLink81[30] , 
        \ScanLink81[29] , \ScanLink146[6] , \Level4Out8[29] , \Level1Out40[5] , 
        \Level1Out43[6] , \Level1Out78[13] , \Level1Out91[0] , 
        \Level1Out101[9] , \Level2Out0[26] , \Level4Out196[3] , 
        \Level1Out192[18] , \ScanLink182[19] , \ScanLink241[4] , 
        \Level4Out144[5] , \Level2Out72[19] , \ScanLink121[1] , 
        \ScanLink122[2] , \ScanLink179[18] , \ScanLink242[7] , 
        \Level2Out24[18] , \Level4Out224[0] , \Level8Out56[13] , 
        \Level32Load160[0] , \Level1Out83[12] , \Level1Out96[26] , 
        \Level2Out170[6] , \ScanLink88[3] , \Level1Out92[3] , 
        \Level1Out169[19] , \Level2Out126[29] , \Level8Out24[7] , 
        \Level2Out170[31] , \ScanLink116[31] , \Level2Out126[30] , 
        \Level2Out170[28] , \Level2Out210[3] , \ScanLink116[28] , 
        \ScanLink135[19] , \ScanLink140[29] , \Level2Out136[3] , 
        \ScanLink140[30] , \ScanLink163[18] , \ScanLink7[25] , 
        \Level1Out106[30] , \Level1Out159[0] , \ScanLink179[8] , 
        \Level1Out196[9] , \ScanLink204[2] , \Level4Out88[8] , 
        \Level1Out125[18] , \Level1Out17[23] , \Level1Out21[26] , 
        \Level1Out54[16] , \Level1Out99[12] , \Level1Out106[29] , 
        \Level1Out150[28] , \Level1Out239[5] , \Level1Out150[31] , 
        \ScanLink164[7] , \Level1Out173[19] , \ScanLink207[1] , 
        \ScanLink59[6] , \Level1Out77[27] , \Level4Out44[2] , 
        \Level32Load32[0] , \Level1Out62[13] , \ScanLink167[4] , 
        \Level1Out188[18] , \Level1Out34[12] , \Level1Out41[22] , 
        \Level4Load112[0] , \Level16Out128[18] , \Level1Out188[5] , 
        \ScanLink198[19] , \ScanLink7[16] , \Level1Load27[0] , \ScanLink44[9] , 
        \Level4Out96[4] , \Level1Out227[9] , \Level2Out68[19] , 
        \ScanLink15[18] , \Level1Out62[4] , \Level1Out99[21] , 
        \ScanLink100[3] , \Level2Out180[1] , \Level16Out240[31] , 
        \Level1Out123[8] , \Level1Load244[0] , \Level2Out152[7] , 
        \Level16Out240[28] , \Level32Out128[4] , \Level2Out232[2] , 
        \ScanLink228[19] , \Level1Out17[10] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink60[28] , \ScanLink43[19] , \ScanLink60[31] , 
        \Level1Out21[15] , \Level1Out34[21] , \Level1Out62[20] , 
        \Level1Out41[11] , \Level4Out20[6] , \Level1Out54[25] , 
        \Level1Out61[7] , \Level1Out77[14] , \ScanLink103[0] , 
        \Level2Out202[18] , \Level2Out254[19] , \Level1Out142[1] , 
        \Level1Out238[18] , \Level2Out114[27] , \Level1Out1[24] , 
        \Level1Out1[17] , \Level1Out5[26] , \Level1Out5[15] , \ScanLink28[11] , 
        \ScanLink41[4] , \Level1Out178[26] , \ScanLink85[11] , 
        \Level1Out87[19] , \Level1Out222[4] , \Level2Out122[22] , 
        \Level2Out142[26] , \Level16Out208[11] , \Level1Out118[22] , 
        \Level2Out174[23] , \Level2Out250[8] , \ScanLink90[25] , 
        \ScanLink93[2] , \ScanLink108[23] , \Level1Out190[7] , 
        \Level2Out98[27] , \ScanLink162[9] , \ScanLink168[27] , 
        \Level2Out74[1] , \ScanLink42[7] , \ScanLink48[15] , \ScanLink90[1] , 
        \ScanLink186[12] , \Level1Out193[4] , \ScanLink200[24] , 
        \Level2Out40[17] , \ScanLink256[25] , \Level2Out16[16] , 
        \ScanLink193[26] , \ScanLink223[15] , \ScanLink236[21] , 
        \ScanLink243[11] , \Level2Out76[12] , \ScanLink215[10] , 
        \Level2Out20[13] , \Level1Out141[2] , \Level1Out183[27] , 
        \Level1Out226[20] , \Level1Out253[10] , \Level4Out88[27] , 
        \Level8Out192[31] , \Level32Out160[27] , \Level1Out205[11] , 
        \Level8Out192[28] , \Level16Out112[0] , \Level1Out210[25] , 
        \Level16Out160[12] , \ScanLink25[0] , \ScanLink85[22] , 
        \ScanLink90[16] , \ScanLink168[14] , \Level1Out196[13] , 
        \Level1Out221[7] , \Level1Out246[24] , \Level1Out233[14] , 
        \ScanLink108[10] , \Level2Out98[14] , \Level2Out10[5] , 
        \ScanLink26[3] , \Level1Out79[5] , \Level1Load89[0] , 
        \Level1Out118[11] , \Level1Out126[5] , \Level2Out122[11] , 
        \Level2Out154[9] , \Level2Out174[10] , \Level1Out125[6] , 
        \Level1Out178[15] , \Level1Out246[0] , \Level2Out114[14] , 
        \Level2Out142[15] , \Level16Out208[22] , \Level1Out210[16] , 
        \Level16Out160[21] , \Level1Out196[20] , \Level16Out176[4] , 
        \Level1Out233[27] , \ScanLink28[22] , \ScanLink48[26] , 
        \ScanLink118[1] , \Level1Out245[3] , \Level1Out246[17] , 
        \Level2Out198[3] , \Level1Out138[9] , \Level1Out183[14] , 
        \Level1Out226[13] , \Level32Out160[14] , \ScanLink193[15] , 
        \Level1Out205[22] , \Level1Out253[23] , \Level4Out88[14] , 
        \ScanLink236[12] , \ScanLink215[23] , \ScanLink243[22] , 
        \Level2Out76[21] , \Level2Out20[20] , \ScanLink200[17] , 
        \Level8Out192[3] , \Level16Out16[1] , \Level1Out67[9] , 
        \ScanLink186[21] , \Level2Out16[25] , \Level2Out40[24] , 
        \ScanLink223[26] , \Level1Out91[9] , \ScanLink256[16] , 
        \Level1Out214[27] , \Level1Out242[26] , \ScanLink8[18] , 
        \Level1Load8[0] , \ScanLink39[27] , \Level1Out101[0] , 
        \Level1Out187[25] , \Level1Out192[11] , \Level1Out222[22] , 
        \Level1Out237[16] , \Level2Out218[22] , \ScanLink121[8] , 
        \ScanLink197[24] , \Level1Out201[13] , \ScanLink232[23] , 
        \ScanLink247[13] , \Level2Out72[10] , \ScanLink59[23] , 
        \ScanLink211[12] , \Level2Out24[11] , \Level2Out44[15] , 
        \Level4Load24[0] , \Level4Out224[9] , \Level16Out32[7] , 
        \ScanLink81[13] , \ScanLink94[27] , \ScanLink182[10] , 
        \ScanLink204[26] , \ScanLink252[27] , \ScanLink227[17] , 
        \Level2Out12[14] , \ScanLink119[15] , \Level2Out34[3] , 
        \Level1Out169[10] , \ScanLink179[11] , \Level2Out126[20] , 
        \Level4Out8[13] , \Level4Out188[6] , \Level2Out170[21] , 
        \Level4Out8[5] , \ScanLink39[14] , \ScanLink59[10] , \Level1Out102[3] , 
        \Level2Out110[25] , \Level1Out109[14] , \Level2Out146[24] , 
        \ScanLink182[23] , \ScanLink204[15] , \Level2Out44[26] , 
        \ScanLink197[17] , \ScanLink227[24] , \ScanLink232[10] , 
        \ScanLink252[14] , \Level2Out12[27] , \ScanLink211[21] , 
        \ScanLink225[9] , \ScanLink247[20] , \Level2Out72[23] , 
        \Level2Out24[22] , \Level4Out120[8] , \ScanLink66[1] , 
        \Level1Out78[30] , \ScanLink158[3] , \Level1Out205[1] , 
        \Level1Out187[16] , \Level1Out222[11] , \Level1Out201[20] , 
        \Level2Out218[11] , \Level1Out78[29] , \Level1Out165[4] , 
        \Level1Out214[14] , \ScanLink238[6] , \Level1Out192[22] , 
        \Level1Out237[25] , \Level1Out242[15] , \Level1Out8[9] , 
        \Level1Out39[7] , \Level1Out109[27] , \Level1Out206[2] , 
        \Level2Out82[1] , \Level2Out110[16] , \ScanLink194[9] , 
        \Level2Out146[17] , \ScanLink11[30] , \ScanLink11[29] , 
        \Level1Out24[8] , \ScanLink65[2] , \Level1Out83[31] , 
        \Level1Out83[28] , \Level1Out169[23] , \Level1Out166[7] , 
        \Level2Out126[13] , \Level2Out170[12] , \ScanLink47[31] , 
        \ScanLink64[19] , \ScanLink81[20] , \ScanLink94[14] , 
        \ScanLink119[26] , \ScanLink179[22] , \Level2Out50[7] , 
        \ScanLink189[6] , \Level4Out8[20] , \Level8Out56[29] , 
        \Level8Out56[30] , \Level1Out97[7] , \ScanLink32[18] , 
        \ScanLink47[28] , \Level1Out13[21] , \Level1Out66[11] , 
        \ScanLink127[6] , \ScanLink19[4] , \Level1Out25[24] , 
        \Level1Out30[10] , \Level1Out45[20] , \Level1Out45[1] , 
        \Level2Out208[8] , \Level1Out50[14] , \Level2Out250[28] , 
        \ScanLink247[3] , \Level2Out206[30] , \Level1Out73[25] , 
        \Level2Load112[0] , \Level2Out250[31] , \ScanLink3[27] , 
        \Level1Out46[2] , \Level1Out249[19] , \Level2Out206[29] , 
        \Level1Out13[12] , \Level1Out21[5] , \Level1Out25[17] , 
        \Level1Out88[24] , \ScanLink124[5] , \Level16Out16[20] , 
        \Level1Out94[4] , \Level1Out119[2] , \ScanLink244[0] , 
        \Level32Out224[28] , \Level32Out224[31] , \Level1Load103[0] , 
        \Level2Out216[4] , \Level2Out176[1] , \Level8Out48[11] , 
        \Level16Out0[25] , \Level1Out50[27] , \Level1Out73[16] , 
        \ScanLink143[2] , \Level32Out0[4] , \Level1Out30[23] , 
        \Level1Out66[22] , \ScanLink223[7] , \Level1Out45[13] , 
        \Level4Out60[4] , \ScanLink131[28] , \ScanLink144[18] , 
        \ScanLink167[30] , \ScanLink191[4] , \Level2Out48[5] , 
        \ScanLink192[7] , \Level1Out0[1] , \ScanLink3[14] , \Level1Out22[6] , 
        \Level1Out88[17] , \ScanLink112[19] , \ScanLink131[31] , 
        \ScanLink167[29] , \ScanLink140[1] , \Level1Out160[9] , 
        \Level16Out0[16] , \Level2Out112[5] , \Level8Out48[22] , 
        \Level2Out56[9] , \Level1Out3[2] , \ScanLink9[21] , \Level1Out34[2] , 
        \Level1Out102[18] , \Level1Out121[30] , \Level1Out121[29] , 
        \Level1Out154[19] , \Level1Out177[31] , \ScanLink220[4] , 
        \Level1Out177[28] , \Level2Out138[18] , \Level16Out16[13] , 
        \ScanLink156[5] , \ScanLink178[31] , \ScanLink68[7] , 
        \ScanLink178[28] , \ScanLink236[0] , \Level2Out88[28] , 
        \Level1Out97[16] , \ScanLink184[3] , \Level2Out88[31] , 
        \Level1Out216[8] , \Level1Load171[0] , \ScanLink9[12] , 
        \Level1Out19[27] , \ScanLink75[8] , \Level1Out168[30] , 
        \Level2Out104[28] , \Level2Out152[30] , \Level4Out40[18] , 
        \Level1Out82[22] , \Level2Out104[31] , \Level2Out152[29] , 
        \ScanLink148[9] , \Level1Out168[29] , \Level4Out16[19] , 
        \ScanLink187[0] , \Level2Out104[1] , \Level8Out232[14] , 
        \Level1Out37[1] , \Level1Out79[23] , \Level1Out193[28] , 
        \Level1Out193[31] , \Level1Out82[11] , \Level1Out82[0] , 
        \ScanLink155[6] , \ScanLink183[29] , \Level1Out208[4] , 
        \Level1Out168[1] , \ScanLink183[30] , \ScanLink235[3] , 
        \Level2Out50[18] , \Level2Load160[0] , \Level4Out76[0] , 
        \Level2Out200[0] , \Level1Out97[25] , \Level2Out160[5] , 
        \Level4Out100[19] , \Level1Out19[14] , \Level1Out50[6] , 
        \Level1Out112[9] , \Level4Out156[18] , \Level1Out53[5] , 
        \ScanLink80[19] , \ScanLink132[1] , \Level2Out24[9] , \ScanLink131[2] , 
        \ScanLink252[4] , \ScanLink210[18] , \ScanLink233[30] , 
        \ScanLink246[19] , \ScanLink58[30] , \ScanLink233[29] , 
        \ScanLink251[7] , \ScanLink58[29] , \Level4Out12[4] , \Level8Out0[28] , 
        \Level1Out79[10] , \Level8Out0[31] , \Level1Out81[3] , 
        \Level4Load196[0] , \Level1Out200[19] , \Level8Out232[27] , 
        \Level1Out223[31] , \Level1Out116[26] , \Level1Out135[17] , 
        \Level1Out140[27] , \Level1Out223[28] , \Level4Out148[20] , 
        \Level1Out163[16] , \Level2Out46[3] , \Level4Out68[16] , 
        \ScanLink10[10] , \ScanLink33[21] , \ScanLink73[6] , 
        \Level1Out103[12] , \Level1Out176[22] , \ScanLink113[13] , 
        \Level1Out120[23] , \Level1Out155[13] , \Level4Out128[24] , 
        \ScanLink166[23] , \ScanLink130[22] , \ScanLink145[12] , 
        \Level2Out94[5] , \Level1Out210[6] , \Level4Out248[5] , 
        \ScanLink106[27] , \ScanLink125[16] , \ScanLink150[26] , 
        \Level1Out170[3] , \ScanLink173[17] , \Level4Out128[0] , 
        \Level1Out213[5] , \Level2Out96[23] , \ScanLink46[11] , 
        \Level16Out240[7] , \Level2Out78[16] , \ScanLink26[15] , 
        \ScanLink65[20] , \ScanLink238[25] , \ScanLink70[14] , 
        \Level1Out173[0] , \ScanLink188[16] , \Level2Out18[12] , 
        \ScanLink53[25] , \ScanLink70[5] , \ScanLink153[8] , 
        \Level1Out248[20] , \Level8Out48[2] , \Level1Out1[30] , 
        \Level1Out1[29] , \ScanLink8[26] , \ScanLink8[0] , \ScanLink10[23] , 
        \Level1Out12[18] , \Level1Out31[29] , \Level1Out198[17] , 
        \Level2Out194[12] , \Level2Out224[21] , \Level4Out216[26] , 
        \Level4Out240[27] , \Level1Out44[19] , \Level1Out67[31] , 
        \Level2Out244[25] , \Level4Load56[0] , \Level4Out220[23] , 
        \ScanLink14[1] , \ScanLink17[2] , \Level1Out31[30] , \Level1Out67[28] , 
        \Level2Out212[24] , \ScanLink106[14] , \ScanLink125[25] , 
        \ScanLink129[0] , \Level1Out228[24] , \Level2Out2[5] , 
        \ScanLink150[15] , \ScanLink113[20] , \ScanLink173[24] , 
        \Level2Out96[10] , \Level1Out114[7] , \ScanLink249[5] , 
        \ScanLink130[11] , \ScanLink166[10] , \ScanLink26[26] , 
        \Level1Out48[4] , \Level1Out56[8] , \Level1Out99[1] , 
        \Level1Out103[21] , \ScanLink145[21] , \Level1Out176[11] , 
        \Level1Out120[10] , \ScanLink70[27] , \Level1Out109[8] , 
        \Level1Out135[24] , \Level1Out155[20] , \Level2Out22[7] , 
        \Level4Out128[17] , \Level4Out148[13] , \Level1Out116[15] , 
        \Level1Out140[14] , \Level1Out163[25] , \Level4Out68[25] , 
        \Level1Out198[24] , \Level1Out228[17] , \Level2Out194[21] , 
        \Level2Out218[2] , \Level2Out244[16] , \Level2Out212[17] , 
        \Level4Out220[10] , \Level32Out96[31] , \Level1Out248[13] , 
        \Level4Out240[14] , \Level2Out178[7] , \Level2Out224[12] , 
        \Level32Out96[28] , \Level4Out152[8] , \Level4Out216[15] , 
        \ScanLink53[16] , \ScanLink188[25] , \Level2Out18[21] , 
        \Level16Out224[3] , \ScanLink33[12] , \ScanLink46[22] , 
        \ScanLink65[13] , \Level1Out117[4] , \ScanLink238[16] , 
        \Level2Out78[25] , \Level16Out144[6] , \ScanLink14[21] , 
        \ScanLink14[12] , \ScanLink22[17] , \ScanLink74[16] , 
        \Level1Load129[0] , \Level1Out189[21] , \Level2Out190[10] , 
        \Level8Out248[19] , \Level2Out216[26] , \Level2Out240[27] , 
        \Level4Out224[21] , \Level1Out239[12] , \Level4Out244[25] , 
        \Level8Out184[7] , \Level2Out220[23] , \Level4Out212[24] , 
        \Level1Out133[2] , \ScanLink229[13] , \Level16Out160[0] , 
        \ScanLink30[7] , \ScanLink37[23] , \ScanLink57[27] , \Level1Out253[7] , 
        \ScanLink42[13] , \ScanLink249[17] , \ScanLink33[4] , \ScanLink61[22] , 
        \ScanLink199[20] , \Level2Load138[0] , \ScanLink37[10] , 
        \ScanLink42[20] , \ScanLink54[3] , \ScanLink102[25] , 
        \ScanLink121[14] , \ScanLink154[24] , \Level1Out130[1] , 
        \ScanLink177[15] , \Level2Out92[21] , \Level4Out168[2] , 
        \Level64Out192[6] , \Level1Out107[10] , \ScanLink117[11] , 
        \ScanLink162[21] , \Level2Out222[8] , \ScanLink134[20] , 
        \ScanLink141[10] , \Level1Out250[4] , \Level1Out172[20] , 
        \Level4Out208[7] , \ScanLink110[9] , \Level1Out124[21] , 
        \Level1Out151[11] , \Level2Out148[20] , \Level1Out131[15] , 
        \Level1Out144[25] , \Level1Out167[14] , \Level1Out112[24] , 
        \Level2Out128[24] , \ScanLink61[11] , \Level1Out157[6] , 
        \ScanLink199[13] , \ScanLink249[24] , \ScanLink22[24] , 
        \ScanLink57[14] , \ScanLink74[25] , \ScanLink229[20] , 
        \Level1Out237[3] , \ScanLink86[5] , \Level1Out239[21] , 
        \Level4Out244[16] , \Level64Out64[18] , \Level1Out185[0] , 
        \Level2Out138[5] , \Level1Out8[4] , \Level1Out10[4] , \Level1Out13[7] , 
        \Level1Out15[9] , \Level2Out220[10] , \Level4Out212[17] , 
        \Level1Out16[30] , \Level1Out35[18] , \Level1Out40[28] , 
        \Level2Out240[14] , \Level2Out190[23] , \Level1Out16[29] , 
        \Level1Out40[31] , \Level1Out63[19] , \Level1Out189[12] , 
        \Level2Out216[15] , \Level16Out64[1] , \ScanLink28[5] , 
        \ScanLink29[31] , \ScanLink57[0] , \ScanLink85[6] , \Level1Out131[26] , 
        \Level1Out186[3] , \ScanLink214[8] , \Level4Out224[12] , 
        \Level1Out144[16] , \Level8Out120[30] , \Level8Out176[28] , 
        \ScanLink98[9] , \Level1Out98[18] , \Level1Out107[23] , 
        \Level1Out112[17] , \Level1Out167[27] , \Level2Out128[17] , 
        \Level8Out120[29] , \Level2Out148[13] , \Level8Out176[31] , 
        \ScanLink117[22] , \Level1Out124[12] , \Level1Out172[13] , 
        \Level1Out151[22] , \Level2Out62[5] , \ScanLink209[7] , 
        \ScanLink134[13] , \Level1Out154[5] , \ScanLink162[12] , 
        \Level1Out77[3] , \ScanLink102[16] , \ScanLink121[27] , 
        \ScanLink141[23] , \Level2Out126[9] , \Level1Out234[0] , 
        \Level8Out72[8] , \ScanLink154[17] , \ScanLink169[2] , 
        \Level2Out92[12] , \Level1Out128[3] , \ScanLink177[26] , 
        \ScanLink214[30] , \ScanLink214[29] , \ScanLink237[18] , 
        \ScanLink242[31] , \ScanLink242[28] , \Level4Out36[2] , 
        \Level4Load160[0] , \ScanLink29[28] , \ScanLink115[4] , 
        \Level1Out248[6] , \ScanLink36[9] , \Level1Load55[0] , 
        \Level8Out200[13] , \Level1Out68[15] , \Level1Out204[28] , 
        \Level2Out188[9] , \Level32Out96[7] , \Level1Out252[30] , 
        \Level1Out255[9] , \Level16Out96[15] , \Level1Out86[20] , 
        \Level1Out204[31] , \Level1Out227[19] , \Level1Out252[29] , 
        \Level1Out93[14] , \Level2Out144[3] , \Level4Out104[28] , 
        \Level4Out152[30] , \Level2Out224[6] , \Level4Out152[29] , 
        \Level8Out168[10] , \Level4Out104[31] , \Level1Out68[26] , 
        \Level1Out74[0] , \ScanLink84[31] , \ScanLink116[7] , 
        \Level2Out196[5] , \ScanLink84[28] , \Level1Out151[8] , 
        \Level1Load236[0] , \Level2Load196[0] , \Level4Out80[0] , 
        \Level16Out96[26] , \ScanLink171[0] , \ScanLink187[18] , 
        \Level1Out197[19] , \ScanLink211[5] , \Level8Out200[20] , 
        \Level4Out52[6] , \Level2Out54[29] , \ScanLink83[8] , 
        \Level2Out54[30] , \ScanLink109[30] , \ScanLink109[29] , 
        \ScanLink212[6] , \Level1Out24[5] , \Level1Out86[13] , 
        \Level1Out93[27] , \ScanLink172[3] , \Level1Load187[0] , 
        \Level1Out119[31] , \Level2Out100[19] , \Level2Out120[7] , 
        \Level4Out12[31] , \Level8Out168[23] , \Level4Out44[29] , 
        \Level2Out240[2] , \Level4Out12[28] , \Level1Out119[28] , 
        \Level2Out156[18] , \Level4Out44[30] , \ScanLink146[2] , 
        \ScanLink78[0] , \ScanLink94[19] , \ScanLink226[7] , 
        \Level16Out128[7] , \Level1Out96[11] , \ScanLink194[4] , 
        \Level8Out56[24] , \Level8Out40[7] , \Level16Out48[2] , 
        \Level1Out18[20] , \Level1Out83[25] , \ScanLink197[7] , 
        \Level2Out114[6] , \Level64Out64[6] , \Level2Out0[11] , 
        \Level1Out78[24] , \Level1Out237[28] , \Level1Out242[18] , 
        \Level1Out165[9] , \Level1Out214[19] , \Level1Out237[31] , 
        \ScanLink3[19] , \ScanLink8[15] , \Level1Out27[6] , \ScanLink39[19] , 
        \ScanLink145[1] , \Level1Out218[3] , \ScanLink227[29] , 
        \ScanLink252[19] , \ScanLink204[18] , \ScanLink227[30] , 
        \Level4Out240[0] , \Level1Out83[16] , \Level1Out92[7] , 
        \Level1Out178[6] , \ScanLink225[4] , \Level4Out120[5] , 
        \Level2Out210[7] , \Level4Out8[8] , \Level1Out96[22] , 
        \Level2Out110[31] , \Level8Out24[3] , \Level1Out109[19] , 
        \Level2Out170[2] , \Level2Out146[29] , \Level1Out18[13] , 
        \Level1Out40[1] , \Level2Out110[28] , \Level2Out146[30] , 
        \Level1Out43[2] , \ScanLink119[18] , \ScanLink121[5] , 
        \ScanLink122[6] , \Level8Out56[17] , \ScanLink242[3] , 
        \ScanLink197[30] , \Level4Out224[4] , \Level1Out78[17] , 
        \ScanLink197[29] , \ScanLink241[0] , \Level2Out12[19] , 
        \Level4Out144[1] , \Level2Out44[18] , \Level1Out91[4] , 
        \Level1Load106[0] , \Level1Out187[31] , \Level4Out196[7] , 
        \Level1Out102[15] , \Level1Out117[21] , \Level1Out134[10] , 
        \Level1Out141[20] , \Level1Out187[28] , \Level2Out0[22] , 
        \Level1Out162[11] , \Level2Out56[4] , \Level32Out224[16] , 
        \Level2Out158[11] , \Level1Out177[25] , \Level2Out138[15] , 
        \ScanLink11[17] , \ScanLink32[26] , \ScanLink63[1] , \ScanLink112[14] , 
        \Level1Out121[24] , \Level1Out154[14] , \ScanLink220[9] , 
        \Level16Out224[23] , \ScanLink167[24] , \Level2Out82[10] , 
        \Level2Load208[0] , \ScanLink131[25] , \ScanLink144[15] , 
        \Level2Out84[2] , \Level1Out200[1] , \ScanLink107[20] , 
        \ScanLink124[11] , \ScanLink151[21] , \Level1Out160[4] , 
        \Level2Out112[8] , \ScanLink172[10] , \ScanLink191[9] , 
        \Level1Out203[2] , \ScanLink47[16] , \ScanLink27[12] , 
        \ScanLink64[27] , \ScanLink239[22] , \ScanLink71[13] , 
        \Level1Out163[7] , \Level2Out48[8] , \ScanLink189[11] , 
        \ScanLink52[22] , \ScanLink60[2] , \Level1Out199[10] , 
        \Level1Out249[27] , \Level2Out206[17] , \Level4Out92[10] , 
        \Level8Load192[0] , \Level32Out0[9] , \ScanLink19[9] , 
        \Level1Out21[8] , \Level2Out180[21] , \Level1Out88[30] , 
        \Level1Out89[6] , \Level1Out94[9] , \ScanLink124[22] , 
        \Level1Load219[0] , \Level2Out230[12] , \Level2Out250[16] , 
        \Level4Out60[9] , \Level4Out184[23] , \Level1Out229[23] , 
        \ScanLink139[7] , \ScanLink151[12] , \Level1Out102[26] , 
        \Level1Out104[0] , \ScanLink107[13] , \ScanLink112[27] , 
        \ScanLink172[23] , \Level2Out82[23] , \Level2Out216[9] , 
        \Level2Load16[0] , \ScanLink124[8] , \ScanLink131[16] , 
        \ScanLink167[17] , \Level16Out0[28] , \ScanLink144[26] , 
        \Level16Out0[31] , \Level1Out177[16] , \Level2Out138[26] , 
        \Level1Out121[17] , \Level1Out134[23] , \Level1Out154[27] , 
        \Level2Out32[0] , \Level16Out224[10] , \Level1Out141[13] , 
        \Level1Out88[29] , \Level1Out117[12] , \Level2Out158[22] , 
        \Level1Out162[22] , \Level32Out224[25] , \Level1Out199[23] , 
        \Level1Out229[10] , \Level2Out208[5] , \Level2Out230[21] , 
        \Level4Out184[10] , \Level1Out73[28] , \ScanLink0[5] , \ScanLink3[6] , 
        \ScanLink5[8] , \ScanLink11[24] , \Level1Out25[30] , 
        \Level1Out249[14] , \Level4Out92[23] , \Level1Out25[29] , 
        \Level1Out50[19] , \Level2Out168[0] , \Level2Out206[24] , 
        \Level1Out73[31] , \Level2Out250[25] , \Level2Out180[12] , 
        \ScanLink27[21] , \ScanLink52[11] , \Level1Out58[3] , \ScanLink71[20] , 
        \ScanLink189[22] , \ScanLink32[15] , \ScanLink47[25] , 
        \ScanLink64[14] , \Level1Out107[3] , \ScanLink239[11] , 
        \ScanLink15[15] , \ScanLink20[0] , \Level1Out21[18] , 
        \Level1Out54[31] , \Level1Out77[19] , \Level1Out188[26] , 
        \Level2Out234[10] , \Level4Out180[21] , \Level16Out128[26] , 
        \Level2Out202[15] , \Level4Out96[12] , \Level1Out238[15] , 
        \ScanLink23[10] , \Level1Out54[28] , \Level2Out184[23] , 
        \Level32Out128[13] , \Level2Out254[14] , \ScanLink75[11] , 
        \Level1Out123[5] , \Level2Out68[27] , \ScanLink228[14] , 
        \Level64Out0[1] , \ScanLink36[24] , \ScanLink56[20] , 
        \Level1Out243[0] , \ScanLink43[14] , \ScanLink248[10] , 
        \ScanLink23[3] , \ScanLink60[25] , \ScanLink198[27] , 
        \Level4Load208[0] , \ScanLink36[17] , \ScanLink43[27] , 
        \ScanLink44[4] , \Level1Out62[9] , \ScanLink103[22] , 
        \ScanLink120[13] , \ScanLink155[23] , \Level32Out128[9] , 
        \Level1Out120[6] , \ScanLink176[12] , \Level1Out106[17] , 
        \ScanLink116[16] , \ScanLink163[26] , \ScanLink135[27] , 
        \ScanLink140[17] , \Level2Out86[12] , \Level1Out240[3] , 
        \Level1Out173[27] , \Level1Out125[26] , \Level1Out150[16] , 
        \Level1Out113[23] , \Level1Out130[12] , \Level1Out145[22] , 
        \Level1Out166[13] , \Level2Out16[6] , \Level16Out240[25] , 
        \ScanLink60[16] , \Level1Out147[1] , \ScanLink198[14] , 
        \Level1Out188[8] , \ScanLink248[23] , \ScanLink7[31] , 
        \ScanLink15[26] , \Level4Out96[9] , \Level1Out18[1] , \ScanLink75[22] , 
        \ScanLink23[23] , \ScanLink56[13] , \ScanLink228[27] , 
        \Level2Out68[14] , \Level1Out227[4] , \ScanLink95[1] , \ScanLink96[2] , 
        \Level1Out238[26] , \Level1Out130[21] , \ScanLink167[9] , 
        \Level1Out195[7] , \Level2Out128[2] , \Level2Out202[26] , 
        \Level4Out96[21] , \Level2Out254[27] , \Level2Out184[10] , 
        \Level2Out234[23] , \Level2Out248[7] , \Level32Out128[20] , 
        \Level1Out188[15] , \Level4Out180[12] , \Level16Out128[15] , 
        \Level16Out240[16] , \Level1Out145[11] , \Level1Out196[4] , 
        \Level4Out88[5] , \Level1Out106[24] , \Level1Out113[10] , 
        \Level1Out166[20] , \Level1Out239[8] , \ScanLink7[28] , 
        \Level1Out125[15] , \Level1Out173[14] , \ScanLink38[2] , 
        \ScanLink47[7] , \ScanLink116[25] , \Level1Out150[25] , 
        \Level2Out72[2] , \ScanLink135[14] , \Level1Out144[2] , 
        \ScanLink219[0] , \Level2Out86[21] , \ScanLink163[15] , 
        \Level1Out67[4] , \ScanLink103[11] , \ScanLink120[20] , 
        \ScanLink140[24] , \ScanLink179[5] , \Level1Out224[7] , 
        \ScanLink155[10] , \Level1Out138[4] , \ScanLink176[21] , 
        \ScanLink193[18] , \Level2Load250[0] , \Level4Out160[7] , 
        \Level1Out69[12] , \ScanLink105[3] , \Level2Out16[28] , 
        \Level2Out40[30] , \Level1Out183[19] , \Level2Out16[31] , 
        \Level2Out40[29] , \Level4Out200[2] , \Level8Out192[16] , 
        \Level16Out176[9] , \Level32Out160[19] , \Level1Out79[8] , 
        \Level1Out87[27] , \Level1Out126[8] , \Level2Out4[13] , 
        \Level4Out88[19] , \Level1Out92[13] , \Level1Load241[0] , 
        \Level2Out142[18] , \Level2Out154[4] , \Level1Out178[18] , 
        \ScanLink168[19] , \Level2Out114[19] , \Level2Out234[1] , 
        \Level1Out64[7] , \ScanLink106[0] , \Level2Out186[2] , 
        \Level8Out32[22] , \Level16Out208[0] , \Level2Out10[8] , 
        \Level2Out98[19] , \Level8Out64[23] , \Level8Out192[25] , 
        \Level1Out5[18] , \Level1Out69[21] , \Level2Out4[20] , 
        \Level1Load22[0] , \ScanLink41[9] , \ScanLink48[18] , \ScanLink161[7] , 
        \Level1Out193[9] , \Level1Out210[31] , \Level1Out233[19] , 
        \Level1Out246[29] , \Level1Out210[28] , \Level1Out246[30] , 
        \ScanLink200[30] , \ScanLink201[2] , \ScanLink256[28] , 
        \ScanLink223[18] , \Level4Out104[3] , \ScanLink200[29] , 
        \ScanLink256[31] , \ScanLink90[31] , \ScanLink90[28] , 
        \ScanLink202[1] , \Level8Out32[11] , \Level8Out64[10] , 
        \Level1Out92[20] , \ScanLink162[4] , \Level2Out130[0] , 
        \ScanLink6[22] , \Level1Out16[7] , \Level1Out87[14] , 
        \Level2Out250[5] , \ScanLink98[4] , \Level1Out222[9] , 
        \Level8Out64[1] , \Level1Out149[7] , \Level1Out154[8] , 
        \Level1Load233[0] , \Level2Out126[4] , \ScanLink214[5] , 
        \Level2Out246[1] , \Level8Out72[5] , \Level8Out120[24] , 
        \Level8Out176[25] , \ScanLink6[11] , \Level1Out15[4] , 
        \Level1Out16[24] , \Level1Out20[21] , \Level1Out55[11] , 
        \Level1Out98[15] , \ScanLink174[0] , \Level1Out229[2] , 
        \Level2Out62[8] , \ScanLink217[6] , \Level4Out112[7] , \ScanLink49[1] , 
        \Level1Out63[14] , \Level1Out76[20] , \ScanLink86[8] , 
        \ScanLink177[3] , \Level2Out138[8] , \Level2Out216[18] , 
        \ScanLink22[30] , \ScanLink22[29] , \Level1Out35[15] , 
        \Level1Out40[25] , \Level2Load222[0] , \Level2Out240[19] , 
        \Level8Out248[27] , \ScanLink57[19] , \Level1Load182[0] , 
        \Level1Out198[2] , \Level8Out80[10] , \ScanLink249[30] , 
        \ScanLink249[29] , \ScanLink74[31] , \ScanLink74[28] , 
        \Level64Out64[15] , \ScanLink33[9] , \Level1Out72[3] , 
        \Level1Out98[26] , \ScanLink110[4] , \Level1Out144[31] , 
        \Level2Out190[6] , \Level1Out112[29] , \Level1Out167[19] , 
        \Level2Out128[29] , \Level1Out144[28] , \Level8Out120[17] , 
        \Level2Out128[30] , \ScanLink102[28] , \Level1Out112[30] , 
        \Level8Out176[16] , \Level1Out131[18] , \ScanLink154[30] , 
        \ScanLink177[18] , \Level1Load50[0] , \ScanLink102[31] , 
        \ScanLink154[29] , \ScanLink121[19] , \Level1Out250[9] , 
        \Level2Out142[0] , \Level8Out16[1] , \Level2Out222[5] , 
        \Level64Out64[26] , \Level1Out0[23] , \Level1Out0[10] , 
        \Level1Out4[21] , \Level1Out4[12] , \Level1Out10[9] , 
        \Level1Out16[17] , \Level2Out18[0] , \Level8Out80[23] , 
        \Level1Out20[12] , \Level1Out35[26] , \Level1Out63[27] , 
        \Level8Out248[14] , \Level1Out40[16] , \Level4Out176[3] , 
        \Level4Out212[29] , \ScanLink51[3] , \Level1Out55[22] , 
        \Level1Out71[0] , \Level1Out76[13] , \ScanLink113[7] , 
        \Level4Out212[30] , \Level4Out244[31] , \Level4Out216[6] , 
        \Level4Out244[28] , \Level1Out152[6] , \Level1Out179[21] , 
        \Level2Out160[10] , \Level4Out24[20] , \Level4Out152[17] , 
        \Level4Out104[16] , \ScanLink83[5] , \ScanLink84[16] , 
        \Level1Out119[25] , \Level1Out232[3] , \Level2Out136[11] , 
        \Level4Out12[25] , \Level4Out72[21] , \Level2Load92[0] , 
        \Level2Out100[14] , \Level2Out156[15] , \Level4Out164[12] , 
        \Level4Out132[13] , \Level4Out44[24] , \ScanLink109[24] , 
        \Level1Out180[0] , \ScanLink169[20] , \Level64Out0[11] , 
        \ScanLink29[16] , \ScanLink91[22] , \Level2Out64[6] , \ScanLink49[12] , 
        \ScanLink80[6] , \Level1Out183[3] , \ScanLink201[23] , 
        \Level2Out34[20] , \ScanLink211[8] , \Level2Out62[21] , 
        \ScanLink187[15] , \ScanLink222[12] , \ScanLink192[21] , 
        \ScanLink242[16] , \Level32Out224[0] , \ScanLink214[17] , 
        \ScanLink237[26] , \Level2Out54[24] , \ScanLink52[0] , 
        \Level1Out151[5] , \Level1Out182[20] , \Level1Out252[17] , 
        \Level1Out227[27] , \Level1Out204[16] , \Level1Out211[22] , 
        \Level1Out247[23] , \ScanLink28[8] , \Level1Out197[14] , 
        \Level1Out231[0] , \Level2Out208[13] , \Level1Out232[13] , 
        \ScanLink35[7] , \ScanLink84[25] , \ScanLink91[11] , \ScanLink169[13] , 
        \Level2Out196[8] , \Level64Out0[22] , \ScanLink109[17] , 
        \Level2Out156[26] , \ScanLink36[4] , \Level1Out69[2] , 
        \Level1Out119[16] , \Level1Out136[2] , \Level4Out12[16] , 
        \Level4Out164[21] , \Level4Out44[17] , \Level2Out100[27] , 
        \Level4Out28[3] , \Level4Out132[20] , \Level1Out93[19] , 
        \Level1Out179[12] , \Level2Out136[22] , \Level2Out160[23] , 
        \Level4Out24[13] , \Level4Out152[24] , \Level4Out72[12] , 
        \Level4Out104[25] , \Level1Out135[1] , \Level1Out211[11] , 
        \Level1Out197[27] , \Level1Out232[20] , \Level1Out247[10] , 
        \Level2Out208[20] , \ScanLink29[25] , \ScanLink49[21] , 
        \Level1Out68[18] , \ScanLink108[6] , \Level1Out255[4] , 
        \Level2Out188[4] , \Level16Out96[18] , \Level1Out182[13] , 
        \ScanLink192[12] , \Level1Out204[25] , \Level1Out227[14] , 
        \Level1Out252[24] , \ScanLink214[24] , \ScanLink237[15] , 
        \ScanLink242[25] , \ScanLink115[9] , \Level2Out54[17] , 
        \ScanLink201[10] , \Level2Out34[13] , \ScanLink187[26] , 
        \ScanLink222[21] , \Level1Out215[20] , \Level2Out62[12] , 
        \Level1Out6[2] , \ScanLink11[1] , \ScanLink12[2] , \Level1Out193[16] , 
        \Level1Out236[11] , \Level1Out243[21] , \Level1Out19[19] , 
        \ScanLink38[20] , \Level1Out53[8] , \Level1Out111[7] , 
        \Level1Out186[22] , \Level1Out223[25] , \Level1Out200[14] , 
        \Level4Out208[13] , \ScanLink196[23] , \ScanLink246[14] , 
        \ScanLink233[24] , \Level2Out50[26] , \ScanLink58[24] , 
        \ScanLink210[15] , \ScanLink80[14] , \ScanLink95[20] , 
        \ScanLink183[17] , \ScanLink205[21] , \ScanLink226[10] , 
        \ScanLink253[20] , \Level2Out30[22] , \Level2Out66[23] , 
        \Level4Out12[9] , \Level8Out0[25] , \ScanLink118[12] , 
        \Level2Out88[16] , \ScanLink252[9] , \Level2Out24[4] , 
        \Level1Out97[31] , \Level1Out168[17] , \ScanLink178[16] , 
        \Level2Out4[6] , \Level4Out16[27] , \Level2Out104[16] , 
        \Level2Out152[17] , \Level4Out160[10] , \Level4Out136[11] , 
        \Level4Out40[26] , \Level1Out97[28] , \Level1Out112[4] , 
        \Level4Out20[22] , \Level2Out164[12] , \Level4Out156[15] , 
        \Level4Out100[14] , \ScanLink58[17] , \Level1Out108[13] , 
        \Level2Out132[13] , \Level2Out160[8] , \Level4Out76[23] , 
        \ScanLink205[12] , \Level1Out208[9] , \Level2Out30[11] , 
        \ScanLink38[13] , \ScanLink183[24] , \ScanLink226[23] , 
        \Level8Out0[16] , \ScanLink196[10] , \ScanLink253[13] , 
        \Level2Out66[10] , \ScanLink210[26] , \ScanLink233[17] , 
        \ScanLink246[27] , \Level2Out50[15] , \Level32Out160[3] , 
        \ScanLink76[6] , \ScanLink148[4] , \Level1Out215[6] , 
        \Level1Out175[3] , \Level1Out186[11] , \Level1Out200[27] , 
        \Level1Out223[16] , \Level8Out232[19] , \Level1Out215[13] , 
        \ScanLink228[1] , \Level4Out208[20] , \Level1Out193[25] , 
        \Level1Out236[22] , \Level1Out0[19] , \Level1Out0[5] , \ScanLink2[20] , 
        \Level1Out5[1] , \Level1Out29[0] , \Level1Out243[12] , \ScanLink75[5] , 
        \Level1Out108[20] , \Level2Out92[6] , \Level2Out164[21] , 
        \Level4Out20[11] , \Level4Out156[26] , \Level1Out216[5] , 
        \Level4Out76[10] , \Level2Out132[20] , \Level2Out152[24] , 
        \Level4Out100[27] , \Level4Out160[23] , \ScanLink80[27] , 
        \Level1Out168[24] , \Level1Out176[0] , \Level4Out16[14] , 
        \Level2Load64[0] , \Level4Out40[15] , \Level2Out104[25] , 
        \Level4Out68[1] , \Level4Out136[22] , \ScanLink156[8] , 
        \ScanLink178[25] , \Level2Out40[0] , \ScanLink199[1] , 
        \Level1Out12[26] , \Level1Out48[9] , \ScanLink95[13] , 
        \ScanLink118[21] , \Level2Out88[25] , \Level128Out128[7] , 
        \ScanLink188[31] , \Level1Out67[16] , \Level1Out87[0] , 
        \ScanLink188[28] , \Level1Out117[9] , \ScanLink137[1] , 
        \Level2Out78[31] , \Level2Out78[28] , \Level4Out180[3] , 
        \Level4Out232[0] , \Level64Out192[22] , \Level1Out24[23] , 
        \Level1Out31[17] , \Level1Out44[27] , \Level1Out55[6] , 
        \Level1Out51[13] , \Level1Out198[30] , \Level4Out0[0] , 
        \Level32Out96[25] , \Level1Out56[5] , \Level1Out72[22] , 
        \Level4Out152[5] , \Level4Out216[18] , \Level1Out198[29] , 
        \Level4Out240[19] , \Level8Out112[23] , \ScanLink2[13] , 
        \Level1Out12[15] , \Level1Out24[10] , \Level1Out84[3] , 
        \Level1Out89[23] , \Level1Out116[18] , \ScanLink134[2] , 
        \Level1Out135[30] , \Level8Out144[22] , \Level4Out68[28] , 
        \Level1Out163[28] , \Level1Out109[5] , \Level1Out135[29] , 
        \ScanLink254[7] , \Level4Out68[31] , \Level1Out140[19] , 
        \Level1Out163[31] , \ScanLink106[19] , \ScanLink125[31] , 
        \ScanLink125[28] , \ScanLink173[29] , \Level2Out206[3] , 
        \Level8Out32[7] , \ScanLink150[18] , \ScanLink173[30] , 
        \Level2Out2[8] , \ScanLink249[8] , \Level2Out166[6] , \Level1Out31[2] , 
        \Level1Out51[20] , \Level32Out96[16] , \Level1Out72[11] , 
        \ScanLink153[5] , \Level2Out212[29] , \Level64Out192[11] , 
        \ScanLink26[18] , \Level1Out31[24] , \Level1Out67[25] , 
        \Level1Out228[29] , \Level2Out244[31] , \ScanLink233[0] , 
        \Level2Out212[30] , \Level1Out44[14] , \Level1Out228[30] , 
        \Level2Out244[28] , \Level4Out136[1] , \Level1Load174[0] , 
        \ScanLink238[28] , \ScanLink181[3] , \Level2Out58[2] , 
        \Level1Out213[8] , \ScanLink238[31] , \Level1Out32[1] , 
        \ScanLink53[31] , \ScanLink53[28] , \ScanLink70[8] , \ScanLink70[19] , 
        \Level1Out89[10] , \ScanLink150[6] , \ScanLink182[0] , 
        \Level2Out94[8] , \Level4Out248[8] , \Level8Out56[3] , 
        \Level2Out102[2] , \Level1Out4[31] , \ScanLink28[1] , \Level1Out74[4] , 
        \ScanLink230[3] , \Level4Out128[30] , \Level4Out128[29] , 
        \Level8Out112[10] , \Level8Out144[11] , \ScanLink116[3] , 
        \Level1Out68[11] , \Level1Out86[24] , \ScanLink91[18] , 
        \Level2Out196[1] , \Level1Out93[10] , \Level2Out224[2] , 
        \Level8Out168[14] , \Level4Out132[30] , \Level4Out164[28] , 
        \Level2Out144[7] , \Level4Out132[29] , \Level4Out164[31] , 
        \Level16Out96[11] , \Level1Out135[8] , \Level1Out211[18] , 
        \Level1Out232[30] , \Level32Out96[3] , \Level1Out4[28] , 
        \Level1Out232[29] , \Level2Out208[30] , \Level8Out200[17] , 
        \ScanLink6[18] , \Level1Out10[0] , \ScanLink49[31] , \Level1Out77[7] , 
        \ScanLink115[0] , \ScanLink201[19] , \Level1Out247[19] , 
        \Level1Load252[0] , \Level1Out248[2] , \Level2Out208[29] , 
        \ScanLink222[31] , \ScanLink222[28] , \ScanLink49[28] , 
        \Level1Out128[7] , \Level4Out36[6] , \Level1Out86[17] , 
        \Level1Out93[23] , \Level1Out179[31] , \Level2Out240[6] , 
        \Level4Out24[29] , \Level8Out168[27] , \Level2Out136[18] , 
        \Level2Out160[19] , \Level4Out72[31] , \Level4Out24[30] , 
        \ScanLink169[30] , \Level1Out179[28] , \Level2Out120[3] , 
        \Level4Out72[28] , \ScanLink169[29] , \ScanLink172[7] , 
        \Level64Out0[18] , \Level1Out13[3] , \Level1Out180[9] , 
        \ScanLink212[2] , \Level1Load31[0] , \ScanLink52[9] , \ScanLink171[4] , 
        \ScanLink192[28] , \Level4Load104[0] , \Level32Out224[9] , 
        \ScanLink192[31] , \ScanLink211[1] , \Level2Out34[29] , 
        \Level2Out62[31] , \Level1Out231[9] , \Level2Out34[30] , 
        \Level2Out62[28] , \Level4Out52[2] , \Level8Out200[24] , 
        \Level1Out182[29] , \Level16Out96[22] , \Level1Out68[22] , 
        \Level1Out112[20] , \Level1Out167[10] , \Level1Out182[30] , 
        \Level4Out80[4] , \Level2Out128[20] , \Level1Out131[11] , 
        \Level1Out144[21] , \ScanLink8[4] , \ScanLink14[16] , \ScanLink33[0] , 
        \ScanLink102[21] , \Level1Out107[14] , \Level1Out124[25] , 
        \Level1Out151[15] , \Level1Out172[24] , \ScanLink117[15] , 
        \ScanLink134[24] , \ScanLink141[14] , \Level2Out148[24] , 
        \Level1Out250[0] , \Level8Out16[8] , \ScanLink162[25] , 
        \Level4Out208[3] , \Level1Out130[5] , \ScanLink177[11] , 
        \Level4Out168[6] , \Level2Out92[25] , \Level64Out192[2] , 
        \ScanLink121[10] , \ScanLink154[20] , \Level2Out142[9] , 
        \ScanLink249[13] , \ScanLink22[13] , \ScanLink37[27] , 
        \ScanLink61[26] , \ScanLink199[24] , \Level2Out18[9] , 
        \Level1Out253[3] , \ScanLink42[17] , \ScanLink30[3] , 
        \Level1Out55[18] , \ScanLink57[23] , \ScanLink57[4] , \Level1Out71[9] , 
        \ScanLink74[12] , \Level1Out133[6] , \ScanLink229[17] , 
        \Level2Out220[27] , \Level4Out212[20] , \Level16Out160[4] , 
        \ScanLink102[12] , \Level1Out189[25] , \Level1Out239[16] , 
        \Level4Out244[21] , \Level8Out184[3] , \Level2Out216[22] , 
        \Level4Out224[25] , \Level2Out190[14] , \Level2Out240[23] , 
        \ScanLink121[23] , \ScanLink169[6] , \ScanLink177[22] , 
        \Level2Out92[16] , \Level2Out246[8] , \Level1Out234[4] , 
        \ScanLink134[17] , \ScanLink154[13] , \ScanLink85[2] , 
        \Level1Out107[27] , \ScanLink117[26] , \ScanLink141[27] , 
        \Level1Out124[16] , \Level1Out154[1] , \ScanLink209[3] , 
        \ScanLink162[16] , \Level1Out151[26] , \Level2Out62[1] , 
        \ScanLink174[9] , \Level2Out148[17] , \Level1Out112[13] , 
        \Level1Out172[17] , \Level1Out131[22] , \Level1Out167[23] , 
        \Level2Out128[13] , \Level1Out144[12] , \Level1Out186[7] , 
        \Level1Out189[16] , \Level2Out190[27] , \Level2Out216[11] , 
        \Level2Out240[10] , \Level4Out224[16] , \Level16Out64[5] , 
        \Level1Out76[30] , \Level1Out185[4] , \ScanLink14[25] , 
        \Level1Out20[31] , \Level1Out20[28] , \Level2Out220[14] , 
        \ScanLink49[8] , \Level1Out76[29] , \Level4Out212[13] , 
        \ScanLink86[1] , \Level1Out239[25] , \Level4Out244[12] , 
        \ScanLink22[20] , \ScanLink57[10] , \Level2Out138[1] , 
        \Level1Out237[7] , \ScanLink61[15] , \ScanLink74[21] , 
        \Level1Out157[2] , \ScanLink199[17] , \ScanLink229[24] , 
        \Level8Out80[19] , \ScanLink249[20] , \Level1Out24[19] , 
        \ScanLink37[14] , \ScanLink42[24] , \ScanLink54[7] , 
        \Level1Out228[20] , \Level2Out212[20] , \Level4Out220[27] , 
        \Level64Out192[18] , \ScanLink233[9] , \Level2Out194[16] , 
        \Level2Out244[21] , \Level4Out136[8] , \Level4Out216[22] , 
        \Level1Out51[29] , \Level2Out224[25] , \Level1Out198[13] , 
        \Level1Out248[24] , \Level8Out48[6] , \Level4Out240[23] , 
        \ScanLink2[30] , \ScanLink2[29] , \Level1Out3[6] , \ScanLink10[14] , 
        \ScanLink26[11] , \Level1Out51[30] , \Level1Out72[18] , 
        \ScanLink53[21] , \ScanLink70[1] , \ScanLink70[10] , \Level1Out173[4] , 
        \ScanLink188[12] , \Level2Out18[16] , \Level2Out78[12] , 
        \ScanLink33[25] , \ScanLink65[24] , \ScanLink238[21] , 
        \Level1Out213[1] , \ScanLink46[15] , \Level16Out240[3] , 
        \ScanLink73[2] , \ScanLink106[23] , \Level1Out170[7] , 
        \ScanLink173[13] , \Level2Out96[27] , \Level4Out128[4] , 
        \Level1Out89[19] , \Level1Out103[16] , \ScanLink113[17] , 
        \ScanLink125[12] , \ScanLink150[22] , \ScanLink130[26] , 
        \ScanLink145[16] , \ScanLink182[9] , \Level1Out210[2] , 
        \ScanLink166[27] , \Level4Out248[1] , \Level1Out120[27] , 
        \Level1Out155[17] , \Level2Out94[1] , \Level4Out128[20] , 
        \Level8Out112[19] , \Level1Out176[26] , \Level8Out144[18] , 
        \Level1Out116[22] , \Level1Out163[12] , \Level4Out68[12] , 
        \ScanLink10[27] , \Level1Out32[8] , \Level1Out140[23] , 
        \ScanLink65[17] , \Level1Out117[0] , \Level1Out135[13] , 
        \Level4Out148[24] , \ScanLink238[12] , \Level2Out46[7] , 
        \Level2Out78[21] , \Level16Out144[2] , \ScanLink14[5] , 
        \ScanLink26[22] , \ScanLink33[16] , \ScanLink46[26] , \ScanLink53[12] , 
        \Level1Out48[0] , \ScanLink70[23] , \Level16Out224[7] , 
        \Level1Load69[0] , \Level1Out87[9] , \Level1Out116[11] , 
        \ScanLink137[8] , \ScanLink188[21] , \Level2Out18[25] , 
        \Level1Out198[20] , \Level2Out224[16] , \Level4Out216[11] , 
        \Level1Out248[17] , \Level4Load32[0] , \Level4Out240[10] , 
        \Level2Out178[3] , \Level1Out228[13] , \Level2Out194[25] , 
        \Level2Out212[13] , \Level2Out218[6] , \Level2Out244[12] , 
        \Level4Out220[14] , \Level4Out232[9] , \Level4Out0[9] , 
        \Level4Out68[21] , \Level1Out99[5] , \Level1Out135[20] , 
        \Level1Out163[21] , \Level4Out148[17] , \Level1Out140[10] , 
        \Level1Out120[14] , \Level1Out103[25] , \Level1Out155[24] , 
        \Level2Out22[3] , \Level4Out128[13] , \Level1Out5[8] , \ScanLink9[25] , 
        \ScanLink17[6] , \ScanLink130[15] , \Level1Out176[15] , 
        \Level1Out19[23] , \Level1Out37[5] , \ScanLink106[10] , 
        \ScanLink113[24] , \ScanLink145[25] , \ScanLink249[1] , 
        \Level1Out114[3] , \ScanLink166[14] , \Level2Out96[14] , 
        \ScanLink125[21] , \ScanLink173[20] , \Level2Out2[1] , 
        \ScanLink129[4] , \ScanLink150[11] , \ScanLink155[2] , 
        \Level1Out168[5] , \ScanLink196[19] , \ScanLink235[7] , 
        \Level1Out208[0] , \Level4Out76[4] , \Level2Out30[18] , 
        \Level1Out79[27] , \ScanLink228[8] , \Level2Out66[19] , 
        \Level1Out186[18] , \ScanLink187[4] , \Level4Out208[30] , 
        \Level1Out29[9] , \Level1Out82[26] , \Level4Out208[29] , 
        \Level8Out232[10] , \Level1Out176[9] , \Level2Out104[5] , 
        \Level4Out68[8] , \Level1Out108[30] , \Level2Out164[28] , 
        \Level1Out34[6] , \ScanLink68[3] , \Level1Out97[12] , 
        \Level1Out108[29] , \ScanLink184[7] , \Level2Out132[30] , 
        \Level4Out20[18] , \Level2Out164[31] , \Level4Out76[19] , 
        \ScanLink118[31] , \Level2Out132[29] , \ScanLink118[28] , 
        \ScanLink236[4] , \ScanLink156[1] , \Level2Out40[9] , \ScanLink199[8] , 
        \Level1Out19[10] , \Level1Out81[7] , \Level1Out243[31] , 
        \Level8Out232[23] , \Level1Out215[29] , \Level1Out243[28] , 
        \ScanLink3[23] , \ScanLink9[16] , \ScanLink38[30] , \Level1Out53[1] , 
        \Level1Out79[14] , \ScanLink205[31] , \ScanLink205[28] , 
        \Level1Out215[30] , \Level1Out236[18] , \ScanLink253[30] , 
        \Level2Load104[0] , \ScanLink226[19] , \ScanLink251[3] , 
        \ScanLink253[29] , \Level4Out12[0] , \ScanLink38[29] , 
        \ScanLink131[6] , \Level1Out50[2] , \ScanLink95[30] , \ScanLink252[0] , 
        \ScanLink95[29] , \ScanLink132[5] , \ScanLink11[8] , \Level1Out46[6] , 
        \Level1Out82[15] , \Level1Out97[21] , \Level2Out160[1] , 
        \Level1Out82[4] , \Level4Out160[19] , \Level1Out88[20] , 
        \Level1Out94[0] , \Level1Out104[9] , \Level1Load115[0] , 
        \Level2Out200[4] , \Level4Out136[18] , \Level2Out176[5] , 
        \Level16Out0[21] , \Level8Out48[15] , \Level1Out119[6] , 
        \ScanLink244[4] , \Level2Out216[0] , \ScanLink124[1] , 
        \Level16Out16[24] , \ScanLink3[10] , \Level1Out13[25] , 
        \ScanLink19[0] , \Level1Out73[21] , \Level2Out32[9] , 
        \Level16Out224[19] , \Level1Out25[20] , \Level1Out50[10] , 
        \Level2Out168[9] , \ScanLink247[7] , \Level1Out30[14] , 
        \Level1Out45[24] , \Level1Out45[5] , \Level2Out230[28] , 
        \Level1Out66[15] , \ScanLink127[2] , \Level1Out229[19] , 
        \Level2Out230[31] , \Level4Out184[19] , \ScanLink27[31] , 
        \ScanLink71[29] , \ScanLink239[18] , \Level4Load180[0] , 
        \Level1Out97[3] , \ScanLink27[28] , \ScanLink52[18] , \ScanLink71[30] , 
        \Level16Out16[17] , \Level1Out22[2] , \ScanLink220[0] , 
        \ScanLink63[8] , \Level1Out88[13] , \Level1Out117[31] , 
        \Level1Out141[29] , \Level1Out134[19] , \ScanLink140[5] , 
        \Level1Out141[30] , \Level1Out162[18] , \Level1Out117[28] , 
        \Level2Out158[18] , \ScanLink107[30] , \ScanLink151[28] , 
        \Level8Out48[26] , \ScanLink107[29] , \ScanLink124[18] , 
        \Level2Out112[1] , \ScanLink151[31] , \ScanLink172[19] , 
        \Level1Out1[20] , \Level1Out1[13] , \Level1Out13[16] , 
        \Level1Out30[27] , \Level1Load167[0] , \ScanLink189[18] , 
        \ScanLink192[3] , \Level2Out82[19] , \Level16Out0[12] , 
        \Level1Out200[8] , \ScanLink191[0] , \ScanLink223[3] , 
        \Level2Out48[1] , \Level1Out45[17] , \Level4Out60[0] , 
        \Level2Load176[0] , \Level1Out21[1] , \Level1Out25[13] , 
        \Level1Out66[26] , \Level1Out73[12] , \ScanLink143[6] , 
        \Level2Out180[31] , \Level4Out92[19] , \Level32Out0[0] , 
        \Level1Out199[19] , \Level2Out180[28] , \ScanLink39[23] , 
        \Level1Out40[8] , \Level1Out50[23] , \ScanLink81[17] , 
        \Level1Out102[7] , \Level1Out109[10] , \Level2Out146[20] , 
        \Level2Out110[21] , \Level1Out169[14] , \Level2Out126[24] , 
        \Level2Out170[25] , \Level4Out8[1] , \Level4Out8[17] , 
        \ScanLink179[15] , \Level4Out188[2] , \ScanLink59[27] , 
        \ScanLink94[23] , \ScanLink119[11] , \ScanLink182[14] , 
        \ScanLink241[9] , \ScanLink252[23] , \Level2Out34[7] , 
        \Level2Out12[10] , \Level4Out144[8] , \ScanLink227[13] , 
        \Level2Out44[11] , \ScanLink204[22] , \Level1Out101[4] , 
        \ScanLink197[20] , \ScanLink211[16] , \ScanLink232[27] , 
        \ScanLink247[17] , \Level2Out24[15] , \Level16Out32[3] , 
        \Level2Out72[14] , \Level1Out187[21] , \Level1Out201[17] , 
        \Level1Out222[26] , \Level2Out218[26] , \Level1Out39[3] , 
        \ScanLink65[6] , \ScanLink78[9] , \ScanLink94[10] , \ScanLink119[22] , 
        \Level1Out192[15] , \Level1Out242[22] , \Level1Out214[23] , 
        \Level1Out237[12] , \ScanLink81[24] , \ScanLink189[2] , 
        \Level4Out8[24] , \Level2Out50[3] , \Level1Out166[3] , 
        \ScanLink179[26] , \Level2Out170[16] , \Level1Out96[18] , 
        \Level1Out109[23] , \Level1Out169[27] , \Level2Out126[17] , 
        \Level1Out206[6] , \Level2Out146[13] , \ScanLink66[5] , 
        \Level1Out192[26] , \Level2Out82[5] , \Level2Out110[12] , 
        \Level1Out237[21] , \Level1Out5[11] , \Level1Out18[30] , 
        \Level1Out165[0] , \Level1Out214[10] , \ScanLink238[2] , 
        \Level1Out242[11] , \Level1Out201[24] , \Level1Out18[29] , 
        \ScanLink158[7] , \Level1Out205[5] , \Level1Out187[12] , 
        \Level1Out222[15] , \ScanLink39[10] , \ScanLink211[25] , 
        \Level2Out0[18] , \Level2Out218[15] , \Level2Out24[26] , 
        \Level4Load40[0] , \ScanLink59[14] , \ScanLink182[27] , 
        \ScanLink197[13] , \ScanLink232[14] , \ScanLink247[24] , 
        \Level2Out12[23] , \Level2Out72[27] , \ScanLink227[20] , 
        \ScanLink252[10] , \ScanLink145[8] , \ScanLink204[11] , 
        \Level1Out246[20] , \Level2Out44[22] , \Level4Out240[9] , 
        \ScanLink42[3] , \Level1Out69[31] , \Level1Out141[6] , 
        \Level1Out196[17] , \Level1Out221[3] , \Level1Out210[21] , 
        \Level1Out233[10] , \Level16Out160[16] , \Level2Out4[30] , 
        \Level16Out112[4] , \Level1Out205[15] , \ScanLink48[11] , 
        \Level1Out69[28] , \Level1Out253[14] , \Level2Out4[29] , 
        \Level4Out88[23] , \Level1Out183[23] , \Level1Out226[24] , 
        \Level32Out160[23] , \ScanLink215[14] , \Level2Out20[17] , 
        \ScanLink243[15] , \Level2Out76[16] , \ScanLink3[21] , \ScanLink5[1] , 
        \Level1Out5[22] , \ScanLink26[7] , \ScanLink28[26] , \ScanLink28[15] , 
        \ScanLink186[16] , \ScanLink193[22] , \ScanLink236[25] , 
        \Level1Out193[0] , \ScanLink256[21] , \ScanLink223[11] , 
        \Level2Out16[12] , \ScanLink41[0] , \ScanLink85[15] , \ScanLink90[21] , 
        \ScanLink90[5] , \ScanLink168[23] , \ScanLink200[20] , 
        \Level2Out40[13] , \ScanLink93[6] , \Level2Out74[5] , 
        \Level8Out32[18] , \ScanLink108[27] , \Level1Out190[3] , 
        \ScanLink202[8] , \Level8Out64[19] , \Level1Out118[26] , 
        \Level1Out222[0] , \Level2Out98[23] , \Level2Out122[26] , 
        \Level2Out174[27] , \Level8Out64[8] , \Level1Out178[22] , 
        \Level1Out92[30] , \Level1Out92[29] , \Level2Out114[23] , 
        \Level2Out130[9] , \Level16Out208[15] , \Level2Out142[22] , 
        \Level1Out142[5] , \ScanLink186[25] , \ScanLink200[13] , 
        \ScanLink223[22] , \ScanLink256[12] , \Level2Out16[21] , 
        \Level8Out192[7] , \Level16Out16[5] , \ScanLink48[22] , 
        \ScanLink215[27] , \Level2Out20[24] , \Level2Out40[20] , 
        \ScanLink118[5] , \ScanLink193[11] , \ScanLink236[16] , 
        \Level1Out205[26] , \ScanLink243[26] , \Level2Out76[25] , 
        \Level1Out245[7] , \Level1Out183[10] , \Level1Out226[17] , 
        \Level32Out160[10] , \Level1Out196[24] , \Level1Out253[27] , 
        \Level4Out88[10] , \Level1Out233[23] , \Level1Out246[13] , 
        \Level1Out18[8] , \ScanLink25[4] , \Level1Out79[1] , \Level1Out125[2] , 
        \Level1Out210[12] , \Level2Out198[7] , \Level16Out160[25] , 
        \Level1Out178[11] , \Level1Out246[4] , \Level16Out176[0] , 
        \Level2Out142[11] , \Level16Out208[26] , \Level1Out118[15] , 
        \Level1Out126[1] , \Level2Out114[10] , \Level2Out234[8] , 
        \Level2Out174[14] , \ScanLink85[26] , \ScanLink106[9] , 
        \Level2Out122[15] , \ScanLink108[14] , \Level16Out208[9] , 
        \Level2Out10[1] , \Level2Out98[10] , \ScanLink90[12] , 
        \ScanLink168[10] , \Level1Out147[8] , \Level1Load220[0] , 
        \Level2Load180[0] , \Level1Out188[1] , \ScanLink6[2] , \ScanLink7[21] , 
        \Level1Out17[27] , \Level1Out34[16] , \Level1Out41[26] , 
        \Level4Out96[0] , \Level1Out62[17] , \ScanLink167[0] , 
        \Level1Out21[22] , \Level1Out54[12] , \ScanLink59[2] , 
        \Level1Out77[23] , \Level4Out96[28] , \Level32Out128[30] , 
        \ScanLink207[5] , \Level32Out128[29] , \Level1Out99[16] , 
        \ScanLink164[3] , \Level1Out239[1] , \Level2Out184[19] , 
        \Level4Out44[6] , \Level4Out96[31] , \Level1Load191[0] , 
        \ScanLink95[8] , \Level1Out130[31] , \Level1Out130[28] , 
        \Level1Out145[18] , \Level1Out159[4] , \ScanLink204[6] , 
        \Level1Out166[30] , \ScanLink103[18] , \Level1Out113[19] , 
        \ScanLink120[30] , \ScanLink120[29] , \Level1Out166[29] , 
        \ScanLink155[19] , \ScanLink176[31] , \ScanLink176[28] , 
        \ScanLink219[9] , \Level2Out86[28] , \ScanLink7[12] , 
        \Level1Out17[14] , \Level1Out21[11] , \Level1Out77[10] , 
        \ScanLink88[7] , \Level2Out86[31] , \ScanLink103[4] , 
        \Level2Out136[7] , \Level4Load176[0] , \Level1Out34[25] , 
        \Level1Out54[21] , \Level1Out61[3] , \Level1Out41[15] , 
        \Level2Out234[19] , \Level4Out20[2] , \Level4Out180[31] , 
        \ScanLink20[9] , \ScanLink23[19] , \ScanLink56[30] , \Level1Out62[24] , 
        \Level4Out180[28] , \ScanLink75[18] , \Level1Out243[9] , 
        \ScanLink248[19] , \Level64Out0[8] , \Level1Load43[0] , 
        \ScanLink56[29] , \Level1Out62[0] , \Level2Out152[3] , 
        \Level2Out232[6] , \Level32Out128[0] , \Level1Out99[25] , 
        \ScanLink100[7] , \Level2Out180[5] , \Level1Out13[27] , 
        \Level1Out30[16] , \Level1Out58[8] , \Level1Out97[1] , 
        \Level1Out107[8] , \ScanLink189[30] , \ScanLink189[29] , 
        \Level1Out45[26] , \Level1Out45[7] , \ScanLink19[2] , 
        \Level1Out66[17] , \ScanLink127[0] , \Level1Out199[28] , 
        \Level4Out92[28] , \Level1Out25[22] , \Level1Out73[23] , 
        \Level2Out180[19] , \Level4Out92[31] , \Level1Out50[12] , 
        \ScanLink124[3] , \Level1Out199[31] , \ScanLink247[5] , 
        \Level16Out16[26] , \Level1Out13[14] , \Level1Out21[3] , 
        \Level1Out25[11] , \Level1Out46[4] , \Level1Out50[21] , 
        \Level1Out73[10] , \Level1Out88[22] , \Level1Out119[4] , 
        \Level1Out134[28] , \Level1Out141[18] , \Level1Out162[30] , 
        \ScanLink244[6] , \Level2Out158[30] , \Level1Out94[2] , 
        \Level1Out117[19] , \Level1Out162[29] , \ScanLink124[29] , 
        \Level1Out134[31] , \Level2Out158[29] , \ScanLink151[19] , 
        \Level8Out48[17] , \ScanLink172[31] , \ScanLink172[28] , 
        \Level2Out216[2] , \ScanLink107[18] , \ScanLink124[30] , 
        \Level2Out82[31] , \Level2Out82[28] , \Level2Out176[7] , 
        \Level16Out0[23] , \ScanLink143[4] , \Level32Out0[2] , 
        \Level4Load136[0] , \Level1Out30[25] , \Level1Out45[15] , 
        \ScanLink223[1] , \Level1Out229[31] , \Level4Out60[2] , 
        \Level2Out230[19] , \Level4Out184[31] , \Level1Out66[24] , 
        \Level1Out229[28] , \ScanLink27[19] , \ScanLink52[30] , 
        \ScanLink191[2] , \Level1Out203[9] , \ScanLink239[30] , 
        \Level4Out184[28] , \ScanLink239[29] , \Level2Out48[3] , 
        \ScanLink52[29] , \ScanLink71[18] , \ScanLink60[9] , \Level2Out84[9] , 
        \Level16Out0[10] , \Level1Out1[22] , \Level1Out1[11] , \ScanLink3[12] , 
        \Level1Out22[0] , \ScanLink192[1] , \Level2Out112[3] , 
        \Level8Out48[24] , \Level1Out88[11] , \ScanLink140[7] , 
        \Level16Out16[15] , \Level16Out224[31] , \Level1Out192[17] , 
        \ScanLink220[2] , \Level16Out224[28] , \Level1Out237[10] , 
        \Level1Out242[20] , \Level1Out18[18] , \Level1Out101[6] , 
        \Level1Out201[15] , \Level1Out214[21] , \Level1Out187[23] , 
        \Level2Out0[30] , \Level1Out222[24] , \ScanLink39[21] , 
        \ScanLink211[14] , \Level2Out0[29] , \Level2Out218[24] , 
        \Level2Out24[17] , \Level16Out32[1] , \ScanLink39[12] , 
        \Level1Out43[9] , \ScanLink197[22] , \ScanLink232[25] , 
        \ScanLink247[15] , \Level2Out72[16] , \ScanLink59[25] , 
        \ScanLink182[16] , \ScanLink227[11] , \ScanLink252[21] , 
        \Level2Out12[12] , \ScanLink59[16] , \ScanLink81[15] , 
        \ScanLink94[21] , \ScanLink119[13] , \ScanLink204[20] , 
        \Level2Out44[13] , \Level2Out34[5] , \ScanLink242[8] , 
        \Level4Out8[15] , \Level4Out188[0] , \Level1Out96[30] , 
        \Level1Out96[29] , \Level1Out109[12] , \Level1Out169[16] , 
        \ScanLink179[17] , \Level2Out170[27] , \Level4Out8[3] , 
        \Level2Out126[26] , \Level8Out24[8] , \Level2Out170[9] , 
        \Level2Out146[22] , \Level1Out102[5] , \ScanLink182[25] , 
        \ScanLink227[22] , \ScanLink252[12] , \Level2Out110[23] , 
        \Level1Out218[8] , \Level2Out12[21] , \Level2Out44[20] , 
        \ScanLink204[13] , \ScanLink158[5] , \Level1Out187[10] , 
        \ScanLink197[11] , \ScanLink211[27] , \Level2Out24[24] , 
        \ScanLink247[26] , \Level2Out72[25] , \Level1Out201[26] , 
        \ScanLink232[16] , \Level1Out205[7] , \Level2Out218[17] , 
        \Level1Out222[17] , \Level1Out242[13] , \Level1Out4[19] , 
        \ScanLink5[3] , \Level1Out5[20] , \Level1Out5[13] , \ScanLink28[17] , 
        \Level1Out39[1] , \ScanLink66[7] , \Level1Out192[24] , 
        \Level1Out237[23] , \Level1Out109[21] , \Level1Out165[2] , 
        \Level1Out214[12] , \ScanLink238[0] , \Level1Out206[4] , 
        \Level2Out146[11] , \Level16Out48[9] , \Level2Out82[7] , 
        \Level2Out110[10] , \ScanLink41[2] , \ScanLink65[4] , 
        \Level1Out166[1] , \Level2Out170[14] , \Level1Out169[25] , 
        \Level2Out126[15] , \ScanLink81[26] , \ScanLink146[9] , 
        \Level8Load8[0] , \ScanLink189[0] , \Level4Out8[26] , \ScanLink94[12] , 
        \ScanLink179[24] , \Level2Out50[1] , \ScanLink119[20] , 
        \Level2Out142[20] , \Level16Load48[0] , \Level16Out208[17] , 
        \ScanLink85[17] , \ScanLink93[4] , \Level1Out118[24] , 
        \Level1Out142[7] , \Level1Out178[20] , \Level2Out114[21] , 
        \Level2Out174[25] , \Level1Out222[2] , \Level1Load238[0] , 
        \Level2Out122[24] , \Level2Load198[0] , \ScanLink108[25] , 
        \Level2Out98[21] , \Level1Out190[1] , \ScanLink90[23] , 
        \ScanLink168[21] , \Level2Out74[7] , \ScanLink186[14] , 
        \ScanLink223[13] , \Level2Out16[10] , \Level4Out104[8] , 
        \Level1Out193[2] , \ScanLink200[22] , \ScanLink201[9] , 
        \ScanLink256[23] , \ScanLink42[1] , \ScanLink48[13] , \ScanLink90[7] , 
        \Level2Out40[11] , \ScanLink215[16] , \Level2Out20[15] , 
        \Level1Out141[4] , \ScanLink193[20] , \Level1Out205[17] , 
        \ScanLink236[27] , \ScanLink243[17] , \Level2Out76[14] , 
        \Level16Out112[6] , \Level1Out183[21] , \Level1Out226[26] , 
        \Level32Out160[21] , \Level1Out196[15] , \Level1Out233[12] , 
        \Level1Out253[16] , \Level4Out88[21] , \ScanLink25[6] , 
        \ScanLink38[9] , \ScanLink90[10] , \ScanLink168[12] , 
        \Level1Load189[0] , \Level1Out210[23] , \Level1Out221[1] , 
        \Level1Out246[22] , \Level16Out160[14] , \Level2Out186[9] , 
        \ScanLink85[24] , \Level8Out32[29] , \Level8Out64[31] , 
        \ScanLink108[16] , \Level2Out10[3] , \Level2Out98[12] , 
        \Level8Out32[30] , \Level8Out64[28] , \Level1Out126[3] , 
        \Level2Out174[16] , \Level2Out122[17] , \Level1Out79[3] , 
        \Level1Out92[18] , \Level1Out118[17] , \Level1Out178[13] , 
        \Level1Out246[6] , \Level2Out142[13] , \Level16Out208[24] , 
        \Level2Out114[12] , \ScanLink6[0] , \ScanLink26[5] , 
        \Level1Out196[26] , \Level1Out233[21] , \Level1Out246[11] , 
        \Level2Out198[5] , \ScanLink28[24] , \ScanLink48[20] , 
        \Level1Out69[19] , \Level1Out125[0] , \Level1Out210[10] , 
        \Level16Out176[2] , \Level16Out160[27] , \Level1Out183[12] , 
        \Level1Out205[24] , \Level1Out245[5] , \Level1Out253[25] , 
        \Level2Out4[18] , \Level4Out88[12] , \Level1Out226[15] , 
        \Level32Out160[12] , \ScanLink118[7] , \ScanLink215[25] , 
        \Level2Out20[26] , \ScanLink186[27] , \ScanLink193[13] , 
        \ScanLink243[24] , \Level2Out76[27] , \ScanLink223[20] , 
        \ScanLink236[14] , \ScanLink256[10] , \Level2Out16[23] , 
        \ScanLink105[8] , \ScanLink200[11] , \Level2Out40[22] , 
        \Level4Out200[9] , \Level16Out16[7] , \Level8Out192[5] , 
        \ScanLink7[23] , \ScanLink88[5] , \Level1Out144[9] , \Level2Out136[5] , 
        \Level1Out99[14] , \Level1Out159[6] , \ScanLink204[4] , 
        \ScanLink164[1] , \Level1Out239[3] , \Level1Out17[25] , 
        \Level1Out21[20] , \ScanLink59[0] , \Level1Out77[21] , 
        \Level2Out72[9] , \Level2Out128[9] , \ScanLink96[9] , \Level4Out44[4] , 
        \Level1Out34[14] , \Level1Out54[10] , \ScanLink207[7] , 
        \Level1Out41[24] , \Level2Out234[28] , \Level4Out180[19] , 
        \Level1Out62[15] , \ScanLink167[2] , \Level2Out234[31] , 
        \ScanLink248[31] , \ScanLink248[28] , \ScanLink7[10] , 
        \ScanLink23[31] , \Level1Out188[3] , \Level4Out96[2] , 
        \ScanLink23[28] , \ScanLink75[29] , \ScanLink56[18] , \ScanLink75[30] , 
        \Level1Out99[27] , \Level2Out180[7] , \Level1Out17[16] , 
        \ScanLink23[8] , \Level1Out62[2] , \Level1Out113[31] , 
        \Level1Out130[19] , \ScanLink100[5] , \Level1Out113[28] , 
        \Level1Out145[29] , \Level1Out166[18] , \ScanLink103[30] , 
        \ScanLink120[18] , \Level1Out145[30] , \Level2Out152[1] , 
        \Level1Out34[27] , \Level1Out41[17] , \ScanLink103[29] , 
        \ScanLink155[28] , \Level32Out128[2] , \Level1Load127[0] , 
        \ScanLink155[31] , \ScanLink176[19] , \Level2Out86[19] , 
        \Level2Out232[4] , \Level1Out240[8] , \Level4Out20[0] , 
        \Level1Out62[26] , \Level1Out21[13] , \Level1Out54[23] , 
        \Level1Out77[12] , \Level2Load136[0] , \ScanLink103[6] , 
        \Level2Out184[31] , \Level4Out96[19] , \ScanLink28[3] , 
        \Level1Out61[1] , \Level2Out184[28] , \Level32Out128[18] , 
        \Level1Out68[13] , \Level1Out77[5] , \Level1Load87[0] , 
        \Level1Out128[5] , \ScanLink192[19] , \Level4Out36[4] , 
        \ScanLink115[2] , \Level1Out248[0] , \Level2Out34[18] , 
        \Level2Out62[19] , \Level8Out200[15] , \Level32Out96[1] , 
        \Level16Out96[13] , \Level1Out69[9] , \Level1Out86[26] , 
        \Level1Out182[18] , \Level1Out136[9] , \Level2Out144[5] , 
        \Level4Out28[8] , \Level2Out136[30] , \Level2Out224[0] , 
        \Level8Out168[16] , \Level4Out24[18] , \Level1Out93[12] , 
        \Level1Out179[19] , \Level2Out136[29] , \Level2Out160[28] , 
        \Level2Out160[31] , \Level2Out196[3] , \Level4Out72[19] , 
        \Level1Out68[20] , \Level1Out74[6] , \ScanLink169[18] , 
        \Level64Out0[29] , \Level64Out0[30] , \ScanLink116[1] , 
        \Level16Out96[20] , \Level1Out211[30] , \Level1Out211[29] , 
        \Level4Out80[6] , \Level1Out247[31] , \Level1Out232[18] , 
        \Level1Out247[28] , \Level8Out200[26] , \Level1Out10[2] , 
        \Level1Out13[1] , \Level1Out183[8] , \ScanLink201[31] , 
        \ScanLink201[28] , \Level2Out208[18] , \Level2Load144[0] , 
        \Level4Out52[0] , \ScanLink211[3] , \ScanLink222[19] , 
        \ScanLink49[19] , \ScanLink91[30] , \ScanLink171[6] , \ScanLink172[5] , 
        \ScanLink212[0] , \Level4Load4[0] , \Level1Out20[19] , \ScanLink51[8] , 
        \ScanLink91[29] , \Level2Out120[1] , \Level8Out168[25] , 
        \Level1Out55[29] , \Level1Out86[15] , \Level1Out93[21] , 
        \Level4Out164[19] , \Level1Load155[0] , \Level1Out232[8] , 
        \Level1Out189[27] , \Level2Out240[4] , \Level4Out132[18] , 
        \Level2Out190[16] , \Level2Out216[20] , \Level2Out240[21] , 
        \Level4Out224[27] , \Level4Out176[8] , \Level2Out220[25] , 
        \Level4Out212[22] , \Level1Out55[30] , \Level1Out76[18] , 
        \Level1Out239[14] , \Level4Out244[23] , \Level8Out184[1] , 
        \Level1Out0[31] , \Level1Out0[7] , \ScanLink2[18] , \Level1Out3[4] , 
        \ScanLink6[30] , \ScanLink6[29] , \ScanLink8[6] , \ScanLink14[27] , 
        \ScanLink14[14] , \ScanLink22[11] , \ScanLink57[21] , \ScanLink30[1] , 
        \ScanLink61[24] , \ScanLink74[10] , \Level1Out133[4] , 
        \ScanLink229[15] , \Level16Out160[6] , \ScanLink199[26] , 
        \Level8Out80[28] , \ScanLink249[11] , \ScanLink33[2] , 
        \ScanLink37[25] , \ScanLink42[15] , \Level1Out253[1] , 
        \Level8Out80[31] , \ScanLink102[23] , \Level2Out92[27] , 
        \Level4Out168[4] , \Level64Out192[0] , \ScanLink121[12] , 
        \Level1Out130[7] , \ScanLink177[13] , \Level1Out72[8] , 
        \Level1Out107[16] , \ScanLink117[17] , \ScanLink134[26] , 
        \ScanLink154[22] , \ScanLink141[16] , \Level4Out208[1] , 
        \Level1Out250[2] , \Level1Out124[27] , \ScanLink162[27] , 
        \Level1Out151[17] , \Level2Out148[26] , \Level1Out112[22] , 
        \Level1Out172[26] , \Level1Out131[13] , \Level1Out167[12] , 
        \Level2Out128[22] , \Level1Out144[23] , \ScanLink249[22] , 
        \ScanLink22[22] , \ScanLink37[16] , \ScanLink61[17] , 
        \Level1Out157[0] , \ScanLink199[15] , \Level1Out198[9] , 
        \ScanLink42[26] , \ScanLink54[5] , \ScanLink57[12] , \ScanLink74[23] , 
        \Level1Out237[5] , \ScanLink229[26] , \Level2Out220[16] , 
        \Level4Out212[11] , \Level1Load29[0] , \ScanLink86[3] , 
        \Level1Out185[6] , \Level1Out239[27] , \Level2Out138[3] , 
        \Level4Load72[0] , \Level4Out244[10] , \ScanLink177[8] , 
        \Level2Out216[13] , \Level4Out224[14] , \Level16Out64[7] , 
        \Level1Out189[14] , \Level2Out190[25] , \Level2Out240[12] , 
        \ScanLink85[0] , \Level1Out167[21] , \Level2Out128[11] , 
        \Level1Out112[11] , \Level1Out131[20] , \Level1Out144[10] , 
        \Level1Out186[5] , \Level1Out124[14] , \Level1Out151[24] , 
        \Level2Out62[3] , \ScanLink57[6] , \Level1Out107[25] , 
        \Level1Out172[15] , \Level1Out229[9] , \ScanLink134[15] , 
        \ScanLink141[25] , \Level2Out148[15] , \ScanLink102[10] , 
        \ScanLink117[24] , \ScanLink162[14] , \ScanLink209[1] , 
        \Level1Out154[3] , \ScanLink177[20] , \Level2Out92[14] , 
        \Level1Out116[20] , \ScanLink121[21] , \ScanLink154[11] , 
        \Level1Out234[6] , \ScanLink169[4] , \Level4Out68[10] , 
        \Level1Out120[25] , \Level1Out135[11] , \Level1Out163[10] , 
        \Level2Out46[5] , \Level1Out140[21] , \Level4Out148[26] , 
        \ScanLink10[16] , \ScanLink65[26] , \ScanLink73[0] , 
        \Level1Out103[14] , \Level1Out155[15] , \ScanLink230[8] , 
        \Level4Out128[22] , \ScanLink106[21] , \ScanLink113[15] , 
        \ScanLink130[24] , \Level1Out176[24] , \ScanLink145[14] , 
        \Level4Out248[3] , \Level1Out210[0] , \Level8Out56[8] , 
        \ScanLink166[25] , \Level2Out94[3] , \Level4Out128[6] , 
        \ScanLink125[10] , \Level1Out170[5] , \Level2Out96[25] , 
        \ScanLink173[11] , \Level2Out102[9] , \ScanLink150[20] , 
        \ScanLink238[23] , \Level2Out58[9] , \Level2Out78[10] , 
        \ScanLink26[13] , \ScanLink33[27] , \ScanLink46[17] , 
        \Level16Out240[1] , \ScanLink181[8] , \Level1Out213[3] , 
        \ScanLink53[23] , \Level1Out31[9] , \ScanLink70[12] , \ScanLink70[3] , 
        \Level4Load84[0] , \Level1Out173[6] , \ScanLink188[10] , 
        \Level2Out18[14] , \Level2Out224[27] , \Level4Out216[20] , 
        \ScanLink9[27] , \ScanLink10[25] , \ScanLink17[4] , \Level1Out84[8] , 
        \ScanLink173[22] , \Level1Out198[11] , \Level4Out240[21] , 
        \Level1Out228[22] , \Level1Out248[26] , \Level8Out48[4] , 
        \Level2Out194[14] , \Level2Out212[22] , \Level2Out244[23] , 
        \Level4Out220[25] , \Level2Out206[8] , \ScanLink106[12] , 
        \ScanLink125[23] , \ScanLink129[6] , \ScanLink150[13] , 
        \Level2Out96[16] , \ScanLink130[17] , \ScanLink145[27] , 
        \Level2Out2[3] , \Level1Out24[31] , \Level1Out24[28] , 
        \Level1Out89[31] , \Level1Out89[28] , \Level1Out99[7] , 
        \ScanLink113[26] , \ScanLink166[16] , \Level1Out114[1] , 
        \ScanLink249[3] , \Level1Out155[26] , \Level8Out144[30] , 
        \Level2Out22[1] , \Level4Out128[11] , \Level1Out103[27] , 
        \Level1Out120[16] , \Level8Out112[28] , \Level1Out176[17] , 
        \Level8Out144[29] , \Level8Out112[31] , \ScanLink134[9] , 
        \Level1Out163[23] , \Level1Out116[13] , \Level4Out68[23] , 
        \Level1Out135[22] , \Level1Out140[12] , \Level1Out228[11] , 
        \Level2Out212[11] , \Level4Out148[15] , \Level4Out220[16] , 
        \Level64Out192[29] , \Level2Out194[27] , \Level2Out218[4] , 
        \Level64Out192[30] , \Level2Out244[10] , \Level1Out51[18] , 
        \Level1Out72[30] , \Level2Out224[14] , \Level4Out216[13] , 
        \ScanLink26[20] , \Level1Out72[29] , \Level1Out248[15] , 
        \Level2Out178[1] , \Level1Out198[22] , \Level4Out240[12] , 
        \Level1Out48[2] , \ScanLink53[10] , \Level16Out224[5] , 
        \ScanLink70[21] , \ScanLink188[23] , \Level2Out18[27] , 
        \Level2Out78[23] , \Level4Out180[8] , \Level16Out144[0] , 
        \ScanLink14[7] , \ScanLink33[14] , \ScanLink65[15] , \Level1Out117[2] , 
        \ScanLink238[10] , \Level1Out34[4] , \ScanLink46[24] , \ScanLink68[1] , 
        \ScanLink156[3] , \ScanLink95[18] , \ScanLink236[6] , 
        \Level1Out19[21] , \Level1Out82[24] , \Level1Out97[10] , 
        \ScanLink184[5] , \Level2Out104[7] , \Level4Out136[30] , 
        \Level4Out136[29] , \Level4Out160[28] , \Level4Out160[31] , 
        \ScanLink187[6] , \Level8Out232[12] , \Level1Out0[28] , 
        \Level1Out175[8] , \Level1Out215[18] , \Level1Out236[30] , 
        \Level1Load212[0] , \ScanLink6[20] , \Level1Load6[0] , \Level1Out6[9] , 
        \Level1Out79[25] , \Level1Out236[29] , \Level1Out243[19] , 
        \ScanLink9[14] , \Level1Out37[7] , \ScanLink155[0] , \ScanLink205[19] , 
        \Level1Out208[2] , \ScanLink226[31] , \ScanLink226[28] , 
        \ScanLink253[18] , \ScanLink38[18] , \Level1Out168[7] , 
        \ScanLink235[5] , \Level4Out76[6] , \Level1Out82[17] , 
        \Level32Out160[8] , \Level1Out82[6] , \Level2Out200[6] , 
        \Level2Out164[19] , \Level4Out76[31] , \Level1Out50[0] , 
        \Level1Out97[23] , \Level1Out108[18] , \Level2Out160[3] , 
        \Level4Out20[29] , \Level4Out76[28] , \ScanLink118[19] , 
        \ScanLink132[7] , \Level2Out132[18] , \Level4Out20[30] , 
        \ScanLink196[28] , \ScanLink252[2] , \ScanLink12[9] , \Level1Out53[3] , 
        \Level1Load71[0] , \Level1Out79[16] , \Level1Out81[5] , 
        \ScanLink131[4] , \ScanLink196[31] , \Level4Load144[0] , 
        \ScanLink251[1] , \Level2Out30[30] , \Level2Out30[29] , 
        \Level2Out66[31] , \Level4Out12[2] , \Level2Out66[28] , 
        \Level32Load64[0] , \Level1Out186[29] , \Level1Out15[6] , 
        \Level1Out16[26] , \Level1Out19[12] , \Level1Out157[9] , 
        \Level1Out186[30] , \Level8Out232[21] , \Level4Out208[18] , 
        \Level64Out64[17] , \Level1Out198[0] , \Level8Out80[12] , 
        \Level1Out35[17] , \Level1Out63[16] , \ScanLink177[1] , 
        \Level8Load80[0] , \Level8Out248[25] , \Level1Out20[23] , 
        \Level1Out40[27] , \ScanLink49[3] , \Level1Out55[13] , 
        \Level4Out112[5] , \Level4Out212[18] , \Level1Out76[22] , 
        \ScanLink217[4] , \Level4Out244[19] , \Level1Out16[15] , 
        \Level1Out16[5] , \Level1Out20[10] , \Level1Out55[20] , 
        \ScanLink85[9] , \Level1Out98[17] , \Level1Out167[28] , 
        \ScanLink174[2] , \Level1Out229[0] , \Level2Out128[18] , 
        \ScanLink98[6] , \ScanLink102[19] , \Level1Out112[18] , 
        \Level1Out131[30] , \Level1Out131[29] , \Level1Out144[19] , 
        \Level8Out120[26] , \Level1Out167[31] , \ScanLink214[7] , 
        \Level8Out176[27] , \Level1Out149[5] , \ScanLink177[29] , 
        \Level2Out246[3] , \ScanLink121[31] , \ScanLink121[28] , 
        \ScanLink154[18] , \ScanLink177[30] , \Level8Out72[7] , 
        \Level2Out126[6] , \ScanLink209[8] , \Level1Out63[25] , 
        \Level1Out71[2] , \Level1Out76[11] , \ScanLink113[5] , 
        \Level4Out216[4] , \Level8Out184[8] , \Level2Out240[31] , 
        \Level1Out35[24] , \Level1Out40[14] , \Level2Out216[29] , 
        \Level4Out176[1] , \Level2Out240[28] , \Level8Out248[16] , 
        \ScanLink57[28] , \Level1Load134[0] , \Level2Out18[2] , 
        \Level2Out216[30] , \ScanLink249[18] , \Level8Out80[21] , 
        \Level1Out253[8] , \Level1Out4[10] , \ScanLink6[13] , \ScanLink22[18] , 
        \ScanLink30[8] , \Level64Out64[24] , \ScanLink57[31] , 
        \Level1Out72[1] , \ScanLink74[19] , \ScanLink110[6] , 
        \Level2Out142[2] , \Level2Out222[7] , \Level4Out208[8] , 
        \Level8Out16[3] , \Level64Out192[9] , \Level8Out120[15] , 
        \Level8Out176[14] , \Level1Out98[24] , \Level2Out190[4] , 
        \Level1Out197[16] , \Level1Out211[20] , \Level1Out232[11] , 
        \Level2Out208[11] , \Level1Out13[8] , \ScanLink52[2] , 
        \Level1Out68[29] , \Level1Out182[22] , \Level1Out227[25] , 
        \Level1Out231[2] , \Level1Out247[21] , \Level16Out96[29] , 
        \Level1Out68[30] , \Level1Out204[14] , \Level1Out252[15] , 
        \Level16Out96[30] , \Level1Out151[7] , \ScanLink192[23] , 
        \ScanLink237[24] , \ScanLink242[14] , \ScanLink29[27] , 
        \ScanLink29[14] , \ScanLink49[10] , \ScanLink214[15] , 
        \Level32Out224[2] , \ScanLink201[21] , \Level2Out54[26] , 
        \Level2Out34[22] , \ScanLink51[1] , \ScanLink80[4] , \ScanLink83[7] , 
        \ScanLink84[14] , \ScanLink91[20] , \ScanLink169[22] , 
        \Level1Out183[1] , \ScanLink187[17] , \Level4Out52[9] , 
        \ScanLink222[10] , \Level2Out62[23] , \Level2Out64[4] , 
        \Level64Out0[13] , \ScanLink109[26] , \Level1Out180[2] , 
        \ScanLink212[9] , \Level1Out93[31] , \Level1Out119[27] , 
        \Level2Out156[17] , \Level4Out164[10] , \Level1Out152[4] , 
        \Level1Out232[1] , \Level2Out100[16] , \Level4Out12[27] , 
        \Level4Out44[26] , \Level2Out160[12] , \Level4Out132[11] , 
        \Level4Out24[22] , \Level4Out152[15] , \Level1Out93[28] , 
        \Level2Out120[8] , \Level2Out136[13] , \Level4Out72[23] , 
        \Level1Out179[23] , \Level4Out104[14] , \ScanLink187[24] , 
        \ScanLink201[12] , \Level1Out248[9] , \Level2Out34[11] , 
        \Level2Out62[10] , \ScanLink222[23] , \ScanLink242[27] , 
        \Level1Out0[21] , \Level1Out0[12] , \Level1Out4[23] , 
        \Level1Load48[0] , \ScanLink192[10] , \ScanLink237[17] , 
        \Level2Out54[15] , \ScanLink49[23] , \ScanLink214[26] , 
        \ScanLink108[4] , \Level1Out182[11] , \Level1Out227[16] , 
        \Level1Out252[26] , \Level1Out255[6] , \Level1Out135[3] , 
        \Level1Out204[27] , \Level1Out211[13] , \Level32Out96[8] , 
        \ScanLink11[3] , \ScanLink35[5] , \ScanLink36[6] , \Level1Out197[25] , 
        \Level1Out247[12] , \Level2Out188[6] , \Level2Out208[22] , 
        \Level1Out232[22] , \Level1Out69[0] , \Level2Out224[9] , 
        \Level4Out24[11] , \Level1Out119[14] , \Level1Out179[10] , 
        \Level2Out160[21] , \Level4Out152[26] , \Level4Out104[27] , 
        \Level2Out136[20] , \Level4Out12[14] , \Level4Out72[10] , 
        \Level4Out164[23] , \ScanLink84[27] , \Level1Out136[0] , 
        \Level2Load24[0] , \Level2Out100[25] , \Level2Out156[24] , 
        \Level4Out132[22] , \Level4Out28[1] , \Level4Out44[15] , 
        \ScanLink91[13] , \ScanLink109[15] , \ScanLink116[8] , 
        \ScanLink169[11] , \Level64Out0[20] , \Level1Out108[11] , 
        \Level1Out112[6] , \Level2Out164[10] , \Level4Out156[17] , 
        \Level4Out20[20] , \Level4Out76[21] , \Level2Out132[11] , 
        \ScanLink12[0] , \ScanLink38[22] , \Level1Out50[9] , \ScanLink80[16] , 
        \Level1Out168[15] , \Level2Out152[15] , \Level4Out100[16] , 
        \Level4Out16[25] , \Level4Out160[12] , \Level2Out4[4] , 
        \Level2Out104[14] , \Level4Out40[24] , \Level4Out136[13] , 
        \ScanLink95[22] , \ScanLink118[10] , \ScanLink178[14] , 
        \Level2Out24[6] , \Level2Out88[14] , \ScanLink58[26] , 
        \ScanLink183[15] , \ScanLink205[23] , \Level2Out30[20] , 
        \Level8Out0[27] , \ScanLink196[21] , \ScanLink226[12] , 
        \ScanLink233[26] , \ScanLink251[8] , \ScanLink253[22] , 
        \Level2Out66[21] , \ScanLink210[17] , \ScanLink246[16] , 
        \Level2Out50[24] , \Level1Out186[20] , \Level1Out223[27] , 
        \Level8Out232[31] , \Level1Out111[5] , \Level1Out200[16] , 
        \Level8Out232[28] , \Level1Out193[14] , \Level1Out215[22] , 
        \Level4Out208[11] , \Level1Out236[13] , \Level1Out243[23] , 
        \Level1Out5[3] , \ScanLink68[8] , \Level128Out128[5] , 
        \ScanLink80[25] , \ScanLink95[11] , \ScanLink118[23] , 
        \Level2Out40[2] , \Level2Out88[27] , \ScanLink178[27] , 
        \Level1Out29[2] , \ScanLink75[7] , \Level1Out168[26] , 
        \ScanLink199[3] , \Level4Out16[16] , \Level1Out176[2] , 
        \Level2Out104[27] , \Level2Out152[26] , \Level4Out160[21] , 
        \Level4Out68[3] , \Level4Out136[20] , \Level4Out40[17] , 
        \Level2Out92[4] , \Level4Out20[13] , \Level1Out97[19] , 
        \Level2Out164[23] , \Level4Out156[24] , \Level4Out100[25] , 
        \Level1Out108[22] , \Level1Out216[7] , \Level2Out132[22] , 
        \Level4Out76[12] , \Level1Out175[1] , \Level1Out215[11] , 
        \ScanLink228[3] , \Level1Out243[10] , \Level1Out1[18] , 
        \ScanLink2[22] , \Level1Out6[0] , \Level1Out19[31] , \Level1Out19[28] , 
        \ScanLink76[4] , \Level1Out193[27] , \Level1Out236[20] , 
        \ScanLink148[6] , \Level1Out186[13] , \Level1Out215[4] , 
        \Level1Out223[14] , \Level4Out208[22] , \ScanLink38[11] , 
        \ScanLink196[12] , \Level1Out200[25] , \ScanLink233[15] , 
        \ScanLink246[25] , \Level2Out50[17] , \ScanLink210[24] , 
        \Level32Out160[1] , \ScanLink58[15] , \Level1Out84[1] , 
        \Level1Out114[8] , \ScanLink155[9] , \ScanLink183[26] , 
        \ScanLink205[10] , \Level2Out30[13] , \ScanLink253[11] , 
        \Level2Out66[12] , \Level8Out0[14] , \ScanLink226[21] , 
        \Level2Out166[4] , \Level2Out206[1] , \Level1Out89[21] , 
        \Level8Out32[5] , \Level1Out109[7] , \ScanLink254[5] , \ScanLink2[11] , 
        \Level1Out12[24] , \Level1Out24[21] , \Level1Out56[7] , 
        \Level2Out22[8] , \Level4Out128[18] , \Level8Out112[21] , 
        \ScanLink134[0] , \Level8Out144[20] , \Level16Load112[0] , 
        \Level4Out152[7] , \Level1Out51[11] , \Level1Out72[20] , 
        \Level2Out178[8] , \Level32Out96[27] , \Level2Out212[18] , 
        \Level64Out192[20] , \ScanLink26[30] , \ScanLink26[29] , 
        \Level1Out31[15] , \Level1Out67[14] , \ScanLink137[3] , 
        \Level4Out232[2] , \Level1Out228[18] , \Level4Out0[2] , 
        \Level1Out44[25] , \Level1Out55[4] , \Level2Out244[19] , 
        \ScanLink238[19] , \Level4Out180[1] , \Level16Out144[9] , 
        \ScanLink53[19] , \ScanLink70[31] , \ScanLink70[28] , \Level1Out87[2] , 
        \Level8Out112[12] , \ScanLink8[24] , \Level1Out8[6] , 
        \Level1Load10[0] , \Level1Out32[3] , \Level1Out89[12] , 
        \Level1Out116[29] , \ScanLink230[1] , \Level8Out144[13] , 
        \Level4Out68[19] , \Level1Out116[30] , \Level1Out135[18] , 
        \Level1Out140[31] , \Level1Out163[19] , \ScanLink150[4] , 
        \Level1Out140[28] , \ScanLink106[31] , \ScanLink106[28] , 
        \ScanLink125[19] , \ScanLink150[30] , \ScanLink173[18] , 
        \Level2Out102[0] , \Level1Out12[17] , \Level1Out67[27] , 
        \ScanLink73[9] , \ScanLink150[29] , \ScanLink181[1] , \ScanLink182[2] , 
        \Level1Out210[9] , \Level8Out56[1] , \ScanLink188[19] , 
        \Level2Out58[0] , \Level2Out78[19] , \Level16Out240[8] , 
        \Level64Out192[13] , \Level1Out18[22] , \Level1Out24[12] , 
        \Level1Out31[26] , \Level1Out44[16] , \ScanLink233[2] , 
        \Level4Out136[3] , \Level1Out51[22] , \Level4Out240[31] , 
        \Level4Out216[29] , \Level32Out96[14] , \Level1Out27[4] , 
        \Level1Out31[0] , \Level1Out72[13] , \Level1Out198[18] , 
        \Level4Out240[28] , \ScanLink153[7] , \Level4Out216[30] , 
        \Level1Out178[4] , \ScanLink197[18] , \ScanLink225[6] , 
        \Level4Out120[7] , \Level2Out12[28] , \Level2Out44[30] , 
        \Level2Load210[0] , \Level1Out78[26] , \ScanLink145[3] , 
        \Level1Out218[1] , \Level2Out44[29] , \Level4Out240[2] , 
        \Level2Out12[31] , \ScanLink238[9] , \Level64Out64[4] , 
        \Level1Out83[27] , \Level1Out166[8] , \Level1Out187[19] , 
        \ScanLink197[5] , \Level2Out0[13] , \Level1Load201[0] , 
        \Level2Out114[4] , \Level1Out96[13] , \Level1Out109[28] , 
        \Level16Out48[0] , \ScanLink194[6] , \Level2Out146[18] , 
        \Level8Out40[5] , \Level1Out18[11] , \Level1Out24[7] , 
        \Level1Out39[8] , \Level2Out110[19] , \ScanLink78[2] , 
        \Level1Out109[31] , \ScanLink119[29] , \Level16Out128[5] , 
        \ScanLink226[5] , \Level8Out56[26] , \ScanLink119[30] , 
        \ScanLink146[0] , \ScanLink189[9] , \Level16Load160[0] , 
        \Level2Out50[8] , \Level2Out0[20] , \Level4Out196[5] , 
        \Level1Out78[15] , \Level1Out214[31] , \Level1Out237[19] , 
        \ScanLink8[17] , \ScanLink39[31] , \ScanLink39[28] , \Level1Out91[6] , 
        \Level1Out214[28] , \Level1Out242[29] , \Level1Out242[30] , 
        \ScanLink121[7] , \ScanLink204[30] , \Level4Out144[3] , 
        \ScanLink204[29] , \ScanLink227[18] , \ScanLink241[2] , 
        \ScanLink252[28] , \ScanLink252[31] , \Level4Out224[6] , 
        \Level16Out32[8] , \Level1Out43[0] , \Level1Out40[3] , 
        \ScanLink242[1] , \Level4Out188[9] , \Level1Load62[0] , 
        \ScanLink94[31] , \ScanLink94[28] , \ScanLink122[4] , 
        \Level8Out56[15] , \Level1Out96[20] , \Level2Out170[0] , 
        \Level1Out50[31] , \Level1Out83[14] , \Level1Out92[5] , 
        \Level2Out210[5] , \Level8Out24[1] , \ScanLink223[8] , 
        \Level1Out229[21] , \Level2Out230[10] , \Level4Out184[21] , 
        \Level1Out73[19] , \Level1Out199[12] , \ScanLink11[26] , 
        \ScanLink11[15] , \Level1Out25[18] , \Level1Out50[28] , 
        \Level1Out249[25] , \Level2Out206[15] , \Level4Out92[12] , 
        \Level2Out180[23] , \Level2Out250[14] , \ScanLink27[10] , 
        \ScanLink52[20] , \ScanLink71[11] , \Level1Out163[5] , 
        \ScanLink189[13] , \ScanLink32[24] , \ScanLink47[14] , \ScanLink60[0] , 
        \Level1Out203[0] , \ScanLink64[25] , \ScanLink239[20] , 
        \Level1Out22[9] , \ScanLink63[3] , \ScanLink124[13] , 
        \Level4Load248[0] , \Level1Out102[17] , \ScanLink107[22] , 
        \ScanLink151[23] , \ScanLink112[16] , \Level1Out160[6] , 
        \ScanLink172[12] , \ScanLink131[27] , \ScanLink167[26] , 
        \Level2Out82[12] , \Level2Out84[0] , \Level16Out0[19] , 
        \ScanLink144[17] , \ScanLink192[8] , \Level1Out200[3] , 
        \Level1Out121[26] , \Level1Out177[27] , \Level2Out138[17] , 
        \Level1Out134[12] , \Level1Out154[16] , \Level16Out224[21] , 
        \Level2Out56[6] , \ScanLink32[17] , \Level1Out88[18] , 
        \Level1Out117[23] , \Level1Out141[22] , \Level1Out162[13] , 
        \Level2Out158[13] , \Level32Out224[14] , \ScanLink47[27] , 
        \ScanLink27[23] , \Level1Out58[1] , \ScanLink64[16] , 
        \Level1Out107[1] , \ScanLink239[13] , \ScanLink71[22] , 
        \Level1Out97[8] , \ScanLink189[20] , \ScanLink52[13] , 
        \Level1Out199[21] , \Level1Out249[16] , \Level2Out206[26] , 
        \Level2Out168[2] , \Level4Out92[21] , \Level1Out0[3] , \ScanLink0[7] , 
        \ScanLink3[31] , \Level1Out117[10] , \ScanLink127[9] , 
        \Level2Out180[10] , \Level2Out208[7] , \Level2Out250[27] , 
        \Level2Out230[23] , \Level4Out184[12] , \Level1Out134[21] , 
        \Level1Out141[11] , \Level1Out229[12] , \Level1Out162[20] , 
        \Level2Out158[20] , \Level32Out224[27] , \ScanLink3[28] , 
        \Level1Out102[24] , \Level1Out177[14] , \Level2Out138[24] , 
        \Level1Out5[30] , \Level1Out5[29] , \ScanLink6[9] , \ScanLink7[19] , 
        \Level1Out89[4] , \Level1Out154[25] , \Level2Out32[2] , 
        \Level16Out224[12] , \Level1Out104[2] , \ScanLink112[25] , 
        \Level1Out121[15] , \ScanLink167[15] , \Level2Out82[21] , 
        \Level1Out106[15] , \ScanLink107[11] , \ScanLink124[20] , 
        \ScanLink131[14] , \ScanLink144[24] , \ScanLink139[5] , 
        \ScanLink151[10] , \ScanLink172[21] , \Level1Out113[21] , 
        \Level1Out130[10] , \Level2Out16[4] , \Level16Out240[27] , 
        \Level1Out145[20] , \Level1Out166[11] , \Level1Out125[24] , 
        \Level1Out173[25] , \ScanLink15[17] , \ScanLink23[1] , 
        \ScanLink116[14] , \Level1Out150[14] , \Level2Out86[10] , 
        \ScanLink120[11] , \ScanLink135[25] , \ScanLink163[24] , 
        \Level2Load248[0] , \ScanLink140[15] , \Level1Out240[1] , 
        \Level2Out152[8] , \ScanLink36[26] , \ScanLink43[16] , 
        \ScanLink103[20] , \ScanLink155[21] , \Level1Out120[4] , 
        \ScanLink176[10] , \Level1Out243[2] , \ScanLink60[27] , 
        \ScanLink198[25] , \ScanLink248[12] , \ScanLink20[2] , 
        \ScanLink23[12] , \ScanLink56[22] , \ScanLink75[13] , 
        \Level1Out123[7] , \ScanLink228[16] , \Level64Out0[3] , 
        \Level2Out68[25] , \Level1Out61[8] , \Level1Out238[17] , 
        \Level2Out184[21] , \Level2Out202[17] , \Level4Out96[10] , 
        \Level2Out254[16] , \Level32Out128[11] , \ScanLink103[13] , 
        \ScanLink120[22] , \ScanLink155[12] , \Level1Out188[24] , 
        \Level2Out234[12] , \Level4Out20[9] , \Level4Out180[23] , 
        \Level16Out128[24] , \Level1Out224[5] , \ScanLink176[23] , 
        \ScanLink179[7] , \ScanLink163[17] , \ScanLink15[24] , 
        \Level1Out18[3] , \Level1Out21[30] , \ScanLink47[5] , 
        \ScanLink116[27] , \ScanLink219[2] , \Level2Out86[23] , 
        \ScanLink135[16] , \ScanLink140[26] , \Level1Out144[0] , 
        \Level2Load56[0] , \ScanLink95[3] , \Level1Out106[26] , 
        \Level1Out173[16] , \Level1Out113[12] , \Level1Out125[17] , 
        \Level1Out150[27] , \ScanLink164[8] , \Level2Out72[0] , 
        \Level1Out130[23] , \Level1Out145[13] , \Level4Out88[7] , 
        \Level1Out196[6] , \Level1Out166[22] , \Level16Out240[14] , 
        \Level1Out188[17] , \Level2Out234[21] , \Level2Out248[5] , 
        \Level4Out180[10] , \Level16Out128[17] , \Level2Out202[24] , 
        \Level1Out21[29] , \ScanLink59[9] , \Level1Out238[24] , 
        \Level2Out128[0] , \Level4Out96[23] , \Level1Out77[28] , 
        \ScanLink96[0] , \Level32Out128[22] , \Level1Out54[19] , 
        \Level1Out77[31] , \Level2Out184[12] , \Level2Out254[25] , 
        \Level1Out195[5] , \Level2Out68[16] , \ScanLink23[21] , 
        \ScanLink75[20] , \ScanLink228[25] , \ScanLink36[15] , 
        \ScanLink56[11] , \Level1Out227[6] , \ScanLink43[25] , \ScanLink44[6] , 
        \ScanLink248[21] , \ScanLink38[0] , \ScanLink60[14] , 
        \Level1Out147[3] , \ScanLink198[16] , \Level1Out64[5] , 
        \ScanLink106[2] , \Level8Out32[20] , \Level16Out208[2] , 
        \Level8Out64[21] , \ScanLink90[19] , \Level1Load94[0] , 
        \Level2Out186[0] , \Level1Out69[10] , \Level1Out87[25] , 
        \Level1Out92[11] , \Level2Out234[3] , \Level2Out4[11] , 
        \Level2Out154[6] , \Level8Out192[14] , \Level1Out246[18] , 
        \Level1Out233[28] , \ScanLink48[30] , \ScanLink48[29] , 
        \Level1Out67[6] , \Level1Out125[9] , \Level1Out210[19] , 
        \Level1Out233[31] , \ScanLink223[29] , \ScanLink256[19] , 
        \ScanLink105[1] , \ScanLink223[30] , \Level4Out200[0] , 
        \ScanLink200[18] , \Level1Out138[6] , \Level4Out160[5] , 
        \Level1Out87[16] , \Level2Out250[7] , \Level8Out64[3] , 
        \Level1Out92[22] , \Level1Out178[29] , \Level2Out130[2] , 
        \Level2Out142[29] , \Level2Out114[31] , \Level2Out142[30] , 
        \ScanLink3[4] , \Level1Load146[0] , \ScanLink161[5] , \ScanLink162[6] , 
        \ScanLink168[31] , \ScanLink168[28] , \Level1Out178[30] , 
        \Level2Out114[28] , \Level1Out190[8] , \ScanLink202[3] , 
        \Level2Out98[31] , \Level8Out32[13] , \Level2Out98[28] , 
        \Level8Out64[12] , \ScanLink193[30] , \ScanLink193[29] , 
        \ScanLink201[0] , \Level2Out16[19] , \Level4Out104[1] , 
        \Level1Out221[8] , \Level2Out40[18] , \ScanLink9[23] , 
        \Level1Load15[0] , \Level1Out37[3] , \ScanLink42[8] , 
        \Level1Out69[23] , \Level1Out183[31] , \Level8Out192[27] , 
        \Level32Out160[31] , \Level4Out88[31] , \Level1Out183[28] , 
        \Level32Out160[28] , \Level1Out168[3] , \ScanLink210[30] , 
        \ScanLink210[29] , \ScanLink246[31] , \Level2Out4[22] , 
        \Level4Out88[28] , \ScanLink246[28] , \Level4Out76[2] , 
        \ScanLink233[18] , \ScanLink235[1] , \Level4Load120[0] , 
        \Level8Out0[19] , \ScanLink58[18] , \ScanLink155[4] , 
        \Level1Out208[6] , \Level1Out19[25] , \ScanLink76[9] , 
        \Level1Out79[21] , \Level1Out200[28] , \Level8Out232[16] , 
        \Level1Out82[20] , \ScanLink187[2] , \Level1Out215[9] , 
        \Level1Out200[31] , \Level1Out223[19] , \Level1Out97[14] , 
        \Level2Out104[3] , \Level4Out100[28] , \ScanLink184[1] , 
        \Level4Out156[30] , \ScanLink9[10] , \Level1Out19[16] , 
        \Level1Out34[0] , \ScanLink68[5] , \ScanLink236[2] , \Level2Out92[9] , 
        \Level4Out100[31] , \Level4Out156[29] , \ScanLink80[31] , 
        \Level128Out128[8] , \ScanLink80[28] , \ScanLink156[7] , 
        \Level1Out111[8] , \Level8Out232[25] , \Level1Out50[4] , 
        \Level1Out53[7] , \Level1Out79[12] , \Level1Out81[1] , 
        \Level1Out193[19] , \ScanLink131[0] , \ScanLink183[18] , 
        \Level4Out12[6] , \ScanLink251[5] , \Level2Out50[29] , 
        \ScanLink178[19] , \ScanLink252[6] , \Level2Out50[30] , 
        \Level2Out88[19] , \Level1Out97[27] , \ScanLink132[3] , 
        \Level2Out160[7] , \Level1Out82[13] , \Level1Out82[2] , 
        \Level2Out200[2] , \Level4Out40[29] , \Level1Out168[18] , 
        \Level2Out104[19] , \Level4Out16[31] , \Level2Out152[18] , 
        \Level4Out40[30] , \Level4Out16[28] , \Level1Out198[15] , 
        \Level1Out228[26] , \Level2Out4[9] , \Level2Out194[10] , 
        \Level2Out244[27] , \Level2Out212[26] , \Level4Out220[21] , 
        \Level4Out240[25] , \Level1Out1[26] , \Level1Out1[15] , \ScanLink3[9] , 
        \Level1Out3[0] , \ScanLink10[12] , \ScanLink26[17] , \ScanLink53[27] , 
        \ScanLink70[16] , \Level1Load169[0] , \Level1Out248[22] , 
        \Level8Out48[0] , \Level32Out96[19] , \Level2Out224[23] , 
        \Level4Out216[24] , \Level1Out173[2] , \ScanLink188[14] , 
        \Level2Out18[10] , \Level16Load208[0] , \ScanLink33[23] , 
        \ScanLink46[13] , \ScanLink70[7] , \Level16Out240[5] , 
        \Level1Out213[7] , \ScanLink65[22] , \ScanLink238[27] , 
        \Level2Out78[14] , \ScanLink73[4] , \ScanLink125[14] , 
        \Level1Out103[10] , \ScanLink106[25] , \ScanLink150[24] , 
        \Level2Load178[0] , \Level2Out96[21] , \Level4Out128[2] , 
        \ScanLink113[11] , \Level1Out170[1] , \ScanLink173[15] , 
        \ScanLink130[20] , \ScanLink166[21] , \Level2Out94[7] , 
        \ScanLink145[10] , \Level4Out248[7] , \Level1Out210[4] , 
        \Level1Out116[24] , \Level1Out120[21] , \Level1Out176[20] , 
        \Level1Out135[15] , \Level1Out155[11] , \Level2Out46[1] , 
        \Level4Out128[26] , \Level1Out140[25] , \Level4Out148[22] , 
        \Level4Out68[14] , \ScanLink5[7] , \ScanLink8[2] , \ScanLink10[21] , 
        \ScanLink14[3] , \ScanLink33[10] , \ScanLink150[9] , 
        \Level1Out163[14] , \ScanLink46[20] , \Level2Out78[27] , 
        \Level16Out144[4] , \Level1Out12[30] , \ScanLink26[24] , 
        \Level1Out48[6] , \ScanLink65[11] , \Level1Out117[6] , 
        \ScanLink238[14] , \ScanLink70[25] , \ScanLink188[27] , 
        \Level2Out18[23] , \ScanLink53[14] , \Level16Out224[1] , 
        \Level1Out198[26] , \Level1Out248[11] , \Level2Out178[5] , 
        \Level4Out240[16] , \Level2Out218[0] , \Level2Out224[10] , 
        \Level4Out216[17] , \Level1Out12[29] , \Level1Out31[18] , 
        \Level2Out194[23] , \Level1Out44[28] , \Level1Out55[9] , 
        \Level2Out244[14] , \ScanLink14[10] , \ScanLink17[0] , 
        \Level1Out44[31] , \Level2Out212[15] , \Level4Out220[12] , 
        \Level1Out67[19] , \Level1Out228[15] , \Level1Out99[3] , 
        \Level1Out103[23] , \Level1Out116[17] , \Level1Out135[26] , 
        \Level1Out140[16] , \Level1Out163[27] , \ScanLink254[8] , 
        \Level4Out148[11] , \Level4Out68[27] , \Level1Out176[13] , 
        \Level1Out155[22] , \Level2Out22[5] , \Level4Out128[15] , 
        \ScanLink113[22] , \Level1Out120[12] , \ScanLink166[12] , 
        \ScanLink249[7] , \Level1Out114[5] , \ScanLink130[13] , 
        \ScanLink145[23] , \Level2Out166[9] , \ScanLink33[6] , 
        \Level1Out98[30] , \Level1Out98[29] , \ScanLink106[16] , 
        \ScanLink125[27] , \ScanLink150[17] , \Level8Out32[8] , 
        \ScanLink129[2] , \Level2Out2[7] , \ScanLink173[26] , 
        \Level2Out96[12] , \Level1Out107[12] , \Level1Out112[26] , 
        \Level1Out131[17] , \Level1Out144[27] , \Level8Out176[19] , 
        \Level1Out167[16] , \Level2Out128[26] , \Level8Out120[18] , 
        \Level2Out148[22] , \Level2Out190[9] , \Level1Out172[22] , 
        \Level1Out124[23] , \ScanLink117[13] , \Level1Out151[13] , 
        \ScanLink121[16] , \ScanLink134[22] , \ScanLink162[23] , 
        \ScanLink141[12] , \Level4Out208[5] , \Level1Out250[6] , 
        \ScanLink37[21] , \ScanLink42[11] , \ScanLink102[27] , 
        \ScanLink154[26] , \Level4Out168[0] , \Level1Out130[3] , 
        \Level2Out92[23] , \Level64Out192[4] , \ScanLink177[17] , 
        \Level1Out253[5] , \ScanLink61[20] , \ScanLink199[22] , 
        \ScanLink249[15] , \Level1Out16[18] , \ScanLink22[15] , 
        \ScanLink57[25] , \ScanLink74[14] , \Level1Out133[0] , 
        \ScanLink229[11] , \Level16Out160[2] , \Level64Out64[30] , 
        \ScanLink30[5] , \Level1Out35[30] , \Level1Out35[29] , 
        \Level1Out40[19] , \Level1Out63[31] , \ScanLink113[8] , 
        \Level1Out239[10] , \Level4Out216[9] , \Level64Out64[29] , 
        \Level4Out244[27] , \Level8Out184[5] , \Level2Out220[21] , 
        \Level4Out212[26] , \Level2Out240[25] , \Level1Out63[28] , 
        \Level2Out190[12] , \Level1Out189[23] , \Level2Out216[24] , 
        \Level4Load16[0] , \Level4Out224[23] , \Level1Out16[8] , 
        \ScanLink57[2] , \ScanLink102[14] , \ScanLink121[25] , 
        \ScanLink154[15] , \ScanLink169[0] , \Level1Out234[2] , 
        \ScanLink177[24] , \ScanLink117[20] , \ScanLink162[10] , 
        \Level2Out92[10] , \ScanLink134[11] , \ScanLink141[21] , 
        \Level1Out154[7] , \ScanLink209[5] , \Level1Out107[21] , 
        \Level1Out172[11] , \Level1Out124[10] , \Level1Out151[20] , 
        \Level2Out148[11] , \Level2Out62[7] , \ScanLink85[4] , 
        \Level1Out112[15] , \Level1Out131[24] , \Level1Out144[14] , 
        \Level1Out149[8] , \Level1Out186[1] , \Level1Out167[25] , 
        \Level2Out128[15] , \ScanLink86[7] , \Level1Out189[10] , 
        \Level2Out190[21] , \Level8Out248[28] , \Level2Out216[17] , 
        \Level2Out240[16] , \Level4Out224[10] , \Level8Out248[31] , 
        \Level16Out64[3] , \Level1Out239[23] , \Level2Out138[7] , 
        \Level4Out244[14] , \Level2Out220[12] , \Level4Out112[8] , 
        \Level4Out212[15] , \Level1Out10[6] , \ScanLink14[23] , 
        \ScanLink22[26] , \ScanLink74[27] , \Level1Out185[2] , 
        \ScanLink217[9] , \ScanLink229[22] , \ScanLink37[12] , 
        \ScanLink57[16] , \Level1Out237[1] , \ScanLink42[22] , \ScanLink54[1] , 
        \ScanLink249[26] , \ScanLink28[7] , \ScanLink61[13] , 
        \Level1Out157[4] , \ScanLink199[11] , \Level1Out74[2] , 
        \ScanLink116[5] , \ScanLink109[18] , \Level2Out196[7] , 
        \ScanLink35[8] , \Level1Out86[22] , \Level1Out93[16] , 
        \Level1Load131[0] , \Level2Out224[4] , \Level8Out168[12] , 
        \Level2Out100[28] , \Level2Out156[30] , \Level4Out44[18] , 
        \Level2Out100[31] , \Level2Out144[1] , \Level4Out12[19] , 
        \Level2Out156[29] , \Level1Out68[17] , \ScanLink108[9] , 
        \Level1Out119[19] , \Level16Out96[17] , \Level1Out77[1] , 
        \ScanLink187[29] , \Level1Out197[31] , \Level1Out197[28] , 
        \Level8Out200[11] , \Level32Out96[5] , \Level1Out86[11] , 
        \ScanLink115[6] , \ScanLink187[30] , \Level1Out248[4] , 
        \Level1Out128[1] , \Level2Out54[18] , \Level2Load120[0] , 
        \Level4Out36[0] , \Level2Out240[0] , \Level1Out93[25] , 
        \Level2Out120[5] , \Level1Out152[9] , \Level4Out104[19] , 
        \Level4Out152[18] , \Level8Out168[21] , \Level2Out64[9] , 
        \Level1Out13[5] , \ScanLink84[19] , \ScanLink172[1] , \ScanLink212[4] , 
        \ScanLink171[2] , \ScanLink214[18] , \ScanLink237[30] , 
        \ScanLink237[29] , \ScanLink29[19] , \ScanLink211[7] , 
        \ScanLink242[19] , \Level4Out52[4] , \Level1Out68[24] , 
        \ScanLink80[9] , \Level1Out204[19] , \Level1Out227[31] , 
        \Level4Out80[2] , \Level8Out200[22] , \Level1Out227[28] , 
        \Level16Out96[24] , \ScanLink228[31] , \Level1Out252[18] , 
        \ScanLink228[28] , \Level1Out5[17] , \ScanLink6[4] , \ScanLink7[27] , 
        \ScanLink15[30] , \ScanLink15[29] , \Level4Out96[6] , \ScanLink43[31] , 
        \ScanLink60[19] , \Level1Out188[7] , \Level1Out17[21] , 
        \ScanLink36[18] , \ScanLink43[28] , \Level1Out21[24] , 
        \Level1Out34[10] , \Level1Out62[11] , \ScanLink167[6] , 
        \Level2Out248[8] , \Level1Out41[20] , \Level4Out44[0] , 
        \Level1Out54[14] , \Level2Out202[30] , \ScanLink59[4] , 
        \Level1Out195[8] , \ScanLink207[3] , \Level1Out238[30] , 
        \Level2Out254[28] , \Level2Load152[0] , \Level2Out202[29] , 
        \Level1Out77[25] , \Level1Out238[29] , \Level2Out254[31] , 
        \ScanLink47[8] , \ScanLink88[1] , \Level1Out99[10] , 
        \Level1Load143[0] , \Level1Out159[2] , \ScanLink164[5] , 
        \Level1Out239[7] , \ScanLink204[0] , \Level16Out240[19] , 
        \Level1Out224[8] , \Level2Out136[1] , \ScanLink7[14] , 
        \Level1Out17[12] , \Level1Out21[17] , \Level1Out54[27] , 
        \Level1Out61[5] , \Level1Out62[22] , \Level1Out77[16] , 
        \Level1Load91[0] , \ScanLink103[2] , \Level1Out188[29] , 
        \Level1Out34[23] , \Level1Out41[13] , \Level16Out128[29] , 
        \Level1Out188[30] , \Level4Out20[4] , \Level16Out128[30] , 
        \Level1Out62[6] , \ScanLink100[1] , \ScanLink116[19] , 
        \ScanLink135[28] , \ScanLink198[31] , \ScanLink198[28] , 
        \Level2Out68[31] , \Level2Out68[28] , \ScanLink140[18] , 
        \ScanLink163[30] , \Level2Out232[0] , \Level1Out120[9] , 
        \ScanLink135[31] , \ScanLink163[29] , \Level2Out152[5] , 
        \Level32Out128[6] , \Level2Out16[9] , \Level1Out125[29] , 
        \Level1Out99[23] , \Level1Out106[18] , \Level1Out150[19] , 
        \Level1Out173[31] , \Level2Out180[3] , \Level1Out125[30] , 
        \Level1Out173[28] , \Level1Out196[11] , \Level1Out210[27] , 
        \Level16Out160[10] , \Level1Out233[16] , \Level1Out246[26] , 
        \ScanLink42[5] , \Level1Out183[25] , \Level1Out221[5] , 
        \Level1Out226[22] , \Level32Out160[25] , \Level1Out253[12] , 
        \Level4Out88[25] , \Level1Out5[24] , \ScanLink28[20] , 
        \ScanLink28[13] , \ScanLink48[17] , \Level1Out141[0] , 
        \Level1Out205[13] , \Level16Out112[2] , \ScanLink193[24] , 
        \ScanLink215[12] , \ScanLink236[23] , \ScanLink243[13] , 
        \Level2Out76[10] , \Level2Out20[11] , \ScanLink161[8] , 
        \ScanLink200[26] , \ScanLink41[6] , \ScanLink85[13] , \ScanLink90[27] , 
        \ScanLink90[3] , \Level2Out40[15] , \Level4Load64[0] , 
        \ScanLink168[25] , \ScanLink186[10] , \ScanLink223[17] , 
        \Level1Out193[6] , \Level2Out16[14] , \ScanLink256[27] , 
        \Level2Out74[3] , \ScanLink108[21] , \Level1Out190[5] , 
        \Level2Out98[25] , \ScanLink93[0] , \Level1Out118[20] , 
        \Level1Out142[3] , \Level1Out222[6] , \Level2Out122[20] , 
        \Level2Out174[21] , \Level2Out114[25] , \Level2Out142[24] , 
        \Level16Out208[13] , \Level1Out178[24] , \ScanLink48[24] , 
        \ScanLink186[23] , \ScanLink200[15] , \Level2Out40[26] , 
        \Level16Out16[3] , \Level8Out192[1] , \ScanLink223[24] , 
        \ScanLink256[14] , \ScanLink193[17] , \ScanLink243[20] , 
        \Level2Out16[27] , \Level2Out76[23] , \Level4Out160[8] , 
        \ScanLink215[21] , \ScanLink236[10] , \Level2Out20[22] , 
        \ScanLink118[3] , \Level1Out183[16] , \Level1Out245[1] , 
        \Level1Out253[21] , \Level4Out88[16] , \Level1Out226[11] , 
        \Level32Out160[16] , \Level1Out125[4] , \Level1Out205[20] , 
        \Level8Out192[19] , \Level1Out210[14] , \Level16Out176[6] , 
        \Level16Out160[23] , \Level1Out246[15] , \ScanLink25[2] , 
        \ScanLink26[1] , \Level1Out196[22] , \Level1Out233[25] , 
        \Level2Out198[1] , \Level1Out79[7] , \Level2Out114[16] , 
        \Level1Out87[28] , \Level1Out178[17] , \Level1Out246[2] , 
        \Level2Out142[17] , \Level16Out208[20] , \Level2Out122[13] , 
        \Level1Out118[13] , \ScanLink39[25] , \ScanLink59[21] , 
        \Level1Out64[8] , \ScanLink85[20] , \Level1Out87[31] , 
        \Level1Out126[7] , \Level2Out174[12] , \Level2Out10[7] , 
        \ScanLink81[11] , \Level1Out83[19] , \ScanLink90[14] , 
        \ScanLink108[12] , \ScanLink168[16] , \Level2Out98[16] , 
        \Level1Out102[1] , \Level1Out109[16] , \Level2Out110[27] , 
        \Level2Out146[26] , \Level1Out92[8] , \Level1Out169[12] , 
        \Level2Out126[22] , \Level2Out170[23] , \Level4Out8[7] , 
        \Level2Out210[8] , \Level4Out188[4] , \ScanLink94[25] , 
        \ScanLink119[17] , \ScanLink122[9] , \ScanLink179[13] , 
        \Level4Out8[11] , \Level8Out56[18] , \Level2Out34[1] , 
        \ScanLink182[12] , \ScanLink204[24] , \ScanLink227[15] , 
        \Level2Out12[16] , \Level2Out44[17] , \ScanLink197[26] , 
        \ScanLink252[25] , \ScanLink211[10] , \ScanLink232[21] , 
        \ScanLink247[11] , \Level2Out72[12] , \Level2Out24[13] , 
        \Level16Out32[5] , \Level1Out78[18] , \Level1Out101[2] , 
        \Level1Out187[27] , \Level1Out201[11] , \Level1Out222[20] , 
        \Level2Out218[20] , \Level4Out196[8] , \Level1Out192[13] , 
        \Level1Out214[25] , \Level1Out237[14] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink65[0] , \ScanLink81[22] , \ScanLink94[16] , 
        \Level1Out242[24] , \Level16Out128[8] , \ScanLink119[24] , 
        \ScanLink226[8] , \Level2Out50[5] , \Level1Out169[21] , 
        \ScanLink179[20] , \ScanLink189[4] , \Level4Out8[22] , 
        \Level2Out126[11] , \Level2Out114[9] , \Level1Out166[5] , 
        \Level2Out170[10] , \Level1Out39[5] , \Level2Out82[3] , 
        \Level2Out110[14] , \Level1Out109[25] , \Level2Out146[15] , 
        \Level8Out40[8] , \Level1Out165[6] , \Level1Out206[0] , 
        \Level1Out214[16] , \ScanLink238[4] , \ScanLink3[25] , 
        \Level1Out27[9] , \ScanLink39[16] , \ScanLink66[3] , 
        \Level1Out192[20] , \Level1Out237[27] , \Level1Out242[17] , 
        \ScanLink158[1] , \Level1Out187[14] , \ScanLink197[8] , 
        \Level2Out218[13] , \Level4Load92[0] , \Level1Out205[3] , 
        \Level1Out222[13] , \Level1Out178[9] , \ScanLink197[15] , 
        \Level1Out201[22] , \Level64Out64[9] , \ScanLink247[22] , 
        \Level2Out72[21] , \ScanLink232[12] , \ScanLink59[12] , 
        \ScanLink211[23] , \Level2Out24[20] , \Level2Out44[24] , 
        \ScanLink204[17] , \ScanLink252[16] , \Level1Out88[26] , 
        \Level1Out94[6] , \ScanLink112[31] , \ScanLink131[19] , 
        \ScanLink144[29] , \ScanLink182[21] , \ScanLink227[26] , 
        \Level2Out12[25] , \Level2Out176[3] , \ScanLink112[28] , 
        \ScanLink144[30] , \ScanLink167[18] , \Level2Out216[6] , 
        \Level16Out0[27] , \ScanLink139[8] , \Level8Out48[13] , 
        \Level1Out119[0] , \ScanLink244[2] , \ScanLink3[16] , 
        \Level1Out13[23] , \ScanLink19[6] , \Level1Out25[26] , 
        \Level1Out46[0] , \Level1Out89[9] , \Level1Out154[28] , 
        \Level2Out138[30] , \Level1Out121[18] , \Level1Out102[30] , 
        \Level1Out102[29] , \ScanLink124[7] , \Level1Out154[31] , 
        \Level1Out177[19] , \Level2Out138[29] , \Level16Out16[22] , 
        \Level1Out50[16] , \Level1Out73[27] , \ScanLink247[1] , 
        \Level1Out30[12] , \Level1Out66[13] , \ScanLink127[4] , 
        \Level1Out45[22] , \Level1Out45[3] , \Level4Load152[0] , 
        \Level1Load67[0] , \Level1Out97[5] , \Level1Out22[4] , 
        \Level1Out88[15] , \ScanLink220[6] , \Level16Out16[11] , 
        \Level32Out224[19] , \ScanLink140[3] , \ScanLink192[5] , 
        \Level2Out112[7] , \Level8Out48[20] , \Level16Out0[14] , 
        \ScanLink11[18] , \ScanLink32[30] , \ScanLink64[28] , 
        \Level1Out163[8] , \Level1Load204[0] , \Level2Out48[7] , 
        \Level1Out13[10] , \ScanLink32[29] , \ScanLink47[19] , 
        \ScanLink64[31] , \ScanLink191[6] , \Level1Out66[20] , 
        \Level1Out30[21] , \Level1Out45[11] , \ScanLink223[5] , 
        \Level4Out60[6] , \Level1Out50[25] , \Level2Out250[19] , 
        \Level1Out21[7] , \Level1Out25[15] , \Level1Out249[31] , 
        \Level1Out73[14] , \Level32Out0[6] , \ScanLink0[3] , \ScanLink3[0] , 
        \ScanLink26[8] , \ScanLink28[30] , \ScanLink28[29] , \Level1Out138[2] , 
        \ScanLink143[0] , \Level1Out249[28] , \Level2Out206[18] , 
        \ScanLink215[31] , \ScanLink243[29] , \Level4Out160[1] , 
        \ScanLink236[19] , \ScanLink215[28] , \ScanLink243[30] , 
        \Level4Out200[4] , \ScanLink105[5] , \Level8Out192[8] , 
        \Level1Out67[2] , \Level2Out198[8] , \ScanLink38[4] , 
        \Level1Out69[14] , \Level1Out205[30] , \Level1Out245[8] , 
        \Level1Out253[28] , \Level2Out4[15] , \Level1Out226[18] , 
        \Level1Out87[21] , \Level1Load122[0] , \Level1Out253[31] , 
        \Level1Out205[29] , \Level8Out192[10] , \Level1Out92[15] , 
        \Level2Out154[2] , \Level2Out234[7] , \Level16Out208[30] , 
        \Level16Out208[29] , \Level2Out186[4] , \Level1Out64[1] , 
        \ScanLink85[29] , \Level8Out64[25] , \Level1Out69[27] , 
        \ScanLink85[30] , \ScanLink106[6] , \Level8Out32[24] , 
        \Level16Out208[6] , \Level2Out4[26] , \Level8Out192[23] , 
        \ScanLink93[9] , \ScanLink108[31] , \ScanLink108[28] , 
        \Level1Out141[9] , \ScanLink161[1] , \ScanLink186[19] , 
        \Level1Out196[18] , \Level16Out160[19] , \Level4Out104[5] , 
        \ScanLink201[4] , \Level2Out20[18] , \Level2Out76[19] , 
        \Level8Load96[0] , \ScanLink202[7] , \Level8Out32[17] , 
        \Level8Out64[16] , \ScanLink162[2] , \ScanLink15[20] , 
        \ScanLink15[13] , \ScanLink20[6] , \ScanLink23[16] , \ScanLink56[26] , 
        \Level1Out87[12] , \Level1Out92[26] , \Level2Out130[6] , 
        \Level1Out118[29] , \Level2Out122[29] , \Level2Out174[31] , 
        \Level8Out64[7] , \Level1Out118[30] , \Level1Out188[20] , 
        \Level2Out122[30] , \Level2Out174[28] , \Level2Out250[3] , 
        \Level1Out238[13] , \Level2Out184[25] , \Level2Out234[16] , 
        \Level4Out180[27] , \Level16Out128[20] , \Level2Out254[12] , 
        \Level32Out128[15] , \Level2Out202[13] , \Level4Out96[14] , 
        \ScanLink60[23] , \ScanLink75[17] , \Level1Out123[3] , 
        \ScanLink228[12] , \Level64Out0[7] , \Level2Out68[21] , 
        \ScanLink198[21] , \ScanLink248[16] , \ScanLink23[5] , 
        \ScanLink36[22] , \ScanLink43[12] , \Level1Out243[6] , 
        \ScanLink103[24] , \ScanLink120[15] , \Level1Out120[0] , 
        \Level2Load32[0] , \ScanLink176[14] , \ScanLink100[8] , 
        \Level1Out106[11] , \ScanLink116[10] , \ScanLink135[21] , 
        \ScanLink155[25] , \ScanLink140[11] , \Level1Out240[5] , 
        \Level1Out125[20] , \ScanLink163[20] , \Level2Out86[14] , 
        \Level2Out232[9] , \Level1Out150[10] , \Level1Out113[25] , 
        \Level1Out173[21] , \Level1Out130[14] , \Level1Out166[15] , 
        \Level2Out16[0] , \Level16Out240[23] , \Level1Out145[24] , 
        \ScanLink248[25] , \Level1Out17[31] , \Level1Out17[28] , 
        \Level1Out18[7] , \ScanLink23[25] , \ScanLink36[11] , \ScanLink60[10] , 
        \Level1Out147[7] , \ScanLink198[12] , \ScanLink43[21] , 
        \ScanLink44[2] , \ScanLink56[15] , \Level1Out227[2] , 
        \Level2Out68[12] , \ScanLink75[24] , \ScanLink96[4] , 
        \Level1Out195[1] , \ScanLink228[21] , \Level2Out184[16] , 
        \Level4Out44[9] , \Level32Out128[26] , \Level2Out254[21] , 
        \Level1Out238[20] , \Level2Out128[4] , \Level2Out202[20] , 
        \Level4Out96[27] , \Level4Out180[14] , \Level1Out41[30] , 
        \Level16Out128[13] , \Level1Out62[18] , \Level1Out188[13] , 
        \Level2Out234[25] , \Level2Out248[1] , \Level1Out34[19] , 
        \Level1Out41[29] , \ScanLink47[1] , \ScanLink88[8] , \ScanLink95[7] , 
        \Level1Out166[26] , \Level1Out99[19] , \Level1Out113[16] , 
        \Level1Out125[13] , \Level1Out130[27] , \Level1Out145[17] , 
        \Level4Out88[3] , \Level1Out150[23] , \Level1Out196[2] , 
        \ScanLink204[9] , \Level16Out240[10] , \Level2Out72[4] , 
        \Level1Out173[12] , \Level1Out106[22] , \ScanLink140[22] , 
        \Level2Out136[8] , \ScanLink135[12] , \Level1Out102[13] , 
        \ScanLink103[17] , \ScanLink116[23] , \ScanLink163[13] , 
        \Level1Out144[4] , \ScanLink219[6] , \Level2Out86[27] , 
        \ScanLink176[27] , \Level1Out117[27] , \ScanLink120[26] , 
        \ScanLink155[16] , \ScanLink179[3] , \Level1Out224[1] , 
        \Level1Out121[22] , \Level1Out134[16] , \Level1Out162[17] , 
        \Level2Out158[17] , \Level2Out56[2] , \Level32Out224[10] , 
        \Level1Out141[26] , \Level1Out154[12] , \Level16Out224[25] , 
        \Level16Out16[18] , \ScanLink112[12] , \ScanLink131[23] , 
        \Level1Out177[23] , \Level2Out138[13] , \ScanLink144[13] , 
        \Level1Out200[7] , \Level2Out82[16] , \Level2Out84[4] , 
        \ScanLink11[11] , \ScanLink63[7] , \ScanLink107[26] , 
        \ScanLink167[22] , \ScanLink124[17] , \Level1Out160[2] , 
        \Level8Out48[30] , \ScanLink172[16] , \ScanLink64[21] , 
        \ScanLink151[27] , \Level8Out48[29] , \ScanLink239[24] , 
        \ScanLink27[14] , \ScanLink32[20] , \ScanLink47[10] , 
        \Level1Out203[4] , \ScanLink52[24] , \ScanLink60[4] , \ScanLink71[15] , 
        \Level1Out163[1] , \ScanLink189[17] , \Level1Out199[16] , 
        \Level2Out180[27] , \Level2Out250[10] , \Level1Out13[19] , 
        \Level1Out30[31] , \Level1Out66[29] , \ScanLink143[9] , 
        \Level1Out249[21] , \Level2Out206[11] , \Level4Out92[16] , 
        \Level1Out229[25] , \Level1Out30[28] , \Level1Out45[18] , 
        \Level1Out66[30] , \Level4Out184[25] , \Level1Out46[9] , 
        \Level1Out89[0] , \Level1Out104[6] , \ScanLink107[15] , 
        \ScanLink172[25] , \Level2Out230[14] , \ScanLink112[21] , 
        \ScanLink124[24] , \ScanLink151[14] , \ScanLink131[10] , 
        \ScanLink139[1] , \ScanLink144[20] , \ScanLink167[11] , 
        \Level2Out82[25] , \Level1Out154[21] , \Level2Out32[6] , 
        \Level16Out224[16] , \Level1Out102[20] , \Level1Out121[11] , 
        \Level1Out177[10] , \Level2Out138[20] , \Level1Out117[14] , 
        \Level1Out162[24] , \Level2Out158[24] , \Level32Out224[23] , 
        \Level1Out119[9] , \Level1Out134[25] , \Level1Out141[15] , 
        \Level1Out199[25] , \Level1Out229[16] , \Level4Out184[16] , 
        \ScanLink247[8] , \Level2Out180[14] , \Level2Out208[3] , 
        \Level2Out230[27] , \Level2Out250[23] , \Level1Out249[12] , 
        \Level2Out206[22] , \Level2Out168[6] , \Level4Out92[25] , 
        \Level1Out0[25] , \Level1Out0[16] , \ScanLink2[26] , \ScanLink8[20] , 
        \ScanLink11[22] , \ScanLink27[27] , \ScanLink52[17] , \Level1Out58[5] , 
        \ScanLink71[26] , \ScanLink189[24] , \Level1Out24[3] , 
        \ScanLink32[13] , \ScanLink64[12] , \Level1Out107[5] , 
        \ScanLink239[17] , \ScanLink47[23] , \ScanLink179[29] , 
        \ScanLink78[6] , \ScanLink146[4] , \ScanLink179[30] , 
        \Level8Out56[22] , \ScanLink226[1] , \Level16Out128[1] , 
        \ScanLink8[13] , \Level1Out8[2] , \Level1Out96[17] , \Level1Out18[26] , 
        \ScanLink65[9] , \Level1Out83[23] , \Level1Out169[28] , 
        \ScanLink194[2] , \Level1Out206[9] , \Level16Out48[4] , 
        \Level8Out40[1] , \Level2Out114[0] , \Level2Out126[18] , 
        \Level1Out169[31] , \Level2Out170[19] , \Level1Out27[0] , 
        \Level1Out78[22] , \ScanLink158[8] , \ScanLink197[1] , 
        \Level2Out0[17] , \Level1Out192[30] , \Level64Out64[0] , 
        \ScanLink145[7] , \ScanLink182[31] , \Level1Out192[29] , 
        \Level1Out218[5] , \Level4Out240[6] , \ScanLink182[28] , 
        \Level1Out83[10] , \Level1Out178[0] , \ScanLink225[2] , 
        \Level2Out24[30] , \Level2Out72[28] , \Level4Out120[3] , 
        \Level2Out24[29] , \Level2Out72[31] , \Level8Out24[5] , 
        \Level1Out92[1] , \Level2Out210[1] , \ScanLink10[31] , 
        \Level1Out18[15] , \Level1Out40[7] , \Level1Out96[24] , 
        \Level1Out102[8] , \Level2Out170[4] , \ScanLink122[0] , 
        \Level2Out34[8] , \Level8Out56[11] , \Level1Out43[4] , 
        \ScanLink81[18] , \ScanLink232[28] , \ScanLink242[5] , 
        \Level4Out8[18] , \ScanLink59[31] , \ScanLink59[28] , \ScanLink121[3] , 
        \ScanLink211[19] , \ScanLink232[31] , \ScanLink247[18] , 
        \Level4Out224[2] , \Level1Out78[11] , \Level1Out91[2] , 
        \ScanLink241[6] , \Level4Out144[7] , \Level1Out222[29] , 
        \Level2Out0[24] , \Level2Out218[29] , \Level1Out87[6] , 
        \Level1Out201[18] , \Level1Out222[30] , \Level2Out218[30] , 
        \Level4Out196[1] , \Level16Out224[8] , \ScanLink10[28] , 
        \ScanLink33[19] , \ScanLink46[29] , \Level1Out12[20] , 
        \Level1Out31[11] , \ScanLink46[30] , \Level4Out180[5] , 
        \ScanLink65[18] , \Level2Out218[9] , \Level1Out44[21] , 
        \Level1Out55[0] , \Level4Out0[6] , \Level4Out232[6] , 
        \Level64Out192[24] , \Level1Out24[25] , \Level1Out67[10] , 
        \ScanLink137[7] , \Level1Out72[24] , \Level1Out248[18] , 
        \Level2Out224[19] , \Level1Out51[15] , \Level4Out152[3] , 
        \Level32Out96[23] , \ScanLink134[4] , \Level2Load18[0] , 
        \Level8Out144[24] , \ScanLink2[15] , \Level1Load3[0] , \Level1Out3[9] , 
        \Level1Out12[13] , \ScanLink17[9] , \Level1Out56[3] , 
        \Level8Out112[25] , \Level1Load74[0] , \Level1Out84[5] , 
        \Level1Out89[25] , \Level1Out109[3] , \ScanLink254[1] , 
        \Level4Out148[18] , \Level2Out206[5] , \Level8Out32[1] , 
        \Level2Out166[0] , \Level1Out24[16] , \Level1Out51[26] , 
        \Level1Out72[17] , \ScanLink153[3] , \Level8Out48[9] , 
        \Level32Out96[10] , \Level1Out31[22] , \Level1Out31[4] , 
        \Level2Load206[0] , \Level1Out44[12] , \Level4Out136[7] , 
        \ScanLink233[6] , \Level2Out194[19] , \Level4Out220[31] , 
        \Level1Out67[23] , \Level4Out220[28] , \Level64Out192[17] , 
        \Level1Out32[7] , \ScanLink113[18] , \ScanLink181[5] , 
        \Level2Out18[19] , \Level2Out58[4] , \ScanLink130[30] , 
        \ScanLink130[29] , \ScanLink166[28] , \ScanLink145[19] , 
        \ScanLink166[31] , \Level1Out170[8] , \ScanLink182[6] , 
        \Level1Load217[0] , \Level2Out102[4] , \Level8Out56[5] , 
        \Level2Out96[31] , \Level2Out96[28] , \Level2Out46[8] , 
        \Level1Out89[16] , \Level1Out103[19] , \ScanLink150[0] , 
        \Level16Load176[0] , \Level1Out120[31] , \Level1Out120[28] , 
        \Level1Out176[29] , \Level8Out144[17] , \Level8Out112[16] , 
        \Level1Out155[18] , \Level1Out176[30] , \Level1Out193[10] , 
        \ScanLink230[5] , \Level1Out236[17] , \ScanLink12[4] , 
        \Level1Out81[8] , \Level1Out215[26] , \Level1Out243[27] , 
        \Level1Out111[1] , \Level1Out200[12] , \Level1Out186[24] , 
        \Level1Out223[23] , \Level4Out208[15] , \ScanLink38[26] , 
        \ScanLink131[9] , \ScanLink210[13] , \Level2Out50[20] , 
        \ScanLink58[22] , \ScanLink183[11] , \ScanLink196[25] , 
        \ScanLink233[22] , \ScanLink246[12] , \Level8Out0[23] , 
        \ScanLink226[16] , \ScanLink253[26] , \Level2Out66[25] , 
        \ScanLink95[26] , \Level1Load108[0] , \ScanLink118[14] , 
        \ScanLink205[27] , \Level2Out30[24] , \Level2Out88[10] , 
        \Level2Out24[2] , \Level1Out6[4] , \ScanLink9[19] , \ScanLink11[7] , 
        \ScanLink80[12] , \Level1Out108[15] , \Level1Out168[11] , 
        \ScanLink178[10] , \Level2Out104[10] , \Level4Out40[20] , 
        \Level2Out152[11] , \Level4Out136[17] , \Level4Out16[21] , 
        \Level4Out160[16] , \Level2Out4[0] , \Level4Out76[25] , 
        \Level2Out132[15] , \Level4Out100[12] , \Level2Out164[14] , 
        \Level4Out156[13] , \Level1Out112[2] , \Level4Out20[24] , 
        \ScanLink183[22] , \ScanLink253[15] , \Level2Out66[16] , 
        \Level8Out0[10] , \ScanLink226[25] , \ScanLink38[15] , 
        \ScanLink58[11] , \ScanLink205[14] , \Level2Out30[17] , 
        \Level2Out50[13] , \ScanLink148[2] , \Level1Out186[17] , 
        \ScanLink196[16] , \ScanLink210[20] , \ScanLink233[11] , 
        \ScanLink235[8] , \ScanLink246[21] , \Level32Out160[5] , 
        \Level1Out200[21] , \Level4Out208[26] , \Level1Out215[0] , 
        \Level1Out223[10] , \Level1Out4[27] , \Level1Out4[14] , 
        \Level1Out5[7] , \Level1Out29[6] , \ScanLink76[0] , \Level1Out79[28] , 
        \Level1Out193[23] , \Level1Out243[14] , \Level1Out236[24] , 
        \Level1Out79[31] , \Level1Out215[15] , \ScanLink228[7] , 
        \Level1Out108[26] , \Level1Out175[5] , \ScanLink184[8] , 
        \Level2Out132[26] , \Level4Out100[21] , \Level4Out76[16] , 
        \Level1Out216[3] , \Level2Out92[0] , \Level4Out20[17] , 
        \ScanLink75[3] , \Level1Out82[30] , \Level2Out164[27] , 
        \Level4Out156[20] , \Level4Out136[24] , \Level1Out82[29] , 
        \Level1Out176[6] , \Level2Out104[23] , \Level4Out68[7] , 
        \Level4Out40[13] , \Level1Out168[22] , \Level4Out16[12] , 
        \Level2Out152[22] , \Level4Out160[25] , \ScanLink29[10] , 
        \Level1Out34[9] , \ScanLink80[21] , \ScanLink199[7] , 
        \ScanLink178[23] , \Level2Out40[6] , \ScanLink51[5] , \ScanLink95[15] , 
        \ScanLink118[27] , \Level2Out88[23] , \Level2Out136[17] , 
        \Level4Out72[27] , \Level128Out128[1] , \Level8Out168[31] , 
        \Level4Out104[10] , \ScanLink83[3] , \Level1Out86[18] , 
        \Level1Out119[23] , \Level1Out152[0] , \Level1Out179[27] , 
        \Level2Out160[16] , \Level4Out152[11] , \Level8Out168[28] , 
        \Level2Load40[0] , \Level4Out24[26] , \Level2Out100[12] , 
        \Level2Out240[9] , \Level4Out44[22] , \Level2Out156[13] , 
        \Level4Out132[15] , \Level4Out164[14] , \Level1Out232[5] , 
        \Level4Out12[23] , \ScanLink84[10] , \ScanLink109[22] , 
        \Level1Out180[6] , \ScanLink91[24] , \ScanLink169[26] , 
        \Level2Out64[0] , \ScanLink172[8] , \Level64Out0[17] , 
        \Level1Out183[5] , \ScanLink187[13] , \ScanLink222[14] , 
        \ScanLink201[25] , \Level2Out34[26] , \Level2Out62[27] , 
        \ScanLink49[14] , \ScanLink80[0] , \ScanLink214[11] , \ScanLink52[6] , 
        \Level1Out151[3] , \ScanLink192[27] , \ScanLink237[20] , 
        \Level2Out54[22] , \Level1Out204[10] , \ScanLink242[10] , 
        \Level32Out224[6] , \Level1Out182[26] , \Level1Out227[21] , 
        \Level1Out197[12] , \Level1Out252[11] , \Level1Out232[15] , 
        \Level1Out247[25] , \Level2Out208[15] , \ScanLink35[1] , 
        \ScanLink84[23] , \ScanLink91[17] , \ScanLink169[15] , 
        \Level1Out211[24] , \Level1Out231[6] , \Level64Out0[24] , 
        \ScanLink109[11] , \Level1Out136[4] , \Level2Out100[21] , 
        \Level4Out28[5] , \Level4Out132[26] , \Level4Out44[11] , 
        \Level2Out144[8] , \Level4Out12[10] , \Level4Out164[27] , 
        \Level1Out69[4] , \Level1Out119[10] , \Level1Out179[14] , 
        \Level2Out156[20] , \Level4Out104[23] , \Level2Out136[24] , 
        \Level4Out24[15] , \Level4Out72[14] , \Level1Out247[16] , 
        \Level2Out160[25] , \Level4Out152[22] , \ScanLink6[24] , 
        \ScanLink29[23] , \ScanLink36[2] , \Level1Out197[21] , 
        \Level2Out188[2] , \Level2Out208[26] , \Level1Out232[26] , 
        \ScanLink49[27] , \ScanLink108[0] , \Level1Out135[7] , 
        \Level1Out211[17] , \Level8Out200[18] , \Level1Out182[15] , 
        \Level1Out204[23] , \Level1Out227[12] , \Level1Out252[22] , 
        \Level1Out255[2] , \ScanLink214[22] , \Level2Out54[11] , 
        \Level1Out77[8] , \Level1Out128[8] , \ScanLink192[14] , 
        \ScanLink237[13] , \ScanLink242[23] , \Level4Out36[9] , 
        \Level2Out62[14] , \ScanLink187[20] , \ScanLink222[27] , 
        \ScanLink98[2] , \ScanLink117[29] , \ScanLink141[31] , 
        \ScanLink162[19] , \ScanLink201[16] , \Level2Out34[15] , 
        \ScanLink134[18] , \ScanLink141[28] , \Level2Out126[2] , 
        \Level1Out98[13] , \ScanLink117[30] , \Level1Out149[1] , 
        \ScanLink169[9] , \Level8Out72[3] , \Level1Out186[8] , 
        \ScanLink214[3] , \Level2Out92[19] , \Level2Out246[7] , 
        \Level8Out176[23] , \Level8Out120[22] , \Level1Out107[28] , 
        \Level1Out151[30] , \Level1Out172[18] , \ScanLink174[6] , 
        \Level1Out229[4] , \Level2Out148[18] , \ScanLink6[17] , 
        \Level1Out15[2] , \Level1Out16[1] , \Level1Out151[29] , 
        \Level1Out20[27] , \ScanLink49[7] , \Level1Out107[31] , 
        \Level1Out124[19] , \Level1Out76[26] , \Level4Out112[1] , 
        \Level1Out35[13] , \Level1Out55[17] , \ScanLink217[0] , 
        \Level8Out248[21] , \Level2Out190[28] , \Level1Out16[22] , 
        \Level1Out40[23] , \ScanLink54[8] , \Level1Out63[12] , 
        \ScanLink177[5] , \Level2Out190[31] , \Level4Out224[19] , 
        \Level1Out189[19] , \Level1Load82[0] , \Level1Load150[0] , 
        \Level1Out198[4] , \ScanLink199[18] , \Level8Out80[16] , 
        \Level1Out237[8] , \Level64Out64[13] , \Level2Out190[0] , 
        \Level1Out98[20] , \Level1Out72[5] , \ScanLink110[2] , 
        \Level8Out120[11] , \Level8Out176[10] , \Level1Out133[9] , 
        \ScanLink229[18] , \Level2Out142[6] , \Level2Out222[3] , 
        \Level4Out168[9] , \Level8Out16[7] , \Level1Out0[2] , \Level1Out3[1] , 
        \ScanLink14[19] , \ScanLink37[31] , \ScanLink37[28] , \ScanLink42[18] , 
        \ScanLink61[30] , \Level64Out64[20] , \ScanLink61[29] , 
        \Level2Out18[6] , \Level8Out80[25] , \Level1Out16[11] , 
        \Level1Out35[20] , \Level1Out40[10] , \Level4Out176[5] , 
        \Level8Out248[12] , \Level1Out63[21] , \Level1Out20[14] , 
        \Level1Out55[24] , \Level1Out76[15] , \Level1Out239[19] , 
        \Level4Out216[0] , \ScanLink113[1] , \Level2Out220[31] , 
        \Level1Out71[6] , \Level2Out220[28] , \ScanLink73[5] , 
        \ScanLink106[24] , \ScanLink113[10] , \ScanLink130[21] , 
        \Level4Out248[6] , \ScanLink145[11] , \Level1Out210[5] , 
        \Level2Out94[6] , \ScanLink166[20] , \ScanLink125[15] , 
        \Level1Out170[0] , \ScanLink173[14] , \Level2Out96[20] , 
        \Level4Out128[3] , \Level2Load62[0] , \ScanLink150[25] , 
        \Level1Out103[11] , \Level1Out116[25] , \Level1Out120[20] , 
        \Level1Out135[14] , \ScanLink150[8] , \Level4Out68[15] , 
        \Level1Out163[15] , \Level2Out46[0] , \Level4Out148[23] , 
        \Level1Out140[24] , \Level1Out155[10] , \Level4Out128[27] , 
        \Level1Out176[21] , \Level2Out224[22] , \Level32Out96[18] , 
        \Level4Out216[25] , \ScanLink3[24] , \ScanLink3[8] , \ScanLink8[3] , 
        \ScanLink9[22] , \ScanLink10[20] , \ScanLink10[13] , \ScanLink65[23] , 
        \Level1Out198[14] , \Level1Out228[27] , \Level1Out248[23] , 
        \Level4Out240[24] , \Level8Out48[1] , \Level2Out194[11] , 
        \Level2Out212[27] , \Level2Out244[26] , \Level4Out220[20] , 
        \ScanLink238[26] , \ScanLink17[1] , \ScanLink26[16] , \ScanLink33[22] , 
        \ScanLink46[12] , \Level2Out78[15] , \Level16Out240[4] , 
        \ScanLink53[26] , \Level1Out213[6] , \ScanLink70[6] , \ScanLink70[17] , 
        \ScanLink188[15] , \Level2Out18[11] , \Level1Out99[2] , 
        \Level1Out120[13] , \Level1Out155[23] , \Level1Out173[3] , 
        \Level4Out128[14] , \Level2Out22[4] , \Level1Out103[22] , 
        \Level1Out176[12] , \ScanLink106[17] , \Level1Out116[16] , 
        \Level1Out163[26] , \Level1Out135[27] , \Level1Out140[17] , 
        \Level4Out68[26] , \Level4Out148[10] , \ScanLink173[27] , 
        \ScanLink254[9] , \ScanLink125[26] , \ScanLink129[3] , 
        \ScanLink150[16] , \Level2Out96[13] , \Level2Out2[6] , 
        \ScanLink145[22] , \Level8Out32[9] , \Level2Out166[8] , 
        \ScanLink26[25] , \ScanLink113[23] , \Level1Out114[4] , 
        \ScanLink130[12] , \ScanLink166[13] , \ScanLink249[6] , 
        \Level16Out224[0] , \Level1Out48[7] , \ScanLink53[15] , 
        \ScanLink188[26] , \Level2Out18[22] , \ScanLink70[24] , 
        \Level1Out12[31] , \Level1Out12[28] , \ScanLink14[2] , 
        \ScanLink33[11] , \ScanLink65[10] , \Level2Out78[26] , 
        \Level16Out144[5] , \Level1Out117[7] , \ScanLink238[15] , 
        \ScanLink46[21] , \Level4Out220[13] , \Level1Out44[30] , 
        \Level2Out212[14] , \Level1Out67[18] , \Level1Out228[14] , 
        \Level2Out194[22] , \Level1Out31[19] , \Level1Out44[29] , 
        \Level2Out218[1] , \Level1Out55[8] , \Level2Out244[15] , 
        \Level1Out198[27] , \Level1Out248[10] , \Level2Out178[4] , 
        \Level2Out224[11] , \Level4Out216[16] , \Level2Out92[8] , 
        \Level4Out100[30] , \Level4Out240[17] , \ScanLink9[11] , 
        \Level1Out19[24] , \Level1Out34[1] , \ScanLink80[29] , 
        \Level1Out82[21] , \Level1Out97[15] , \Level4Out156[28] , 
        \ScanLink184[0] , \Level4Out100[29] , \Level2Out104[2] , 
        \Level4Out156[31] , \Level1Out37[2] , \ScanLink58[19] , 
        \ScanLink68[4] , \ScanLink80[30] , \ScanLink156[6] , \ScanLink155[5] , 
        \ScanLink236[3] , \Level128Out128[9] , \Level1Out208[7] , 
        \Level1Out168[2] , \ScanLink246[29] , \Level4Out76[3] , 
        \Level8Out0[18] , \ScanLink210[31] , \ScanLink210[28] , 
        \ScanLink233[19] , \ScanLink235[0] , \ScanLink246[30] , 
        \Level1Out50[5] , \ScanLink76[8] , \Level1Load172[0] , 
        \ScanLink187[3] , \Level1Out200[30] , \Level1Out215[8] , 
        \Level1Out223[18] , \Level1Out200[29] , \Level8Out232[17] , 
        \Level1Out79[20] , \ScanLink132[2] , \Level2Out88[18] , 
        \Level1Out82[12] , \ScanLink178[18] , \ScanLink252[7] , 
        \Level2Out4[8] , \Level2Out152[19] , \Level4Out40[31] , 
        \Level1Out82[3] , \Level1Out168[19] , \Level4Out16[29] , 
        \Level2Out200[3] , \Level4Out40[28] , \Level2Out104[18] , 
        \Level4Out16[30] , \Level1Out10[7] , \Level1Out13[4] , 
        \Level1Out19[17] , \Level1Out79[13] , \Level1Out81[0] , 
        \Level1Out97[26] , \Level2Out160[6] , \Level1Out193[18] , 
        \ScanLink28[6] , \Level1Out53[6] , \Level1Out111[9] , 
        \Level8Out232[24] , \Level2Out50[31] , \Level1Out68[16] , 
        \ScanLink108[8] , \ScanLink131[1] , \ScanLink183[19] , 
        \Level2Out50[28] , \Level4Load224[0] , \Level1Out197[30] , 
        \ScanLink251[4] , \Level4Out12[7] , \Level32Out96[4] , 
        \Level1Out197[29] , \Level8Out200[10] , \Level1Out77[0] , 
        \ScanLink115[7] , \Level1Out128[0] , \Level4Out36[1] , 
        \Level16Out96[16] , \ScanLink187[31] , \Level2Out54[19] , 
        \ScanLink187[28] , \Level1Out248[5] , \Level2Out196[6] , 
        \ScanLink29[18] , \ScanLink35[9] , \Level1Load56[0] , \Level1Out74[3] , 
        \ScanLink109[19] , \ScanLink116[4] , \Level2Out144[0] , 
        \Level1Out86[23] , \Level2Out100[30] , \Level4Out12[18] , 
        \Level1Out119[18] , \Level2Out156[28] , \ScanLink80[8] , 
        \Level1Out93[17] , \Level2Out100[29] , \Level2Out156[31] , 
        \Level4Out44[19] , \Level2Out224[5] , \Level8Out168[13] , 
        \Level1Load184[0] , \ScanLink211[6] , \Level4Out52[5] , 
        \ScanLink237[28] , \Level2Load224[0] , \Level1Out68[25] , 
        \ScanLink171[3] , \ScanLink214[19] , \ScanLink237[31] , 
        \ScanLink242[18] , \ScanLink84[18] , \Level1Out86[10] , 
        \Level1Out93[24] , \Level1Out152[8] , \Level1Out204[18] , 
        \Level1Out227[30] , \Level1Out227[29] , \Level1Out252[19] , 
        \Level16Out96[25] , \Level4Out80[3] , \Level4Out152[19] , 
        \Level8Out200[23] , \Level1Load235[0] , \Level8Out168[20] , 
        \Level2Out120[4] , \Level4Out104[18] , \Level2Out240[1] , 
        \ScanLink172[0] , \ScanLink212[5] , \Level2Out64[8] , \ScanLink14[11] , 
        \ScanLink22[14] , \ScanLink30[4] , \ScanLink57[24] , 
        \Level64Out64[28] , \ScanLink61[21] , \ScanLink74[15] , 
        \ScanLink229[10] , \Level16Out160[3] , \Level1Out133[1] , 
        \Level64Out64[31] , \ScanLink199[23] , \Level1Out16[19] , 
        \Level1Out35[31] , \ScanLink37[20] , \ScanLink42[10] , 
        \ScanLink249[14] , \Level1Out63[29] , \Level1Out189[22] , 
        \Level1Out253[4] , \Level2Out216[25] , \ScanLink33[7] , 
        \Level1Out35[28] , \Level1Out40[18] , \Level1Out63[30] , 
        \Level2Out240[24] , \Level4Out224[22] , \Level1Out98[31] , 
        \ScanLink113[9] , \Level1Out239[11] , \Level2Out190[13] , 
        \Level2Out220[20] , \Level4Out212[27] , \Level4Out244[26] , 
        \Level4Out216[8] , \Level1Out124[22] , \Level8Out184[4] , 
        \Level1Out98[28] , \Level1Out107[13] , \Level1Out151[12] , 
        \Level2Out148[23] , \Level2Out190[8] , \ScanLink102[26] , 
        \Level1Out112[27] , \Level1Out172[23] , \Level8Out120[19] , 
        \Level1Out131[16] , \Level1Out167[17] , \Level2Out128[27] , 
        \Level1Out144[26] , \Level8Out176[18] , \Level2Out92[22] , 
        \Level64Out192[5] , \ScanLink121[17] , \Level1Out130[2] , 
        \ScanLink177[16] , \Level4Out168[1] , \ScanLink154[27] , 
        \ScanLink117[12] , \ScanLink134[23] , \Level4Out208[4] , 
        \ScanLink141[13] , \Level1Out250[7] , \ScanLink162[22] , 
        \Level4Out112[9] , \Level4Out212[14] , \ScanLink14[22] , 
        \ScanLink86[6] , \Level1Out185[3] , \Level2Out220[13] , 
        \ScanLink217[8] , \Level2Out138[6] , \Level1Out189[11] , 
        \Level1Out239[22] , \Level4Out244[15] , \Level2Out216[16] , 
        \Level4Out224[11] , \Level16Out64[2] , \Level8Out248[30] , 
        \Level2Out190[20] , \Level2Out240[17] , \Level8Out248[29] , 
        \Level1Out16[9] , \ScanLink22[27] , \ScanLink37[13] , \ScanLink61[12] , 
        \ScanLink249[27] , \Level1Out157[5] , \ScanLink199[10] , 
        \ScanLink42[23] , \ScanLink54[0] , \ScanLink57[17] , \Level1Out237[0] , 
        \ScanLink57[3] , \ScanLink74[26] , \ScanLink229[23] , 
        \Level32Load128[0] , \ScanLink141[20] , \ScanLink85[5] , 
        \ScanLink102[15] , \ScanLink117[21] , \ScanLink134[10] , 
        \Level1Out154[6] , \ScanLink162[11] , \ScanLink209[4] , 
        \ScanLink177[25] , \Level2Out92[11] , \ScanLink121[24] , 
        \ScanLink154[14] , \Level1Out167[24] , \ScanLink169[1] , 
        \Level1Out234[3] , \Level2Out128[14] , \Level1Out112[14] , 
        \Level1Out131[25] , \Level1Out144[15] , \Level1Out149[9] , 
        \Level1Out186[0] , \Level1Out151[21] , \Level2Load94[0] , 
        \Level2Out62[6] , \ScanLink41[7] , \ScanLink85[12] , \ScanLink93[1] , 
        \Level1Out107[20] , \Level1Out124[11] , \Level1Out172[10] , 
        \Level2Out148[10] , \ScanLink108[20] , \Level2Out98[24] , 
        \Level1Out190[4] , \ScanLink90[26] , \Level1Load158[0] , 
        \Level2Out74[2] , \ScanLink168[24] , \Level1Out178[25] , 
        \Level2Out142[25] , \Level16Out208[12] , \Level1Out118[21] , 
        \Level1Out142[2] , \Level2Out114[24] , \Level2Out174[20] , 
        \Level1Out205[12] , \Level1Out222[7] , \Level2Out122[21] , 
        \ScanLink5[6] , \Level1Out5[25] , \Level1Out5[16] , \ScanLink42[4] , 
        \Level1Out141[1] , \Level16Out112[3] , \Level1Out183[24] , 
        \Level1Out226[23] , \Level32Out160[24] , \Level1Out253[13] , 
        \Level4Out88[24] , \Level1Out196[10] , \Level1Out221[4] , 
        \Level1Out233[17] , \ScanLink25[3] , \ScanLink28[12] , \ScanLink90[2] , 
        \ScanLink186[11] , \Level1Out210[26] , \Level1Out246[27] , 
        \Level16Out160[11] , \Level2Out16[15] , \Level1Out193[7] , 
        \ScanLink223[16] , \ScanLink200[27] , \ScanLink256[26] , 
        \Level2Out40[14] , \ScanLink48[16] , \Level1Out87[30] , 
        \ScanLink161[9] , \ScanLink215[13] , \Level2Out20[10] , 
        \ScanLink193[25] , \ScanLink236[22] , \ScanLink243[12] , 
        \Level2Out76[11] , \Level1Out87[29] , \Level1Out126[6] , 
        \Level2Out174[13] , \Level2Out122[12] , \ScanLink28[21] , 
        \ScanLink48[25] , \Level1Out64[9] , \Level1Out79[6] , 
        \Level1Out118[12] , \Level1Out178[16] , \Level1Out246[3] , 
        \Level2Out142[16] , \Level16Out208[21] , \Level2Out114[17] , 
        \ScanLink85[21] , \ScanLink90[15] , \ScanLink168[17] , 
        \ScanLink108[13] , \Level2Out10[6] , \Level2Out98[17] , 
        \ScanLink186[22] , \ScanLink193[16] , \ScanLink215[20] , 
        \ScanLink236[11] , \ScanLink243[21] , \Level2Out20[23] , 
        \Level4Out160[9] , \Level2Out76[22] , \ScanLink256[15] , 
        \Level2Out16[26] , \ScanLink223[25] , \Level2Out40[27] , 
        \ScanLink200[14] , \Level16Out16[2] , \Level2Out198[0] , 
        \Level8Out192[0] , \ScanLink6[5] , \ScanLink7[26] , \ScanLink26[0] , 
        \Level1Out246[14] , \Level1Out99[11] , \ScanLink118[2] , 
        \Level1Out125[5] , \Level1Out196[23] , \Level1Out233[24] , 
        \Level16Out176[7] , \Level1Out183[17] , \Level1Out205[21] , 
        \Level1Out210[15] , \Level16Out160[22] , \Level1Out226[10] , 
        \Level1Out253[20] , \Level8Out192[18] , \Level4Out88[17] , 
        \Level32Out160[17] , \Level1Out159[3] , \Level1Out245[0] , 
        \ScanLink204[1] , \Level16Out240[18] , \ScanLink164[4] , 
        \Level1Out239[6] , \ScanLink15[31] , \Level1Load24[0] , 
        \ScanLink47[9] , \Level2Out136[0] , \ScanLink88[0] , \Level1Out224[9] , 
        \ScanLink15[28] , \ScanLink36[19] , \ScanLink43[29] , \Level4Out96[7] , 
        \ScanLink7[15] , \Level1Out17[20] , \Level1Out21[25] , 
        \ScanLink43[30] , \Level1Out188[6] , \ScanLink59[5] , \ScanLink60[18] , 
        \Level1Out77[24] , \ScanLink228[30] , \ScanLink228[29] , 
        \Level2Out202[28] , \Level1Out238[28] , \Level2Out254[30] , 
        \Level2Out202[31] , \Level4Out44[1] , \Level1Out34[11] , 
        \Level1Out54[15] , \Level1Out195[9] , \ScanLink207[2] , 
        \Level1Out238[31] , \Level2Out254[29] , \Level2Load48[0] , 
        \Level1Out41[21] , \Level2Out248[9] , \Level1Out62[10] , 
        \Level1Out99[22] , \Level1Out106[19] , \ScanLink116[18] , 
        \Level1Out120[8] , \ScanLink167[7] , \Level1Load247[0] , 
        \Level2Out152[4] , \Level32Out128[7] , \ScanLink135[30] , 
        \Level2Out232[1] , \ScanLink135[29] , \ScanLink163[28] , 
        \ScanLink140[19] , \ScanLink163[31] , \Level1Out125[31] , 
        \Level1Out173[29] , \Level2Out180[2] , \Level1Out125[28] , 
        \Level1Out150[18] , \Level1Out173[30] , \Level1Out13[22] , 
        \Level1Out17[13] , \Level1Out34[22] , \Level1Out41[12] , 
        \Level1Out62[7] , \Level2Out16[8] , \ScanLink100[0] , 
        \Level1Out188[31] , \Level4Out20[5] , \Level1Out62[23] , 
        \Level16Out128[31] , \Level1Out188[28] , \Level1Out21[16] , 
        \Level1Out54[26] , \Level1Out77[17] , \Level16Out128[28] , 
        \ScanLink103[3] , \Level1Out61[4] , \Level1Out30[13] , 
        \ScanLink198[30] , \Level2Out68[30] , \Level2Out68[29] , 
        \ScanLink198[29] , \Level1Out45[23] , \Level1Out45[2] , 
        \ScanLink19[7] , \Level1Out66[12] , \ScanLink127[5] , 
        \Level1Out25[27] , \Level1Out73[26] , \Level1Out50[17] , 
        \ScanLink247[0] , \Level1Out94[7] , \Level1Out97[4] , 
        \Level1Load100[0] , \ScanLink139[9] , \Level8Out48[12] , 
        \Level2Out216[7] , \Level1Out102[28] , \ScanLink112[30] , 
        \ScanLink112[29] , \ScanLink144[31] , \ScanLink167[19] , 
        \Level16Out0[26] , \ScanLink131[18] , \ScanLink144[28] , 
        \Level2Out176[2] , \ScanLink124[6] , \Level1Out154[30] , 
        \Level1Out177[18] , \Level2Out138[28] , \Level1Out154[29] , 
        \Level16Out16[23] , \Level2Out138[31] , \ScanLink11[19] , 
        \ScanLink32[31] , \ScanLink32[28] , \Level1Out46[1] , \ScanLink47[18] , 
        \ScanLink64[30] , \Level1Out88[27] , \Level1Out89[8] , 
        \Level1Out102[31] , \Level1Out121[19] , \Level1Out119[1] , 
        \ScanLink244[3] , \ScanLink64[29] , \ScanLink191[7] , \Level2Out48[6] , 
        \Level1Out163[9] , \Level1Out73[15] , \ScanLink143[1] , 
        \Level32Out0[7] , \Level1Out249[29] , \Level2Out206[19] , 
        \ScanLink3[17] , \Level1Out13[11] , \Level1Out21[6] , 
        \Level1Out50[24] , \Level2Out250[18] , \Level1Out25[14] , 
        \Level1Out30[20] , \Level1Out45[10] , \Level1Out249[30] , 
        \Level4Out60[7] , \Level1Out66[21] , \ScanLink223[4] , 
        \Level1Out22[5] , \Level1Out88[14] , \ScanLink140[2] , 
        \Level32Out224[18] , \ScanLink220[7] , \Level16Out16[10] , 
        \Level16Out0[15] , \ScanLink0[2] , \Level1Out1[27] , \Level1Out1[14] , 
        \ScanLink39[24] , \ScanLink192[4] , \ScanLink211[11] , 
        \Level2Out24[12] , \Level2Out112[6] , \Level8Out48[21] , 
        \Level16Out32[4] , \ScanLink59[20] , \ScanLink182[13] , 
        \ScanLink197[27] , \ScanLink232[20] , \ScanLink247[10] , 
        \Level2Out72[13] , \ScanLink204[25] , \ScanLink227[14] , 
        \ScanLink252[24] , \Level2Out12[17] , \Level1Out78[19] , 
        \Level2Out44[16] , \Level1Out192[12] , \Level1Out237[15] , 
        \Level1Out242[25] , \ScanLink81[10] , \Level1Out83[18] , 
        \Level1Out92[9] , \Level1Out101[3] , \Level1Out201[10] , 
        \Level1Out214[24] , \Level4Out196[9] , \Level1Out187[26] , 
        \Level1Out222[21] , \Level2Out170[22] , \Level2Out210[9] , 
        \Level2Out218[21] , \Level4Out8[6] , \Level1Out169[13] , 
        \ScanLink94[24] , \Level1Out102[0] , \Level1Out109[17] , 
        \Level2Out126[23] , \Level2Out146[27] , \ScanLink119[16] , 
        \Level2Load10[0] , \Level2Out34[0] , \Level2Out110[26] , 
        \ScanLink122[8] , \Level8Out56[19] , \ScanLink179[12] , 
        \Level4Out8[10] , \Level4Out188[5] , \ScanLink158[0] , 
        \Level1Out187[15] , \Level1Out201[23] , \Level64Out64[8] , 
        \Level1Out222[12] , \Level2Out218[12] , \ScanLink197[9] , 
        \Level1Out205[2] , \Level1Out242[16] , \ScanLink8[31] , 
        \Level1Out27[8] , \ScanLink66[2] , \Level1Out165[7] , 
        \Level1Out192[21] , \Level1Out237[26] , \Level1Out214[17] , 
        \ScanLink238[5] , \ScanLink252[17] , \ScanLink39[17] , 
        \ScanLink59[13] , \ScanLink182[20] , \ScanLink204[16] , 
        \ScanLink227[27] , \Level2Out12[24] , \Level2Out44[25] , 
        \ScanLink81[23] , \Level1Out178[8] , \ScanLink211[22] , 
        \Level2Out24[21] , \ScanLink247[23] , \Level2Out72[20] , 
        \ScanLink179[21] , \ScanLink189[5] , \ScanLink197[14] , 
        \ScanLink232[13] , \Level4Out8[23] , \Level16Load0[0] , 
        \ScanLink94[17] , \Level2Out50[4] , \ScanLink119[25] , 
        \ScanLink226[9] , \Level16Out128[9] , \ScanLink8[28] , 
        \Level1Out109[24] , \Level1Out206[1] , \Level2Out146[14] , 
        \Level8Out40[9] , \Level2Out82[2] , \Level2Out110[15] , 
        \ScanLink15[21] , \ScanLink15[12] , \ScanLink23[4] , \Level1Out39[4] , 
        \ScanLink65[1] , \Level1Out166[4] , \Level2Out170[11] , 
        \Level1Out169[20] , \Level2Out114[8] , \Level2Out126[10] , 
        \ScanLink116[11] , \Level2Out86[15] , \Level2Out232[8] , 
        \ScanLink120[14] , \ScanLink135[20] , \ScanLink163[21] , 
        \ScanLink140[10] , \Level1Out240[4] , \ScanLink155[24] , 
        \ScanLink36[23] , \ScanLink43[13] , \ScanLink100[9] , 
        \ScanLink103[25] , \Level2Load128[0] , \Level1Out113[24] , 
        \Level1Out120[1] , \ScanLink176[15] , \Level1Out130[15] , 
        \Level2Out16[1] , \Level16Out240[22] , \Level1Out145[25] , 
        \Level1Out106[10] , \Level1Out166[14] , \Level1Out125[21] , 
        \Level1Out173[20] , \Level1Load139[0] , \Level1Out150[11] , 
        \Level1Out238[12] , \Level2Out202[12] , \Level4Out96[15] , 
        \Level1Out188[21] , \Level2Out184[24] , \Level2Out254[13] , 
        \Level2Out234[17] , \Level32Out128[14] , \Level4Out180[26] , 
        \Level16Out128[21] , \ScanLink60[22] , \Level1Out243[7] , 
        \ScanLink198[20] , \Level1Out18[6] , \ScanLink20[7] , \ScanLink56[27] , 
        \ScanLink75[16] , \ScanLink228[13] , \ScanLink248[17] , 
        \Level64Out0[6] , \Level1Out123[2] , \Level2Out68[20] , 
        \ScanLink23[17] , \ScanLink47[0] , \ScanLink95[6] , \Level1Out99[18] , 
        \Level1Out106[23] , \Level1Out173[13] , \Level1Out113[17] , 
        \Level1Out125[12] , \Level1Out150[22] , \Level2Out72[5] , 
        \Level1Out130[26] , \Level1Out145[16] , \Level4Out88[2] , 
        \Level1Out196[3] , \Level1Out166[27] , \ScanLink204[8] , 
        \Level16Out240[11] , \ScanLink103[16] , \ScanLink120[27] , 
        \ScanLink155[17] , \ScanLink176[26] , \ScanLink179[2] , 
        \Level1Out224[0] , \ScanLink116[22] , \Level1Out144[5] , 
        \ScanLink163[12] , \ScanLink219[7] , \Level2Out86[26] , 
        \ScanLink140[23] , \Level2Out136[9] , \ScanLink88[9] , 
        \ScanLink135[13] , \ScanLink228[20] , \Level2Out68[13] , 
        \ScanLink23[24] , \ScanLink75[25] , \ScanLink36[10] , \ScanLink56[14] , 
        \Level1Out227[3] , \ScanLink43[20] , \ScanLink44[3] , 
        \Level1Out17[30] , \ScanLink60[11] , \ScanLink248[24] , 
        \Level1Out147[6] , \ScanLink198[13] , \Level1Out17[29] , 
        \Level1Out34[18] , \Level2Out234[24] , \Level1Out41[28] , 
        \Level2Out248[0] , \ScanLink26[9] , \ScanLink28[31] , \ScanLink38[5] , 
        \Level1Out41[31] , \Level4Out180[15] , \Level16Out128[12] , 
        \Level1Out62[19] , \Level1Out188[12] , \Level1Out64[0] , 
        \ScanLink85[31] , \Level1Out87[20] , \Level1Out92[14] , 
        \ScanLink96[5] , \Level2Out128[5] , \Level2Out202[21] , 
        \Level4Out96[26] , \Level1Out195[0] , \Level1Out238[21] , 
        \Level2Out184[17] , \Level32Out128[27] , \Level4Out44[8] , 
        \Level2Out254[20] , \Level16Out208[28] , \Level2Out154[3] , 
        \Level2Out234[6] , \Level16Out208[31] , \Level16Out208[7] , 
        \ScanLink85[28] , \ScanLink106[7] , \Level8Out32[25] , 
        \Level8Out64[24] , \Level2Out186[5] , \Level32Load224[0] , 
        \ScanLink28[28] , \Level1Out67[3] , \Level4Out200[5] , 
        \Level1Load45[0] , \Level1Out69[15] , \ScanLink105[4] , 
        \Level1Out138[3] , \ScanLink215[29] , \ScanLink243[31] , 
        \Level8Out192[9] , \ScanLink243[28] , \Level4Out160[0] , 
        \Level1Out205[31] , \Level1Out205[28] , \ScanLink215[30] , 
        \ScanLink236[18] , \Level1Out253[30] , \Level1Out253[29] , 
        \Level8Out192[11] , \Level2Out4[14] , \Level1Out226[19] , 
        \Level1Out245[9] , \Level2Out198[9] , \Level1Out87[13] , 
        \ScanLink93[8] , \ScanLink108[30] , \ScanLink162[3] , 
        \Level1Load197[0] , \Level8Out32[16] , \ScanLink108[29] , 
        \Level1Out118[31] , \ScanLink202[6] , \Level2Out174[29] , 
        \Level2Out250[2] , \Level8Out64[17] , \Level1Out118[28] , 
        \Level2Out122[31] , \Level2Out174[30] , \Level2Out122[28] , 
        \Level8Out64[6] , \Level1Out92[27] , \Level2Out130[7] , \ScanLink3[1] , 
        \Level1Out196[19] , \Level16Out160[18] , \ScanLink8[21] , 
        \Level1Out8[3] , \Level1Out18[27] , \Level1Out69[26] , 
        \Level1Out141[8] , \Level8Out192[22] , \Level1Load226[0] , 
        \Level1Out78[23] , \ScanLink161[0] , \Level2Out4[27] , 
        \Level2Load186[0] , \Level2Out20[19] , \ScanLink186[18] , 
        \Level2Out76[18] , \Level1Out192[28] , \ScanLink201[5] , 
        \Level4Out104[4] , \Level1Out192[31] , \Level64Out64[1] , 
        \Level1Out24[2] , \Level1Out27[1] , \ScanLink158[9] , \Level2Out0[16] , 
        \Level1Out178[1] , \ScanLink197[0] , \Level2Out24[28] , 
        \Level2Out72[30] , \Level2Load170[0] , \Level2Out72[29] , 
        \Level4Out120[2] , \ScanLink182[29] , \ScanLink225[3] , 
        \Level2Out24[31] , \ScanLink78[7] , \ScanLink145[6] , 
        \ScanLink182[30] , \Level4Out240[7] , \Level1Out218[4] , 
        \ScanLink226[0] , \Level16Out128[0] , \Level8Out56[23] , 
        \ScanLink146[5] , \ScanLink179[31] , \ScanLink179[28] , 
        \ScanLink65[8] , \Level1Out83[22] , \Level1Out169[30] , 
        \Level2Out114[1] , \Level2Out170[18] , \Level1Out169[29] , 
        \Level2Out126[19] , \Level16Out48[5] , \Level1Out96[16] , 
        \Level1Load161[0] , \ScanLink194[3] , \Level1Out206[8] , 
        \Level8Out40[0] , \ScanLink8[12] , \Level1Out18[14] , \Level1Out43[5] , 
        \ScanLink59[30] , \Level4Out144[6] , \ScanLink59[29] , 
        \ScanLink241[7] , \ScanLink121[2] , \ScanLink211[18] , 
        \ScanLink232[30] , \Level4Out224[3] , \ScanLink232[29] , 
        \Level1Out201[19] , \Level1Out222[31] , \ScanLink247[19] , 
        \Level4Out196[0] , \Level1Out222[28] , \Level2Out218[31] , 
        \Level2Out0[25] , \Level2Out218[28] , \Level1Out78[10] , 
        \Level1Out91[3] , \Level1Out96[25] , \Level2Out170[5] , 
        \Level1Out102[9] , \ScanLink11[10] , \ScanLink27[15] , 
        \Level1Out40[6] , \ScanLink81[19] , \Level1Out83[11] , 
        \Level1Out92[0] , \Level2Out210[0] , \Level8Out24[4] , 
        \ScanLink242[4] , \Level4Out8[19] , \Level2Out34[9] , \ScanLink52[25] , 
        \ScanLink71[14] , \ScanLink122[1] , \ScanLink189[16] , 
        \Level8Out56[10] , \Level1Out163[0] , \ScanLink60[5] , 
        \ScanLink32[21] , \ScanLink47[11] , \ScanLink64[20] , 
        \Level1Out203[5] , \ScanLink239[25] , \Level1Out13[18] , 
        \Level1Out30[30] , \Level1Out30[29] , \Level1Out45[19] , 
        \Level1Out66[31] , \Level1Out66[28] , \Level2Out230[15] , 
        \Level1Out229[24] , \Level4Out184[24] , \ScanLink63[6] , 
        \Level1Out102[12] , \ScanLink143[8] , \Level1Out199[17] , 
        \Level1Out249[20] , \Level4Out92[17] , \Level2Out180[26] , 
        \Level2Out206[10] , \Level2Out250[11] , \Level1Out117[26] , 
        \Level1Out121[23] , \Level1Out177[22] , \Level16Out16[19] , 
        \Level2Out138[12] , \Level1Out134[17] , \Level1Out154[13] , 
        \Level16Out224[24] , \Level2Out56[3] , \Level1Out141[27] , 
        \ScanLink124[16] , \Level1Out162[16] , \Level2Out158[16] , 
        \Level32Out224[11] , \ScanLink151[26] , \Level8Out48[28] , 
        \ScanLink107[27] , \ScanLink112[13] , \Level1Out160[3] , 
        \ScanLink172[17] , \Level8Out48[31] , \Level2Out84[5] , 
        \ScanLink167[23] , \Level2Out82[17] , \Level4Load128[0] , 
        \ScanLink131[22] , \ScanLink144[12] , \Level1Out200[6] , 
        \Level1Out249[13] , \Level2Out168[7] , \Level2Out206[23] , 
        \Level4Out92[24] , \Level1Out0[24] , \Level1Out0[17] , \ScanLink9[18] , 
        \ScanLink11[23] , \ScanLink32[12] , \Level1Out199[24] , 
        \Level1Out229[17] , \ScanLink247[9] , \Level2Out180[15] , 
        \Level2Out208[2] , \Level2Out230[26] , \Level2Out250[22] , 
        \Level4Out184[17] , \ScanLink47[22] , \ScanLink27[26] , 
        \Level1Out58[4] , \ScanLink64[13] , \Level1Out107[4] , 
        \ScanLink189[25] , \ScanLink239[16] , \ScanLink71[27] , 
        \Level1Out46[8] , \ScanLink52[16] , \Level1Out102[21] , 
        \Level1Out104[7] , \ScanLink167[10] , \ScanLink107[14] , 
        \ScanLink112[20] , \ScanLink124[25] , \ScanLink131[11] , 
        \ScanLink144[21] , \Level2Out82[24] , \ScanLink139[0] , 
        \ScanLink151[15] , \ScanLink172[24] , \Level1Out117[15] , 
        \Level1Out119[8] , \Level1Out141[14] , \Level1Out134[24] , 
        \Level1Out162[25] , \Level32Out224[22] , \Level2Out158[25] , 
        \Level1Out177[11] , \Level2Out138[21] , \Level1Out121[10] , 
        \Level1Out154[20] , \Level2Out32[7] , \Level16Out224[17] , 
        \ScanLink80[13] , \Level1Out89[1] , \ScanLink178[11] , 
        \ScanLink95[27] , \ScanLink118[15] , \Level2Out24[3] , 
        \Level2Out88[11] , \Level1Out112[3] , \Level2Out164[15] , 
        \Level4Out156[12] , \Level4Out20[25] , \ScanLink11[6] , 
        \Level1Out108[14] , \Level2Out132[14] , \Level4Out76[24] , 
        \ScanLink12[5] , \Level1Out168[10] , \Level2Out4[1] , 
        \Level2Out152[10] , \Level4Out100[13] , \Level4Out160[17] , 
        \Level1Out186[25] , \Level2Out104[11] , \Level4Out16[20] , 
        \Level4Out40[21] , \Level4Out136[16] , \Level1Out223[22] , 
        \Level1Out81[9] , \Level1Out111[0] , \Level1Out200[13] , 
        \Level4Out208[14] , \Level1Out215[27] , \Level1Out193[11] , 
        \Level1Out236[16] , \Level1Out243[26] , \Level1Out5[6] , 
        \Level1Out29[7] , \ScanLink38[27] , \ScanLink58[23] , 
        \ScanLink205[26] , \Level2Out30[25] , \ScanLink183[10] , 
        \ScanLink226[17] , \ScanLink196[24] , \ScanLink253[27] , 
        \Level2Out66[24] , \Level8Out0[22] , \ScanLink210[12] , 
        \ScanLink233[23] , \ScanLink246[13] , \ScanLink75[2] , 
        \Level1Out82[28] , \ScanLink131[8] , \Level2Out50[21] , 
        \Level1Out168[23] , \Level4Out16[13] , \Level4Out160[24] , 
        \Level1Out82[31] , \Level2Out104[22] , \Level2Out152[23] , 
        \Level4Out68[6] , \Level4Out136[25] , \Level1Out176[7] , 
        \Level4Out40[12] , \Level2Out92[1] , \Level2Out164[26] , 
        \Level4Out20[16] , \Level4Out156[21] , \Level1Out34[8] , 
        \ScanLink80[20] , \ScanLink95[14] , \Level1Out108[27] , 
        \ScanLink184[9] , \Level2Out132[27] , \Level4Out100[20] , 
        \Level1Out216[2] , \Level4Out76[17] , \Level128Out128[0] , 
        \ScanLink118[26] , \ScanLink178[22] , \Level2Out88[22] , 
        \Level2Out40[7] , \Level1Out6[5] , \ScanLink38[14] , \ScanLink196[17] , 
        \ScanLink199[6] , \ScanLink246[20] , \ScanLink233[10] , 
        \ScanLink235[9] , \ScanLink210[21] , \Level2Out50[12] , 
        \Level32Out160[4] , \ScanLink58[10] , \ScanLink205[15] , 
        \Level2Out30[16] , \Level1Out79[30] , \Level1Out175[4] , 
        \ScanLink183[23] , \ScanLink226[24] , \ScanLink253[14] , 
        \Level2Out66[17] , \Level8Out0[11] , \Level1Out215[14] , 
        \ScanLink228[6] , \Level1Out243[15] , \ScanLink2[27] , \ScanLink76[1] , 
        \Level1Out79[29] , \Level1Out89[24] , \ScanLink148[3] , 
        \Level1Out186[16] , \Level1Out193[22] , \Level1Out236[25] , 
        \Level1Out223[11] , \Level1Out200[20] , \Level1Out215[1] , 
        \Level4Out208[27] , \Level1Out109[2] , \ScanLink254[0] , 
        \Level4Out148[19] , \ScanLink2[14] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink17[8] , \Level1Out56[2] , \ScanLink134[5] , 
        \Level8Out112[24] , \Level8Out144[25] , \Level2Out166[1] , 
        \Level1Out84[4] , \Level1Load113[0] , \Level2Out206[4] , 
        \Level8Out32[0] , \ScanLink46[31] , \Level4Out180[4] , 
        \ScanLink65[19] , \Level1Out12[21] , \Level1Out24[24] , 
        \ScanLink33[18] , \ScanLink46[28] , \Level1Out87[7] , 
        \Level16Out224[9] , \Level2Out224[18] , \Level4Out152[2] , 
        \Level1Out51[14] , \Level1Out72[25] , \Level1Out248[19] , 
        \Level32Out96[22] , \Level2Load102[0] , \Level1Out31[10] , 
        \Level1Out67[11] , \Level4Out232[7] , \Level64Out192[25] , 
        \ScanLink137[6] , \Level4Out0[7] , \Level1Out44[20] , 
        \Level2Out218[8] , \Level1Out55[1] , \ScanLink113[19] , 
        \ScanLink130[28] , \Level1Out170[9] , \Level2Out96[29] , 
        \Level2Out96[30] , \Level2Out102[5] , \ScanLink145[18] , 
        \ScanLink182[7] , \Level8Out56[4] , \ScanLink166[30] , 
        \Level1Out120[29] , \ScanLink130[31] , \ScanLink166[29] , 
        \Level1Out155[19] , \Level8Out112[17] , \Level1Out176[31] , 
        \ScanLink230[4] , \Level1Out3[8] , \Level1Out103[18] , 
        \Level1Out120[30] , \Level1Out176[28] , \Level8Out144[16] , 
        \ScanLink6[25] , \Level1Out12[12] , \Level1Out32[6] , 
        \Level1Out89[17] , \ScanLink150[1] , \Level2Out46[9] , 
        \Level1Out67[22] , \Level1Out15[3] , \Level1Out16[23] , 
        \Level1Out24[17] , \Level1Out31[23] , \Level1Out44[13] , 
        \Level4Out220[29] , \Level64Out192[16] , \Level2Out194[18] , 
        \Level4Out136[6] , \Level4Out220[30] , \Level1Out31[5] , 
        \Level1Out51[27] , \ScanLink233[7] , \Level32Out96[11] , 
        \Level1Out72[16] , \ScanLink153[2] , \ScanLink181[4] , 
        \Level2Out18[18] , \Level8Out48[8] , \Level2Out58[5] , 
        \Level2Out190[30] , \Level4Out224[18] , \Level1Out35[12] , 
        \Level1Out63[13] , \ScanLink177[4] , \Level1Out189[18] , 
        \Level1Out40[22] , \Level2Out190[29] , \Level8Out248[20] , 
        \Level1Out20[26] , \Level1Load37[0] , \ScanLink49[6] , 
        \Level1Out55[16] , \ScanLink217[1] , \Level4Out112[0] , 
        \Level1Out76[27] , \Level1Out198[5] , \Level1Out237[9] , 
        \Level64Out64[12] , \ScanLink199[19] , \Level8Out80[17] , 
        \ScanLink54[9] , \ScanLink98[3] , \ScanLink117[31] , \ScanLink134[19] , 
        \ScanLink141[29] , \ScanLink169[8] , \Level2Out92[18] , 
        \Level2Out246[6] , \Level8Out72[2] , \Level2Out126[3] , 
        \ScanLink117[28] , \ScanLink141[30] , \ScanLink162[18] , 
        \Level1Out151[28] , \ScanLink14[18] , \Level1Out16[0] , 
        \Level1Out124[18] , \ScanLink37[30] , \ScanLink61[28] , 
        \Level1Out98[12] , \Level1Out107[30] , \Level1Out172[19] , 
        \Level1Out107[29] , \Level1Out151[31] , \ScanLink174[7] , 
        \Level2Out148[19] , \Level1Out149[0] , \Level1Out229[5] , 
        \Level8Out120[23] , \Level8Out176[22] , \Level1Out186[9] , 
        \ScanLink214[2] , \Level2Out18[7] , \Level8Out80[24] , 
        \ScanLink37[29] , \ScanLink42[19] , \ScanLink61[31] , 
        \Level1Load254[0] , \Level1Out1[23] , \Level1Out1[10] , 
        \Level1Out4[26] , \Level1Out4[15] , \ScanLink6[16] , \Level1Out16[10] , 
        \Level1Out20[15] , \Level1Out55[25] , \Level1Out133[8] , 
        \ScanLink229[19] , \Level64Out64[21] , \Level1Out71[7] , 
        \Level1Out63[20] , \Level1Out76[14] , \Level2Out220[29] , 
        \ScanLink113[0] , \Level1Out239[18] , \Level4Out216[1] , 
        \Level2Out220[30] , \Level1Out35[21] , \Level1Out40[11] , 
        \Level4Out176[4] , \Level1Out72[4] , \ScanLink110[3] , 
        \Level8Out120[10] , \Level8Out248[13] , \Level8Out176[11] , 
        \ScanLink29[11] , \ScanLink49[15] , \Level1Out98[21] , 
        \Level2Out190[1] , \ScanLink192[26] , \Level2Out142[7] , 
        \Level2Out222[2] , \Level8Out16[6] , \Level4Out168[8] , 
        \ScanLink237[21] , \ScanLink242[11] , \Level32Out224[7] , 
        \ScanLink80[1] , \ScanLink201[24] , \ScanLink214[10] , 
        \Level2Out54[23] , \Level2Out34[27] , \Level1Out183[4] , 
        \ScanLink187[12] , \ScanLink222[15] , \Level1Out197[13] , 
        \Level1Out211[25] , \Level2Out62[26] , \Level1Out232[14] , 
        \Level1Out231[7] , \Level2Out208[14] , \ScanLink51[4] , 
        \ScanLink52[7] , \Level1Out182[27] , \Level1Out247[24] , 
        \Level1Out227[20] , \Level1Out252[10] , \Level1Out86[19] , 
        \Level1Out119[22] , \Level1Out151[2] , \Level1Out204[11] , 
        \Level2Out156[12] , \Level4Out164[15] , \Level1Out152[1] , 
        \Level1Out232[4] , \Level2Out100[13] , \Level2Out240[8] , 
        \Level4Out12[22] , \Level4Out44[23] , \Level2Out160[17] , 
        \Level4Out132[14] , \Level4Out24[27] , \Level4Out152[10] , 
        \Level1Out179[26] , \Level2Out136[16] , \Level4Out72[26] , 
        \Level8Out168[29] , \ScanLink83[2] , \ScanLink84[11] , 
        \ScanLink91[25] , \ScanLink172[9] , \Level4Out104[11] , 
        \Level8Out168[30] , \Level64Out0[16] , \Level2Out64[1] , 
        \ScanLink109[23] , \ScanLink169[27] , \Level1Out180[7] , 
        \ScanLink108[1] , \Level1Out182[14] , \Level1Out252[23] , 
        \Level1Out227[13] , \Level1Out135[6] , \Level1Out204[22] , 
        \Level1Out255[3] , \Level64Load192[0] , \Level1Out211[16] , 
        \Level2Out188[3] , \Level1Out18[19] , \ScanLink29[22] , 
        \ScanLink36[3] , \Level1Out247[17] , \Level2Out208[27] , 
        \Level1Out197[20] , \Level1Out232[27] , \Level8Out200[19] , 
        \ScanLink35[0] , \ScanLink49[26] , \Level1Out77[9] , \ScanLink201[17] , 
        \Level2Out34[14] , \Level2Out62[15] , \Level1Out128[9] , 
        \ScanLink187[21] , \ScanLink222[26] , \ScanLink242[22] , 
        \Level4Out36[8] , \ScanLink192[15] , \ScanLink237[12] , 
        \Level2Out54[10] , \Level1Out69[5] , \ScanLink84[22] , 
        \ScanLink214[23] , \ScanLink91[16] , \ScanLink109[10] , 
        \Level64Out0[25] , \ScanLink169[14] , \Level2Out160[24] , 
        \Level4Out24[14] , \Level4Out152[23] , \Level1Load99[0] , 
        \Level1Out179[15] , \Level2Out136[25] , \Level4Out104[22] , 
        \Level2Out144[9] , \Level4Out72[15] , \Level1Out119[11] , 
        \Level4Out12[11] , \ScanLink81[14] , \Level1Out136[5] , 
        \Level2Out100[20] , \Level2Out156[21] , \Level4Out164[26] , 
        \Level4Out132[27] , \Level4Out28[4] , \ScanLink179[16] , 
        \Level4Out44[10] , \Level4Out188[1] , \ScanLink94[20] , 
        \ScanLink119[12] , \ScanLink242[9] , \Level2Out34[4] , 
        \Level4Out8[14] , \Level1Out96[31] , \Level1Out102[4] , 
        \Level2Out110[22] , \Level1Out96[28] , \Level1Out109[13] , 
        \Level2Out146[23] , \Level2Out170[8] , \Level1Out169[17] , 
        \Level1Out187[22] , \Level1Out222[25] , \Level2Out126[27] , 
        \Level2Out170[26] , \Level4Out8[2] , \Level8Out24[9] , 
        \Level1Out101[7] , \Level1Out201[14] , \Level2Out0[28] , 
        \Level2Out218[25] , \Level2Out0[31] , \Level1Out192[16] , 
        \Level1Out214[20] , \Level1Out237[11] , \Level1Load18[0] , 
        \ScanLink39[20] , \Level1Out43[8] , \ScanLink59[24] , 
        \ScanLink204[21] , \Level1Out242[21] , \ScanLink182[17] , 
        \Level2Out12[13] , \Level2Out44[12] , \ScanLink197[23] , 
        \ScanLink227[10] , \ScanLink232[24] , \ScanLink252[20] , 
        \ScanLink247[14] , \Level2Out72[17] , \ScanLink211[15] , 
        \Level16Out32[0] , \Level2Out24[16] , \ScanLink39[13] , 
        \Level1Out39[0] , \ScanLink65[5] , \Level1Out169[24] , 
        \Level2Out126[14] , \Level1Out166[0] , \Level2Load74[0] , 
        \Level2Out170[15] , \Level2Out82[6] , \Level2Out110[11] , 
        \ScanLink81[27] , \ScanLink94[13] , \Level1Out109[20] , 
        \Level2Out146[10] , \Level16Out48[8] , \Level1Out206[5] , 
        \ScanLink119[21] , \ScanLink179[25] , \Level2Out50[0] , 
        \ScanLink146[8] , \ScanLink189[1] , \Level4Out8[27] , 
        \ScanLink197[10] , \ScanLink232[17] , \ScanLink247[27] , 
        \Level2Out72[24] , \ScanLink59[17] , \ScanLink204[12] , 
        \ScanLink211[26] , \Level2Out24[25] , \Level2Out44[21] , 
        \Level1Out218[9] , \Level1Out165[3] , \ScanLink182[24] , 
        \ScanLink252[13] , \Level2Out12[20] , \ScanLink227[23] , 
        \Level2Load6[0] , \Level1Out214[13] , \ScanLink238[1] , 
        \ScanLink3[20] , \ScanLink66[6] , \Level1Out242[12] , 
        \Level1Out88[23] , \ScanLink158[4] , \Level1Out187[11] , 
        \Level1Out192[25] , \Level1Out222[16] , \Level1Out237[22] , 
        \Level2Out218[16] , \Level1Out162[28] , \Level1Out201[27] , 
        \Level1Out205[6] , \Level1Out117[18] , \Level1Out119[5] , 
        \Level1Out134[30] , \Level1Out141[19] , \Level2Out158[28] , 
        \Level1Out162[31] , \Level1Out134[29] , \ScanLink244[7] , 
        \Level2Out158[31] , \Level1Out13[26] , \ScanLink19[3] , 
        \Level1Out25[23] , \Level1Out46[5] , \Level1Out58[9] , 
        \Level1Out94[3] , \ScanLink107[19] , \ScanLink124[2] , 
        \ScanLink172[29] , \Level2Out82[30] , \Level2Out176[6] , 
        \Level16Out16[27] , \Level2Out82[29] , \Level16Out0[22] , 
        \Level2Out216[3] , \ScanLink124[31] , \Level1Out97[0] , 
        \Level1Out107[9] , \ScanLink124[28] , \ScanLink151[18] , 
        \ScanLink172[30] , \Level8Out48[16] , \ScanLink189[31] , 
        \ScanLink189[28] , \Level2Out180[18] , \Level4Out92[30] , 
        \Level1Out50[13] , \ScanLink247[4] , \Level1Out73[22] , 
        \Level1Out199[30] , \Level4Out92[29] , \Level4Load232[0] , 
        \Level1Out199[29] , \Level1Out30[17] , \Level1Out66[16] , 
        \ScanLink127[1] , \Level1Out45[27] , \Level1Out45[6] , 
        \ScanLink192[0] , \Level2Out112[2] , \Level8Out48[25] , 
        \Level2Out84[8] , \Level16Out0[11] , \ScanLink3[13] , \ScanLink220[3] , 
        \Level16Out224[29] , \ScanLink5[2] , \Level1Out13[15] , 
        \Level1Out22[1] , \Level1Out88[10] , \Level16Out16[14] , 
        \Level16Out224[30] , \ScanLink140[6] , \Level1Out66[25] , 
        \Level1Out229[29] , \Level4Out184[29] , \Level1Out17[24] , 
        \Level1Out21[2] , \Level1Out30[24] , \Level1Out45[14] , 
        \Level1Out229[30] , \Level2Out230[18] , \Level4Out60[3] , 
        \Level4Out184[30] , \Level1Out50[20] , \ScanLink223[0] , 
        \Level1Out25[10] , \ScanLink27[18] , \ScanLink52[28] , 
        \Level1Out73[11] , \ScanLink143[5] , \Level32Out0[3] , \ScanLink60[8] , 
        \ScanLink52[31] , \ScanLink71[19] , \Level1Load164[0] , 
        \Level2Out48[2] , \ScanLink191[3] , \Level1Out203[8] , 
        \ScanLink239[31] , \ScanLink239[28] , \Level2Out234[30] , 
        \Level1Out21[21] , \Level1Out34[15] , \Level1Out62[14] , 
        \Level4Out180[18] , \ScanLink167[3] , \Level1Load192[0] , 
        \Level1Out41[25] , \Level2Load232[0] , \Level2Out234[29] , 
        \Level4Out44[5] , \ScanLink23[30] , \ScanLink23[29] , 
        \Level1Out54[11] , \ScanLink207[6] , \ScanLink59[1] , \ScanLink96[8] , 
        \Level2Out128[8] , \Level1Out77[20] , \ScanLink56[19] , 
        \ScanLink75[31] , \ScanLink75[28] , \Level4Out96[3] , \Level1Out5[21] , 
        \Level1Out5[12] , \ScanLink6[1] , \ScanLink88[4] , \Level1Out188[2] , 
        \ScanLink248[29] , \Level1Load223[0] , \ScanLink248[30] , 
        \Level2Out136[4] , \ScanLink7[22] , \Level1Out144[8] , 
        \Level2Out72[8] , \ScanLink7[11] , \Level1Out17[17] , 
        \Level1Out21[12] , \Level1Out54[22] , \Level1Out99[15] , 
        \Level1Out159[7] , \ScanLink164[0] , \Level1Out239[2] , 
        \ScanLink204[5] , \Level1Out61[0] , \Level32Out128[19] , 
        \Level1Out62[27] , \Level1Out77[13] , \Level2Out184[29] , 
        \ScanLink103[7] , \Level2Out184[30] , \Level4Out96[18] , 
        \Level1Out34[26] , \Level1Out41[16] , \Level4Out20[1] , 
        \Level1Out62[3] , \ScanLink100[4] , \Level1Out113[29] , 
        \Level1Out145[31] , \Level1Out166[19] , \Level1Out113[30] , 
        \Level1Out130[18] , \Level1Out145[28] , \ScanLink23[9] , 
        \Level1Load40[0] , \Level1Out99[26] , \Level2Out180[6] , 
        \ScanLink103[31] , \ScanLink103[28] , \Level1Out240[9] , 
        \Level2Out86[18] , \Level2Out232[5] , \ScanLink120[19] , 
        \ScanLink155[30] , \ScanLink176[18] , \Level2Out152[0] , 
        \ScanLink155[29] , \Level32Out128[3] , \ScanLink28[16] , 
        \ScanLink48[12] , \ScanLink193[21] , \ScanLink236[26] , 
        \ScanLink243[16] , \Level2Out76[15] , \ScanLink90[6] , 
        \ScanLink200[23] , \ScanLink215[17] , \Level2Out20[14] , 
        \Level2Out40[10] , \ScanLink186[15] , \Level1Out193[3] , 
        \ScanLink223[12] , \Level2Out16[11] , \Level4Out104[9] , 
        \Level1Out196[14] , \ScanLink201[8] , \Level1Out210[22] , 
        \ScanLink256[22] , \Level16Out160[15] , \Level1Out221[0] , 
        \Level1Out233[13] , \Level1Out246[23] , \ScanLink41[3] , 
        \ScanLink42[0] , \Level1Out183[20] , \Level1Out226[27] , 
        \Level32Out160[20] , \Level1Out253[17] , \Level4Out88[20] , 
        \Level1Out118[25] , \Level1Out141[5] , \Level1Out205[16] , 
        \Level16Out112[7] , \Level1Out142[6] , \Level1Out222[3] , 
        \Level2Out122[25] , \Level2Out174[24] , \Level8Load88[0] , 
        \Level1Out178[21] , \Level2Out114[20] , \Level2Out142[21] , 
        \Level16Out208[16] , \Level1Out69[18] , \ScanLink85[16] , 
        \ScanLink90[22] , \Level2Out74[6] , \ScanLink108[24] , 
        \ScanLink168[20] , \Level1Out190[0] , \Level2Out98[20] , 
        \Level2Load82[0] , \ScanLink93[5] , \Level1Out253[24] , 
        \Level2Out4[19] , \Level4Out88[13] , \ScanLink118[6] , 
        \Level1Out183[13] , \Level1Out226[14] , \Level32Out160[13] , 
        \Level1Out125[1] , \Level1Out205[25] , \Level1Out245[4] , 
        \Level16Out176[3] , \Level1Out210[11] , \Level1Out246[10] , 
        \Level2Out198[4] , \Level16Out160[26] , \ScanLink14[15] , 
        \Level1Out20[18] , \ScanLink25[7] , \ScanLink26[4] , \ScanLink28[25] , 
        \Level1Out196[27] , \Level1Out233[20] , \Level2Out40[23] , 
        \ScanLink38[8] , \ScanLink48[21] , \ScanLink105[9] , \Level4Out200[8] , 
        \Level16Out16[6] , \ScanLink186[26] , \ScanLink200[10] , 
        \ScanLink256[11] , \Level8Out192[4] , \ScanLink193[12] , 
        \ScanLink223[21] , \ScanLink236[15] , \ScanLink243[25] , 
        \Level2Out16[22] , \Level2Out76[26] , \ScanLink85[25] , 
        \ScanLink215[24] , \Level2Out20[27] , \Level2Out10[2] , 
        \ScanLink108[17] , \Level8Out64[29] , \Level2Out98[13] , 
        \Level2Out186[8] , \Level8Out32[31] , \Level8Out32[28] , 
        \Level8Out64[30] , \Level1Out79[2] , \ScanLink90[11] , 
        \ScanLink168[13] , \Level2Out114[13] , \Level1Out92[19] , 
        \Level1Out178[12] , \Level1Out118[16] , \Level1Out246[7] , 
        \Level2Out142[12] , \Level16Out208[25] , \Level2Out122[16] , 
        \ScanLink33[3] , \ScanLink117[16] , \Level1Out126[2] , 
        \Level2Out174[17] , \ScanLink121[13] , \ScanLink134[27] , 
        \ScanLink162[26] , \Level4Out208[0] , \ScanLink141[17] , 
        \Level1Out250[3] , \ScanLink154[23] , \Level1Out55[31] , 
        \Level1Out72[9] , \ScanLink102[22] , \Level1Out130[6] , 
        \ScanLink177[12] , \Level2Out92[26] , \Level64Out192[1] , 
        \Level4Out168[5] , \Level1Out131[12] , \Level1Out107[17] , 
        \Level1Out112[23] , \Level1Out144[22] , \Level1Out167[13] , 
        \Level2Out128[23] , \Level2Out148[27] , \Level1Out124[26] , 
        \Level1Out172[27] , \Level1Out151[16] , \Level1Out55[28] , 
        \Level1Out76[19] , \Level1Out239[15] , \Level4Out244[22] , 
        \Level8Out184[0] , \Level2Out220[24] , \ScanLink37[24] , 
        \ScanLink42[14] , \Level1Out189[26] , \Level2Out190[17] , 
        \Level2Out240[20] , \Level4Out212[23] , \Level4Out176[9] , 
        \Level2Out216[21] , \Level4Out224[26] , \Level8Out80[30] , 
        \ScanLink61[25] , \Level1Out253[0] , \Level8Out80[29] , 
        \ScanLink199[27] , \ScanLink74[11] , \ScanLink229[14] , 
        \ScanLink249[10] , \Level16Out160[7] , \Level1Out133[5] , 
        \Level1Out0[30] , \Level1Out0[29] , \Level1Out4[18] , \ScanLink6[31] , 
        \ScanLink22[10] , \ScanLink30[0] , \ScanLink57[20] , 
        \Level1Out172[14] , \ScanLink6[28] , \Level1Out107[24] , 
        \Level1Out151[25] , \Level1Out229[8] , \Level2Out148[14] , 
        \Level2Out62[2] , \ScanLink8[7] , \ScanLink14[26] , \ScanLink22[23] , 
        \ScanLink57[7] , \ScanLink85[1] , \Level1Out112[10] , 
        \Level1Out124[15] , \Level1Out131[21] , \Level1Out144[11] , 
        \Level1Out167[20] , \Level1Out186[4] , \Level2Out128[10] , 
        \ScanLink102[11] , \ScanLink121[20] , \ScanLink154[10] , 
        \ScanLink169[5] , \ScanLink177[21] , \Level1Out234[7] , 
        \ScanLink117[25] , \Level1Out154[2] , \ScanLink162[15] , 
        \Level2Out92[15] , \ScanLink141[24] , \ScanLink209[0] , 
        \ScanLink74[22] , \ScanLink134[14] , \ScanLink229[27] , 
        \ScanLink37[17] , \ScanLink57[13] , \Level1Out237[4] , 
        \ScanLink42[27] , \ScanLink54[4] , \ScanLink61[16] , \ScanLink249[23] , 
        \ScanLink86[2] , \Level1Out157[1] , \Level1Out198[8] , 
        \ScanLink177[9] , \Level1Out189[15] , \ScanLink199[14] , 
        \Level2Out190[24] , \Level2Out216[12] , \Level2Out240[13] , 
        \Level4Out224[15] , \Level16Out64[6] , \Level2Out138[2] , 
        \Level1Out239[26] , \Level4Out244[11] , \Level4Out212[10] , 
        \Level1Out10[3] , \ScanLink28[2] , \Level1Out69[8] , \Level1Out93[13] , 
        \Level1Out185[7] , \Level2Out220[17] , \Level2Out136[28] , 
        \Level1Out179[18] , \Level2Out136[31] , \Level2Out160[30] , 
        \Level4Out72[18] , \Level4Out24[19] , \Level2Out160[29] , 
        \Level2Out224[1] , \Level8Out168[17] , \Level1Out74[7] , 
        \Level1Out86[27] , \Level1Out136[8] , \Level4Out28[9] , 
        \Level1Load251[0] , \Level2Out144[4] , \ScanLink116[0] , 
        \ScanLink169[19] , \Level2Out196[2] , \Level64Out0[31] , 
        \Level1Out68[12] , \Level1Out77[4] , \Level2Out62[18] , 
        \Level64Out0[28] , \ScanLink115[3] , \Level2Out34[19] , 
        \Level2Load240[0] , \Level1Out128[4] , \Level1Out248[1] , 
        \Level4Out36[5] , \Level1Out182[19] , \ScanLink192[18] , 
        \Level8Out200[14] , \Level16Out96[12] , \Level32Out96[0] , 
        \Level1Load32[0] , \Level1Out86[14] , \ScanLink91[31] , 
        \ScanLink91[28] , \ScanLink172[4] , \ScanLink212[1] , 
        \Level1Out232[9] , \Level2Out240[5] , \Level4Out132[19] , 
        \Level4Out164[18] , \ScanLink51[9] , \Level1Out93[20] , 
        \Level2Out120[0] , \Level1Out211[31] , \Level8Out168[24] , 
        \Level8Out200[27] , \Level1Out232[19] , \Level1Out13[0] , 
        \ScanLink49[18] , \Level1Out68[21] , \Level1Out211[28] , 
        \Level1Out247[29] , \Level2Out208[19] , \Level1Out247[30] , 
        \Level4Out80[7] , \Level16Out96[21] , \ScanLink171[7] , 
        \Level1Out183[9] , \ScanLink201[30] , \ScanLink211[2] , 
        \ScanLink222[18] , \Level4Out52[1] , \ScanLink201[29] , 
        \Level1Out243[18] , \Level1Out79[24] , \Level1Out236[28] , 
        \Level1Out0[6] , \Level1Out6[8] , \Level1Out19[20] , \Level1Out175[9] , 
        \Level1Out215[19] , \Level1Out236[31] , \Level8Out232[13] , 
        \Level1Out37[6] , \ScanLink38[19] , \ScanLink187[7] , 
        \Level1Out168[6] , \Level4Out76[7] , \Level4Load240[0] , 
        \Level32Out160[9] , \ScanLink226[29] , \ScanLink235[4] , 
        \ScanLink253[19] , \ScanLink9[26] , \Level1Out34[5] , \ScanLink68[0] , 
        \ScanLink95[19] , \ScanLink155[1] , \ScanLink226[30] , 
        \ScanLink205[18] , \Level1Out208[3] , \ScanLink236[7] , 
        \ScanLink156[2] , \Level1Out82[25] , \Level2Out104[6] , 
        \Level4Out136[28] , \Level4Out160[30] , \Level1Out97[11] , 
        \Level4Out136[31] , \Level4Out160[29] , \ScanLink184[4] , 
        \ScanLink9[15] , \ScanLink12[8] , \Level1Out19[13] , \Level1Out53[2] , 
        \ScanLink131[5] , \ScanLink196[30] , \ScanLink251[0] , 
        \Level2Out30[31] , \Level2Out66[29] , \Level4Out12[3] , 
        \Level2Out30[28] , \Level2Out66[30] , \ScanLink196[29] , 
        \Level1Out186[31] , \Level1Out186[28] , \Level4Out208[19] , 
        \Level8Out232[20] , \Level1Out79[17] , \Level1Out81[4] , 
        \Level1Load116[0] , \Level1Out97[22] , \Level1Out108[19] , 
        \Level4Out76[29] , \Level2Out160[2] , \Level2Out132[19] , 
        \Level2Out164[18] , \Level4Out20[31] , \Level4Out20[28] , 
        \Level4Out76[30] , \ScanLink10[17] , \ScanLink26[12] , 
        \Level1Out50[1] , \Level1Out82[16] , \Level1Out82[7] , 
        \Level2Out200[7] , \ScanLink118[18] , \ScanLink252[3] , 
        \ScanLink53[22] , \ScanLink70[13] , \ScanLink132[6] , 
        \ScanLink188[11] , \Level2Out18[15] , \Level1Out173[7] , 
        \ScanLink70[2] , \ScanLink33[26] , \ScanLink46[16] , 
        \Level16Out240[0] , \ScanLink65[27] , \ScanLink181[9] , 
        \Level1Out213[2] , \Level2Out58[8] , \ScanLink238[22] , 
        \Level1Out198[10] , \Level1Load209[0] , \Level1Out228[23] , 
        \Level2Out78[11] , \Level2Out194[15] , \Level2Out244[22] , 
        \Level2Out212[23] , \Level4Out220[24] , \Level4Out240[20] , 
        \ScanLink2[19] , \Level1Out31[8] , \Level1Out248[27] , 
        \Level8Out48[5] , \Level1Out103[15] , \Level2Out224[26] , 
        \Level4Out216[21] , \Level1Out120[24] , \Level1Out176[25] , 
        \Level1Out155[14] , \ScanLink230[9] , \Level4Out128[23] , 
        \Level1Out3[5] , \Level1Out135[10] , \Level2Out46[4] , 
        \Level4Out148[27] , \Level1Out140[20] , \Level1Out4[22] , 
        \Level1Out4[11] , \ScanLink10[24] , \ScanLink14[6] , \Level1Out24[30] , 
        \ScanLink73[1] , \Level1Out116[21] , \ScanLink125[11] , 
        \Level1Out163[11] , \Level4Out68[11] , \ScanLink150[21] , 
        \Level2Out102[8] , \ScanLink106[20] , \Level2Out96[24] , 
        \ScanLink113[14] , \Level1Out170[4] , \ScanLink173[10] , 
        \Level4Out128[7] , \Level2Out94[2] , \ScanLink130[25] , 
        \ScanLink166[24] , \Level2Load218[0] , \Level4Out248[2] , 
        \ScanLink145[15] , \Level1Out210[1] , \Level8Out56[9] , 
        \Level2Out178[0] , \Level1Out24[29] , \Level1Out72[28] , 
        \Level1Out198[23] , \Level1Out248[14] , \Level4Out240[13] , 
        \Level4Out216[12] , \ScanLink33[15] , \Level1Out51[19] , 
        \Level1Out72[31] , \Level2Out224[15] , \Level1Out228[10] , 
        \Level2Out194[26] , \Level2Out212[10] , \Level2Out218[5] , 
        \Level64Out192[31] , \Level2Out244[11] , \Level4Out220[17] , 
        \Level64Out192[28] , \ScanLink46[25] , \Level4Out180[9] , 
        \ScanLink17[5] , \ScanLink26[21] , \Level1Out48[3] , \ScanLink65[14] , 
        \Level2Out78[22] , \Level16Out144[1] , \Level1Out117[3] , 
        \ScanLink188[22] , \ScanLink238[11] , \Level2Out18[26] , 
        \ScanLink70[20] , \Level16Out224[4] , \ScanLink53[11] , 
        \ScanLink113[27] , \Level1Out114[0] , \ScanLink166[17] , 
        \ScanLink249[2] , \ScanLink145[26] , \ScanLink51[0] , \ScanLink83[6] , 
        \Level1Out84[9] , \ScanLink106[13] , \ScanLink125[22] , 
        \ScanLink130[16] , \ScanLink150[12] , \Level2Out2[2] , 
        \ScanLink129[7] , \ScanLink173[23] , \Level2Out96[17] , 
        \Level2Out206[9] , \Level1Out89[30] , \Level1Out89[29] , 
        \Level1Out135[23] , \Level1Out140[13] , \Level4Out148[14] , 
        \Level1Out99[6] , \Level1Out103[26] , \Level1Out116[12] , 
        \Level1Out163[22] , \Level1Out176[16] , \Level4Out68[22] , 
        \Level8Out144[28] , \Level1Out120[17] , \ScanLink134[8] , 
        \Level1Out155[27] , \Level4Out128[10] , \Level8Out112[30] , 
        \Level2Out22[0] , \Level8Out144[31] , \Level8Out112[29] , 
        \ScanLink84[15] , \ScanLink109[27] , \Level1Out180[3] , 
        \ScanLink212[8] , \ScanLink91[21] , \Level2Out64[5] , 
        \ScanLink169[23] , \Level1Out179[22] , \Level2Out120[9] , 
        \Level4Out72[22] , \Level64Out0[12] , \Level2Out136[12] , 
        \Level4Out104[15] , \ScanLink52[3] , \Level1Out68[31] , 
        \Level1Out93[30] , \Level1Out93[29] , \Level1Out152[5] , 
        \Level2Out160[13] , \Level4Out152[14] , \Level4Out24[23] , 
        \Level1Out119[26] , \Level2Out100[17] , \Level4Out44[27] , 
        \Level2Out156[16] , \Level4Out132[10] , \Level1Out204[15] , 
        \Level1Out232[0] , \Level4Out12[26] , \Level4Out164[11] , 
        \Level1Out68[28] , \Level1Out151[6] , \Level16Out96[31] , 
        \Level1Out182[23] , \Level1Out227[24] , \Level1Out252[14] , 
        \Level16Out96[28] , \Level1Out197[17] , \Level1Out232[10] , 
        \Level1Out231[3] , \Level1Out247[20] , \Level2Out208[10] , 
        \Level1Out13[9] , \ScanLink29[15] , \ScanLink80[5] , \Level1Out183[0] , 
        \ScanLink187[16] , \Level1Out211[21] , \ScanLink222[11] , 
        \Level4Out52[8] , \ScanLink201[20] , \Level2Out34[23] , 
        \Level2Out62[22] , \ScanLink49[11] , \ScanLink192[22] , 
        \ScanLink214[14] , \Level2Out54[27] , \ScanLink237[25] , 
        \ScanLink242[15] , \Level32Out224[3] , \ScanLink29[26] , 
        \ScanLink35[4] , \Level1Out136[1] , \Level2Out100[24] , 
        \Level4Out28[0] , \Level4Out132[23] , \Level4Out44[14] , 
        \Level4Out12[15] , \ScanLink49[22] , \Level1Out69[1] , 
        \Level1Out119[15] , \Level1Out179[11] , \Level2Out156[25] , 
        \Level4Out164[22] , \Level2Out136[21] , \Level4Out104[26] , 
        \Level2Out160[20] , \Level2Out224[8] , \Level4Out24[10] , 
        \Level4Out72[11] , \Level4Out152[27] , \ScanLink84[26] , 
        \ScanLink91[12] , \ScanLink116[9] , \ScanLink169[10] , 
        \Level64Out0[21] , \ScanLink109[14] , \Level2Out54[14] , 
        \ScanLink187[25] , \ScanLink192[11] , \ScanLink214[27] , 
        \ScanLink242[26] , \ScanLink222[22] , \ScanLink237[16] , 
        \Level2Out62[11] , \ScanLink201[13] , \Level2Out34[10] , 
        \Level1Out247[13] , \Level1Out248[8] , \Level2Out188[7] , 
        \ScanLink6[21] , \ScanLink36[7] , \Level2Out208[23] , \ScanLink85[8] , 
        \ScanLink108[5] , \Level1Out135[2] , \Level1Out197[24] , 
        \Level1Out232[23] , \Level32Out96[9] , \Level1Out182[10] , 
        \Level1Out204[26] , \Level1Out211[12] , \Level1Out252[27] , 
        \Level1Out227[17] , \Level1Out112[19] , \Level1Out131[28] , 
        \Level1Out144[18] , \Level1Out255[7] , \Level8Out176[26] , 
        \Level1Out149[4] , \Level1Out167[30] , \ScanLink214[6] , 
        \Level1Out167[29] , \Level2Out128[19] , \Level8Out120[27] , 
        \Level1Out98[16] , \Level1Out131[31] , \ScanLink174[3] , 
        \Level1Load181[0] , \Level1Out229[1] , \ScanLink6[12] , 
        \Level1Out15[7] , \Level1Out16[4] , \Level1Out20[22] , \ScanLink49[2] , 
        \ScanLink98[7] , \ScanLink209[9] , \Level2Out126[7] , 
        \ScanLink102[18] , \ScanLink121[29] , \ScanLink154[19] , 
        \ScanLink177[31] , \ScanLink177[28] , \Level8Out72[6] , 
        \Level2Out246[2] , \ScanLink121[30] , \Level1Out157[8] , 
        \Level1Out198[1] , \Level1Load230[0] , \Level2Load190[0] , 
        \Level8Out80[13] , \Level4Out244[18] , \Level64Out64[16] , 
        \Level1Out76[23] , \Level4Out112[4] , \Level4Out212[19] , 
        \Level1Out35[16] , \Level1Out55[12] , \ScanLink217[5] , 
        \Level1Out40[26] , \Level8Out248[24] , \Level1Out16[27] , 
        \Level1Out63[17] , \Level1Out98[25] , \ScanLink177[0] , 
        \Level2Out142[3] , \Level2Out190[5] , \Level2Out222[6] , 
        \Level64Out192[8] , \Level4Out208[9] , \Level8Out16[2] , 
        \Level1Out16[14] , \Level1Out35[25] , \Level1Out40[15] , 
        \Level1Out72[0] , \Level8Out176[15] , \ScanLink110[7] , 
        \Level8Out120[14] , \Level2Out216[31] , \Level2Out240[29] , 
        \Level4Out176[0] , \Level1Out63[24] , \Level8Out248[17] , 
        \Level2Out240[30] , \Level1Out20[11] , \Level1Out55[21] , 
        \Level1Out76[10] , \Level2Out216[28] , \Level4Out216[5] , 
        \ScanLink113[4] , \Level8Out184[9] , \Level1Out71[3] , 
        \ScanLink57[30] , \ScanLink57[29] , \ScanLink74[18] , \Level1Out0[20] , 
        \Level1Out0[13] , \ScanLink2[23] , \Level1Out12[25] , \ScanLink22[19] , 
        \ScanLink30[9] , \Level1Load53[0] , \Level64Out64[25] , 
        \Level1Out31[14] , \ScanLink249[19] , \Level1Out253[9] , 
        \Level2Out18[3] , \Level8Out80[20] , \Level1Out44[24] , 
        \Level2Out244[18] , \Level4Out0[3] , \Level1Out55[5] , 
        \Level2Out212[19] , \Level4Out232[3] , \Level1Out24[20] , 
        \Level1Out67[15] , \Level64Out192[21] , \Level1Out72[21] , 
        \ScanLink137[2] , \Level1Out228[19] , \Level2Out178[9] , 
        \ScanLink26[31] , \Level1Out51[10] , \Level4Out152[6] , 
        \Level32Out96[26] , \ScanLink26[28] , \ScanLink70[29] , 
        \Level1Out87[3] , \ScanLink53[18] , \ScanLink70[30] , \Level1Out84[0] , 
        \ScanLink238[18] , \Level4Out180[0] , \Level16Out144[8] , 
        \Level2Out206[0] , \Level8Out32[4] , \Level1Out114[9] , 
        \ScanLink134[1] , \Level2Out166[5] , \Level8Out144[21] , 
        \Level2Out22[9] , \Level4Out128[19] , \ScanLink2[10] , 
        \Level1Out12[16] , \Level1Out24[13] , \Level1Out31[1] , 
        \Level1Out51[23] , \Level1Out56[6] , \Level1Out72[12] , 
        \Level1Out89[20] , \Level1Out109[6] , \Level8Out112[20] , 
        \ScanLink254[4] , \ScanLink181[0] , \Level8Load0[0] , 
        \Level16Out240[9] , \ScanLink188[18] , \Level2Out58[1] , 
        \Level2Out78[18] , \ScanLink153[6] , \Level1Out198[19] , 
        \Level4Out240[29] , \Level4Out216[31] , \Level4Out240[30] , 
        \Level32Out96[15] , \Level1Out31[27] , \Level1Out44[17] , 
        \Level4Out136[2] , \Level4Out216[28] , \Level1Out67[26] , 
        \ScanLink233[3] , \Level1Out32[2] , \Level1Out116[31] , 
        \Level1Out135[19] , \Level2Load166[0] , \Level64Out192[12] , 
        \Level1Out89[13] , \Level1Out116[28] , \Level1Out140[29] , 
        \Level4Out68[18] , \Level1Out163[18] , \Level1Out140[30] , 
        \ScanLink150[5] , \ScanLink230[0] , \Level8Out112[13] , 
        \Level8Out144[12] , \ScanLink38[23] , \ScanLink73[8] , 
        \ScanLink106[30] , \ScanLink125[18] , \Level1Load177[0] , 
        \ScanLink182[3] , \Level1Out210[8] , \Level2Out102[1] , 
        \Level8Out56[0] , \ScanLink150[28] , \ScanLink106[29] , 
        \ScanLink150[31] , \ScanLink173[19] , \ScanLink210[16] , 
        \ScanLink58[27] , \ScanLink183[14] , \ScanLink196[20] , 
        \Level2Out50[25] , \ScanLink226[13] , \ScanLink233[27] , 
        \ScanLink246[17] , \ScanLink205[22] , \ScanLink251[9] , 
        \ScanLink253[23] , \Level8Out0[26] , \Level2Out66[20] , 
        \Level2Out30[21] , \Level1Out193[15] , \Level1Out236[12] , 
        \ScanLink11[2] , \ScanLink12[1] , \Level1Out111[4] , 
        \Level1Out200[17] , \Level1Out215[23] , \Level1Out243[22] , 
        \Level4Out208[10] , \Level8Out232[29] , \Level1Out186[21] , 
        \Level1Out223[26] , \Level8Out232[30] , \Level1Out108[10] , 
        \Level1Out168[14] , \Level2Out4[5] , \Level2Out104[15] , 
        \Level4Out40[25] , \Level2Out152[14] , \Level4Out136[12] , 
        \Level4Out160[13] , \Level4Out16[24] , \Level2Out132[10] , 
        \Level4Out76[20] , \Level4Out100[17] , \Level1Out19[30] , 
        \Level1Out50[8] , \ScanLink95[23] , \Level1Out112[7] , 
        \Level2Out164[11] , \Level4Out20[21] , \Level4Out156[16] , 
        \ScanLink118[11] , \Level2Out24[7] , \Level2Out88[15] , 
        \ScanLink80[17] , \ScanLink178[15] , \Level4Out208[23] , 
        \Level1Out19[29] , \Level1Out200[24] , \ScanLink148[7] , 
        \Level1Out186[12] , \Level1Out223[15] , \Level1Out215[5] , 
        \Level1Out5[2] , \Level1Out6[1] , \ScanLink76[5] , \Level1Out243[11] , 
        \Level1Out175[0] , \Level1Out193[26] , \Level1Out236[21] , 
        \ScanLink183[27] , \Level1Out215[10] , \ScanLink226[20] , 
        \ScanLink228[2] , \ScanLink253[10] , \Level2Out66[13] , 
        \Level8Out0[15] , \ScanLink38[10] , \ScanLink58[14] , \ScanLink155[8] , 
        \ScanLink205[11] , \Level2Out30[12] , \ScanLink196[13] , 
        \ScanLink210[25] , \Level2Out50[16] , \Level32Out160[0] , 
        \ScanLink246[24] , \ScanLink233[14] , \Level1Out22[8] , 
        \Level1Out29[3] , \ScanLink68[9] , \ScanLink80[24] , \ScanLink178[26] , 
        \ScanLink199[2] , \ScanLink95[10] , \Level2Out40[3] , 
        \ScanLink118[22] , \Level2Out88[26] , \Level128Out128[4] , 
        \Level1Out97[18] , \Level1Out108[23] , \Level2Out132[23] , 
        \Level4Out100[24] , \Level1Out216[6] , \Level4Out76[13] , 
        \Level2Out92[5] , \Level2Out164[22] , \Level4Out20[12] , 
        \Level4Out156[25] , \ScanLink63[2] , \ScanLink75[6] , 
        \Level1Out168[27] , \Level1Out176[3] , \Level2Out104[26] , 
        \Level4Out136[21] , \Level4Out68[2] , \Level4Out40[16] , 
        \Level4Out16[17] , \Level4Out160[20] , \ScanLink107[23] , 
        \ScanLink112[17] , \ScanLink131[26] , \Level2Out152[27] , 
        \ScanLink144[16] , \ScanLink192[9] , \Level1Out200[2] , 
        \Level2Out82[13] , \Level2Out84[1] , \Level16Out0[18] , 
        \ScanLink167[27] , \ScanLink124[12] , \Level1Out160[7] , 
        \ScanLink172[13] , \ScanLink151[22] , \Level1Out88[19] , 
        \Level1Out117[22] , \Level2Out158[12] , \Level1Out134[13] , 
        \Level1Out162[12] , \Level32Out224[15] , \Level2Out56[7] , 
        \Level1Out141[23] , \Level1Out25[19] , \Level1Out50[29] , 
        \Level1Out102[16] , \Level1Out121[27] , \Level1Out154[17] , 
        \Level16Out224[20] , \Level1Out177[26] , \Level2Out138[16] , 
        \Level2Out180[22] , \Level2Out250[15] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink11[14] , \Level1Out50[30] , \ScanLink64[24] , 
        \Level1Out73[18] , \Level1Out199[13] , \ScanLink223[9] , 
        \Level1Out229[20] , \Level1Out249[24] , \Level4Out92[13] , 
        \Level2Out206[14] , \Level2Out230[11] , \Level4Out184[20] , 
        \ScanLink239[21] , \ScanLink27[11] , \ScanLink32[25] , 
        \ScanLink47[15] , \ScanLink52[21] , \Level1Out203[1] , \ScanLink60[1] , 
        \ScanLink71[10] , \ScanLink189[12] , \Level1Out154[24] , 
        \Level1Out163[4] , \Level2Out32[3] , \Level16Out224[13] , 
        \Level1Out89[5] , \Level1Out121[14] , \Level1Out177[15] , 
        \Level2Out138[25] , \ScanLink11[27] , \ScanLink27[22] , 
        \Level1Load79[0] , \Level1Out102[25] , \Level1Out104[3] , 
        \ScanLink107[10] , \Level1Out117[11] , \Level1Out162[21] , 
        \Level32Out224[26] , \Level2Out158[21] , \Level1Out134[20] , 
        \Level1Out141[10] , \ScanLink172[20] , \ScanLink124[21] , 
        \ScanLink151[11] , \ScanLink131[15] , \ScanLink139[4] , 
        \ScanLink144[25] , \ScanLink167[14] , \ScanLink112[24] , 
        \Level2Out82[20] , \ScanLink52[12] , \Level1Out58[0] , 
        \Level1Out97[9] , \ScanLink189[21] , \ScanLink71[23] , 
        \ScanLink32[16] , \ScanLink64[17] , \Level1Out107[0] , 
        \ScanLink239[12] , \ScanLink47[26] , \ScanLink127[8] , 
        \Level1Out229[13] , \Level4Out184[13] , \Level1Out249[17] , 
        \Level2Out168[3] , \Level2Out180[11] , \Level2Out208[6] , 
        \Level2Out230[22] , \Level2Out250[26] , \Level2Out206[27] , 
        \Level4Out92[20] , \ScanLink0[6] , \Level1Out1[19] , \ScanLink8[25] , 
        \Level1Out199[20] , \Level2Out110[18] , \ScanLink8[16] , 
        \Level1Out8[7] , \Level1Out39[9] , \Level1Out109[30] , 
        \Level1Out96[12] , \Level16Out48[1] , \Level1Out18[23] , 
        \Level1Out24[6] , \Level1Out83[26] , \Level1Out109[29] , 
        \ScanLink194[7] , \Level2Out114[5] , \Level2Out146[19] , 
        \Level8Out40[4] , \Level1Out166[9] , \Level2Out50[9] , 
        \Level1Out27[5] , \ScanLink78[3] , \ScanLink119[31] , \ScanLink146[1] , 
        \ScanLink189[8] , \Level8Out56[27] , \ScanLink119[28] , 
        \ScanLink226[4] , \Level16Out128[4] , \ScanLink145[2] , 
        \Level2Out12[30] , \Level2Out44[28] , \Level4Out240[3] , 
        \Level1Out218[0] , \Level2Out12[29] , \Level2Out44[31] , 
        \Level1Out178[5] , \Level4Out120[6] , \ScanLink197[19] , 
        \ScanLink225[7] , \Level1Out40[2] , \Level1Out78[27] , 
        \Level1Out187[18] , \Level2Out0[12] , \ScanLink197[4] , 
        \ScanLink238[8] , \Level64Out64[5] , \ScanLink94[30] , 
        \ScanLink122[5] , \Level8Out56[14] , \Level1Out83[15] , 
        \ScanLink94[29] , \ScanLink242[0] , \Level4Out188[8] , 
        \Level8Out24[0] , \Level1Out92[4] , \Level1Load105[0] , 
        \Level2Out210[4] , \Level1Out78[14] , \Level1Out91[7] , 
        \Level1Out96[21] , \Level2Out170[1] , \Level1Out214[29] , 
        \Level1Out214[30] , \Level1Out242[31] , \Level1Out237[18] , 
        \Level1Out242[28] , \ScanLink3[5] , \Level1Out5[31] , 
        \Level1Out18[10] , \Level2Out0[21] , \Level16Load32[0] , 
        \ScanLink39[30] , \Level4Out196[4] , \ScanLink39[29] , 
        \Level1Out43[1] , \Level4Out224[7] , \Level16Out32[9] , 
        \ScanLink121[6] , \ScanLink204[31] , \ScanLink204[28] , 
        \ScanLink252[30] , \Level2Load114[0] , \ScanLink227[19] , 
        \ScanLink241[3] , \Level4Out144[2] , \ScanLink252[29] , 
        \Level1Out5[28] , \Level1Out125[8] , \Level1Out210[18] , 
        \Level1Out233[30] , \Level1Load242[0] , \Level1Load21[0] , 
        \ScanLink38[1] , \ScanLink48[31] , \Level1Out69[11] , 
        \Level1Out233[29] , \Level1Out246[19] , \Level2Out4[10] , 
        \Level4Out160[4] , \Level8Out192[15] , \ScanLink48[28] , 
        \Level1Out138[7] , \Level1Out67[7] , \ScanLink105[0] , 
        \ScanLink200[19] , \ScanLink223[31] , \Level4Out200[1] , 
        \ScanLink223[28] , \ScanLink256[18] , \Level2Out186[1] , 
        \Level1Out64[4] , \ScanLink90[18] , \Level8Out64[20] , 
        \Level1Out87[24] , \ScanLink106[3] , \Level8Out32[21] , 
        \Level16Out208[3] , \Level2Out154[7] , \Level1Out92[10] , 
        \Level2Out234[2] , \ScanLink161[4] , \ScanLink193[31] , 
        \ScanLink193[28] , \ScanLink201[1] , \Level2Out16[18] , 
        \Level2Out40[19] , \Level4Out104[0] , \Level1Out183[29] , 
        \Level32Out160[29] , \ScanLink42[9] , \Level1Out69[22] , 
        \Level2Out4[23] , \Level4Out88[29] , \Level1Out183[30] , 
        \Level8Out192[26] , \Level32Out160[30] , \Level1Out221[9] , 
        \Level4Out88[30] , \Level2Out142[31] , \ScanLink6[8] , \ScanLink7[18] , 
        \ScanLink15[16] , \ScanLink20[3] , \ScanLink56[23] , \Level1Out87[17] , 
        \Level1Out92[23] , \Level1Out178[31] , \Level2Out114[29] , 
        \Level2Out114[30] , \Level2Out130[3] , \Level2Out142[28] , 
        \Level1Out178[28] , \Level8Out64[2] , \ScanLink162[7] , 
        \Level1Out190[9] , \ScanLink202[2] , \Level2Out98[29] , 
        \Level2Out250[6] , \Level2Out98[30] , \Level8Out64[13] , 
        \Level8Out32[12] , \ScanLink168[30] , \ScanLink168[29] , 
        \ScanLink23[13] , \ScanLink60[26] , \ScanLink75[12] , 
        \ScanLink228[17] , \Level64Out0[2] , \Level1Out123[6] , 
        \Level2Out68[24] , \ScanLink198[24] , \ScanLink36[27] , 
        \ScanLink43[17] , \ScanLink248[13] , \Level1Out61[9] , 
        \Level1Out188[25] , \Level1Out243[3] , \Level2Out234[13] , 
        \Level4Out20[8] , \Level4Out180[22] , \Level16Out128[25] , 
        \Level2Out254[17] , \Level1Out125[25] , \Level1Out238[16] , 
        \Level2Out184[20] , \Level32Out128[10] , \Level2Out202[16] , 
        \Level4Out96[11] , \Level1Out150[15] , \ScanLink15[25] , 
        \Level1Out21[31] , \Level1Out21[28] , \ScanLink23[0] , 
        \ScanLink103[21] , \Level1Out106[14] , \Level1Out113[20] , 
        \Level1Out173[24] , \Level1Out130[11] , \Level1Out166[10] , 
        \Level2Out16[5] , \Level16Out240[26] , \Level1Out145[21] , 
        \ScanLink120[10] , \Level1Out120[5] , \ScanLink176[11] , 
        \Level2Out152[9] , \ScanLink155[20] , \ScanLink116[15] , 
        \ScanLink135[24] , \ScanLink140[14] , \Level1Out240[0] , 
        \ScanLink163[25] , \Level2Out86[11] , \Level1Out54[18] , 
        \Level1Out77[30] , \Level1Out195[4] , \Level2Out184[13] , 
        \Level32Out128[23] , \Level2Out254[24] , \Level2Out128[1] , 
        \ScanLink59[8] , \Level1Out77[29] , \ScanLink96[1] , 
        \Level2Out202[25] , \Level4Out96[22] , \Level1Out188[16] , 
        \Level1Out238[25] , \Level4Out180[11] , \Level16Out128[16] , 
        \Level2Out234[20] , \Level2Out248[4] , \Level1Out18[2] , 
        \ScanLink23[20] , \ScanLink36[14] , \ScanLink60[15] , 
        \ScanLink248[20] , \Level1Out147[2] , \ScanLink198[17] , 
        \ScanLink43[24] , \ScanLink44[7] , \ScanLink56[10] , \Level1Out227[7] , 
        \ScanLink228[24] , \Level2Out68[17] , \ScanLink47[4] , 
        \ScanLink75[21] , \ScanLink140[27] , \ScanLink135[17] , 
        \ScanLink11[16] , \ScanLink27[13] , \ScanLink60[3] , \ScanLink95[2] , 
        \ScanLink103[12] , \ScanLink116[26] , \Level1Out144[1] , 
        \ScanLink163[16] , \ScanLink176[22] , \ScanLink219[3] , 
        \Level2Out86[22] , \ScanLink120[23] , \ScanLink155[13] , 
        \ScanLink179[6] , \Level1Out166[23] , \Level1Out224[4] , 
        \Level1Out106[27] , \Level1Out113[13] , \Level1Out125[16] , 
        \Level1Out130[22] , \Level1Out145[12] , \Level4Out88[6] , 
        \Level1Out150[26] , \Level1Out196[7] , \Level16Out240[15] , 
        \Level2Out72[1] , \Level1Out173[17] , \ScanLink164[9] , 
        \ScanLink52[23] , \ScanLink71[12] , \Level1Out163[6] , 
        \ScanLink189[10] , \Level1Out21[9] , \ScanLink32[27] , 
        \ScanLink64[26] , \Level2Out48[9] , \ScanLink239[23] , 
        \ScanLink47[17] , \ScanLink191[8] , \Level1Out203[3] , 
        \Level1Out229[22] , \Level4Out184[22] , \Level2Out230[13] , 
        \Level4Out60[8] , \Level1Out249[26] , \Level2Out180[20] , 
        \Level2Out206[16] , \Level2Out250[17] , \Level4Out92[11] , 
        \ScanLink3[18] , \Level1Out154[15] , \Level1Out199[11] , 
        \Level32Out0[8] , \ScanLink220[8] , \Level16Out224[22] , 
        \Level1Out25[28] , \Level1Out50[18] , \ScanLink63[0] , 
        \Level1Out102[14] , \Level1Out121[25] , \Level1Out177[24] , 
        \Level2Out138[14] , \ScanLink107[21] , \Level1Out117[20] , 
        \Level1Out162[10] , \Level2Out158[10] , \Level32Out224[17] , 
        \Level1Out134[11] , \Level1Out141[21] , \Level1Out160[5] , 
        \ScanLink172[11] , \Level2Out56[5] , \ScanLink151[20] , 
        \ScanLink112[15] , \ScanLink124[10] , \Level2Out112[9] , 
        \ScanLink131[24] , \ScanLink144[14] , \Level1Out200[0] , 
        \ScanLink167[25] , \Level2Out84[3] , \Level2Out82[11] , 
        \Level1Out73[30] , \Level2Out180[13] , \Level2Out250[24] , 
        \ScanLink0[4] , \Level1Out1[31] , \ScanLink11[25] , \ScanLink19[8] , 
        \Level1Out73[29] , \Level1Out25[31] , \Level1Out199[22] , 
        \Level1Out249[15] , \Level2Out168[1] , \Level2Out206[25] , 
        \Level4Out92[22] , \ScanLink64[15] , \Level1Out229[11] , 
        \Level2Out208[4] , \Level2Out230[20] , \Level4Out184[11] , 
        \Level1Out107[2] , \ScanLink239[10] , \ScanLink27[20] , 
        \ScanLink32[14] , \ScanLink47[24] , \ScanLink52[10] , \Level1Out58[2] , 
        \ScanLink71[21] , \ScanLink189[23] , \Level1Out88[31] , 
        \Level1Out88[28] , \Level1Out94[8] , \Level1Out104[1] , 
        \ScanLink131[17] , \Level16Out0[30] , \ScanLink144[27] , 
        \Level16Out0[29] , \ScanLink107[12] , \ScanLink112[26] , 
        \ScanLink167[16] , \Level2Out82[22] , \Level1Out117[13] , 
        \ScanLink124[23] , \ScanLink139[6] , \ScanLink172[22] , 
        \Level2Out216[8] , \ScanLink151[13] , \Level1Out162[23] , 
        \Level2Out158[23] , \Level32Out224[24] , \Level1Out134[22] , 
        \Level1Out141[12] , \Level1Out89[7] , \Level1Out121[16] , 
        \Level1Out102[27] , \ScanLink124[9] , \Level1Out154[26] , 
        \Level2Out32[1] , \Level16Out224[11] , \Level1Out165[8] , 
        \Level1Out177[17] , \Level2Out138[27] , \Level1Out214[18] , 
        \Level1Out237[30] , \Level1Out1[28] , \Level1Out78[25] , 
        \Level1Out237[29] , \ScanLink8[27] , \Level1Out18[21] , 
        \ScanLink197[6] , \Level1Load202[0] , \Level1Out242[19] , 
        \Level2Out0[10] , \Level1Out24[4] , \Level1Out27[7] , \ScanLink39[18] , 
        \Level1Out178[7] , \Level64Out64[7] , \ScanLink225[5] , 
        \Level4Out120[4] , \ScanLink145[0] , \ScanLink204[19] , 
        \Level1Out218[2] , \ScanLink227[31] , \Level4Out240[1] , 
        \ScanLink78[1] , \ScanLink227[28] , \ScanLink252[18] , 
        \ScanLink94[18] , \ScanLink226[6] , \Level8Out56[25] , 
        \Level16Out128[6] , \Level1Out83[24] , \ScanLink146[3] , 
        \Level2Out114[7] , \ScanLink8[14] , \Level1Out8[5] , \ScanLink194[5] , 
        \Level8Out40[6] , \Level1Out18[12] , \Level1Out43[3] , 
        \Level1Out96[10] , \ScanLink241[1] , \Level2Out44[19] , 
        \Level16Out48[3] , \Level2Out12[18] , \Level4Out144[0] , 
        \ScanLink121[4] , \ScanLink197[28] , \ScanLink197[31] , 
        \Level4Out224[5] , \Level1Load61[0] , \Level1Out187[29] , 
        \Level2Out0[23] , \Level1Out78[16] , \Level1Out91[5] , 
        \Level1Out187[30] , \Level4Out196[6] , \Level2Out110[29] , 
        \ScanLink38[3] , \Level1Out40[0] , \Level1Out83[17] , 
        \Level1Out96[23] , \Level2Out146[31] , \Level1Out109[18] , 
        \Level2Out110[30] , \Level2Out146[28] , \Level2Out170[3] , 
        \Level1Out92[6] , \Level8Out24[2] , \ScanLink122[7] , \ScanLink242[2] , 
        \Level2Out210[6] , \Level4Out8[9] , \Level8Out56[16] , 
        \Level1Out64[6] , \Level1Out79[9] , \ScanLink119[19] , 
        \Level1Out87[26] , \Level1Out92[12] , \Level1Out178[19] , 
        \Level2Out114[18] , \Level2Out142[19] , \Level2Out234[0] , 
        \Level2Out154[5] , \Level1Out126[9] , \Level2Out98[18] , 
        \ScanLink106[1] , \Level2Out10[9] , \Level8Out64[22] , 
        \Level8Out32[23] , \Level16Out208[1] , \Level1Out67[5] , 
        \ScanLink105[2] , \ScanLink168[18] , \Level2Out186[3] , 
        \Level2Out16[30] , \Level2Out40[28] , \Level4Out200[3] , 
        \Level1Out69[13] , \Level1Load97[0] , \Level1Out138[5] , 
        \Level2Out16[29] , \Level2Out40[31] , \ScanLink193[19] , 
        \Level4Out160[6] , \Level1Out87[15] , \ScanLink90[30] , 
        \Level1Out183[18] , \Level32Out160[18] , \Level2Out4[12] , 
        \Level4Out88[18] , \Level8Out192[17] , \Level16Out176[8] , 
        \ScanLink90[29] , \ScanLink162[5] , \ScanLink202[0] , 
        \Level8Out64[11] , \Level16Load224[0] , \Level1Out222[8] , 
        \Level8Out32[10] , \Level1Load145[0] , \Level2Out250[4] , 
        \Level8Out64[0] , \ScanLink3[7] , \Level1Out5[19] , \ScanLink41[8] , 
        \Level1Out92[21] , \Level1Out210[29] , \Level1Out246[31] , 
        \Level2Out130[1] , \Level1Out246[28] , \Level1Out69[20] , 
        \Level1Out210[30] , \Level1Out233[18] , \Level2Out4[21] , 
        \Level1Out4[20] , \Level1Out4[13] , \ScanLink5[9] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink15[14] , \Level1Out21[19] , \ScanLink23[2] , 
        \ScanLink48[19] , \ScanLink161[6] , \Level8Out192[24] , 
        \ScanLink103[23] , \ScanLink116[17] , \ScanLink135[26] , 
        \ScanLink140[16] , \Level1Out193[8] , \ScanLink200[28] , 
        \ScanLink256[30] , \Level2Load154[0] , \ScanLink200[31] , 
        \ScanLink201[3] , \ScanLink223[19] , \ScanLink256[29] , 
        \Level1Out240[2] , \Level4Out104[2] , \ScanLink163[27] , 
        \Level2Out86[13] , \Level1Out120[7] , \ScanLink176[13] , 
        \ScanLink155[22] , \Level32Out128[8] , \Level1Out62[8] , 
        \Level1Out113[22] , \ScanLink120[12] , \Level1Out166[12] , 
        \Level1Out145[23] , \Level1Out106[16] , \Level1Out125[27] , 
        \Level1Out130[13] , \Level1Out150[17] , \Level2Out16[7] , 
        \Level16Out240[24] , \Level1Out173[26] , \Level32Out128[12] , 
        \Level1Out54[30] , \Level1Out54[29] , \Level2Out184[22] , 
        \Level2Out254[15] , \Level1Out77[18] , \Level1Out238[14] , 
        \Level2Out202[14] , \Level4Out96[13] , \Level1Out188[27] , 
        \Level4Out180[20] , \Level16Out128[27] , \Level2Out234[11] , 
        \ScanLink20[1] , \ScanLink36[25] , \ScanLink60[24] , \ScanLink248[11] , 
        \ScanLink198[26] , \ScanLink43[15] , \Level1Out243[1] , 
        \ScanLink23[11] , \ScanLink56[21] , \ScanLink75[10] , 
        \Level1Out123[4] , \ScanLink228[15] , \Level2Out68[26] , 
        \Level64Out0[0] , \Level1Out125[14] , \Level1Out150[24] , 
        \Level2Out72[3] , \Level1Out106[25] , \Level1Out173[15] , 
        \Level1Out239[9] , \ScanLink15[27] , \Level1Out18[0] , 
        \ScanLink23[22] , \Level1Load39[0] , \ScanLink95[0] , 
        \Level1Out113[11] , \ScanLink47[6] , \ScanLink103[10] , 
        \Level1Out130[20] , \Level1Out166[21] , \Level1Out196[5] , 
        \Level16Out240[17] , \Level1Out145[10] , \Level4Out88[4] , 
        \ScanLink120[21] , \ScanLink176[20] , \ScanLink155[11] , 
        \ScanLink179[4] , \Level1Out224[6] , \ScanLink56[12] , 
        \ScanLink116[24] , \ScanLink135[15] , \ScanLink140[25] , 
        \Level1Out144[3] , \ScanLink219[1] , \Level2Out86[20] , 
        \ScanLink163[14] , \Level1Out227[5] , \ScanLink75[23] , 
        \ScanLink228[26] , \ScanLink60[17] , \Level1Out188[9] , 
        \Level2Out68[15] , \Level1Out147[0] , \ScanLink198[15] , 
        \Level4Out96[8] , \ScanLink29[17] , \ScanLink36[16] , \ScanLink43[26] , 
        \ScanLink248[22] , \ScanLink44[5] , \ScanLink49[13] , \ScanLink96[3] , 
        \ScanLink167[8] , \Level1Out188[14] , \Level1Out195[6] , 
        \Level2Out234[22] , \Level4Out180[13] , \Level16Out128[14] , 
        \Level2Out248[6] , \Level2Out184[11] , \Level2Out254[26] , 
        \Level32Out128[21] , \Level1Out238[27] , \Level2Out54[25] , 
        \Level2Out128[3] , \Level2Out202[27] , \Level4Out96[20] , 
        \ScanLink80[7] , \Level1Out183[2] , \ScanLink192[20] , 
        \ScanLink214[16] , \ScanLink237[27] , \ScanLink242[17] , 
        \Level32Out224[1] , \ScanLink211[9] , \Level2Out62[20] , 
        \ScanLink187[14] , \ScanLink222[13] , \ScanLink201[22] , 
        \Level1Out231[1] , \Level2Out34[21] , \Level1Out10[8] , 
        \ScanLink51[2] , \ScanLink52[1] , \Level1Out151[4] , 
        \Level1Out197[15] , \Level1Out247[22] , \Level2Out208[12] , 
        \Level1Load199[0] , \Level1Out232[12] , \Level1Out211[23] , 
        \Level1Out204[17] , \Level1Out252[16] , \Level1Out119[24] , 
        \Level1Out182[21] , \Level1Out227[26] , \Level1Out232[2] , 
        \Level2Out100[15] , \Level4Out132[12] , \Level4Out44[25] , 
        \Level4Out12[24] , \Level4Out164[13] , \Level2Out156[14] , 
        \Level1Out152[7] , \Level1Out179[20] , \Level4Out104[17] , 
        \Level2Out136[10] , \Level4Out24[21] , \Level4Out72[20] , 
        \Level2Out160[11] , \Level4Out152[16] , \ScanLink36[5] , 
        \Level1Out68[19] , \ScanLink83[4] , \ScanLink91[23] , 
        \ScanLink169[21] , \Level2Out64[7] , \Level64Out0[10] , 
        \ScanLink84[17] , \Level1Load228[0] , \Level2Load188[0] , 
        \ScanLink108[7] , \ScanLink109[25] , \Level1Out180[1] , 
        \Level1Out204[24] , \Level1Out182[12] , \Level1Out227[15] , 
        \Level1Out252[25] , \Level1Out255[5] , \Level16Out96[19] , 
        \Level1Out197[26] , \Level1Out232[21] , \Level2Out188[5] , 
        \Level2Out208[21] , \ScanLink6[23] , \Level1Out15[5] , \ScanLink28[9] , 
        \ScanLink29[24] , \ScanLink115[8] , \Level1Out135[0] , 
        \Level1Out247[11] , \ScanLink187[27] , \Level1Out211[10] , 
        \ScanLink201[11] , \ScanLink222[20] , \Level2Out62[13] , 
        \Level2Out34[12] , \ScanLink49[20] , \ScanLink84[24] , 
        \ScanLink109[16] , \ScanLink192[13] , \ScanLink214[25] , 
        \ScanLink237[14] , \Level2Out54[16] , \ScanLink242[24] , 
        \ScanLink91[10] , \ScanLink169[12] , \ScanLink35[6] , \Level1Out69[3] , 
        \Level1Out93[18] , \Level2Out136[23] , \Level2Out196[9] , 
        \Level64Out0[23] , \Level4Out72[13] , \Level1Out179[13] , 
        \Level4Out104[24] , \Level2Out160[22] , \Level4Out152[25] , 
        \Level1Out119[17] , \Level1Out136[3] , \Level4Out24[12] , 
        \Level2Out100[26] , \Level4Out44[16] , \Level2Out156[27] , 
        \Level4Out28[2] , \Level4Out132[21] , \Level4Out164[20] , 
        \Level1Out40[24] , \Level4Out12[17] , \Level2Out240[18] , 
        \Level1Out16[25] , \Level1Out35[14] , \Level1Out63[15] , 
        \Level8Out248[26] , \ScanLink177[2] , \Level1Out16[6] , 
        \Level1Out20[20] , \ScanLink49[0] , \Level1Out76[21] , \ScanLink86[9] , 
        \Level2Out216[19] , \Level1Out55[10] , \ScanLink217[7] , 
        \Level2Out138[9] , \ScanLink22[31] , \ScanLink74[29] , 
        \Level4Out112[6] , \ScanLink22[28] , \ScanLink57[18] , 
        \ScanLink74[30] , \Level64Out64[14] , \ScanLink98[5] , 
        \Level1Out154[9] , \Level1Out198[3] , \ScanLink249[31] , 
        \ScanLink249[28] , \Level8Out80[11] , \Level2Out246[0] , 
        \Level8Out72[4] , \Level1Out98[14] , \ScanLink174[1] , 
        \Level2Out126[5] , \Level1Out229[3] , \Level2Out62[9] , 
        \Level1Out149[6] , \ScanLink214[4] , \Level2Out18[1] , 
        \Level8Out80[22] , \Level8Out120[25] , \Level8Out176[24] , 
        \Level64Out64[27] , \Level1Out0[22] , \Level1Out0[11] , 
        \ScanLink2[21] , \ScanLink6[10] , \Level1Out16[16] , \Level1Out20[13] , 
        \Level1Out71[1] , \Level1Out76[12] , \ScanLink113[6] , 
        \Level4Out212[31] , \Level4Out216[7] , \Level4Out244[29] , 
        \Level1Out35[27] , \Level1Out55[23] , \Level4Out212[28] , 
        \Level4Out244[30] , \Level1Out40[17] , \Level4Out176[2] , 
        \Level8Out248[15] , \Level2Load126[0] , \Level1Out63[26] , 
        \Level1Out72[2] , \Level8Out176[17] , \Level1Out98[27] , 
        \ScanLink110[5] , \Level1Out112[31] , \Level1Out144[29] , 
        \Level2Out128[31] , \Level1Out131[19] , \Level2Out128[28] , 
        \Level1Out112[28] , \Level1Out144[30] , \Level1Out167[18] , 
        \Level8Out120[16] , \Level2Out190[7] , \ScanLink33[8] , 
        \Level1Load137[0] , \ScanLink154[28] , \Level1Out250[8] , 
        \Level2Out222[4] , \Level8Out16[0] , \Level1Out56[4] , 
        \Level1Out89[22] , \ScanLink102[30] , \ScanLink102[29] , 
        \ScanLink121[18] , \Level2Out142[1] , \ScanLink154[31] , 
        \ScanLink177[19] , \Level1Out109[4] , \Level1Out116[19] , 
        \Level1Out135[31] , \Level1Out135[28] , \Level1Out140[18] , 
        \Level1Out163[30] , \ScanLink254[6] , \Level4Out68[30] , 
        \Level4Out68[29] , \ScanLink134[3] , \Level1Out163[29] , 
        \Level8Out144[23] , \Level8Out112[22] , \ScanLink2[12] , 
        \Level1Out12[27] , \Level1Out24[22] , \Level1Out48[8] , 
        \Level1Out84[2] , \ScanLink106[18] , \ScanLink125[30] , 
        \ScanLink125[29] , \ScanLink249[9] , \Level2Out2[9] , 
        \Level2Out166[7] , \ScanLink150[19] , \ScanLink173[31] , 
        \Level8Out32[6] , \Level1Out87[1] , \Level1Out117[8] , 
        \ScanLink173[28] , \Level2Out78[30] , \Level2Out206[2] , 
        \ScanLink188[29] , \Level2Out78[29] , \Level4Out180[2] , 
        \Level1Out51[12] , \Level1Out72[23] , \ScanLink188[30] , 
        \Level1Out198[28] , \Level4Out240[18] , \Level1Out198[31] , 
        \Level4Out152[4] , \Level4Out216[19] , \Level32Out96[24] , 
        \Level1Out31[16] , \Level1Out44[26] , \Level1Out55[7] , 
        \Level4Out0[1] , \Level1Out67[17] , \ScanLink137[0] , \ScanLink182[1] , 
        \Level2Out94[9] , \Level2Out102[3] , \Level4Load48[0] , 
        \Level4Out232[1] , \Level64Out192[23] , \Level8Out56[2] , 
        \ScanLink230[2] , \Level4Out128[31] , \Level4Out248[9] , 
        \Level8Out144[10] , \Level4Out128[28] , \ScanLink11[0] , 
        \Level1Out12[14] , \Level1Out31[25] , \Level1Out32[0] , 
        \Level8Out112[11] , \Level1Out89[11] , \ScanLink150[7] , 
        \Level1Out44[15] , \Level1Out228[31] , \ScanLink233[1] , 
        \Level2Out212[31] , \Level2Out244[29] , \Level2Out212[28] , 
        \Level4Out136[0] , \Level1Load13[0] , \Level1Out24[11] , 
        \Level1Out31[3] , \Level1Out67[24] , \Level1Out228[28] , 
        \Level64Out192[10] , \Level2Out244[30] , \Level1Out72[10] , 
        \ScanLink153[4] , \ScanLink26[19] , \Level1Out51[21] , 
        \ScanLink53[30] , \ScanLink70[18] , \Level32Out96[17] , 
        \ScanLink70[9] , \ScanLink53[29] , \ScanLink80[15] , \ScanLink178[17] , 
        \ScanLink181[2] , \Level1Out213[9] , \ScanLink238[30] , 
        \ScanLink238[29] , \Level2Out58[3] , \ScanLink95[21] , 
        \ScanLink252[8] , \Level4Load188[0] , \ScanLink118[13] , 
        \Level2Out24[5] , \Level2Out88[17] , \ScanLink12[3] , 
        \Level1Out19[18] , \Level1Out97[30] , \Level1Out97[29] , 
        \Level4Out100[15] , \Level1Out108[12] , \Level2Out132[12] , 
        \Level4Out76[22] , \Level2Out160[9] , \Level1Out111[6] , 
        \Level1Out112[5] , \Level1Out168[16] , \Level2Out4[7] , 
        \Level2Out104[17] , \Level2Out164[13] , \Level4Out20[23] , 
        \Level4Out156[14] , \Level4Out136[10] , \Level4Out40[27] , 
        \Level4Out16[26] , \Level2Out152[16] , \Level4Out160[11] , 
        \Level4Out208[12] , \Level1Out200[15] , \Level1Out186[23] , 
        \Level1Out223[24] , \Level1Out243[20] , \Level1Out5[0] , 
        \Level1Out29[1] , \ScanLink38[21] , \ScanLink58[25] , 
        \ScanLink183[16] , \Level1Out193[17] , \Level1Out215[21] , 
        \Level1Out236[10] , \ScanLink253[21] , \Level2Out66[22] , 
        \ScanLink205[20] , \ScanLink226[11] , \Level2Out30[23] , 
        \Level4Out12[8] , \Level8Out0[24] , \Level1Out53[9] , 
        \ScanLink210[14] , \Level2Out50[27] , \ScanLink75[4] , 
        \Level1Out176[1] , \ScanLink196[22] , \ScanLink233[25] , 
        \ScanLink246[15] , \Level4Out40[14] , \Level2Out104[24] , 
        \Level4Out68[0] , \Level2Out152[25] , \Level4Out136[23] , 
        \Level1Out108[21] , \Level1Out168[25] , \Level4Out16[15] , 
        \Level4Out160[22] , \Level1Out216[4] , \Level4Out76[11] , 
        \Level2Out132[21] , \Level2Out164[20] , \Level4Out100[26] , 
        \Level4Out156[27] , \ScanLink95[12] , \ScanLink118[20] , 
        \Level2Out92[7] , \Level4Out20[10] , \Level2Out88[24] , 
        \ScanLink156[9] , \ScanLink199[0] , \Level128Out128[6] , 
        \Level1Out6[3] , \ScanLink38[12] , \ScanLink80[26] , \ScanLink178[24] , 
        \Level2Out40[1] , \ScanLink210[27] , \Level32Out160[2] , 
        \ScanLink58[16] , \ScanLink183[25] , \ScanLink196[11] , 
        \ScanLink233[16] , \Level2Out50[14] , \ScanLink246[26] , 
        \ScanLink205[13] , \ScanLink226[22] , \ScanLink253[12] , 
        \Level2Out66[11] , \Level8Out0[17] , \Level2Out30[10] , 
        \Level1Out208[8] , \ScanLink76[7] , \Level1Out193[24] , 
        \Level1Out236[23] , \Level1Out243[13] , \Level1Out0[18] , 
        \Level1Out4[30] , \Level1Out4[29] , \ScanLink6[19] , \ScanLink14[17] , 
        \ScanLink22[12] , \ScanLink30[2] , \ScanLink74[13] , \Level1Out133[7] , 
        \ScanLink148[5] , \Level1Out175[2] , \Level1Out200[26] , 
        \Level1Out215[12] , \ScanLink228[0] , \Level4Out208[21] , 
        \Level8Out232[18] , \Level1Out186[10] , \Level1Out223[17] , 
        \Level1Out215[7] , \ScanLink229[16] , \Level16Out160[5] , 
        \ScanLink37[26] , \ScanLink57[22] , \Level16Load128[0] , 
        \ScanLink42[16] , \Level1Out253[2] , \ScanLink61[27] , 
        \ScanLink249[12] , \Level1Out71[8] , \Level1Out189[24] , 
        \ScanLink199[25] , \Level2Out18[8] , \Level2Out190[15] , 
        \Level2Out216[23] , \Level2Out240[22] , \Level4Out224[24] , 
        \Level1Out239[17] , \Level1Load249[0] , \Level8Out184[2] , 
        \Level4Out244[20] , \Level1Out107[15] , \Level1Out172[25] , 
        \Level2Out220[26] , \Level4Out212[21] , \Level1Out151[14] , 
        \Level2Out148[25] , \ScanLink8[5] , \Level1Out20[30] , \ScanLink33[1] , 
        \Level1Out112[21] , \Level1Out124[24] , \Level1Out131[10] , 
        \Level1Out144[20] , \Level1Out167[11] , \Level2Out128[21] , 
        \ScanLink154[21] , \ScanLink49[9] , \ScanLink86[0] , \ScanLink102[20] , 
        \ScanLink121[11] , \Level1Out130[4] , \ScanLink177[10] , 
        \Level2Out142[8] , \Level2Out92[24] , \Level64Out192[3] , 
        \ScanLink117[14] , \ScanLink162[24] , \Level4Out168[7] , 
        \ScanLink134[25] , \ScanLink141[15] , \Level1Out250[1] , 
        \Level8Out16[9] , \Level4Out208[2] , \Level1Out239[24] , 
        \Level4Out244[13] , \Level1Out76[28] , \Level2Out138[0] , 
        \Level1Out55[19] , \Level1Out185[5] , \Level1Out76[31] , 
        \Level2Out220[15] , \ScanLink14[24] , \Level1Out20[29] , 
        \Level4Out212[12] , \ScanLink37[15] , \ScanLink42[25] , 
        \Level1Out189[17] , \Level2Out190[26] , \Level2Out240[11] , 
        \Level2Out216[10] , \Level4Out224[17] , \Level16Out64[4] , 
        \ScanLink54[6] , \ScanLink61[14] , \Level8Out80[18] , 
        \Level1Out157[3] , \ScanLink199[16] , \ScanLink22[21] , 
        \ScanLink57[11] , \ScanLink74[20] , \ScanLink229[25] , 
        \ScanLink249[21] , \Level1Out237[6] , \ScanLink57[5] , 
        \ScanLink117[27] , \Level1Out154[0] , \Level2Load46[0] , 
        \ScanLink209[2] , \ScanLink162[17] , \ScanLink85[3] , 
        \ScanLink102[13] , \ScanLink121[22] , \ScanLink134[16] , 
        \ScanLink141[26] , \ScanLink154[12] , \ScanLink169[7] , 
        \Level1Out234[5] , \Level2Out92[17] , \Level1Out131[23] , 
        \ScanLink177[23] , \Level1Out186[6] , \Level2Out246[9] , 
        \Level1Out144[13] , \Level1Out107[26] , \Level1Out112[12] , 
        \Level1Out167[22] , \Level2Out128[12] , \ScanLink174[8] , 
        \Level2Out148[16] , \Level1Out124[17] , \Level1Out172[16] , 
        \Level1Out151[27] , \Level2Out62[0] , \Level1Out232[28] , 
        \Level8Out200[16] , \Level1Out247[18] , \Level1Out135[9] , 
        \Level2Out208[28] , \Level32Out96[2] , \Level1Out211[19] , 
        \Level1Out232[31] , \Level1Load5[0] , \Level1Out5[9] , \ScanLink9[24] , 
        \Level1Out10[1] , \Level1Out13[2] , \ScanLink28[0] , \ScanLink49[30] , 
        \ScanLink49[29] , \Level1Out68[10] , \Level2Out208[31] , 
        \Level16Out96[10] , \Level1Out128[6] , \Level4Load200[0] , 
        \Level1Out77[6] , \Level4Out36[7] , \ScanLink91[19] , \ScanLink115[1] , 
        \ScanLink222[29] , \ScanLink201[18] , \ScanLink222[30] , 
        \Level1Out248[3] , \Level1Out74[5] , \Level1Load84[0] , 
        \ScanLink116[2] , \Level2Out196[0] , \Level1Out86[25] , 
        \Level2Out144[6] , \Level4Out132[28] , \Level4Out164[30] , 
        \Level4Out164[29] , \Level4Out132[31] , \Level1Out93[11] , 
        \ScanLink171[5] , \ScanLink211[0] , \Level2Out224[3] , 
        \Level8Out168[15] , \Level2Out34[31] , \Level2Out62[29] , 
        \Level2Out34[28] , \Level2Out62[30] , \Level4Out52[3] , 
        \ScanLink192[30] , \Level32Out224[8] , \ScanLink52[8] , 
        \Level1Out182[31] , \ScanLink192[29] , \Level4Out80[5] , 
        \Level1Out68[23] , \Level1Out86[16] , \Level1Out93[22] , 
        \Level1Load156[0] , \Level1Out182[28] , \Level1Out231[8] , 
        \Level16Out96[23] , \Level8Out200[25] , \Level1Out179[29] , 
        \Level2Out136[19] , \Level4Out24[31] , \Level1Out179[30] , 
        \Level2Out120[2] , \Level4Out72[29] , \Level4Out24[28] , 
        \Level2Out160[18] , \Level8Out168[26] , \Level2Out240[7] , 
        \Level4Out72[30] , \Level1Out180[8] , \ScanLink212[3] , 
        \Level1Out29[8] , \Level1Out97[13] , \Level1Out108[28] , 
        \ScanLink169[31] , \ScanLink169[28] , \ScanLink172[6] , 
        \ScanLink184[6] , \Level64Out0[19] , \Level2Out164[30] , 
        \Level4Out76[18] , \Level1Out108[31] , \Level2Out132[28] , 
        \Level2Out164[29] , \Level2Out132[31] , \Level4Out20[19] , 
        \Level1Out82[27] , \Level1Out176[8] , \Level1Load211[0] , 
        \Level4Out68[9] , \Level2Out104[4] , \ScanLink156[0] , 
        \ScanLink199[9] , \Level1Out19[22] , \Level1Out34[7] , 
        \Level1Out37[4] , \ScanLink68[2] , \ScanLink118[29] , \ScanLink236[5] , 
        \Level2Out40[8] , \ScanLink118[30] , \ScanLink155[3] , 
        \Level2Out30[19] , \Level2Out66[18] , \Level2Load200[0] , 
        \Level1Out168[4] , \Level1Out208[1] , \Level1Out186[19] , 
        \ScanLink196[18] , \ScanLink235[6] , \Level4Out76[5] , 
        \Level4Out208[28] , \Level8Out232[11] , \ScanLink187[5] , 
        \Level4Out208[31] , \Level1Out50[3] , \Level1Out79[26] , 
        \ScanLink95[28] , \ScanLink228[9] , \ScanLink9[17] , \ScanLink11[9] , 
        \Level1Out82[14] , \Level1Out82[5] , \ScanLink95[31] , 
        \ScanLink132[4] , \ScanLink252[1] , \Level4Out136[19] , 
        \Level2Out200[5] , \Level1Out97[20] , \Level4Out160[18] , 
        \Level1Load72[0] , \Level2Out160[0] , \Level1Out0[4] , \Level1Out3[7] , 
        \Level1Out19[11] , \Level1Out79[15] , \Level1Out236[19] , 
        \Level1Out243[29] , \Level1Out81[6] , \Level1Out215[31] , 
        \Level1Out215[28] , \Level1Out243[30] , \Level8Out232[22] , 
        \Level1Out32[9] , \ScanLink38[31] , \ScanLink38[28] , \ScanLink131[7] , 
        \Level1Out53[0] , \ScanLink73[3] , \ScanLink113[16] , 
        \ScanLink166[26] , \ScanLink205[30] , \ScanLink226[18] , 
        \ScanLink251[2] , \ScanLink253[28] , \ScanLink205[29] , 
        \ScanLink253[31] , \Level4Out12[1] , \Level2Out94[0] , 
        \ScanLink130[27] , \ScanLink145[17] , \ScanLink182[8] , 
        \Level1Out210[3] , \Level4Out248[0] , \ScanLink150[23] , 
        \ScanLink106[22] , \ScanLink125[13] , \Level1Out170[6] , 
        \ScanLink173[12] , \Level2Out96[26] , \Level4Out128[5] , 
        \Level1Out89[18] , \Level1Out135[12] , \Level1Out140[22] , 
        \Level1Out163[13] , \Level2Out46[6] , \Level4Out148[25] , 
        \Level1Out103[17] , \Level1Out116[23] , \Level4Out68[13] , 
        \Level1Out176[27] , \Level8Out144[19] , \Level1Out120[26] , 
        \Level1Out155[16] , \Level4Out128[21] , \Level1Out248[25] , 
        \Level8Out48[7] , \Level8Out112[18] , \Level1Out1[12] , 
        \ScanLink2[31] , \ScanLink10[15] , \Level1Out24[18] , 
        \Level1Out51[31] , \Level1Out72[19] , \Level1Out198[12] , 
        \Level4Out240[22] , \ScanLink33[24] , \Level1Out51[28] , 
        \Level2Out224[24] , \Level4Out216[23] , \Level1Out228[21] , 
        \ScanLink233[8] , \Level2Out194[17] , \Level2Out212[21] , 
        \Level2Out244[20] , \Level4Out136[9] , \Level4Out220[26] , 
        \Level64Out192[19] , \ScanLink46[14] , \Level1Out213[0] , 
        \Level16Out240[2] , \ScanLink26[10] , \ScanLink65[25] , 
        \Level2Out78[13] , \ScanLink70[11] , \Level1Out173[5] , 
        \ScanLink238[20] , \ScanLink188[13] , \Level2Out18[17] , 
        \ScanLink70[0] , \ScanLink53[20] , \Level1Out103[24] , 
        \Level1Out176[14] , \ScanLink2[28] , \Level1Out99[4] , 
        \Level1Out120[15] , \Level1Out155[25] , \Level2Out22[2] , 
        \Level4Out128[12] , \ScanLink10[26] , \ScanLink14[4] , \ScanLink17[7] , 
        \ScanLink106[11] , \Level1Out116[10] , \Level1Out135[21] , 
        \Level1Out140[11] , \Level4Out148[16] , \Level4Out68[20] , 
        \ScanLink125[20] , \ScanLink129[5] , \Level1Out163[20] , 
        \ScanLink150[10] , \Level2Out2[0] , \ScanLink113[25] , 
        \Level1Out114[2] , \ScanLink173[21] , \Level2Out96[15] , 
        \ScanLink166[15] , \ScanLink249[0] , \ScanLink26[23] , 
        \Level1Out48[1] , \ScanLink70[22] , \Level1Out87[8] , 
        \ScanLink130[14] , \ScanLink145[24] , \ScanLink188[20] , 
        \Level2Out18[24] , \ScanLink53[13] , \Level16Out224[6] , 
        \ScanLink46[27] , \ScanLink33[17] , \ScanLink65[16] , 
        \Level1Out117[1] , \ScanLink238[13] , \ScanLink39[22] , 
        \ScanLink137[9] , \Level1Out228[12] , \Level2Out78[20] , 
        \Level16Out144[3] , \Level2Out194[24] , \Level2Out244[13] , 
        \Level4Out0[8] , \Level2Out218[7] , \ScanLink197[21] , 
        \Level1Out198[21] , \Level2Out212[12] , \Level4Out220[15] , 
        \Level4Out232[8] , \Level4Out240[11] , \ScanLink247[16] , 
        \Level1Out248[16] , \Level2Out178[2] , \Level2Out72[15] , 
        \Level2Out224[17] , \Level4Out216[10] , \ScanLink232[26] , 
        \ScanLink59[26] , \ScanLink204[23] , \ScanLink211[17] , 
        \Level2Out24[14] , \Level16Out32[2] , \Level2Out44[10] , 
        \ScanLink182[15] , \ScanLink227[12] , \ScanLink241[8] , 
        \ScanLink252[22] , \Level1Out214[22] , \Level2Out12[11] , 
        \Level4Out144[9] , \Level1Out242[23] , \Level1Out101[5] , 
        \Level1Out187[20] , \Level1Out192[14] , \Level1Out237[13] , 
        \Level2Out218[27] , \Level1Out222[27] , \Level1Out102[6] , 
        \Level1Out169[15] , \Level1Out201[16] , \Level2Out126[25] , 
        \Level2Out110[20] , \Level2Out170[24] , \Level4Out8[0] , 
        \Level1Out109[11] , \Level2Out146[21] , \Level1Out1[21] , 
        \Level1Out18[31] , \Level1Out18[28] , \Level1Out40[9] , 
        \ScanLink81[16] , \ScanLink94[22] , \ScanLink119[10] , 
        \Level2Out34[6] , \ScanLink179[14] , \ScanLink158[6] , 
        \Level4Out8[16] , \Level4Out188[3] , \Level1Out187[13] , 
        \Level1Out205[4] , \Level1Out222[14] , \Level1Out201[25] , 
        \Level2Out0[19] , \Level2Out218[14] , \ScanLink66[4] , 
        \Level1Out165[1] , \Level1Out214[11] , \ScanLink238[3] , 
        \Level1Out192[27] , \Level1Out237[20] , \Level1Out242[10] , 
        \ScanLink3[22] , \Level1Out13[24] , \ScanLink39[11] , \ScanLink59[15] , 
        \ScanLink145[9] , \ScanLink204[10] , \ScanLink182[26] , 
        \ScanLink227[21] , \Level2Out44[23] , \Level4Out240[8] , 
        \ScanLink197[12] , \ScanLink252[11] , \Level2Out12[22] , 
        \ScanLink211[24] , \ScanLink232[15] , \ScanLink247[25] , 
        \Level2Out72[26] , \Level2Out24[27] , \Level1Out39[2] , 
        \ScanLink78[8] , \ScanLink81[25] , \ScanLink179[27] , \ScanLink189[3] , 
        \Level2Out50[2] , \Level4Out8[25] , \ScanLink94[11] , 
        \ScanLink119[23] , \ScanLink65[7] , \Level1Out96[19] , 
        \Level1Out109[22] , \Level1Out206[7] , \Level2Out82[4] , 
        \Level2Out110[13] , \Level2Out146[12] , \Level1Out66[14] , 
        \Level1Out166[2] , \Level1Out169[26] , \Level2Out126[16] , 
        \Level1Out229[18] , \Level2Out170[17] , \ScanLink127[3] , 
        \ScanLink19[1] , \Level1Out25[21] , \Level1Out30[15] , 
        \Level1Out45[25] , \Level2Out230[30] , \Level4Out184[18] , 
        \Level1Out45[4] , \Level2Out230[29] , \Level1Out50[11] , 
        \ScanLink247[6] , \ScanLink27[30] , \ScanLink27[29] , \ScanLink52[19] , 
        \Level1Out73[20] , \Level2Out168[8] , \ScanLink71[31] , 
        \ScanLink71[28] , \Level1Out97[2] , \Level1Out46[7] , \Level1Out94[1] , 
        \ScanLink239[19] , \Level1Out104[8] , \Level2Out176[4] , 
        \Level2Out216[1] , \Level8Out48[14] , \Level16Out0[20] , 
        \Level2Out32[8] , \Level16Out224[18] , \ScanLink3[11] , 
        \Level1Out13[17] , \Level1Out21[0] , \Level1Out88[21] , 
        \ScanLink124[0] , \Level16Out16[25] , \Level1Out119[7] , 
        \ScanLink189[19] , \ScanLink191[1] , \ScanLink244[5] , 
        \Level2Out48[0] , \Level1Out25[12] , \Level2Out180[29] , 
        \Level1Out50[22] , \Level1Out73[13] , \ScanLink143[7] , 
        \Level1Out199[18] , \Level2Out180[30] , \Level4Out92[18] , 
        \Level32Out0[1] , \Level1Out22[3] , \Level1Out30[26] , 
        \Level1Out66[27] , \Level1Out45[16] , \ScanLink223[2] , 
        \Level4Out60[1] , \Level1Out88[12] , \ScanLink140[4] , 
        \Level1Out141[31] , \Level1Out117[29] , \Level1Out162[19] , 
        \Level1Out141[28] , \Level2Out158[19] , \Level1Out117[30] , 
        \Level1Out134[18] , \ScanLink220[1] , \ScanLink192[2] , 
        \Level16Out16[16] , \Level1Out200[9] , \Level1Load0[0] , 
        \Level1Out0[26] , \Level1Out0[15] , \ScanLink5[0] , \ScanLink6[3] , 
        \ScanLink7[20] , \ScanLink63[9] , \ScanLink107[28] , \ScanLink151[30] , 
        \Level2Out82[18] , \Level16Out0[13] , \ScanLink172[18] , 
        \ScanLink151[29] , \Level8Out48[27] , \ScanLink95[9] , 
        \ScanLink107[31] , \Level1Out113[18] , \ScanLink124[19] , 
        \Level1Out130[30] , \Level2Out112[0] , \Level1Out130[29] , 
        \Level1Out159[5] , \Level1Out166[28] , \Level1Out145[19] , 
        \Level1Out166[31] , \ScanLink204[7] , \ScanLink88[6] , 
        \Level1Out99[17] , \ScanLink164[2] , \Level1Out239[0] , 
        \ScanLink219[8] , \Level2Out86[30] , \Level2Out136[6] , 
        \Level2Out86[29] , \ScanLink103[19] , \ScanLink120[31] , 
        \ScanLink120[28] , \ScanLink176[29] , \Level1Out147[9] , 
        \ScanLink155[18] , \ScanLink176[30] , \Level1Out188[0] , 
        \Level4Out96[1] , \Level1Out5[23] , \Level1Out5[10] , \ScanLink7[13] , 
        \Level1Out17[26] , \Level1Out18[9] , \Level1Out21[23] , 
        \Level1Out54[13] , \ScanLink207[4] , \ScanLink59[3] , 
        \Level1Out77[22] , \Level2Out184[18] , \Level4Out44[7] , 
        \Level32Out128[28] , \Level4Out96[30] , \Level1Out62[16] , 
        \Level4Out96[29] , \Level32Out128[31] , \ScanLink167[1] , 
        \Level1Out34[17] , \Level1Out41[27] , \Level2Out152[2] , 
        \Level32Out128[1] , \Level2Out232[7] , \Level1Out17[15] , 
        \Level1Out62[1] , \Level1Out99[24] , \ScanLink100[6] , 
        \Level2Out180[4] , \Level4Out180[29] , \ScanLink20[8] , 
        \Level1Out21[10] , \Level1Out34[24] , \Level1Out62[25] , 
        \Level1Out41[14] , \Level2Out234[18] , \Level4Out180[30] , 
        \Level4Out20[3] , \Level1Out61[2] , \Level1Out54[20] , 
        \Level1Out77[11] , \ScanLink103[5] , \ScanLink23[18] , \ScanLink41[1] , 
        \ScanLink56[31] , \ScanLink56[28] , \ScanLink75[19] , \Level64Out0[9] , 
        \ScanLink85[14] , \Level1Load124[0] , \ScanLink248[18] , 
        \ScanLink202[9] , \Level1Out243[8] , \ScanLink90[20] , \ScanLink93[7] , 
        \ScanLink108[26] , \Level1Out190[2] , \Level2Out98[22] , 
        \Level8Out64[18] , \Level8Out32[19] , \Level1Out92[31] , 
        \ScanLink168[22] , \Level2Out74[4] , \Level1Out92[28] , 
        \Level1Out142[4] , \Level2Out114[22] , \ScanLink42[2] , 
        \Level1Out118[27] , \Level1Out178[23] , \Level1Out222[1] , 
        \Level2Out122[27] , \Level2Out130[8] , \Level2Out142[23] , 
        \Level16Out208[14] , \Level8Out64[9] , \Level1Out253[15] , 
        \Level2Out4[28] , \Level2Out174[26] , \Level4Out88[22] , 
        \Level1Out69[30] , \Level1Out69[29] , \Level1Out183[22] , 
        \Level1Out226[25] , \Level32Out160[22] , \Level1Out141[7] , 
        \Level2Out4[31] , \Level1Out205[14] , \Level1Out210[20] , 
        \Level16Out112[5] , \Level1Out221[2] , \Level16Out160[17] , 
        \ScanLink25[5] , \ScanLink28[14] , \ScanLink90[4] , \Level1Out196[16] , 
        \Level1Out233[11] , \Level1Out246[21] , \Level2Out40[12] , 
        \ScanLink48[10] , \ScanLink186[17] , \Level1Out193[1] , 
        \ScanLink200[21] , \ScanLink256[20] , \ScanLink223[10] , 
        \Level2Out16[13] , \ScanLink193[23] , \ScanLink243[14] , 
        \Level2Out76[17] , \ScanLink236[24] , \ScanLink215[15] , 
        \Level2Out20[16] , \ScanLink26[6] , \ScanLink28[27] , \ScanLink48[23] , 
        \Level1Out79[0] , \Level1Out118[14] , \Level1Out126[0] , 
        \Level2Out122[14] , \Level2Load34[0] , \Level2Out174[15] , 
        \ScanLink85[27] , \ScanLink90[13] , \Level1Out178[10] , 
        \Level1Out246[5] , \Level2Out114[11] , \Level2Out234[9] , 
        \Level2Out142[10] , \Level16Out208[27] , \ScanLink108[15] , 
        \ScanLink168[11] , \Level2Out98[11] , \ScanLink106[8] , 
        \Level2Out10[0] , \ScanLink193[10] , \Level16Out208[8] , 
        \ScanLink236[17] , \ScanLink243[27] , \Level2Out76[24] , 
        \Level1Load58[0] , \ScanLink215[26] , \Level2Out20[25] , 
        \ScanLink200[12] , \Level2Out40[21] , \Level8Out192[6] , 
        \Level16Out16[4] , \Level1Out125[3] , \ScanLink186[24] , 
        \ScanLink223[23] , \Level2Out16[20] , \ScanLink256[13] , 
        \Level1Out210[13] , \Level16Out160[24] , \Level16Out176[1] , 
        \Level1Out196[25] , \Level1Out233[22] , \Level2Out198[6] , 
        \ScanLink38[25] , \ScanLink118[4] , \Level1Out246[12] , 
        \Level1Out183[11] , \ScanLink196[26] , \Level1Out205[27] , 
        \Level1Out226[16] , \Level1Out245[6] , \Level32Out160[11] , 
        \Level1Out253[26] , \Level4Out88[11] , \ScanLink233[21] , 
        \ScanLink246[11] , \ScanLink58[21] , \ScanLink205[24] , 
        \ScanLink210[10] , \Level2Out50[23] , \Level2Out30[27] , 
        \ScanLink183[12] , \ScanLink253[25] , \Level2Out66[26] , 
        \Level1Out215[25] , \ScanLink226[15] , \Level8Out0[20] , 
        \ScanLink11[4] , \ScanLink12[7] , \Level1Out79[18] , 
        \Level1Out193[13] , \Level1Out243[24] , \Level1Out236[14] , 
        \Level1Out82[19] , \Level1Out111[2] , \Level1Out186[27] , 
        \Level1Out223[20] , \Level4Out208[16] , \Level1Out200[11] , 
        \Level2Out4[3] , \Level1Out82[8] , \Level1Out168[12] , 
        \Level4Out16[22] , \Level2Out152[12] , \Level4Out160[15] , 
        \Level4Out136[14] , \Level1Out112[1] , \Level2Out104[13] , 
        \Level2Out200[8] , \Level4Out20[27] , \Level4Out40[23] , 
        \Level2Out164[17] , \Level4Out156[10] , \Level4Out100[11] , 
        \ScanLink76[3] , \ScanLink80[11] , \ScanLink95[25] , 
        \Level1Out108[16] , \Level2Out132[16] , \Level4Out76[26] , 
        \ScanLink132[9] , \ScanLink118[17] , \Level2Out24[1] , 
        \Level2Out88[13] , \ScanLink178[13] , \ScanLink148[1] , 
        \Level1Out175[6] , \Level1Out186[14] , \Level1Out223[13] , 
        \ScanLink187[8] , \Level1Out215[3] , \Level1Out200[22] , 
        \Level4Out208[25] , \Level1Out215[16] , \ScanLink228[4] , 
        \Level1Out193[20] , \Level1Out236[27] , \Level1Out5[4] , 
        \Level1Out6[7] , \ScanLink58[12] , \ScanLink205[17] , 
        \Level1Out243[17] , \Level2Out30[14] , \Level1Out37[9] , 
        \ScanLink183[21] , \ScanLink226[26] , \ScanLink38[16] , 
        \Level1Out168[9] , \ScanLink253[16] , \Level8Out0[13] , 
        \Level2Out66[15] , \ScanLink196[15] , \ScanLink233[12] , 
        \ScanLink210[23] , \ScanLink246[22] , \Level4Out76[8] , 
        \Level32Out160[6] , \ScanLink80[22] , \ScanLink178[20] , 
        \Level2Out50[10] , \ScanLink199[4] , \Level2Out40[5] , \ScanLink9[30] , 
        \ScanLink9[29] , \Level1Out29[5] , \ScanLink95[16] , \ScanLink118[24] , 
        \ScanLink236[8] , \Level128Out128[2] , \Level2Out88[20] , 
        \Level2Out164[24] , \Level4Out156[23] , \Level2Out92[3] , 
        \Level4Out20[14] , \Level1Out108[25] , \Level4Out76[15] , 
        \Level1Out216[0] , \Level2Out132[25] , \Level4Out100[22] , 
        \Level1Out12[23] , \Level1Out67[13] , \ScanLink75[0] , 
        \Level2Out152[21] , \Level1Out168[21] , \Level2Out104[9] , 
        \Level4Out160[26] , \Level4Out16[11] , \Level1Out176[5] , 
        \Level2Out104[20] , \Level4Out40[10] , \Level4Out68[4] , 
        \Level4Out136[27] , \ScanLink137[4] , \Level4Out220[18] , 
        \Level4Out232[5] , \Level1Out31[12] , \Level1Out44[22] , 
        \Level2Out194[30] , \Level64Out192[27] , \Level1Out55[3] , 
        \Level2Out194[29] , \Level4Out0[5] , \Level1Out0[9] , \ScanLink2[25] , 
        \ScanLink14[9] , \Level1Out24[26] , \Level1Out51[16] , 
        \Level32Out96[20] , \Level1Out72[27] , \Level4Out152[0] , 
        \Level1Out87[5] , \Level2Out18[30] , \Level2Out18[29] , 
        \Level4Out180[6] , \Level1Out56[0] , \Level1Load77[0] , 
        \Level1Out84[6] , \Level2Out96[18] , \Level1Out103[30] , 
        \ScanLink113[31] , \ScanLink129[8] , \Level2Out206[6] , 
        \Level8Out32[2] , \ScanLink113[28] , \ScanLink130[19] , 
        \ScanLink145[29] , \Level2Out166[3] , \ScanLink145[30] , 
        \ScanLink166[18] , \Level1Out120[18] , \Level1Out99[9] , 
        \Level1Out155[28] , \Level8Out112[26] , \ScanLink10[18] , 
        \Level1Out89[26] , \Level1Out103[29] , \ScanLink134[7] , 
        \Level1Out155[31] , \Level1Out176[19] , \Level8Out144[27] , 
        \Level1Out109[0] , \ScanLink254[2] , \Level1Out24[15] , 
        \Level1Out31[7] , \ScanLink33[30] , \ScanLink33[29] , \ScanLink65[28] , 
        \Level2Out58[7] , \ScanLink46[19] , \ScanLink181[6] , \ScanLink65[31] , 
        \Level1Out173[8] , \Level1Load214[0] , \Level1Out248[31] , 
        \Level2Out224[29] , \Level1Out51[25] , \Level32Out96[13] , 
        \ScanLink153[0] , \Level1Out248[28] , \Level2Out224[30] , 
        \ScanLink2[16] , \Level1Out12[10] , \Level1Out72[14] , 
        \Level1Out31[21] , \Level1Out67[20] , \Level64Out192[14] , 
        \Level1Out32[4] , \Level1Out44[11] , \ScanLink233[5] , 
        \Level4Out136[4] , \Level1Out89[15] , \ScanLink150[3] , 
        \Level4Out148[31] , \ScanLink230[6] , \Level4Out148[28] , 
        \ScanLink6[27] , \Level1Out16[2] , \Level1Out149[2] , \ScanLink182[5] , 
        \Level8Out112[15] , \Level8Out144[14] , \Level2Out102[7] , 
        \Level4Out128[8] , \Level8Out56[6] , \Level8Out120[21] , 
        \ScanLink214[0] , \Level8Out176[20] , \ScanLink6[14] , \ScanLink8[8] , 
        \ScanLink14[30] , \ScanLink14[29] , \ScanLink42[31] , \ScanLink57[8] , 
        \Level1Out98[10] , \ScanLink174[5] , \Level1Out229[7] , 
        \ScanLink61[19] , \ScanLink98[1] , \Level1Load153[0] , 
        \Level2Out126[1] , \Level2Out246[4] , \Level1Out234[8] , 
        \Level8Out72[0] , \Level8Out80[15] , \Level1Out198[7] , 
        \ScanLink37[18] , \ScanLink42[28] , \Level16Load64[0] , 
        \Level1Out20[24] , \Level1Out55[14] , \Level1Out185[8] , 
        \ScanLink229[31] , \ScanLink229[28] , \Level64Out64[10] , 
        \ScanLink217[3] , \Level1Out239[30] , \Level4Out112[2] , 
        \Level1Out15[1] , \Level1Out16[21] , \ScanLink49[4] , 
        \Level2Out220[18] , \Level1Out63[11] , \Level1Out76[25] , 
        \Level1Out239[29] , \Level2Load142[0] , \ScanLink177[6] , 
        \Level1Out40[20] , \Level16Out64[9] , \Level1Out35[10] , 
        \ScanLink117[19] , \Level1Out130[9] , \Level8Out248[22] , 
        \ScanLink134[31] , \ScanLink134[28] , \ScanLink141[18] , 
        \ScanLink162[30] , \Level2Out92[30] , \Level2Out92[29] , 
        \Level2Out142[5] , \Level8Out16[4] , \ScanLink162[29] , 
        \Level2Out222[0] , \Level1Out151[19] , \Level1Out172[31] , 
        \Level1Out16[12] , \Level1Out72[6] , \Level1Out98[23] , 
        \Level1Out124[29] , \Level2Out148[31] , \Level1Out107[18] , 
        \Level1Out124[30] , \Level1Out172[28] , \Level2Out148[28] , 
        \ScanLink110[1] , \Level2Out190[3] , \Level8Out120[12] , 
        \Level8Out176[13] , \Level1Out20[17] , \Level1Out35[23] , 
        \Level1Out63[22] , \Level1Load81[0] , \Level1Out189[29] , 
        \Level4Out224[29] , \Level1Out40[13] , \Level1Out189[30] , 
        \Level2Out190[18] , \Level4Out224[30] , \Level8Out248[11] , 
        \Level1Out71[5] , \Level4Out176[6] , \Level1Out55[27] , 
        \Level1Out76[16] , \ScanLink113[2] , \Level4Out216[3] , 
        \Level64Out64[23] , \ScanLink0[0] , \ScanLink3[3] , \Level1Out4[24] , 
        \Level1Out4[17] , \ScanLink51[6] , \ScanLink83[0] , \ScanLink84[13] , 
        \ScanLink199[31] , \ScanLink199[28] , \Level2Out18[5] , 
        \Level8Out80[26] , \Level16Out160[8] , \ScanLink109[21] , 
        \Level1Out180[5] , \ScanLink91[27] , \Level64Out0[14] , 
        \Level1Out152[3] , \ScanLink169[25] , \Level2Out64[3] , 
        \Level2Out160[15] , \Level4Out24[25] , \Level4Out152[12] , 
        \Level4Out104[13] , \ScanLink52[5] , \Level1Out119[20] , 
        \Level1Out179[24] , \Level1Out232[6] , \Level2Out136[14] , 
        \Level4Out12[20] , \Level4Out72[24] , \Level4Out164[17] , 
        \Level1Out252[12] , \Level2Out100[11] , \Level2Out156[10] , 
        \Level4Out132[16] , \Level4Out44[21] , \Level1Out151[0] , 
        \Level1Out182[25] , \Level1Out227[22] , \Level1Out204[13] , 
        \Level4Out80[8] , \Level1Out211[27] , \Level8Out200[31] , 
        \Level1Out231[5] , \Level1Out247[26] , \ScanLink29[20] , 
        \ScanLink29[13] , \ScanLink80[3] , \Level1Out197[11] , 
        \Level2Out208[16] , \Level8Out200[28] , \Level1Out232[16] , 
        \ScanLink35[2] , \ScanLink49[17] , \ScanLink171[8] , \Level1Out183[6] , 
        \ScanLink201[26] , \Level2Out34[25] , \Level2Out62[24] , 
        \ScanLink187[10] , \ScanLink192[24] , \ScanLink222[17] , 
        \ScanLink237[23] , \ScanLink242[13] , \Level32Out224[5] , 
        \Level2Out54[21] , \ScanLink214[12] , \Level2Out156[23] , 
        \Level4Out164[24] , \ScanLink49[24] , \Level1Out69[7] , 
        \Level1Out86[31] , \Level1Out86[28] , \Level1Out119[13] , 
        \Level4Out12[13] , \Level1Out136[7] , \Level4Out44[12] , 
        \Level4Out28[6] , \Level2Out100[22] , \Level2Out160[26] , 
        \Level4Out132[25] , \Level4Out152[21] , \Level1Out74[8] , 
        \ScanLink91[14] , \Level1Out179[17] , \Level2Out136[27] , 
        \Level4Out24[16] , \Level4Out72[17] , \Level8Out168[18] , 
        \Level4Out104[20] , \Level64Out0[27] , \ScanLink109[12] , 
        \ScanLink169[16] , \ScanLink84[20] , \ScanLink192[17] , 
        \ScanLink237[10] , \ScanLink242[20] , \ScanLink201[15] , 
        \ScanLink214[21] , \Level2Out34[16] , \Level2Out54[12] , 
        \ScanLink36[1] , \Level1Out135[4] , \ScanLink187[23] , 
        \ScanLink222[24] , \Level2Out62[17] , \Level1Out211[14] , 
        \Level1Out197[22] , \Level1Out232[25] , \Level1Out247[15] , 
        \Level2Out188[1] , \Level2Out208[25] , \ScanLink15[23] , 
        \ScanLink15[10] , \ScanLink20[5] , \ScanLink75[14] , \ScanLink108[3] , 
        \Level1Out123[0] , \Level1Out182[16] , \Level1Out227[11] , 
        \Level1Out204[20] , \Level1Out252[21] , \Level1Out255[1] , 
        \ScanLink228[11] , \Level2Out68[22] , \Level64Out0[4] , 
        \ScanLink23[15] , \ScanLink36[21] , \ScanLink56[25] , \ScanLink43[11] , 
        \Level1Out243[5] , \Level1Out17[18] , \Level1Out34[29] , 
        \ScanLink60[20] , \ScanLink248[15] , \ScanLink198[22] , 
        \Level2Out234[15] , \Level1Out41[19] , \Level1Out62[31] , 
        \Level4Out180[24] , \ScanLink23[6] , \Level1Out34[30] , 
        \Level1Out62[28] , \Level16Out128[23] , \Level1Out99[30] , 
        \Level1Out99[29] , \ScanLink103[8] , \Level1Out188[23] , 
        \Level1Out173[22] , \Level1Out238[10] , \Level2Out202[10] , 
        \Level4Out96[17] , \Level2Out184[26] , \Level32Out128[16] , 
        \Level2Out254[11] , \Level1Out106[12] , \Level1Out150[13] , 
        \Level2Out180[9] , \Level1Out113[26] , \Level1Out125[23] , 
        \Level1Out130[17] , \Level1Out145[27] , \Level1Out166[16] , 
        \Level2Out16[3] , \Level16Out240[20] , \ScanLink155[26] , 
        \ScanLink36[12] , \ScanLink43[22] , \ScanLink96[7] , \ScanLink103[27] , 
        \ScanLink120[16] , \Level1Out120[3] , \ScanLink176[17] , 
        \ScanLink116[13] , \ScanLink163[23] , \Level4Load168[0] , 
        \ScanLink135[22] , \ScanLink140[12] , \Level1Out240[6] , 
        \Level2Out86[17] , \Level1Out188[10] , \Level1Out195[2] , 
        \ScanLink207[9] , \Level1Out238[23] , \Level2Out128[7] , 
        \Level2Out202[23] , \Level4Out96[24] , \Level2Out184[15] , 
        \Level2Out254[22] , \Level2Out234[26] , \Level32Out128[25] , 
        \Level2Out248[2] , \Level4Out180[17] , \Level16Out128[10] , 
        \ScanLink44[1] , \ScanLink60[13] , \Level1Out147[4] , 
        \ScanLink198[11] , \Level1Out18[4] , \ScanLink75[27] , 
        \ScanLink228[22] , \ScanLink248[26] , \ScanLink23[26] , 
        \ScanLink56[16] , \Level1Out227[1] , \Level2Out68[11] , 
        \ScanLink25[8] , \ScanLink38[7] , \ScanLink47[2] , \ScanLink116[20] , 
        \Level1Out144[7] , \ScanLink163[10] , \ScanLink219[5] , 
        \Level2Out86[24] , \Level1Out67[1] , \Level1Out69[17] , 
        \ScanLink95[4] , \ScanLink103[14] , \ScanLink120[25] , 
        \ScanLink135[11] , \ScanLink140[21] , \ScanLink179[0] , 
        \ScanLink155[15] , \Level1Out224[2] , \Level1Out130[24] , 
        \Level1Out159[8] , \ScanLink176[24] , \Level16Out240[13] , 
        \Level1Out145[14] , \Level1Out196[1] , \Level4Out88[0] , 
        \Level1Out106[21] , \Level1Out113[15] , \Level1Out166[25] , 
        \Level1Out125[10] , \Level1Out173[11] , \Level1Out150[20] , 
        \Level2Out72[7] , \Level1Out196[31] , \Level1Out196[28] , 
        \Level16Load16[0] , \Level16Out160[30] , \Level8Out192[13] , 
        \Level16Out160[29] , \ScanLink118[9] , \Level1Out138[1] , 
        \Level2Out4[16] , \Level2Out20[28] , \Level2Load130[0] , 
        \Level2Out76[30] , \Level2Out20[31] , \Level2Out76[29] , 
        \Level4Out160[2] , \ScanLink105[6] , \ScanLink186[29] , 
        \ScanLink186[30] , \Level4Out200[7] , \Level16Out16[9] , 
        \Level16Load240[0] , \Level1Out64[2] , \ScanLink106[5] , 
        \Level2Out186[7] , \ScanLink108[18] , \Level8Out32[27] , 
        \Level16Out208[5] , \Level1Out118[19] , \Level2Out174[18] , 
        \Level8Out64[26] , \ScanLink28[19] , \Level1Out87[22] , 
        \Level2Out122[19] , \Level2Out154[1] , \ScanLink90[9] , 
        \Level1Out92[16] , \Level1Out246[8] , \Level1Load121[0] , 
        \ScanLink201[7] , \Level2Out234[4] , \Level4Out104[6] , 
        \ScanLink161[2] , \Level1Out205[19] , \ScanLink215[18] , 
        \ScanLink236[30] , \ScanLink236[29] , \ScanLink243[19] , 
        \Level1Out226[31] , \Level8Out192[20] , \Level1Out69[24] , 
        \Level1Out226[28] , \Level1Out253[18] , \Level16Out112[8] , 
        \Level2Out4[25] , \Level1Out92[25] , \Level16Out208[19] , 
        \Level1Out142[9] , \Level2Out130[5] , \ScanLink8[23] , \Level1Out8[1] , 
        \ScanLink85[19] , \Level1Out87[11] , \Level2Out250[0] , 
        \Level8Out32[14] , \Level8Out64[4] , \Level8Out64[15] , 
        \Level1Out96[14] , \ScanLink162[1] , \ScanLink202[4] , 
        \Level2Out74[9] , \ScanLink194[1] , \Level8Out40[2] , \Level2Out82[9] , 
        \Level16Out48[7] , \ScanLink8[10] , \Level1Out18[25] , 
        \Level1Out24[0] , \ScanLink81[31] , \Level1Out83[20] , 
        \Level2Out114[3] , \ScanLink146[7] , \Level4Out8[28] , 
        \Level1Out27[3] , \ScanLink78[5] , \ScanLink81[28] , \Level4Out8[31] , 
        \ScanLink226[2] , \Level16Out128[2] , \Level8Out56[21] , 
        \ScanLink59[18] , \ScanLink145[4] , \Level1Out218[6] , 
        \Level1Out178[3] , \ScanLink211[29] , \Level4Out240[5] , 
        \ScanLink247[31] , \ScanLink197[2] , \Level1Out201[31] , 
        \Level1Out201[28] , \ScanLink211[30] , \ScanLink225[1] , 
        \ScanLink232[18] , \ScanLink247[28] , \Level4Out120[0] , 
        \Level1Out222[19] , \Level64Out64[3] , \Level1Out205[9] , 
        \Level2Out0[14] , \Level2Out218[19] , \Level1Out40[4] , 
        \ScanLink66[9] , \Level1Out78[21] , \Level1Out83[13] , 
        \Level1Out92[2] , \ScanLink122[3] , \Level8Out56[12] , 
        \ScanLink179[19] , \ScanLink242[6] , \Level2Out126[31] , 
        \Level1Out169[18] , \Level2Out170[29] , \Level2Out210[2] , 
        \Level1Out96[27] , \Level2Out126[28] , \Level2Out170[30] , 
        \Level8Out24[6] , \Level2Out170[7] , \Level1Out18[16] , 
        \Level1Out78[12] , \Level1Out91[1] , \Level1Out192[19] , 
        \Level1Out101[8] , \Level4Out196[2] , \Level1Out43[7] , 
        \ScanLink121[0] , \Level2Out0[27] , \Level2Out24[19] , 
        \Level4Out224[1] , \Level2Out72[18] , \ScanLink63[4] , 
        \ScanLink112[11] , \ScanLink167[21] , \ScanLink182[18] , 
        \ScanLink241[5] , \Level4Out144[4] , \Level2Out82[15] , 
        \Level2Out84[7] , \ScanLink131[20] , \ScanLink144[10] , 
        \Level1Out200[4] , \ScanLink151[24] , \Level2Load168[0] , 
        \Level1Out102[10] , \ScanLink107[25] , \ScanLink124[14] , 
        \Level1Out160[1] , \ScanLink172[15] , \Level1Out117[24] , 
        \Level1Out134[15] , \Level1Out141[25] , \ScanLink140[9] , 
        \Level1Out162[14] , \Level2Out56[1] , \Level32Out224[13] , 
        \Level2Out158[14] , \Level1Out177[20] , \Level2Out138[10] , 
        \Level1Out121[21] , \Level1Out154[11] , \Level16Out224[26] , 
        \Level1Out249[22] , \Level2Out206[12] , \Level4Out92[15] , 
        \ScanLink11[21] , \ScanLink11[12] , \ScanLink32[23] , 
        \Level1Load179[0] , \Level1Out199[15] , \Level2Out180[24] , 
        \Level1Out229[26] , \Level2Out230[17] , \Level2Out250[13] , 
        \Level4Out184[26] , \ScanLink47[13] , \Level1Out203[7] , 
        \ScanLink27[24] , \ScanLink27[17] , \ScanLink60[7] , \ScanLink64[22] , 
        \ScanLink71[16] , \Level1Out163[2] , \ScanLink239[27] , 
        \ScanLink189[14] , \ScanLink52[27] , \ScanLink52[14] , 
        \Level1Out58[6] , \ScanLink71[25] , \Level1Out89[3] , 
        \Level1Out102[23] , \Level1Out121[12] , \Level1Out177[13] , 
        \Level16Out16[28] , \Level2Out138[23] , \Level16Out16[31] , 
        \Level1Out104[5] , \ScanLink107[16] , \Level1Out117[17] , 
        \Level1Out134[26] , \Level1Out154[22] , \Level2Out32[5] , 
        \Level16Out224[15] , \ScanLink244[8] , \Level1Out141[16] , 
        \ScanLink124[27] , \Level1Out162[27] , \Level2Out158[27] , 
        \Level32Out224[20] , \ScanLink139[2] , \ScanLink151[17] , 
        \Level8Out48[19] , \ScanLink172[26] , \ScanLink112[22] , 
        \Level2Out82[26] , \ScanLink131[13] , \ScanLink167[12] , 
        \ScanLink144[23] , \Level2Out176[9] , \ScanLink189[27] , 
        \ScanLink32[10] , \ScanLink47[20] , \ScanLink64[11] , 
        \Level1Out107[6] , \ScanLink239[14] , \Level1Out13[30] , 
        \Level1Out30[18] , \Level1Out45[28] , \Level1Out45[9] , 
        \Level2Out230[24] , \Level1Out13[29] , \Level1Out45[31] , 
        \Level1Out66[19] , \Level1Out229[15] , \Level2Out208[0] , 
        \Level4Out184[15] , \ScanLink0[9] , \Level1Out5[14] , \ScanLink28[10] , 
        \ScanLink48[14] , \Level1Out199[26] , \Level1Out249[11] , 
        \Level2Out168[5] , \Level2Out180[17] , \Level2Out206[21] , 
        \Level4Out92[26] , \Level2Out250[20] , \ScanLink90[0] , 
        \ScanLink186[13] , \ScanLink193[27] , \ScanLink215[11] , 
        \Level2Out20[12] , \ScanLink243[10] , \Level2Out76[13] , 
        \Level1Out193[5] , \ScanLink236[20] , \ScanLink256[24] , 
        \ScanLink223[14] , \Level2Out16[17] , \Level2Out40[16] , 
        \ScanLink200[25] , \Level1Out221[6] , \Level1Out246[25] , 
        \ScanLink41[5] , \ScanLink42[6] , \Level1Out141[3] , 
        \Level1Out196[12] , \Level1Out233[15] , \Level1Out210[24] , 
        \Level16Out160[13] , \Level1Out205[10] , \Level1Out253[11] , 
        \Level4Out88[26] , \Level8Out192[29] , \Level16Out112[1] , 
        \Level1Out87[18] , \Level1Out183[26] , \Level1Out226[21] , 
        \Level2Out122[23] , \Level2Out174[22] , \Level2Out250[9] , 
        \Level8Out192[30] , \Level32Out160[26] , \Level1Out118[23] , 
        \Level1Out222[5] , \Level1Out142[0] , \Level1Out178[27] , 
        \Level2Load50[0] , \Level2Out142[27] , \Level16Out208[10] , 
        \Level2Out114[26] , \ScanLink3[26] , \ScanLink5[4] , \Level1Out5[27] , 
        \ScanLink26[2] , \ScanLink85[10] , \ScanLink90[24] , \ScanLink93[3] , 
        \ScanLink162[8] , \ScanLink168[26] , \Level2Out74[0] , 
        \ScanLink108[22] , \Level1Out190[6] , \ScanLink118[0] , 
        \Level1Out205[23] , \Level2Out98[26] , \Level1Out183[15] , 
        \Level1Out226[12] , \Level1Out245[2] , \Level32Out160[15] , 
        \Level1Out253[22] , \Level4Out88[15] , \Level1Out196[21] , 
        \Level1Out233[26] , \Level1Out246[16] , \Level2Out198[2] , 
        \Level1Out17[22] , \ScanLink25[1] , \ScanLink28[23] , \Level1Out67[8] , 
        \Level1Out125[7] , \ScanLink186[20] , \Level1Out210[17] , 
        \Level16Out160[20] , \ScanLink223[27] , \Level16Out176[5] , 
        \Level2Out16[24] , \ScanLink200[16] , \ScanLink256[17] , 
        \Level2Out40[25] , \Level8Out192[2] , \Level16Out16[0] , 
        \ScanLink48[27] , \Level1Out79[4] , \ScanLink85[23] , 
        \ScanLink108[11] , \Level1Out138[8] , \ScanLink215[22] , 
        \Level2Out20[21] , \ScanLink193[14] , \ScanLink236[13] , 
        \ScanLink243[23] , \Level2Out76[20] , \Level2Out10[4] , 
        \Level2Out98[15] , \ScanLink90[17] , \ScanLink168[15] , 
        \Level1Out178[14] , \Level1Out246[1] , \Level2Out142[14] , 
        \Level16Out208[23] , \Level1Out118[10] , \Level1Out126[4] , 
        \Level2Out114[15] , \Level2Out174[11] , \Level1Out34[13] , 
        \Level1Out41[23] , \Level2Out122[10] , \Level2Out154[8] , 
        \Level1Out62[12] , \Level1Out188[19] , \ScanLink167[5] , 
        \Level1Out21[27] , \Level1Out54[17] , \ScanLink59[7] , 
        \Level16Out128[19] , \Level1Out77[26] , \ScanLink207[0] , 
        \ScanLink44[8] , \Level1Load140[0] , \Level2Out68[18] , 
        \Level4Out44[3] , \Level1Out227[8] , \Level1Out188[4] , 
        \ScanLink198[18] , \Level4Out96[5] , \ScanLink6[7] , \ScanLink116[29] , 
        \ScanLink179[9] , \ScanLink7[24] , \ScanLink88[2] , \ScanLink140[31] , 
        \ScanLink163[19] , \Level1Out99[13] , \Level1Out106[28] , 
        \ScanLink116[30] , \ScanLink135[18] , \ScanLink140[28] , 
        \Level2Out136[2] , \Level1Out150[30] , \ScanLink164[6] , 
        \Level1Out239[4] , \Level1Out106[31] , \Level1Out173[18] , 
        \Level1Out125[19] , \Level1Out150[29] , \ScanLink7[17] , 
        \ScanLink15[19] , \ScanLink36[28] , \Level1Out159[1] , 
        \Level1Out196[8] , \ScanLink204[3] , \Level4Out88[9] , 
        \ScanLink43[18] , \ScanLink60[30] , \Level1Out17[11] , 
        \Level1Out21[14] , \ScanLink36[31] , \ScanLink60[29] , 
        \Level1Out61[6] , \Level1Out77[15] , \ScanLink103[1] , 
        \Level1Out123[9] , \ScanLink228[18] , \Level1Out238[19] , 
        \Level2Out202[19] , \Level1Out34[20] , \Level1Out54[24] , 
        \Level2Out254[18] , \Level1Out41[10] , \Level4Out20[7] , 
        \Level1Out62[21] , \Level4Load216[0] , \Level1Out62[5] , 
        \Level1Load92[0] , \Level1Out99[20] , \ScanLink100[2] , 
        \Level16Out240[29] , \Level16Out240[30] , \Level2Out180[0] , 
        \Level1Out46[3] , \Level1Out88[25] , \Level1Out119[3] , 
        \Level2Out152[6] , \Level2Out232[3] , \Level32Out128[5] , 
        \ScanLink244[1] , \Level32Out224[30] , \Level32Out224[29] , 
        \ScanLink124[4] , \Level16Out16[21] , \ScanLink11[31] , 
        \ScanLink32[19] , \ScanLink47[29] , \Level1Load64[0] , 
        \Level2Out176[0] , \Level16Out0[24] , \Level1Out94[5] , 
        \Level8Out48[10] , \Level2Out216[5] , \ScanLink11[28] , 
        \ScanLink47[30] , \ScanLink64[18] , \Level1Out97[6] , 
        \Level1Out13[20] , \ScanLink19[5] , \Level1Out73[24] , 
        \Level2Out250[30] , \Level1Out25[25] , \Level1Out50[15] , 
        \ScanLink247[2] , \Level1Out249[18] , \Level2Out206[28] , 
        \Level2Out250[29] , \Level1Out30[11] , \Level1Out45[21] , 
        \Level2Out206[31] , \Level1Out45[0] , \Level1Out66[10] , 
        \Level2Out208[9] , \ScanLink127[7] , \Level1Out160[8] , 
        \Level1Load207[0] , \Level8Out48[23] , \Level2Out112[4] , 
        \ScanLink167[28] , \Level1Out0[0] , \Level1Out1[25] , \Level1Out1[16] , 
        \ScanLink3[15] , \Level1Out102[19] , \ScanLink112[18] , 
        \ScanLink131[30] , \Level16Out0[17] , \Level1Out121[31] , 
        \ScanLink131[29] , \ScanLink144[19] , \ScanLink167[31] , 
        \ScanLink192[6] , \Level1Out177[29] , \Level2Out138[19] , 
        \Level1Out154[18] , \Level1Out177[30] , \Level16Out16[12] , 
        \ScanLink220[5] , \ScanLink8[19] , \Level1Out13[13] , \Level1Out22[7] , 
        \Level1Out121[28] , \Level1Out30[22] , \Level1Out88[16] , 
        \ScanLink140[0] , \Level2Out56[8] , \Level1Out45[12] , 
        \ScanLink223[6] , \Level4Out60[5] , \Level1Out21[4] , 
        \Level1Out66[23] , \Level1Out73[17] , \ScanLink143[3] , 
        \Level32Out0[5] , \Level1Out25[16] , \Level2Load216[0] , 
        \Level1Out50[26] , \ScanLink81[12] , \ScanLink179[10] , 
        \ScanLink191[5] , \Level2Out48[4] , \Level4Out8[12] , \ScanLink94[26] , 
        \Level4Out188[7] , \Level1Out102[2] , \Level1Out109[15] , 
        \Level1Load118[0] , \Level2Out34[2] , \ScanLink119[14] , 
        \Level2Out146[25] , \Level2Out110[24] , \Level1Out101[1] , 
        \Level1Out169[11] , \Level2Out126[21] , \Level2Out170[20] , 
        \Level4Out8[4] , \Level1Out187[24] , \Level1Out201[12] , 
        \Level2Out218[23] , \Level1Out222[23] , \Level1Out8[8] , 
        \ScanLink39[26] , \ScanLink59[22] , \Level1Out91[8] , 
        \Level1Out192[10] , \Level1Out237[17] , \Level1Out242[27] , 
        \ScanLink182[11] , \Level1Out214[26] , \ScanLink227[16] , 
        \ScanLink252[26] , \Level2Out12[15] , \ScanLink204[27] , 
        \Level2Out44[14] , \ScanLink65[3] , \Level1Out83[30] , 
        \ScanLink121[9] , \Level1Out166[6] , \ScanLink197[25] , 
        \ScanLink211[13] , \Level4Out224[8] , \Level16Out32[6] , 
        \ScanLink247[12] , \Level2Out24[10] , \Level2Out72[11] , 
        \ScanLink232[22] , \Level2Out170[13] , \Level1Out83[29] , 
        \Level1Out109[26] , \Level1Out169[22] , \Level2Out126[12] , 
        \ScanLink194[8] , \Level1Out206[3] , \Level2Out146[16] , 
        \Level1Out24[9] , \Level1Out39[6] , \ScanLink94[15] , 
        \ScanLink119[27] , \Level2Out82[0] , \Level2Out110[17] , 
        \ScanLink189[7] , \Level8Out56[31] , \Level8Out56[28] , 
        \Level4Out8[21] , \ScanLink39[15] , \ScanLink81[21] , 
        \ScanLink179[23] , \Level2Out50[6] , \ScanLink211[20] , 
        \Level2Out24[23] , \ScanLink59[11] , \ScanLink182[22] , 
        \ScanLink197[16] , \ScanLink225[8] , \ScanLink227[25] , 
        \ScanLink232[11] , \ScanLink247[21] , \Level4Out120[9] , 
        \Level2Out12[26] , \Level2Out72[22] , \ScanLink204[14] , 
        \ScanLink252[15] , \ScanLink66[0] , \Level2Out44[27] , 
        \Level1Out78[28] , \Level1Out192[23] , \Level1Out237[24] , 
        \ScanLink10[11] , \ScanLink26[14] , \ScanLink70[4] , \Level1Out78[31] , 
        \Level1Out165[5] , \Level1Out242[14] , \ScanLink238[7] , 
        \ScanLink158[2] , \Level1Out201[21] , \Level1Out214[15] , 
        \Level1Out187[17] , \Level1Out205[0] , \Level1Out222[10] , 
        \Level2Out218[10] , \ScanLink53[24] , \ScanLink70[15] , 
        \Level1Out173[1] , \ScanLink188[17] , \Level2Out18[13] , 
        \Level1Out12[19] , \ScanLink33[20] , \ScanLink65[21] , 
        \Level2Out78[17] , \ScanLink238[24] , \ScanLink46[10] , 
        \Level1Out213[4] , \Level16Out240[6] , \Level1Out31[31] , 
        \Level2Out212[25] , \Level4Out220[22] , \Level1Out31[28] , 
        \Level1Out67[29] , \Level1Out228[25] , \Level2Out194[13] , 
        \Level1Out44[18] , \Level1Out67[30] , \ScanLink153[9] , 
        \Level2Out224[20] , \Level2Out244[24] , \Level4Out216[27] , 
        \Level1Out198[16] , \Level1Out248[21] , \Level8Out48[3] , 
        \Level4Out240[26] , \ScanLink0[19] , \Level1Out3[3] , 
        \Level1Out103[13] , \Level1Out120[22] , \Level1Out155[12] , 
        \Level4Out128[25] , \Level1Out176[23] , \Level1Out163[17] , 
        \ScanLink8[1] , \ScanLink9[20] , \ScanLink10[22] , \ScanLink65[12] , 
        \ScanLink73[7] , \ScanLink106[26] , \Level1Out116[27] , 
        \Level4Out68[17] , \Level1Out135[16] , \Level1Out140[26] , 
        \Level1Out170[2] , \ScanLink173[16] , \Level2Out46[2] , 
        \Level4Out148[21] , \Level2Out96[22] , \ScanLink150[27] , 
        \Level4Out128[1] , \ScanLink113[12] , \ScanLink125[17] , 
        \ScanLink130[23] , \ScanLink145[13] , \Level1Out210[7] , 
        \Level4Out248[4] , \ScanLink166[22] , \Level2Out94[4] , 
        \Level1Out198[25] , \Level2Out224[13] , \Level32Out96[29] , 
        \Level4Out152[9] , \Level4Out216[14] , \Level4Out240[15] , 
        \Level32Out96[30] , \Level1Out228[16] , \Level1Out248[12] , 
        \Level2Out178[6] , \Level2Out194[20] , \Level2Out212[16] , 
        \Level2Out244[17] , \Level4Out220[11] , \Level2Out218[3] , 
        \Level1Out117[5] , \ScanLink238[17] , \ScanLink14[0] , 
        \ScanLink46[23] , \Level2Out78[24] , \Level16Out144[7] , 
        \Level1Load16[0] , \ScanLink17[3] , \ScanLink26[27] , \ScanLink33[13] , 
        \ScanLink53[17] , \Level16Out224[2] , \Level1Out48[5] , 
        \ScanLink70[26] , \ScanLink188[24] , \Level2Out18[20] , 
        \Level1Out19[26] , \Level1Out56[9] , \ScanLink106[15] , 
        \ScanLink113[21] , \Level1Out114[6] , \ScanLink130[10] , 
        \ScanLink145[20] , \ScanLink249[4] , \ScanLink166[11] , 
        \Level2Out96[11] , \Level1Out109[9] , \Level1Out116[14] , 
        \ScanLink125[24] , \ScanLink173[25] , \ScanLink129[1] , 
        \Level2Out2[4] , \ScanLink150[14] , \Level4Out68[24] , 
        \Level1Out163[24] , \Level1Out135[25] , \Level1Out140[15] , 
        \Level4Out148[12] , \Level1Out79[22] , \Level1Out99[0] , 
        \Level1Out120[11] , \Level1Out103[20] , \Level1Out155[21] , 
        \Level2Out22[6] , \Level4Out128[16] , \Level1Out176[10] , 
        \Level1Out193[30] , \ScanLink148[8] , \Level1Out193[29] , 
        \ScanLink187[1] , \Level1Out34[3] , \Level1Out37[0] , \ScanLink155[7] , 
        \Level1Out168[0] , \Level8Out232[15] , \ScanLink235[2] , 
        \Level2Out50[19] , \Level4Out76[1] , \ScanLink183[31] , 
        \Level1Out208[5] , \ScanLink68[6] , \ScanLink183[28] , 
        \Level2Out88[30] , \ScanLink236[1] , \Level2Out88[29] , 
        \ScanLink75[9] , \ScanLink156[4] , \ScanLink178[29] , 
        \ScanLink178[30] , \Level2Out152[28] , \Level1Out82[23] , 
        \Level1Out168[28] , \Level2Out104[0] , \Level4Out16[18] , 
        \Level1Out168[31] , \Level2Out104[30] , \Level2Out152[31] , 
        \Level4Out40[19] , \Level2Load8[0] , \Level2Out104[29] , 
        \ScanLink9[13] , \Level1Out19[15] , \Level1Out53[4] , \ScanLink58[31] , 
        \ScanLink58[28] , \Level1Out97[17] , \ScanLink184[2] , 
        \Level1Out216[9] , \ScanLink251[6] , \Level8Out0[30] , 
        \ScanLink246[18] , \Level4Out12[5] , \Level8Out0[29] , 
        \ScanLink131[3] , \ScanLink233[28] , \ScanLink210[19] , 
        \ScanLink233[31] , \Level1Out79[11] , \Level1Out81[2] , 
        \Level1Out200[18] , \Level1Out223[29] , \Level1Out223[30] , 
        \Level8Out232[26] , \Level1Out112[8] , \Level1Out10[5] , 
        \ScanLink28[4] , \Level1Out50[7] , \ScanLink80[18] , \Level1Out82[10] , 
        \Level1Out97[24] , \Level4Out100[18] , \Level4Out156[19] , 
        \Level2Out160[4] , \Level1Out82[1] , \ScanLink252[5] , 
        \Level2Out200[1] , \ScanLink132[0] , \Level1Out74[1] , 
        \Level1Out86[21] , \Level1Out93[15] , \Level2Out24[8] , 
        \Level2Out224[7] , \Level4Out104[30] , \Level4Out152[28] , 
        \Level4Out152[31] , \Level8Out168[11] , \Level2Out144[2] , 
        \Level4Out104[29] , \ScanLink84[30] , \ScanLink84[29] , 
        \ScanLink116[6] , \ScanLink29[30] , \ScanLink29[29] , \ScanLink115[5] , 
        \Level2Out196[4] , \Level1Out248[7] , \Level1Out77[2] , 
        \ScanLink36[8] , \Level1Out68[14] , \Level1Out128[2] , 
        \ScanLink214[31] , \ScanLink237[19] , \ScanLink214[28] , 
        \ScanLink242[29] , \Level4Out36[3] , \Level1Out227[18] , 
        \ScanLink242[30] , \Level1Load132[0] , \Level1Out204[30] , 
        \Level1Out204[29] , \Level1Out252[28] , \Level1Out255[8] , 
        \Level16Out96[14] , \Level1Out252[31] , \Level32Out96[6] , 
        \ScanLink172[2] , \Level2Out188[8] , \Level8Out200[12] , 
        \Level1Out13[6] , \Level1Out68[27] , \ScanLink83[9] , 
        \ScanLink109[28] , \ScanLink212[7] , \Level1Out86[12] , 
        \ScanLink109[31] , \Level1Out93[26] , \Level1Out119[30] , 
        \Level1Out119[29] , \Level2Out156[19] , \Level4Out12[29] , 
        \Level4Out44[31] , \Level2Out100[18] , \Level2Out240[3] , 
        \Level4Out12[30] , \Level4Out44[28] , \Level8Out168[22] , 
        \Level1Out197[18] , \Level2Out120[6] , \Level8Out200[21] , 
        \Level1Out151[9] , \Level16Out96[27] , \Level2Out54[31] , 
        \Level4Out80[1] , \ScanLink14[20] , \ScanLink14[13] , \ScanLink33[5] , 
        \ScanLink102[24] , \ScanLink117[10] , \ScanLink134[21] , 
        \ScanLink141[11] , \ScanLink171[1] , \Level2Out54[28] , 
        \ScanLink187[19] , \ScanLink211[4] , \Level1Out250[5] , 
        \Level4Out52[7] , \Level4Out208[6] , \ScanLink162[20] , 
        \Level1Out130[0] , \ScanLink177[14] , \Level2Out222[9] , 
        \Level2Load22[0] , \ScanLink154[25] , \Level2Out92[20] , 
        \Level64Out192[7] , \Level4Out168[3] , \Level1Out107[11] , 
        \ScanLink110[8] , \ScanLink121[15] , \Level1Out167[15] , 
        \Level2Out128[25] , \Level1Out112[25] , \Level1Out124[20] , 
        \Level1Out131[14] , \Level1Out144[24] , \Level1Out151[10] , 
        \Level1Out172[21] , \Level1Out189[20] , \Level1Out239[13] , 
        \Level2Out148[21] , \Level2Out220[22] , \Level4Out212[25] , 
        \Level8Out184[6] , \Level2Out216[27] , \Level4Out224[20] , 
        \Level4Out244[24] , \Level2Out190[11] , \Level2Out240[26] , 
        \Level8Out248[18] , \ScanLink22[25] , \ScanLink22[16] , 
        \ScanLink30[6] , \ScanLink37[22] , \ScanLink61[23] , \ScanLink249[16] , 
        \ScanLink199[21] , \ScanLink42[12] , \Level1Out253[6] , 
        \ScanLink57[26] , \ScanLink57[15] , \ScanLink57[1] , \ScanLink74[17] , 
        \Level1Out133[3] , \ScanLink229[12] , \Level16Out160[1] , 
        \ScanLink85[7] , \Level1Out98[19] , \Level1Out107[22] , 
        \Level1Out124[13] , \Level1Out151[23] , \Level2Out62[4] , 
        \Level2Out148[12] , \Level1Out172[12] , \Level1Out112[16] , 
        \Level8Out120[28] , \ScanLink102[17] , \Level1Out131[27] , 
        \Level1Out167[26] , \Level2Out128[16] , \Level8Out176[30] , 
        \ScanLink214[9] , \Level8Out120[31] , \Level1Out144[17] , 
        \Level1Out186[2] , \Level8Out176[29] , \ScanLink121[26] , 
        \ScanLink169[3] , \ScanLink177[27] , \Level2Out92[13] , 
        \ScanLink154[16] , \Level1Out234[1] , \Level8Out72[9] , 
        \ScanLink98[8] , \ScanLink134[12] , \ScanLink117[23] , 
        \ScanLink141[22] , \Level1Out154[4] , \Level2Out126[8] , 
        \ScanLink162[13] , \ScanLink209[6] , \Level1Out237[2] , 
        \Level64Out64[19] , \ScanLink61[10] , \ScanLink74[24] , 
        \ScanLink229[21] , \Level1Out157[7] , \ScanLink199[12] , 
        \Level1Out15[8] , \Level1Out16[28] , \ScanLink37[11] , 
        \ScanLink42[21] , \ScanLink249[25] , \ScanLink54[2] , 
        \Level1Out40[30] , \Level1Out63[18] , \Level1Out189[13] , 
        \Level2Out216[14] , \Level4Out224[13] , \Level1Out40[29] , 
        \Level2Out240[15] , \Level16Out64[0] , \Level1Out16[31] , 
        \Level1Out35[19] , \Level1Out185[1] , \Level2Out190[22] , 
        \Level2Out220[11] , \Level1Out9[25] , \Level1Out26[30] , 
        \Level1Out26[29] , \Level1Out53[19] , \Level1Out70[31] , 
        \ScanLink86[4] , \Level4Out212[16] , \Level1Out209[21] , 
        \Level1Out239[20] , \Level2Out138[4] , \Level4Out244[17] , 
        \Level2Out210[10] , \Level4Out84[17] , \Level2Out196[26] , 
        \Level2Out238[5] , \Level2Out246[11] , \ScanLink29[9] , 
        \Level2Out226[15] , \Level1Out70[28] , \Level1Out9[16] , 
        \Level1Out11[8] , \ScanLink12[24] , \ScanLink24[21] , \ScanLink51[11] , 
        \Level2Out158[0] , \Level4Out192[24] , \Level8Out152[0] , 
        \ScanLink67[14] , \Level1Out68[3] , \ScanLink72[20] , 
        \Level1Out137[3] , \Level8Out232[5] , \ScanLink12[17] , 
        \ScanLink31[15] , \ScanLink34[6] , \ScanLink219[20] , \ScanLink44[25] , 
        \ScanLink37[5] , \ScanLink89[21] , \ScanLink104[13] , 
        \Level2Out94[17] , \ScanLink109[7] , \ScanLink127[22] , 
        \ScanLink171[23] , \Level1Out254[5] , \Level2Out226[9] , 
        \Level4Out0[21] , \ScanLink132[16] , \ScanLink152[12] , 
        \Level1Out101[26] , \ScanLink111[27] , \ScanLink147[26] , 
        \Level1Out122[17] , \Level1Out134[0] , \ScanLink164[17] , 
        \Level2Load26[0] , \Level1Out157[27] , \Level2Out118[17] , 
        \ScanLink114[8] , \Level1Out114[12] , \Level1Out174[16] , 
        \Level1Out137[23] , \Level1Out161[22] , \Level1Out142[13] , 
        \Level2Out178[13] , \ScanLink24[12] , \ScanLink31[26] , 
        \ScanLink67[27] , \Level1Out233[2] , \Level2Out78[8] , 
        \Level8Out136[4] , \ScanLink44[16] , \ScanLink219[13] , 
        \ScanLink50[2] , \ScanLink51[22] , \ScanLink72[13] , \Level1Out153[7] , 
        \Level2Out226[26] , \ScanLink82[4] , \Level4Out192[17] , 
        \Level1Out114[21] , \Level1Out161[11] , \Level1Out181[1] , 
        \Level1Load229[0] , \Level2Out210[23] , \Level4Out84[24] , 
        \Level1Out209[12] , \Level2Out196[15] , \Level2Out246[22] , 
        \Level8Out128[8] , \Level1Out137[10] , \Level1Out142[20] , 
        \Level2Out66[4] , \Level2Out178[20] , \Level1Out2[30] , 
        \ScanLink32[8] , \ScanLink53[1] , \ScanLink81[7] , \Level1Out122[24] , 
        \Level1Out157[14] , \ScanLink210[9] , \Level2Out118[24] , 
        \Level1Out182[2] , \Level1Out174[25] , \ScanLink89[12] , 
        \Level1Out101[15] , \ScanLink111[14] , \ScanLink132[25] , 
        \ScanLink147[15] , \Level1Out230[1] , \ScanLink164[24] , 
        \Level2Load238[0] , \Level1Load198[0] , \ScanLink104[20] , 
        \Level1Out150[4] , \ScanLink171[10] , \Level2Out94[24] , 
        \Level4Out108[7] , \Level1Out58[26] , \Level1Out73[2] , 
        \ScanLink127[11] , \ScanLink152[21] , \Level4Out0[12] , 
        \Level2Out122[8] , \ScanLink111[5] , \ScanLink194[29] , 
        \ScanLink194[30] , \Level2Out32[31] , \Level2Out32[28] , 
        \Level2Out64[30] , \Level2Out64[29] , \Level4Out32[3] , 
        \Level1Load136[0] , \Level1Out251[8] , \Level1Out38[22] , 
        \Level1Out184[28] , \Level1Out38[11] , \Level1Out70[1] , 
        \Level1Out80[16] , \Level1Out184[31] , \Level1Out95[22] , 
        \Level1Out129[28] , \Level2Out220[7] , \Level32Out32[10] , 
        \Level32Out64[11] , \Level128Out0[23] , \Level16Out48[13] , 
        \Level2Out166[18] , \ScanLink112[6] , \Level1Out129[31] , 
        \Level2Out130[19] , \Level2Out140[2] , \ScanLink139[29] , 
        \ScanLink139[30] , \Level2Out192[4] , \Level8Out16[22] , 
        \Level8Out40[23] , \Level1Out58[15] , \Level1Out217[19] , 
        \Level1Out234[31] , \Level2Load88[0] , \Level1Out155[9] , 
        \Level4Out84[1] , \Level1Out2[29] , \ScanLink99[5] , 
        \Level1Out234[28] , \Level1Out241[18] , \ScanLink4[31] , 
        \ScanLink4[28] , \Level1Out6[18] , \Level1Load12[0] , \Level1Out14[5] , 
        \Level1Out17[6] , \ScanLink175[1] , \ScanLink224[30] , 
        \Level1Out228[3] , \ScanLink207[18] , \ScanLink224[29] , 
        \ScanLink19[31] , \ScanLink19[28] , \Level1Out148[6] , 
        \ScanLink215[4] , \ScanLink251[19] , \Level4Out56[7] , 
        \Level1Out30[3] , \ScanLink48[0] , \ScanLink176[2] , \Level8Out16[11] , 
        \Level8Out40[10] , \Level1Out80[25] , \ScanLink87[9] , 
        \Level1Out95[11] , \ScanLink97[19] , \ScanLink216[7] , 
        \Level2Out244[3] , \Level16Out48[20] , \Level32Out32[23] , 
        \Level128Out0[10] , \ScanLink93[31] , \ScanLink152[4] , 
        \Level1Out199[3] , \Level2Out124[6] , \ScanLink232[1] , 
        \Level32Out64[22] , \Level8Out24[25] , \ScanLink71[9] , 
        \Level1Out91[20] , \ScanLink93[28] , \Level8Out72[24] , 
        \Level1Out29[14] , \Level1Out49[10] , \Level1Out84[14] , 
        \ScanLink180[2] , \Level2Out100[0] , \Level1Out212[9] , 
        \Level1Out245[30] , \Level1Out213[28] , \Level8Out184[11] , 
        \Level1Out29[27] , \Level1Out33[0] , \ScanLink183[1] , 
        \Level1Out245[29] , \ScanLink203[30] , \ScanLink203[29] , 
        \Level1Out213[31] , \Level1Out230[19] , \ScanLink255[31] , 
        \ScanLink231[2] , \ScanLink255[28] , \Level4Out72[1] , 
        \ScanLink220[18] , \Level1Out49[8] , \ScanLink68[30] , 
        \ScanLink68[29] , \ScanLink151[7] , \Level2Out88[6] , 
        \Level1Out84[27] , \Level1Out116[8] , \Level2Out164[4] , 
        \Level1Out54[7] , \Level1Out86[1] , \Level2Out162[29] , 
        \Level1Out91[13] , \Level1Out158[30] , \Level1Out158[29] , 
        \Level2Out204[1] , \Level2Out134[31] , \Level2Out162[30] , 
        \Level2Out134[28] , \ScanLink148[31] , \ScanLink148[28] , 
        \Level8Out24[16] , \ScanLink256[5] , \Level8Out72[17] , 
        \Level1Out57[4] , \Level1Out108[4] , \ScanLink136[0] , 
        \Level2Out20[8] , \ScanLink190[18] , \ScanLink255[6] , 
        \Level32Out64[6] , \ScanLink135[3] , \Level2Out36[19] , 
        \Level4Out16[5] , \ScanLink248[9] , \Level2Out60[18] , 
        \Level8Out184[22] , \Level1Out49[23] , \Level1Out85[2] , 
        \Level1Out180[19] , \Level1Out110[10] , \Level16Out176[18] , 
        \Level1Out126[15] , \Level1Out133[21] , \Level1Out165[20] , 
        \Level1Out146[11] , \Level1Out7[3] , \Level1Out105[24] , 
        \Level1Out153[25] , \Level1Out209[8] , \Level2Out42[2] , 
        \Level8Out80[9] , \Level1Out4[0] , \ScanLink16[26] , \ScanLink63[16] , 
        \ScanLink77[7] , \ScanLink136[14] , \Level1Out170[14] , 
        \ScanLink98[17] , \ScanLink115[25] , \ScanLink143[24] , 
        \ScanLink160[15] , \Level1Out174[2] , \ScanLink229[0] , 
        \ScanLink100[11] , \ScanLink123[20] , \ScanLink149[5] , 
        \ScanLink175[21] , \Level2Out90[15] , \Level2Out90[4] , 
        \Level1Out214[7] , \Level4Out4[23] , \ScanLink156[10] , 
        \Level1Out177[1] , \ScanLink20[23] , \ScanLink35[17] , 
        \ScanLink40[27] , \ScanLink74[4] , \Level2Out28[21] , \ScanLink55[13] , 
        \ScanLink208[16] , \Level1Out217[4] , \Level8Out112[2] , 
        \Level16Out96[0] , \Level1Out28[1] , \Level2Out48[25] , 
        \ScanLink76[22] , \ScanLink157[9] , \Level1Out218[17] , 
        \Level2Out118[2] , \Level2Out222[17] , \Level4Out196[26] , 
        \ScanLink198[0] , \Level4Out80[15] , \Level4Out252[8] , 
        \ScanLink13[3] , \ScanLink100[22] , \Level1Out110[6] , 
        \Level2Out192[24] , \Level2Out214[12] , \Level2Out242[13] , 
        \ScanLink175[12] , \Level4Out148[5] , \Level2Out90[26] , 
        \ScanLink1[20] , \ScanLink1[13] , \ScanLink2[7] , \ScanLink5[22] , 
        \ScanLink5[11] , \Level1Out7[21] , \ScanLink10[0] , \ScanLink20[10] , 
        \Level1Out22[18] , \Level1Out52[9] , \ScanLink98[24] , 
        \ScanLink123[13] , \ScanLink156[23] , \Level4Out4[10] , 
        \ScanLink136[27] , \ScanLink143[17] , \Level2Out6[4] , 
        \ScanLink160[26] , \Level4Out228[0] , \Level1Out105[17] , 
        \ScanLink115[16] , \Level1Out126[26] , \Level1Out153[16] , 
        \Level1Out170[27] , \Level1Out110[23] , \Level1Out165[13] , 
        \Level1Out133[12] , \Level1Out146[22] , \Level2Out26[6] , 
        \ScanLink253[8] , \Level2Out214[21] , \Level4Out80[26] , 
        \Level2Out192[17] , \Level2Out222[24] , \Level2Out242[20] , 
        \Level16Out192[1] , \Level4Out156[9] , \Level1Out57[31] , 
        \Level1Out57[28] , \Level1Out218[24] , \Level4Out196[15] , 
        \Level1Out74[19] , \ScanLink16[15] , \ScanLink55[20] , 
        \Level2Out48[16] , \ScanLink76[11] , \Level1Out113[5] , 
        \ScanLink208[25] , \Level8Out216[3] , \ScanLink35[24] , 
        \ScanLink63[25] , \Level8Out176[6] , \ScanLink40[14] , 
        \Level2Out28[12] , \Level1Out194[27] , \Level1Out231[20] , 
        \Level1Out244[10] , \Level1Out7[12] , \ScanLink18[8] , 
        \Level1Out48[30] , \Level1Out48[29] , \Level1Out95[8] , 
        \Level1Out105[1] , \Level1Out212[11] , \Level8Out200[7] , 
        \Level2Out228[11] , \Level1Out207[25] , \Level2Out248[15] , 
        \ScanLink138[6] , \Level1Out181[13] , \Level2Out198[22] , 
        \Level1Out224[14] , \Level8Out160[2] , \ScanLink69[10] , 
        \ScanLink191[12] , \ScanLink217[24] , \Level1Out251[24] , 
        \Level2Out6[19] , \Level2Out22[27] , \ScanLink234[15] , 
        \Level1Out88[7] , \ScanLink241[25] , \Level2Out74[26] , 
        \ScanLink92[11] , \ScanLink125[9] , \ScanLink184[26] , 
        \ScanLink221[21] , \ScanLink254[11] , \Level2Out14[22] , 
        \ScanLink202[10] , \Level2Out42[23] , \Level4Out220[8] , 
        \Level1Out59[2] , \ScanLink87[25] , \ScanLink129[26] , 
        \ScanLink149[22] , \Level1Out90[19] , \Level1Out106[2] , 
        \Level1Out139[27] , \Level2Out30[2] , \Level2Out176[17] , 
        \Level4Out144[10] , \Level2Out120[16] , \Level4Out32[27] , 
        \Level8Out128[31] , \Level4Out64[26] , \Level8Out128[28] , 
        \Level2Out140[12] , \Level4Out112[11] , \Level4Out172[15] , 
        \ScanLink62[0] , \ScanLink69[23] , \Level1Out159[23] , 
        \Level2Out116[13] , \Level4Out52[23] , \Level4Out124[14] , 
        \ScanLink184[15] , \ScanLink221[12] , \ScanLink221[8] , 
        \ScanLink254[22] , \Level4Out124[9] , \ScanLink191[21] , 
        \ScanLink202[23] , \Level2Out14[11] , \Level2Out42[10] , 
        \ScanLink217[17] , \Level2Out22[14] , \Level128Out128[19] , 
        \ScanLink241[16] , \Level2Out74[15] , \ScanLink234[26] , 
        \Level1Out161[5] , \Level1Out207[16] , \Level2Out198[11] , 
        \Level8Out240[18] , \Level2Out248[26] , \Level1Out181[20] , 
        \Level1Out251[17] , \Level8Out216[19] , \Level1Out224[27] , 
        \Level1Out244[23] , \Level8Out88[1] , \Level8Out104[6] , 
        \Level1Out15[17] , \Level1Out20[9] , \ScanLink61[3] , 
        \Level1Out194[14] , \Level1Out201[0] , \Level1Out231[13] , 
        \Level16Out80[4] , \Level1Out212[22] , \Level2Out228[22] , 
        \ScanLink87[16] , \ScanLink129[15] , \Level1Out139[14] , 
        \Level1Out159[10] , \Level1Out162[6] , \Level2Out140[21] , 
        \Level4Out172[26] , \Level4Out124[27] , \Level2Out116[20] , 
        \Level4Out32[14] , \Level4Out52[10] , \Level4Out144[23] , 
        \ScanLink190[8] , \Level1Out202[3] , \Level2Out86[0] , 
        \Level2Out176[24] , \Level4Out112[22] , \Level2Out120[25] , 
        \Level4Out64[15] , \ScanLink92[22] , \Level1Out36[26] , 
        \Level1Out93[6] , \ScanLink149[11] , \Level2Out54[6] , 
        \Level8Out96[17] , \ScanLink243[2] , \Level2Out28[0] , 
        \Level1Out43[16] , \Level1Out23[12] , \Level1Out60[27] , 
        \Level1Out75[13] , \ScanLink123[7] , \Level2Out8[2] , 
        \Level2Out186[30] , \Level4Out232[18] , \Level8Out208[21] , 
        \Level1Out41[0] , \Level2Out186[29] , \Level1Out56[22] , 
        \Level8Out136[23] , \Level8Out160[22] , \Level1Out9[5] , 
        \Level1Out15[24] , \Level1Out23[21] , \Level1Out42[3] , 
        \Level1Out147[28] , \ScanLink240[1] , \Level2Out108[18] , 
        \Level16Out192[18] , \Level1Out56[11] , \Level1Load60[0] , 
        \ScanLink101[31] , \Level1Out111[30] , \Level1Out132[18] , 
        \Level1Out111[29] , \ScanLink120[4] , \Level1Out147[31] , 
        \Level1Out164[19] , \ScanLink122[19] , \ScanLink157[29] , 
        \Level2Out172[0] , \Level1Out75[20] , \ScanLink79[1] , 
        \Level1Out90[5] , \ScanLink101[28] , \ScanLink157[30] , 
        \ScanLink174[18] , \Level2Out84[18] , \Level2Out212[5] , 
        \Level2Out108[8] , \Level8Out208[12] , \ScanLink227[6] , 
        \Level4Out64[5] , \Level1Out25[4] , \Level1Out36[15] , 
        \Level1Out43[25] , \Level2Load212[0] , \Level1Out60[14] , 
        \ScanLink147[3] , \Level2Out236[29] , \ScanLink21[30] , 
        \ScanLink77[28] , \Level2Out236[30] , \Level8Out96[24] , 
        \ScanLink21[29] , \ScanLink54[19] , \ScanLink77[31] , \ScanLink195[5] , 
        \Level1Out26[7] , \ScanLink144[0] , \Level1Out164[8] , 
        \Level1Out179[7] , \ScanLink196[6] , \Level1Load203[0] , 
        \Level2Out116[4] , \ScanLink224[5] , \Level1Out219[2] , 
        \Level8Out136[10] , \ScanLink88[18] , \Level2Out52[8] , 
        \Level8Out160[11] , \Level2Out132[2] , \Level2Out252[7] , 
        \ScanLink160[6] , \Level8Out104[24] , \Level4Out108[18] , 
        \Level8Out152[25] , \ScanLink1[4] , \Level1Out11[15] , 
        \Level1Out27[10] , \Level1Out71[11] , \ScanLink163[5] , 
        \Level1Out192[8] , \ScanLink200[3] , \Level1Out32[24] , 
        \Level1Out52[20] , \ScanLink203[0] , \Level2Out232[18] , 
        \Level32Out32[0] , \Level1Out47[14] , \Level1Out208[18] , 
        \Level4Out40[3] , \ScanLink50[31] , \Level1Out64[25] , 
        \Level1Load144[0] , \ScanLink218[19] , \Level1Out223[8] , 
        \Level2Out68[2] , \ScanLink73[19] , \Level4Out92[5] , \Level8Out8[29] , 
        \ScanLink25[18] , \ScanLink40[8] , \ScanLink50[28] , \Level1Out66[5] , 
        \ScanLink104[2] , \Level8Out8[30] , \Level1Out3[23] , \ScanLink4[9] , 
        \Level1Out11[26] , \Level1Out32[17] , \Level1Out47[27] , 
        \Level1Out65[6] , \Level1Out78[9] , \Level1Load96[0] , 
        \Level1Out115[18] , \Level1Out136[29] , \Level1Out139[5] , 
        \Level4Out48[19] , \Level1Out143[19] , \Level8Out104[17] , 
        \Level1Out160[31] , \Level1Out136[30] , \Level1Out160[28] , 
        \ScanLink105[19] , \ScanLink126[28] , \Level2Out184[0] , 
        \Level8Out152[16] , \ScanLink153[18] , \ScanLink170[30] , 
        \ScanLink126[31] , \ScanLink170[29] , \Level2Out236[3] , 
        \Level2Out80[30] , \Level2Out80[29] , \Level2Out156[6] , 
        \Level1Out127[9] , \Level2Out58[19] , \Level1Out64[16] , 
        \ScanLink107[1] , \Level1Out19[0] , \Level1Out27[23] , \ScanLink39[3] , 
        \Level1Out71[22] , \Level4Load212[0] , \Level1Out52[13] , 
        \Level4Out236[29] , \Level2Out182[18] , \Level4Out24[7] , 
        \Level4Out236[30] , \Level1Out226[5] , \Level2Out144[10] , 
        \Level4Out176[17] , \Level32Out0[22] , \Level1Out128[11] , 
        \Level4Out56[21] , \Level1Out146[0] , \Level2Load54[0] , 
        \Level2Out112[11] , \Level2Out254[9] , \Level4Out120[16] , 
        \Level2Out172[15] , \Level1Out148[15] , \Level1Out189[9] , 
        \Level4Out140[12] , \Level4Out36[25] , \ScanLink18[22] , 
        \Level1Load38[0] , \ScanLink45[5] , \Level4Out60[24] , 
        \ScanLink78[26] , \ScanLink83[27] , \ScanLink158[14] , 
        \ScanLink166[8] , \Level2Out124[14] , \Level4Out116[13] , 
        \ScanLink96[13] , \Level1Out194[6] , \Level2Out70[0] , \ScanLink97[3] , 
        \ScanLink138[10] , \ScanLink94[0] , \ScanLink180[24] , 
        \ScanLink225[23] , \Level2Out10[20] , \ScanLink206[12] , 
        \Level1Out238[9] , \ScanLink250[13] , \Level2Out46[21] , 
        \ScanLink213[26] , \Level2Out26[25] , \ScanLink195[10] , 
        \Level1Out197[5] , \ScanLink230[17] , \ScanLink245[27] , 
        \Level2Out70[24] , \ScanLink46[6] , \ScanLink178[4] , 
        \Level1Out185[11] , \Level1Out203[27] , \Level1Out225[6] , 
        \Level1Out220[16] , \Level8Out120[0] , \Level1Out190[25] , 
        \Level1Out235[22] , \Level1Out255[26] , \Level4Out228[11] , 
        \Level4Out248[15] , \Level1Out3[19] , \Level1Out3[10] , 
        \ScanLink21[1] , \ScanLink83[14] , \ScanLink96[20] , \Level1Out145[3] , 
        \Level1Out216[13] , \Level1Out240[12] , \Level8Out240[5] , 
        \ScanLink218[1] , \ScanLink138[23] , \Level2Out14[4] , 
        \ScanLink158[27] , \Level1Out94[28] , \Level1Out148[26] , 
        \Level4Out36[16] , \Level1Out242[1] , \Level2Out172[26] , 
        \Level4Out140[21] , \Level2Out124[27] , \Level4Out116[20] , 
        \Level4Out60[17] , \Level32Out0[11] , \Level1Out94[31] , 
        \Level1Out122[4] , \Level2Out144[23] , \Level2Out150[8] , 
        \Level4Out176[24] , \Level4Out120[25] , \Level1Out128[22] , 
        \Level2Out112[22] , \Level4Out56[12] , \ScanLink5[18] , 
        \ScanLink17[25] , \ScanLink18[11] , \ScanLink22[2] , \Level1Out39[28] , 
        \Level1Out121[7] , \Level1Out190[16] , \Level1Out235[11] , 
        \Level1Out240[21] , \Level1Out241[2] , \Level8Out144[4] , 
        \Level4Out248[26] , \Level1Out216[20] , \Level8Out0[4] , 
        \Level2Out2[31] , \Level8Out224[1] , \Level1Out203[14] , 
        \Level1Out39[31] , \Level1Out255[15] , \Level4Out228[22] , 
        \Level2Out2[28] , \Level1Out63[8] , \Level1Out185[22] , 
        \ScanLink213[15] , \Level1Out220[25] , \ScanLink245[14] , 
        \Level2Out26[16] , \Level2Out70[17] , \ScanLink21[20] , 
        \Level1Out23[31] , \Level1Out75[29] , \ScanLink78[15] , 
        \ScanLink195[23] , \ScanLink230[24] , \ScanLink250[20] , 
        \ScanLink180[17] , \ScanLink225[10] , \Level2Out10[13] , 
        \ScanLink188[3] , \ScanLink206[21] , \Level2Out46[12] , 
        \Level2Out236[20] , \Level4Out204[27] , \Level4Out252[26] , 
        \ScanLink79[8] , \Level2Out200[25] , \Level1Out23[28] , 
        \Level1Out56[18] , \Level1Out75[30] , \Level2Out108[1] , 
        \Level4Out232[22] , \Level1Out219[14] , \Level1Out38[2] , 
        \Level2Out186[13] , \ScanLink54[10] , \ScanLink77[21] , 
        \Level1Out207[7] , \ScanLink209[15] , \ScanLink34[14] , 
        \ScanLink41[24] , \ScanLink64[7] , \ScanLink62[15] , \Level1Out167[2] , 
        \ScanLink17[16] , \ScanLink34[27] , \ScanLink67[4] , \ScanLink99[14] , 
        \ScanLink101[12] , \ScanLink122[23] , \ScanLink159[6] , 
        \Level1Out204[4] , \ScanLink157[13] , \ScanLink114[26] , 
        \ScanLink174[22] , \Level2Out80[7] , \ScanLink161[16] , 
        \Level1Out164[1] , \ScanLink239[3] , \Level2Out84[22] , 
        \ScanLink137[17] , \Level1Out104[27] , \ScanLink142[27] , 
        \Level8Out136[19] , \Level1Out111[13] , \Level1Out127[16] , 
        \ScanLink144[9] , \Level1Out171[17] , \Level32Out192[17] , 
        \Level2Out168[26] , \Level1Out132[22] , \Level1Out152[26] , 
        \Level8Out160[18] , \Level2Out52[1] , \Level1Out147[12] , 
        \Level2Out108[22] , \Level16Out192[22] , \Level1Out164[23] , 
        \ScanLink41[17] , \ScanLink21[13] , \ScanLink62[26] , \Level2Out28[9] , 
        \ScanLink77[12] , \Level1Out103[6] , \Level1Out41[9] , 
        \ScanLink54[23] , \ScanLink209[26] , \Level2Out186[20] , 
        \Level2Out200[16] , \Level4Out232[11] , \Level8Out208[28] , 
        \Level1Out104[14] , \Level1Out111[20] , \Level1Out132[11] , 
        \Level1Out147[21] , \Level1Out219[27] , \Level2Out236[13] , 
        \Level4Out204[14] , \Level8Out208[31] , \Level4Out252[15] , 
        \Level2Out36[5] , \Level2Out108[11] , \Level16Out192[11] , 
        \Level1Out164[10] , \Level1Out171[24] , \Level32Out192[24] , 
        \Level1Out7[31] , \Level1Out7[28] , \Level1Out20[0] , \Level1Out23[3] , 
        \ScanLink99[27] , \Level1Out127[25] , \Level1Out152[15] , 
        \ScanLink240[8] , \ScanLink161[25] , \Level2Out168[15] , 
        \Level1Out100[5] , \ScanLink114[15] , \ScanLink122[10] , 
        \ScanLink137[24] , \ScanLink142[14] , \Level2Out84[11] , 
        \ScanLink157[20] , \Level2Out172[9] , \ScanLink101[21] , 
        \ScanLink174[11] , \ScanLink141[4] , \ScanLink191[31] , 
        \Level128Out128[10] , \Level4Out244[5] , \Level1Out28[17] , 
        \ScanLink191[28] , \ScanLink193[2] , \ScanLink221[1] , 
        \Level2Out98[5] , \Level8Out88[26] , \Level2Out14[18] , 
        \Level4Out124[0] , \Level2Out42[19] , \Level8Out88[8] , 
        \Level1Out201[9] , \Level16Out80[16] , \Level1Out48[13] , 
        \Level1Out181[30] , \Level2Out198[18] , \Level8Out240[11] , 
        \ScanLink62[9] , \Level1Out85[17] , \Level1Out181[29] , 
        \Level2Out6[23] , \Level8Out216[10] , \ScanLink190[1] , 
        \Level2Out86[9] , \Level1Out90[23] , \Level8Out128[12] , 
        \Level1Out159[19] , \Level2Out110[3] , \Level2Out116[30] , 
        \Level2Out116[29] , \Level2Out140[28] , \Level2Out140[31] , 
        \Level4Out52[19] , \Level1Out48[20] , \Level1Out95[1] , 
        \ScanLink142[7] , \ScanLink149[18] , \Level8Out96[4] , 
        \ScanLink222[2] , \Level1Out231[29] , \Level2Out6[10] , 
        \Level8Out216[23] , \Level8Out240[22] , \Level16Out80[25] , 
        \Level1Out28[24] , \Level1Out105[8] , \Level1Out212[18] , 
        \Level1Out231[30] , \Level1Out244[19] , \Level4Out192[2] , 
        \ScanLink18[1] , \Level1Out44[4] , \Level1Out47[7] , \ScanLink221[28] , 
        \Level2Out228[18] , \ScanLink69[19] , \ScanLink125[0] , 
        \ScanLink202[19] , \ScanLink221[31] , \ScanLink254[18] , 
        \ScanLink245[5] , \Level4Out220[1] , \Level128Out128[23] , 
        \Level1Out118[7] , \Level8Out88[15] , \ScanLink126[3] , 
        \Level4Out140[4] , \ScanLink92[18] , \ScanLink246[6] , \ScanLink21[8] , 
        \Level1Out60[2] , \Level1Out85[24] , \Level1Out90[10] , 
        \Level1Out96[2] , \Level2Out214[2] , \Level4Out144[19] , 
        \Level8Out128[21] , \Level2Out174[7] , \Level4Out112[18] , 
        \Level2Out182[7] , \ScanLink96[30] , \ScanLink96[29] , 
        \ScanLink102[5] , \Level32Out0[18] , \Level1Out39[21] , 
        \Level1Out81[15] , \Level1Out94[21] , \Level1Load125[0] , 
        \Level2Out150[1] , \Level4Out116[30] , \Level4Out140[28] , 
        \Level1Out242[8] , \Level2Out230[4] , \Level4Out116[29] , 
        \Level4Out140[31] , \Level1Out240[28] , \Level2Out2[21] , 
        \Level8Out224[8] , \ScanLink4[0] , \ScanLink18[18] , \Level1Out59[25] , 
        \Level1Out216[30] , \Level1Out216[29] , \Level1Out235[18] , 
        \Level1Out240[31] , \Level1Out63[1] , \ScanLink101[6] , 
        \ScanLink206[31] , \ScanLink250[29] , \Level8Out224[17] , 
        \Level4Out164[2] , \ScanLink206[28] , \ScanLink225[19] , 
        \ScanLink250[30] , \Level2Load134[0] , \Level4Out204[7] , 
        \Level1Out146[9] , \Level1Out189[0] , \ScanLink1[30] , \ScanLink7[3] , 
        \Level1Out19[9] , \Level1Out81[26] , \Level1Out94[12] , 
        \Level2Out134[5] , \Level2Out144[19] , \Level4Out56[31] , 
        \ScanLink58[3] , \Level1Out128[18] , \ScanLink206[4] , 
        \Level2Out112[18] , \Level2Out254[0] , \Level4Out56[28] , 
        \Level1Out59[16] , \ScanLink89[6] , \ScanLink94[9] , \ScanLink138[19] , 
        \ScanLink166[1] , \Level2Out70[9] , \Level1Out158[5] , 
        \ScanLink195[19] , \ScanLink205[7] , \ScanLink165[2] , 
        \Level1Out238[0] , \Level2Out10[29] , \Level4Out100[6] , 
        \Level2Out46[31] , \Level2Out10[30] , \Level2Out46[28] , 
        \ScanLink218[8] , \Level8Out224[24] , \Level1Out39[12] , 
        \Level64Out128[4] , \Level1Load59[0] , \Level1Out115[11] , 
        \Level1Out136[20] , \Level1Out185[18] , \Level2Out2[12] , 
        \Level4Out228[18] , \Level8Out120[9] , \Level4Out48[10] , 
        \Level1Out143[10] , \Level4Out168[26] , \Level1Out100[25] , 
        \Level1Out160[21] , \Level2Out184[9] , \ScanLink1[29] , 
        \Level1Out123[14] , \Level1Out175[15] , \Level4Out108[22] , 
        \Level1Out2[20] , \Level1Out8[26] , \ScanLink13[27] , \ScanLink24[5] , 
        \ScanLink27[6] , \ScanLink110[24] , \Level1Out156[24] , 
        \Level4Out28[14] , \Level2Out12[3] , \Level2Out80[20] , 
        \Level1Out124[3] , \ScanLink133[15] , \ScanLink165[14] , 
        \ScanLink88[22] , \ScanLink105[10] , \ScanLink119[4] , 
        \ScanLink126[21] , \ScanLink146[25] , \Level1Out244[6] , 
        \ScanLink153[11] , \ScanLink170[20] , \ScanLink218[23] , 
        \ScanLink30[16] , \ScanLink45[26] , \Level2Out58[10] , 
        \ScanLink66[17] , \Level1Out127[0] , \ScanLink25[22] , 
        \ScanLink50[12] , \ScanLink73[23] , \Level1Out78[0] , \Level8Out8[13] , 
        \Level1Out247[5] , \Level2Out38[14] , \Level2Out204[27] , 
        \Level1Out8[15] , \ScanLink43[2] , \ScanLink107[8] , 
        \Level1Out208[22] , \Level2Out148[3] , \Level4Out236[20] , 
        \Level2Out182[11] , \Level2Out252[26] , \Level2Out228[6] , 
        \Level2Out232[22] , \Level4Out200[25] , \ScanLink88[11] , 
        \ScanLink126[12] , \ScanLink153[22] , \ScanLink91[4] , 
        \ScanLink105[23] , \Level1Out140[7] , \ScanLink170[13] , 
        \ScanLink110[17] , \ScanLink165[27] , \Level2Out80[13] , 
        \ScanLink133[26] , \ScanLink146[16] , \Level1Out220[2] , 
        \Level1Out175[26] , \ScanLink92[7] , \Level1Out100[16] , 
        \Level4Out108[11] , \Level1Out115[22] , \Level1Out123[27] , 
        \Level1Out156[17] , \Level4Out28[27] , \Level1Out192[1] , 
        \Level1Out136[13] , \Level1Out143[23] , \Level2Out76[7] , 
        \Level4Out48[23] , \Level1Out160[12] , \Level1Out191[2] , 
        \ScanLink203[9] , \Level4Out168[15] , \Level32Out32[9] , 
        \Level1Out208[11] , \Level2Out232[11] , \Level4Out200[16] , 
        \ScanLink13[14] , \ScanLink25[11] , \Level1Out27[19] , 
        \Level1Out52[30] , \Level2Out204[14] , \Level4Out236[13] , 
        \Level1Out71[18] , \Level2Out182[22] , \Level1Out52[29] , 
        \ScanLink73[10] , \Level1Out143[4] , \Level2Out252[15] , 
        \Level8Load200[0] , \Level8Out8[20] , \ScanLink30[25] , 
        \ScanLink40[1] , \ScanLink50[21] , \Level1Out223[1] , 
        \Level2Out38[27] , \Level2Out58[23] , \Level16Out0[5] , 
        \ScanLink45[15] , \ScanLink218[10] , \ScanLink56[5] , \ScanLink66[24] , 
        \Level1Out155[0] , \ScanLink208[2] , \Level1Out217[10] , 
        \Level1Out191[26] , \Level2Out188[17] , \Level4Out84[8] , 
        \Level16Out112[17] , \Level16Out144[16] , \Level1Out234[21] , 
        \Level32Out192[6] , \Level1Out2[13] , \ScanLink9[5] , \ScanLink19[21] , 
        \Level1Out38[18] , \ScanLink168[7] , \Level1Out184[12] , 
        \Level1Out221[15] , \Level1Out235[5] , \Level1Out241[11] , 
        \Level1Out202[24] , \Level1Out254[25] , \Level1Out187[6] , 
        \ScanLink194[13] , \ScanLink231[14] , \Level2Out238[24] , 
        \ScanLink244[24] , \ScanLink48[9] , \ScanLink79[25] , \ScanLink84[3] , 
        \ScanLink175[8] , \ScanLink207[11] , \ScanLink212[25] , 
        \Level2Out52[16] , \Level2Out32[12] , \ScanLink139[13] , 
        \ScanLink181[27] , \ScanLink224[20] , \ScanLink251[10] , 
        \Level2Out64[13] , \ScanLink87[0] , \Level1Out184[5] , 
        \ScanLink19[12] , \ScanLink55[6] , \ScanLink82[24] , \ScanLink97[10] , 
        \Level2Out60[3] , \Level8Out16[18] , \ScanLink159[17] , 
        \Level8Out40[19] , \ScanLink79[16] , \Level1Out95[18] , 
        \Level1Out129[12] , \Level1Out149[16] , \Level1Out156[3] , 
        \Level2Out150[27] , \Level128Out0[19] , \Level2Out106[26] , 
        \Level4Out48[2] , \Level1Out236[6] , \Level2Out166[22] , 
        \Level16Out48[29] , \Level16Out48[30] , \ScanLink207[22] , 
        \Level2Out130[23] , \ScanLink251[23] , \Level2Out32[21] , 
        \Level2Out64[20] , \ScanLink181[14] , \ScanLink224[13] , 
        \ScanLink244[17] , \ScanLink32[1] , \ScanLink194[20] , 
        \ScanLink231[27] , \ScanLink212[16] , \Level2Out52[25] , 
        \Level1Out131[4] , \Level1Out184[21] , \Level1Out221[26] , 
        \Level1Out254[16] , \Level1Out202[17] , \Level2Out238[17] , 
        \Level1Out217[23] , \Level2Out188[24] , \Level16Out112[24] , 
        \Level1Out10[16] , \ScanLink31[2] , \Level1Out129[21] , 
        \Level1Out132[7] , \Level1Out191[15] , \Level1Out241[22] , 
        \Level1Out251[1] , \Level1Out234[12] , \Level16Out144[25] , 
        \Level2Out166[11] , \Level2Out130[10] , \Level1Out70[8] , 
        \ScanLink82[17] , \Level1Out149[25] , \Level1Out252[2] , 
        \Level2Out106[15] , \Level2Out150[14] , \Level32Out32[19] , 
        \Level32Out64[18] , \ScanLink97[23] , \ScanLink139[20] , 
        \ScanLink159[24] , \Level1Load248[0] , \Level2Out78[1] , 
        \Level1Out11[1] , \Level1Out26[13] , \Level1Out33[27] , 
        \Level1Out65[26] , \Level2Out8[27] , \Level2Load146[0] , 
        \Level1Out181[8] , \ScanLink213[3] , \Level1Out46[17] , 
        \Level4Out116[2] , \ScanLink0[10] , \Level1Out53[23] , 
        \Level1Out70[12] , \ScanLink173[6] , \Level1Out12[2] , 
        \Level1Out114[28] , \Level1Out142[30] , \Level1Out161[18] , 
        \ScanLink210[0] , \Level8Out248[4] , \Level8Out128[1] , 
        \ScanLink170[5] , \Level2Out178[30] , \ScanLink53[8] , 
        \ScanLink104[29] , \Level1Out114[31] , \Level1Out137[19] , 
        \Level1Out142[29] , \Level64Out128[26] , \Level2Out178[29] , 
        \ScanLink152[31] , \ScanLink171[19] , \Level1Out53[10] , 
        \ScanLink104[30] , \ScanLink127[18] , \ScanLink152[28] , 
        \Level2Out122[1] , \Level1Load157[0] , \Level1Out230[8] , 
        \Level2Out242[4] , \ScanLink0[23] , \Level1Out10[25] , 
        \Level1Out26[20] , \ScanLink29[0] , \Level1Out70[21] , 
        \Level4Out172[6] , \Level1Out65[15] , \Level1Load85[0] , 
        \ScanLink117[2] , \Level2Out158[9] , \Level1Out209[31] , 
        \Level2Out8[14] , \Level2Out210[19] , \Level4Out212[3] , 
        \ScanLink24[31] , \ScanLink24[28] , \Level1Out33[14] , 
        \Level1Out46[24] , \Level1Out75[5] , \Level1Out209[28] , 
        \Level2Out246[18] , \ScanLink51[18] , \ScanLink72[30] , 
        \ScanLink219[30] , \ScanLink219[29] , \Level8Out152[9] , 
        \ScanLink72[29] , \Level1Out76[6] , \ScanLink89[31] , \ScanLink89[28] , 
        \Level1Out134[9] , \Level2Out146[5] , \Level4Out0[31] , 
        \Level2Out226[0] , \Level4Out0[28] , \Level1Out129[6] , 
        \Level2Out194[3] , \Level8Out8[5] , \Level64Out128[15] , 
        \ScanLink1[24] , \ScanLink1[17] , \ScanLink1[0] , \Level1Out1[4] , 
        \ScanLink4[21] , \ScanLink4[12] , \Level1Out52[0] , \Level1Out80[6] , 
        \ScanLink114[1] , \Level1Out249[3] , \Level4Out228[9] , 
        \ScanLink130[7] , \Level2Out162[3] , \Level2Out202[6] , 
        \Level4Out4[19] , \Level4Load28[0] , \Level8Out168[3] , 
        \Level1Load4[0] , \Level1Out22[11] , \ScanLink250[2] , 
        \Level8Out208[6] , \Level16Out32[24] , \Level16Out64[25] , 
        \Level128Out0[6] , \Level1Out51[3] , \Level1Out57[21] , 
        \ScanLink10[9] , \Level1Out14[14] , \Level1Out74[10] , 
        \ScanLink133[4] , \Level4Out4[5] , \Level4Out236[5] , \ScanLink20[19] , 
        \Level1Out37[25] , \Level1Out61[24] , \Level2Out214[28] , 
        \Level2Out242[30] , \ScanLink253[1] , \Level1Out42[15] , 
        \Level2Out214[31] , \Level16Out192[8] , \Level1Out83[5] , 
        \Level2Out242[29] , \Level4Out156[0] , \Level2Out38[3] , 
        \Level1Out36[4] , \ScanLink55[30] , \ScanLink55[29] , 
        \Level1Load73[0] , \Level4Out184[6] , \ScanLink76[18] , 
        \Level16Out32[17] , \Level1Out4[9] , \Level1Out28[8] , 
        \ScanLink100[18] , \Level1Out110[19] , \ScanLink154[3] , 
        \Level1Out209[1] , \Level8Out80[0] , \Level16Out64[16] , 
        \Level1Out133[31] , \Level1Out133[28] , \Level1Out165[29] , 
        \ScanLink234[6] , \Level1Out146[18] , \Level1Out169[4] , 
        \Level1Out165[30] , \ScanLink123[30] , \ScanLink123[29] , 
        \ScanLink175[28] , \ScanLink186[5] , \ScanLink156[19] , 
        \ScanLink175[31] , \ScanLink185[6] , \ScanLink229[9] , 
        \Level2Out106[7] , \Level16Out96[9] , \Level1Out61[17] , 
        \ScanLink157[0] , \Level1Out177[8] , \Level1Load210[0] , 
        \Level2Out28[31] , \Level2Out28[28] , \ScanLink198[9] , 
        \Level1Out6[22] , \Level1Out14[27] , \ScanLink15[4] , 
        \Level1Out22[22] , \Level1Out35[7] , \Level4Out252[1] , 
        \Level1Out37[16] , \Level1Out42[26] , \Level1Out57[12] , 
        \ScanLink237[5] , \Level4Out132[4] , \Level1Out49[1] , \ScanLink69[2] , 
        \Level16Load96[0] , \Level1Out74[23] , \Level1Out86[8] , 
        \Level1Out158[20] , \Level2Out162[20] , \Level2Out204[8] , 
        \Level2Out0[3] , \Level2Out134[21] , \ScanLink16[7] , \ScanLink68[13] , 
        \ScanLink86[26] , \Level1Out116[1] , \Level1Out138[24] , 
        \Level2Out154[25] , \Level2Out20[1] , \Level2Out102[24] , 
        \ScanLink93[12] , \ScanLink128[25] , \ScanLink136[9] , 
        \ScanLink148[21] , \Level1Out98[4] , \ScanLink203[13] , 
        \Level2Out36[10] , \ScanLink185[25] , \ScanLink190[11] , 
        \ScanLink220[22] , \ScanLink235[16] , \ScanLink255[12] , 
        \Level2Out60[11] , \Level1Out115[2] , \ScanLink128[5] , 
        \Level1Out180[10] , \ScanLink216[27] , \ScanLink240[26] , 
        \Level1Out225[17] , \Level2Out56[14] , \Level1Out206[26] , 
        \Level1Out250[27] , \Level4Out188[17] , \Level16Out176[11] , 
        \Level1Out213[12] , \ScanLink248[0] , \Level1Out195[24] , 
        \Level1Out230[23] , \Level1Out245[13] , \ScanLink148[12] , 
        \Level1Out2[7] , \Level1Out6[11] , \ScanLink71[0] , \ScanLink86[15] , 
        \ScanLink93[21] , \Level2Out44[5] , \Level1Out91[30] , 
        \ScanLink128[16] , \ScanLink232[8] , \Level1Out138[17] , 
        \Level1Out212[0] , \Level2Out102[17] , \Level2Out154[16] , 
        \Level1Out158[13] , \Level1Out172[5] , \Level2Out96[3] , 
        \Level2Out134[12] , \Level2Out162[13] , \Level1Out91[29] , 
        \Level1Out213[21] , \Level2Out100[9] , \Level1Out245[20] , 
        \Level8Out184[18] , \Level1Out33[9] , \Level1Out49[19] , 
        \ScanLink72[3] , \ScanLink183[8] , \Level1Out211[3] , 
        \Level1Out195[17] , \Level1Out230[10] , \Level1Out171[6] , 
        \Level1Out180[23] , \Level1Out225[24] , \Level1Out250[14] , 
        \Level4Out188[24] , \Level1Out206[15] , \ScanLink240[15] , 
        \Level16Out176[22] , \ScanLink68[20] , \ScanLink190[22] , 
        \ScanLink235[25] , \ScanLink216[14] , \Level2Out56[27] , 
        \Level1Out3[27] , \ScanLink46[2] , \Level1Out145[7] , 
        \ScanLink185[16] , \ScanLink203[20] , \Level2Out36[23] , 
        \ScanLink255[21] , \Level2Out60[22] , \Level4Out72[8] , 
        \Level1Out216[17] , \ScanLink220[11] , \ScanLink218[5] , 
        \Level8Out240[1] , \Level8Out224[29] , \Level1Out190[21] , 
        \Level1Out235[26] , \Level4Out248[11] , \Level64Out128[9] , 
        \Level1Out240[16] , \Level8Out224[30] , \Level1Out3[14] , 
        \ScanLink18[26] , \Level1Out158[8] , \ScanLink178[0] , 
        \Level1Out185[15] , \Level1Out225[2] , \Level8Out120[4] , 
        \Level1Out220[12] , \ScanLink195[14] , \Level1Out203[23] , 
        \Level1Out255[22] , \Level4Out228[15] , \Level1Out197[1] , 
        \ScanLink230[13] , \ScanLink245[23] , \Level2Out70[20] , 
        \ScanLink18[15] , \Level1Out19[4] , \ScanLink45[1] , \ScanLink78[22] , 
        \ScanLink94[4] , \ScanLink206[16] , \ScanLink213[22] , 
        \Level2Out26[21] , \Level2Out46[25] , \ScanLink83[23] , 
        \ScanLink96[17] , \ScanLink97[7] , \ScanLink138[14] , 
        \ScanLink180[20] , \ScanLink225[27] , \ScanLink250[17] , 
        \Level2Out10[24] , \Level1Out194[2] , \ScanLink206[9] , 
        \Level2Out70[4] , \ScanLink158[10] , \Level4Out60[20] , 
        \Level1Out146[4] , \Level2Out124[10] , \Level2Out134[8] , 
        \Level4Out116[17] , \Level2Out172[11] , \Level4Out140[16] , 
        \Level1Out148[11] , \Level4Out36[21] , \ScanLink78[11] , 
        \Level1Out128[15] , \Level4Out56[25] , \ScanLink206[25] , 
        \Level1Out226[1] , \Level2Out112[15] , \Level2Out144[14] , 
        \Level4Out120[12] , \Level2Out46[16] , \Level4Out176[13] , 
        \Level32Out0[26] , \ScanLink250[24] , \ScanLink180[13] , 
        \ScanLink225[14] , \ScanLink245[10] , \Level2Out10[17] , 
        \Level2Out70[13] , \ScanLink22[6] , \ScanLink195[27] , 
        \ScanLink213[11] , \ScanLink230[20] , \Level2Out26[12] , 
        \Level1Out59[28] , \Level1Out121[3] , \Level1Out185[26] , 
        \Level1Out255[11] , \Level4Out228[26] , \Level1Out220[21] , 
        \Level1Out203[10] , \Level8Out224[5] , \Level1Out216[24] , 
        \Level8Out0[0] , \Level1Out240[25] , \Level8Out144[0] , 
        \ScanLink21[5] , \Level1Out59[31] , \Level1Out190[12] , 
        \Level1Out235[15] , \Level1Out241[6] , \Level4Out248[22] , 
        \Level1Out122[0] , \Level1Out128[26] , \Level2Load30[0] , 
        \Level4Out120[21] , \Level2Out112[26] , \Level4Out56[16] , 
        \Level32Out0[15] , \Level1Out81[18] , \Level2Out144[27] , 
        \Level4Out176[20] , \Level4Out116[24] , \ScanLink83[10] , 
        \Level1Out148[22] , \Level1Out242[5] , \Level2Out124[23] , 
        \Level4Out36[12] , \Level4Out60[13] , \Level2Out172[22] , 
        \Level4Out140[25] , \Level2Out230[9] , \ScanLink96[24] , 
        \ScanLink102[8] , \ScanLink158[23] , \ScanLink138[27] , 
        \Level1Out143[9] , \Level2Out14[0] , \Level4Out92[1] , 
        \Level1Out8[18] , \Level1Out11[11] , \ScanLink13[19] , 
        \ScanLink30[31] , \ScanLink30[28] , \ScanLink66[29] , \Level2Out68[6] , 
        \Level16Out0[8] , \ScanLink45[18] , \ScanLink66[30] , 
        \Level1Out27[14] , \Level1Out32[20] , \Level1Out64[21] , 
        \ScanLink203[4] , \Level32Out32[4] , \Level1Out47[10] , 
        \Level4Out40[7] , \Level1Out52[24] , \Level2Out252[18] , 
        \Level2Out204[19] , \Level1Out71[15] , \ScanLink163[1] , 
        \ScanLink2[3] , \ScanLink91[9] , \ScanLink200[7] , \ScanLink160[2] , 
        \Level4Out168[18] , \Level8Out152[21] , \Level8Out104[20] , 
        \Level1Out11[22] , \Level1Out27[27] , \Level1Out52[17] , 
        \Level2Out132[6] , \Level2Out252[3] , \Level4Out24[3] , 
        \ScanLink39[7] , \Level1Out64[12] , \Level1Out71[26] , 
        \ScanLink107[5] , \Level4Out200[31] , \ScanLink24[8] , 
        \Level1Out32[13] , \Level1Out47[23] , \Level1Out65[2] , 
        \Level4Out200[28] , \Level1Out66[1] , \ScanLink110[30] , 
        \Level1Load120[0] , \Level1Out247[8] , \Level2Out38[19] , 
        \ScanLink133[18] , \ScanLink110[29] , \ScanLink146[28] , 
        \Level2Out156[2] , \ScanLink119[9] , \ScanLink146[31] , 
        \ScanLink165[19] , \Level2Out236[7] , \Level1Out139[1] , 
        \Level2Out184[4] , \Level8Out152[12] , \Level8Out104[13] , 
        \Level32Load0[0] , \Level1Out100[31] , \Level1Out123[19] , 
        \Level1Out4[4] , \ScanLink5[26] , \ScanLink5[15] , \Level1Out42[7] , 
        \Level1Out90[1] , \Level1Out100[28] , \ScanLink104[6] , 
        \Level1Out156[29] , \Level4Out28[19] , \ScanLink137[29] , 
        \ScanLink142[19] , \Level1Out156[30] , \Level1Out175[18] , 
        \ScanLink161[31] , \ScanLink161[28] , \Level1Out100[8] , 
        \ScanLink114[18] , \ScanLink137[30] , \Level2Out212[1] , 
        \ScanLink120[0] , \Level2Out172[4] , \Level2Out36[8] , 
        \Level8Out160[26] , \Level1Out15[13] , \Level1Out23[16] , 
        \Level1Out104[19] , \Level1Out127[28] , \Level1Out152[18] , 
        \Level1Out171[30] , \ScanLink240[5] , \Level2Out168[18] , 
        \Level32Out192[30] , \Level1Out171[29] , \Level8Out136[27] , 
        \Level32Out192[29] , \Level1Out127[31] , \Level1Out41[4] , 
        \Level1Out56[26] , \Level1Out75[17] , \ScanLink123[3] , 
        \Level2Out8[6] , \Level8Out208[25] , \Level1Out26[3] , 
        \Level1Out36[22] , \Level1Out60[23] , \ScanLink243[6] , 
        \Level4Out252[18] , \Level1Out43[12] , \Level4Out204[19] , 
        \Level1Out93[2] , \Level2Out28[4] , \Level8Out96[13] , 
        \Level1Out7[25] , \Level1Out9[1] , \ScanLink67[9] , \ScanLink144[4] , 
        \Level1Out219[6] , \Level8Out160[15] , \Level8Out136[14] , 
        \Level1Out179[3] , \ScanLink224[1] , \ScanLink196[2] , 
        \Level1Out204[9] , \ScanLink99[19] , \Level2Out116[0] , 
        \ScanLink195[1] , \ScanLink209[18] , \Level1Out15[20] , 
        \ScanLink17[31] , \ScanLink17[28] , \ScanLink41[30] , 
        \Level8Out96[20] , \ScanLink62[18] , \ScanLink41[29] , 
        \ScanLink34[19] , \Level1Out60[10] , \ScanLink147[7] , 
        \Level1Out23[25] , \Level1Out25[0] , \Level1Out36[11] , 
        \Level1Out43[21] , \Level1Out56[15] , \Level1Out219[19] , 
        \ScanLink227[2] , \Level2Load68[0] , \Level4Out64[1] , 
        \Level1Out28[29] , \Level1Out44[9] , \Level1Out59[6] , 
        \Level1Out75[24] , \Level2Out200[31] , \ScanLink79[5] , 
        \Level2Out200[28] , \Level8Out208[16] , \Level1Out85[30] , 
        \Level1Out85[29] , \Level1Out159[27] , \Level2Out116[17] , 
        \Level4Out52[27] , \Level4Out124[10] , \Level2Out120[12] , 
        \Level2Out140[16] , \Level4Out64[22] , \Level4Out172[11] , 
        \Level1Out106[6] , \Level2Out176[13] , \Level4Out112[15] , 
        \Level1Out139[23] , \Level4Out144[14] , \Level4Out32[23] , 
        \ScanLink69[14] , \ScanLink87[21] , \Level2Out30[6] , \Level1Out88[3] , 
        \ScanLink92[15] , \ScanLink129[22] , \ScanLink149[26] , 
        \ScanLink202[14] , \Level2Out42[27] , \ScanLink184[22] , 
        \ScanLink221[25] , \Level2Out14[26] , \ScanLink191[16] , 
        \ScanLink245[8] , \ScanLink254[15] , \ScanLink234[11] , 
        \Level8Out88[18] , \Level1Out105[5] , \ScanLink138[2] , 
        \Level1Out181[17] , \ScanLink217[20] , \ScanLink241[21] , 
        \Level2Out74[22] , \Level4Out140[9] , \Level2Out22[23] , 
        \Level8Out160[6] , \Level1Out224[10] , \Level1Out207[21] , 
        \Level1Out251[20] , \Level2Out248[11] , \Level1Out212[15] , 
        \Level2Out198[26] , \Level8Out200[3] , \Level16Out80[31] , 
        \Level2Out228[15] , \Level1Out194[23] , \Level1Out231[24] , 
        \Level16Out80[28] , \Level1Out7[16] , \Level1Out28[30] , 
        \Level1Out244[14] , \ScanLink61[7] , \ScanLink87[12] , 
        \ScanLink92[26] , \ScanLink149[15] , \Level8Out96[9] , 
        \Level1Load178[0] , \Level2Out54[2] , \ScanLink129[11] , 
        \Level1Out139[10] , \Level1Out202[7] , \Level2Out120[21] , 
        \Level4Out112[26] , \Level4Out32[10] , \Level4Out64[11] , 
        \Level4Out144[27] , \Level1Out159[14] , \Level2Out86[4] , 
        \Level2Out176[20] , \Level4Out124[23] , \Level1Out162[2] , 
        \Level2Out116[24] , \Level4Out52[14] , \Level1Out212[26] , 
        \Level2Out140[25] , \Level4Out172[22] , \Level2Out228[26] , 
        \Level8Out88[5] , \ScanLink62[4] , \Level1Out194[10] , 
        \Level1Out201[4] , \Level1Out244[27] , \Level8Out104[2] , 
        \Level1Out231[17] , \Level16Out80[0] , \ScanLink69[27] , 
        \Level1Out161[1] , \Level1Out181[24] , \Level1Out251[13] , 
        \Level1Out224[23] , \ScanLink191[25] , \Level1Out207[12] , 
        \Level2Out198[15] , \ScanLink241[12] , \Level2Out248[22] , 
        \Level2Out74[11] , \ScanLink234[22] , \ScanLink141[9] , 
        \Level2Out98[8] , \ScanLink184[11] , \ScanLink202[27] , 
        \ScanLink217[13] , \Level2Out22[10] , \Level2Out42[14] , 
        \Level4Out244[8] , \ScanLink221[16] , \ScanLink254[26] , 
        \Level2Out14[15] , \ScanLink198[4] , \Level2Out192[20] , 
        \Level2Out242[17] , \Level1Out7[7] , \ScanLink16[22] , 
        \ScanLink20[27] , \Level1Out28[5] , \Level1Out218[13] , 
        \Level2Out118[6] , \Level2Out214[16] , \Level4Out80[11] , 
        \Level4Out196[22] , \ScanLink237[8] , \Level2Out222[13] , 
        \Level4Out132[9] , \ScanLink55[17] , \ScanLink76[26] , 
        \ScanLink208[12] , \Level1Out217[0] , \Level8Out112[6] , 
        \Level16Out96[4] , \ScanLink35[13] , \ScanLink40[23] , \ScanLink74[0] , 
        \Level2Out28[25] , \Level2Out48[21] , \ScanLink63[12] , 
        \Level1Out177[5] , \ScanLink77[3] , \ScanLink98[13] , 
        \ScanLink100[15] , \ScanLink123[24] , \ScanLink186[8] , 
        \Level1Out214[3] , \Level4Out4[27] , \ScanLink149[1] , 
        \ScanLink156[14] , \Level2Out90[11] , \ScanLink115[21] , 
        \ScanLink175[25] , \Level2Out90[0] , \ScanLink229[4] , 
        \ScanLink160[11] , \Level1Out174[6] , \ScanLink136[10] , 
        \Level1Out105[20] , \ScanLink143[20] , \ScanLink10[4] , 
        \ScanLink16[11] , \ScanLink35[20] , \Level1Out36[9] , 
        \Level1Out170[10] , \Level1Out110[14] , \Level1Out126[11] , 
        \Level1Out133[25] , \Level1Out153[21] , \Level2Out42[6] , 
        \Level1Out146[15] , \Level1Out169[9] , \Level1Out165[24] , 
        \Level8Out176[2] , \ScanLink40[10] , \Level2Out28[16] , 
        \Level1Out83[8] , \ScanLink20[14] , \ScanLink63[21] , \ScanLink76[15] , 
        \Level1Out113[1] , \Level8Out216[7] , \ScanLink13[7] , 
        \Level1Out14[19] , \Level1Out37[31] , \Level1Out37[28] , 
        \ScanLink55[24] , \Level2Out48[12] , \ScanLink133[9] , 
        \ScanLink208[21] , \Level4Out196[11] , \Level1Out218[20] , 
        \Level2Out222[20] , \Level4Out236[8] , \Level4Out4[8] , 
        \Level1Out42[18] , \Level1Out61[30] , \Level2Out192[13] , 
        \Level16Out192[5] , \Level2Out242[24] , \Level2Out214[25] , 
        \Level1Out61[29] , \Level4Out80[22] , \ScanLink98[20] , 
        \Level1Out105[13] , \Level1Out110[27] , \Level1Out133[16] , 
        \Level1Out146[26] , \Level2Out26[2] , \Level1Out165[17] , 
        \Level1Out170[23] , \Level16Out64[28] , \Level16Out32[30] , 
        \Level1Out126[22] , \Level1Out153[12] , \Level16Out64[31] , 
        \Level16Out32[29] , \ScanLink160[22] , \ScanLink115[12] , 
        \ScanLink136[23] , \ScanLink143[13] , \Level2Out6[0] , 
        \Level4Out228[4] , \Level1Load1[0] , \Level1Out1[9] , 
        \Level1Out29[10] , \Level1Out33[4] , \ScanLink100[26] , 
        \Level1Out110[2] , \ScanLink123[17] , \ScanLink156[27] , 
        \Level4Out4[14] , \ScanLink175[16] , \Level2Out90[22] , 
        \Level4Out148[1] , \ScanLink151[3] , \ScanLink216[19] , 
        \ScanLink235[31] , \ScanLink183[5] , \ScanLink231[6] , 
        \ScanLink235[28] , \ScanLink240[18] , \Level2Load204[0] , 
        \Level2Out88[2] , \Level4Out72[5] , \Level1Out30[7] , 
        \Level1Out49[14] , \Level1Out206[18] , \Level1Out225[30] , 
        \Level4Out188[30] , \Level8Out184[15] , \Level1Out84[10] , 
        \ScanLink180[6] , \Level1Out225[29] , \Level1Out250[19] , 
        \Level4Out188[29] , \Level1Out91[24] , \Level1Out172[8] , 
        \Level1Load215[0] , \Level2Out100[4] , \Level8Out72[20] , 
        \ScanLink152[0] , \Level2Out44[8] , \Level1Out29[23] , 
        \Level1Out49[27] , \Level1Out85[6] , \ScanLink86[18] , 
        \ScanLink232[5] , \Level8Out24[21] , \ScanLink128[8] , 
        \Level1Out195[30] , \Level1Out195[29] , \Level128Load128[0] , 
        \Level8Out184[26] , \Level1Out54[3] , \Level1Out57[0] , 
        \Level1Out98[9] , \ScanLink185[28] , \Level1Out108[0] , 
        \ScanLink135[7] , \ScanLink185[31] , \ScanLink255[2] , 
        \Level2Out56[19] , \Level32Out64[2] , \ScanLink128[28] , 
        \ScanLink136[4] , \Level4Out16[1] , \ScanLink128[31] , \ScanLink9[8] , 
        \ScanLink15[9] , \Level1Out86[5] , \Level1Out91[17] , \ScanLink256[1] , 
        \Level8Out24[12] , \Level8Out72[13] , \Level1Out138[30] , 
        \Level1Out138[29] , \Level2Out204[5] , \Level2Out102[29] , 
        \Level2Out154[31] , \Level2Out154[28] , \Level1Out38[26] , 
        \Level1Out70[5] , \Level1Load76[0] , \Level1Out84[23] , 
        \Level2Out102[30] , \Level2Out164[0] , \Level1Load80[0] , 
        \ScanLink159[29] , \Level8Out40[27] , \ScanLink159[30] , 
        \Level2Out192[0] , \Level8Out16[26] , \Level1Out80[12] , 
        \Level1Out95[26] , \ScanLink112[2] , \Level1Out149[31] , 
        \Level1Out149[28] , \Level2Out140[6] , \Level16Out48[17] , 
        \Level32Out64[15] , \Level2Out106[18] , \Level2Out220[3] , 
        \Level1Out131[9] , \Level2Out150[19] , \Level32Out32[14] , 
        \Level128Out0[27] , \Level1Out58[22] , \Level1Out191[18] , 
        \Level2Out188[30] , \Level16Out112[30] , \Level16Out144[28] , 
        \Level2Out188[29] , \Level16Out112[29] , \Level1Out73[6] , 
        \ScanLink111[1] , \ScanLink181[19] , \Level4Out32[7] , 
        \Level16Out144[31] , \Level4Load204[0] , \Level2Out52[31] , 
        \Level2Out52[28] , \Level1Out80[21] , \Level1Out199[7] , 
        \Level32Out32[27] , \Level32Out64[26] , \Level128Out0[14] , 
        \Level1Out95[15] , \Level2Out124[2] , \Level1Out184[8] , 
        \Level2Out244[7] , \Level16Out48[24] , \ScanLink216[3] , 
        \Level1Out9[21] , \ScanLink12[20] , \Level1Out14[1] , \ScanLink48[4] , 
        \ScanLink82[30] , \ScanLink176[6] , \Level8Out40[14] , 
        \Level8Load168[0] , \Level8Out16[15] , \Level1Out17[2] , 
        \ScanLink79[28] , \ScanLink82[29] , \Level1Out148[2] , 
        \ScanLink212[31] , \ScanLink212[28] , \ScanLink244[30] , 
        \ScanLink215[0] , \ScanLink231[19] , \ScanLink244[29] , 
        \Level4Out56[3] , \ScanLink31[11] , \ScanLink34[2] , \ScanLink37[1] , 
        \Level1Out38[15] , \ScanLink56[8] , \ScanLink79[31] , 
        \Level1Out228[7] , \ScanLink99[1] , \ScanLink175[5] , 
        \Level1Out58[11] , \Level1Load152[0] , \Level1Out202[29] , 
        \Level4Out84[5] , \Level1Out254[31] , \Level2Out238[29] , 
        \Level1Out101[22] , \Level1Out114[16] , \Level1Out137[27] , 
        \Level1Out202[30] , \Level1Out235[8] , \Level1Out221[18] , 
        \Level1Out254[28] , \Level2Out238[30] , \Level1Out142[17] , 
        \Level2Out178[17] , \Level64Out128[18] , \Level1Out161[26] , 
        \ScanLink111[23] , \Level1Out122[13] , \Level1Out174[12] , 
        \Level8Out8[8] , \Level1Out157[23] , \Level2Out118[13] , 
        \ScanLink132[12] , \Level1Out134[4] , \ScanLink164[13] , 
        \ScanLink89[25] , \ScanLink104[17] , \ScanLink109[3] , 
        \ScanLink147[22] , \Level1Out254[1] , \Level2Out146[8] , 
        \Level4Out0[25] , \ScanLink127[26] , \ScanLink152[16] , 
        \Level2Out94[13] , \ScanLink171[27] , \ScanLink219[24] , 
        \ScanLink44[21] , \ScanLink67[10] , \Level1Out137[7] , 
        \Level8Out232[1] , \ScanLink24[25] , \ScanLink51[15] , 
        \Level1Out68[7] , \ScanLink72[24] , \Level8Out152[4] , 
        \Level4Out192[20] , \Level1Out9[12] , \Level1Out10[31] , 
        \Level1Out46[29] , \Level1Out75[8] , \Level2Out158[4] , 
        \Level2Out226[11] , \Level1Out209[25] , \Level2Out238[1] , 
        \Level2Out246[15] , \Level1Out10[28] , \Level1Out33[19] , 
        \Level2Out196[22] , \Level1Out46[30] , \Level1Out65[18] , 
        \Level4Out84[13] , \ScanLink53[5] , \Level2Out8[19] , 
        \Level2Out210[14] , \ScanLink81[3] , \ScanLink89[16] , 
        \ScanLink127[15] , \ScanLink152[25] , \Level4Out0[16] , 
        \Level2Load42[0] , \ScanLink104[24] , \Level1Out150[0] , 
        \ScanLink171[14] , \Level4Out108[3] , \ScanLink111[10] , 
        \ScanLink164[20] , \Level2Out94[20] , \ScanLink132[21] , 
        \ScanLink147[11] , \Level2Out242[9] , \Level1Out230[5] , 
        \Level1Out174[21] , \ScanLink82[0] , \Level1Out101[11] , 
        \Level1Out114[25] , \Level1Out122[20] , \Level1Out157[10] , 
        \Level1Out182[6] , \Level2Out118[20] , \Level8Out248[9] , 
        \Level1Out137[14] , \Level1Out142[24] , \Level2Out66[0] , 
        \Level2Out178[24] , \Level1Out161[15] , \ScanLink170[8] , 
        \Level8Load48[0] , \Level1Out181[5] , \Level1Out209[16] , 
        \Level2Out196[11] , \Level2Out246[26] , \Level2Out210[27] , 
        \Level4Out84[20] , \Level4Out192[13] , \Level2Out226[22] , 
        \ScanLink0[14] , \Level1Out1[0] , \Level1Out2[3] , \Level1Out6[26] , 
        \ScanLink12[13] , \ScanLink24[16] , \ScanLink72[17] , 
        \Level1Out153[3] , \ScanLink31[22] , \ScanLink50[6] , \ScanLink51[26] , 
        \Level1Out233[6] , \Level8Out136[0] , \ScanLink44[12] , 
        \ScanLink219[17] , \ScanLink16[3] , \ScanLink67[23] , 
        \Level1Out195[20] , \Level1Out230[27] , \ScanLink15[0] , 
        \Level1Out57[9] , \ScanLink68[17] , \Level1Out108[9] , 
        \Level1Out115[6] , \Level1Out213[16] , \Level1Out245[17] , 
        \ScanLink248[4] , \ScanLink128[1] , \Level1Out180[14] , 
        \Level1Out206[22] , \Level16Out176[15] , \Level1Out225[13] , 
        \ScanLink190[15] , \ScanLink216[23] , \Level1Out250[23] , 
        \Level4Out188[13] , \ScanLink235[12] , \Level2Out56[10] , 
        \Level1Out98[0] , \ScanLink240[22] , \Level4Out16[8] , 
        \ScanLink86[22] , \ScanLink93[16] , \ScanLink185[21] , 
        \ScanLink203[17] , \ScanLink220[26] , \ScanLink255[16] , 
        \Level2Out60[15] , \ScanLink256[8] , \Level2Out36[14] , 
        \ScanLink128[21] , \ScanLink148[25] , \Level1Out116[5] , 
        \Level2Out20[5] , \Level1Out138[20] , \Level2Out102[20] , 
        \Level1Out49[5] , \Level2Out0[7] , \Level2Out154[21] , 
        \Level2Out164[9] , \Level2Out134[25] , \Level1Out158[24] , 
        \Level2Out162[24] , \ScanLink185[12] , \ScanLink255[25] , 
        \Level2Out60[26] , \ScanLink203[24] , \ScanLink220[15] , 
        \ScanLink216[10] , \Level2Out36[27] , \Level2Out56[23] , 
        \Level1Out6[15] , \ScanLink68[24] , \ScanLink190[26] , 
        \ScanLink235[21] , \ScanLink240[11] , \ScanLink72[7] , 
        \Level1Out171[2] , \Level1Out206[11] , \Level16Out176[26] , 
        \Level1Out180[27] , \Level1Out225[20] , \Level1Out250[10] , 
        \Level4Out188[20] , \Level1Out29[19] , \Level1Out195[13] , 
        \Level1Out211[7] , \Level1Out245[24] , \Level1Out230[14] , 
        \ScanLink71[4] , \Level1Out213[25] , \Level2Out134[16] , 
        \Level1Out84[19] , \Level1Out138[13] , \Level1Out158[17] , 
        \Level1Out172[1] , \Level2Out102[13] , \Level2Out162[17] , 
        \Level1Out212[4] , \Level2Out96[7] , \ScanLink86[11] , 
        \ScanLink128[12] , \Level2Out154[12] , \ScanLink93[25] , 
        \ScanLink148[16] , \Level2Out44[1] , \Level8Out72[29] , 
        \Level8Out24[31] , \ScanLink152[9] , \Level8Out72[30] , 
        \ScanLink4[25] , \ScanLink4[16] , \Level1Out14[10] , \ScanLink16[18] , 
        \ScanLink35[30] , \ScanLink35[29] , \Level1Out113[8] , 
        \Level8Out24[28] , \ScanLink208[31] , \Level4Out184[2] , 
        \ScanLink208[28] , \ScanLink40[19] , \ScanLink63[31] , 
        \Level1Out83[1] , \Level1Out37[21] , \ScanLink63[28] , 
        \Level2Out38[7] , \ScanLink253[5] , \Level1Out42[11] , 
        \Level4Out156[4] , \Level1Out22[15] , \Level1Out61[20] , 
        \Level1Out74[14] , \ScanLink133[0] , \Level2Out222[30] , 
        \Level4Out196[18] , \Level1Out218[30] , \Level4Out236[1] , 
        \Level1Out51[7] , \Level2Out222[29] , \Level1Out57[25] , 
        \Level1Out218[29] , \Level4Out4[1] , \Level16Out64[21] , 
        \Level128Out0[2] , \Level1Out14[23] , \Level1Out22[26] , 
        \Level1Out52[4] , \ScanLink250[6] , \Level8Out208[2] , 
        \Level16Out32[20] , \Level1Out57[16] , \ScanLink69[6] , 
        \Level1Out74[27] , \Level1Out80[2] , \ScanLink98[29] , 
        \ScanLink130[3] , \Level8Out168[7] , \Level2Out162[7] , 
        \Level4Out148[8] , \ScanLink98[30] , \Level2Out6[9] , 
        \Level2Out202[2] , \ScanLink237[1] , \Level1Out35[3] , 
        \Level4Out132[0] , \Level1Out37[12] , \Level1Out42[22] , 
        \Level1Out61[13] , \ScanLink157[4] , \Level2Out192[29] , 
        \Level4Out80[18] , \Level4Out252[5] , \Level1Load17[0] , 
        \ScanLink74[9] , \Level2Out192[30] , \Level1Out36[0] , 
        \Level1Out105[29] , \ScanLink115[31] , \ScanLink115[28] , 
        \ScanLink185[2] , \Level2Out48[31] , \Level1Out217[9] , 
        \Level2Out48[28] , \ScanLink136[19] , \ScanLink143[30] , 
        \ScanLink160[18] , \ScanLink143[29] , \ScanLink149[8] , 
        \ScanLink186[1] , \Level2Out106[3] , \ScanLink154[7] , 
        \Level1Out169[0] , \ScanLink234[2] , \Level2Out90[18] , 
        \Level2Out90[9] , \Level1Out209[5] , \Level8Out80[4] , 
        \Level1Out126[18] , \Level1Out153[31] , \Level1Out170[19] , 
        \Level16Out64[12] , \Level16Out32[13] , \Level1Out105[30] , 
        \Level1Out12[6] , \ScanLink111[19] , \Level1Out153[28] , 
        \ScanLink164[29] , \Level2Out242[0] , \ScanLink132[31] , 
        \ScanLink132[28] , \ScanLink147[18] , \ScanLink164[30] , 
        \Level1Out150[9] , \Level2Out94[30] , \Level2Out122[5] , 
        \Level2Out94[29] , \Level1Out101[18] , \ScanLink170[1] , 
        \Level2Out66[9] , \Level64Out128[22] , \Level8Out128[5] , 
        \Level1Out174[28] , \Level2Out118[30] , \Level1Out122[30] , 
        \Level1Out11[5] , \Level1Out26[17] , \Level1Out70[16] , 
        \Level1Out122[29] , \Level1Out157[19] , \Level8Out248[0] , 
        \Level1Out174[31] , \ScanLink210[4] , \Level2Out118[29] , 
        \ScanLink173[2] , \ScanLink0[27] , \Level1Out10[12] , 
        \Level1Out33[23] , \Level1Out53[27] , \ScanLink213[7] , 
        \Level2Out196[18] , \Level4Out84[30] , \Level1Out46[13] , 
        \ScanLink82[9] , \Level4Out116[6] , \Level1Out65[22] , 
        \Level2Out8[23] , \Level4Out84[29] , \Level1Out76[2] , 
        \ScanLink114[5] , \Level1Out249[7] , \Level2Out78[5] , 
        \Level8Out136[9] , \Level8Out8[1] , \Level1Out9[28] , 
        \Level1Out10[21] , \ScanLink12[30] , \ScanLink37[8] , 
        \Level1Out129[2] , \Level1Load133[0] , \Level1Out254[8] , 
        \Level2Out194[7] , \Level64Out128[11] , \Level2Out226[4] , 
        \ScanLink44[28] , \Level2Out146[1] , \ScanLink12[29] , 
        \ScanLink31[18] , \ScanLink44[31] , \Level8Out232[8] , 
        \ScanLink67[19] , \Level1Out33[10] , \Level1Out46[20] , 
        \Level1Out75[1] , \Level2Out238[8] , \Level1Out65[11] , 
        \ScanLink117[6] , \Level2Out8[10] , \ScanLink29[4] , 
        \Level2Load122[0] , \Level4Out212[7] , \Level1Out70[25] , 
        \Level1Out53[14] , \Level4Out192[29] , \ScanLink1[9] , 
        \Level1Out2[24] , \ScanLink9[1] , \Level1Out9[31] , \Level2Out226[18] , 
        \Level1Out14[8] , \Level1Out26[24] , \Level4Out172[2] , 
        \Level4Out192[30] , \ScanLink55[2] , \Level1Out80[31] , 
        \Level1Out129[16] , \Level1Out236[2] , \Level2Out130[27] , 
        \Level1Out149[12] , \Level1Out156[7] , \Level2Out166[26] , 
        \Level4Out48[6] , \Level2Out106[22] , \Level1Out80[28] , 
        \Level2Out150[23] , \ScanLink159[13] , \ScanLink82[20] , 
        \Level1Out184[1] , \Level2Out60[7] , \ScanLink19[25] , 
        \ScanLink79[21] , \ScanLink87[4] , \ScanLink97[14] , \ScanLink139[17] , 
        \ScanLink84[7] , \ScanLink181[23] , \ScanLink207[15] , 
        \ScanLink224[24] , \ScanLink251[14] , \Level2Out64[17] , 
        \Level2Out32[16] , \Level1Out187[2] , \ScanLink194[17] , 
        \ScanLink212[21] , \ScanLink231[10] , \Level2Out52[12] , 
        \ScanLink215[9] , \ScanLink244[20] , \ScanLink56[1] , \ScanLink99[8] , 
        \ScanLink168[3] , \Level1Out184[16] , \Level1Out202[20] , 
        \Level1Out221[11] , \Level1Out235[1] , \Level2Out238[20] , 
        \Level1Out254[21] , \Level16Out144[12] , \Level1Out191[22] , 
        \Level32Out192[2] , \Level1Out234[25] , \Level1Out241[15] , 
        \Level1Out2[17] , \ScanLink31[6] , \Level1Out58[18] , 
        \Level1Out217[14] , \ScanLink82[13] , \ScanLink97[27] , 
        \Level1Out155[4] , \ScanLink208[6] , \Level8Load216[0] , 
        \Level2Out188[13] , \Level16Out112[13] , \ScanLink139[24] , 
        \ScanLink159[20] , \Level2Out192[9] , \Level1Out149[21] , 
        \Level2Out106[11] , \Level1Out252[6] , \Level2Out130[14] , 
        \Level2Out150[10] , \Level1Out129[25] , \Level1Out132[3] , 
        \Level2Out166[15] , \Level1Out241[26] , \Level1Out8[22] , 
        \ScanLink19[16] , \ScanLink32[5] , \Level1Out131[0] , 
        \Level1Out191[11] , \Level1Out251[5] , \Level1Out217[27] , 
        \Level1Out234[16] , \Level2Out188[20] , \Level16Out112[20] , 
        \Level16Out144[21] , \Level1Out202[13] , \Level2Out238[13] , 
        \ScanLink111[8] , \Level1Out184[25] , \Level1Out221[22] , 
        \Level1Out254[12] , \Level2Out52[21] , \ScanLink212[12] , 
        \ScanLink244[13] , \ScanLink79[12] , \ScanLink194[24] , 
        \ScanLink231[23] , \ScanLink251[27] , \Level2Out64[24] , 
        \ScanLink181[10] , \ScanLink207[26] , \ScanLink224[17] , 
        \Level2Out32[25] , \Level1Out208[26] , \Level2Out182[15] , 
        \Level2Out228[2] , \Level2Out232[26] , \Level2Out252[22] , 
        \Level4Out200[21] , \Level2Out204[23] , \Level4Out236[24] , 
        \ScanLink13[23] , \ScanLink25[26] , \ScanLink50[16] , 
        \Level2Out148[7] , \Level1Out247[1] , \Level2Out38[10] , 
        \ScanLink66[13] , \ScanLink73[27] , \Level1Out78[4] , 
        \Level1Out127[4] , \Level8Out8[17] , \ScanLink13[10] , \ScanLink24[1] , 
        \ScanLink218[27] , \ScanLink27[2] , \ScanLink30[12] , \ScanLink45[22] , 
        \Level2Out58[14] , \ScanLink88[26] , \ScanLink105[14] , 
        \ScanLink119[0] , \ScanLink170[24] , \Level1Out244[2] , 
        \ScanLink126[25] , \ScanLink133[11] , \ScanLink153[15] , 
        \Level1Out66[8] , \ScanLink110[20] , \ScanLink146[21] , 
        \Level1Out123[10] , \Level1Out124[7] , \Level2Out80[24] , 
        \ScanLink165[10] , \Level1Out100[21] , \Level1Out156[20] , 
        \Level4Out28[10] , \Level2Out12[7] , \Level1Out115[15] , 
        \Level1Out175[11] , \Level4Out108[26] , \Level1Out136[24] , 
        \Level1Out160[25] , \Level4Out168[22] , \Level4Out48[14] , 
        \Level1Out139[8] , \Level1Out143[14] , \ScanLink25[15] , 
        \ScanLink30[21] , \ScanLink66[20] , \Level1Out223[5] , 
        \Level2Out58[27] , \ScanLink45[11] , \ScanLink218[14] , 
        \Level16Out0[1] , \ScanLink40[5] , \ScanLink50[25] , \ScanLink73[14] , 
        \Level1Out143[0] , \Level2Out38[23] , \Level4Out92[8] , 
        \Level8Out8[24] , \ScanLink4[4] , \ScanLink7[7] , \Level1Out8[11] , 
        \Level2Out182[26] , \Level2Out252[11] , \Level4Out236[17] , 
        \Level1Out11[18] , \Level1Out32[30] , \ScanLink92[3] , 
        \ScanLink163[8] , \Level2Out204[10] , \Level1Out32[29] , 
        \Level1Out64[28] , \Level1Out191[6] , \Level1Out39[25] , 
        \ScanLink43[6] , \Level1Out47[19] , \Level1Out64[31] , 
        \Level2Out232[15] , \Level4Out200[12] , \Level1Out208[15] , 
        \ScanLink88[15] , \ScanLink91[0] , \Level1Out115[26] , 
        \Level1Out160[16] , \Level8Out152[28] , \Level1Out123[23] , 
        \Level1Out136[17] , \Level1Out143[27] , \Level4Out168[11] , 
        \Level8Out104[30] , \Level2Out76[3] , \Level8Out152[31] , 
        \Level4Out48[27] , \Level1Out156[13] , \Level1Out192[5] , 
        \Level8Out104[29] , \Level4Out28[23] , \Level1Out175[22] , 
        \Level4Out108[15] , \Level1Out100[12] , \ScanLink110[13] , 
        \ScanLink133[22] , \ScanLink146[12] , \Level1Out220[6] , 
        \ScanLink165[23] , \Level4Load108[0] , \Level2Out80[17] , 
        \ScanLink105[27] , \Level1Out140[3] , \ScanLink170[17] , 
        \Level1Out59[21] , \Level1Out63[5] , \ScanLink126[16] , 
        \ScanLink153[26] , \ScanLink78[18] , \Level1Load93[0] , 
        \ScanLink101[2] , \ScanLink230[29] , \ScanLink245[19] , 
        \ScanLink213[18] , \ScanLink230[30] , \Level4Out204[3] , 
        \Level4Out164[6] , \Level8Out0[9] , \Level1Out220[28] , 
        \Level1Out255[18] , \Level2Out2[25] , \Level8Out144[9] , 
        \Level8Out224[13] , \Level1Out39[16] , \Level1Out60[6] , 
        \Level1Out81[11] , \Level1Out203[19] , \Level1Out220[31] , 
        \Level1Out94[25] , \Level1Out122[9] , \Level2Out230[0] , 
        \Level4Out120[28] , \Level4Out176[30] , \ScanLink102[1] , 
        \Level2Out150[5] , \Level4Out120[31] , \Level4Out176[29] , 
        \ScanLink83[19] , \Level2Out14[9] , \ScanLink178[9] , 
        \Level2Out182[3] , \Level2Out2[16] , \Level1Out59[12] , 
        \Level1Out190[31] , \Level8Out224[20] , \Level8Out240[8] , 
        \Level64Out128[0] , \ScanLink45[8] , \ScanLink58[7] , \ScanLink89[2] , 
        \Level1Out190[28] , \Level4Out248[18] , \ScanLink158[19] , 
        \Level1Out158[1] , \ScanLink165[6] , \ScanLink180[30] , 
        \Level1Out238[4] , \ScanLink180[29] , \Level1Out197[8] , 
        \ScanLink205[3] , \Level2Out26[31] , \ScanLink166[5] , 
        \Level2Out26[28] , \Level2Out70[29] , \Level4Out100[2] , 
        \Level2Out70[30] , \Level2Load150[0] , \Level1Out94[16] , 
        \Level1Load141[0] , \ScanLink206[0] , \Level2Out254[4] , 
        \Level1Out226[8] , \Level1Out81[22] , \Level4Out60[29] , 
        \Level1Out189[4] , \Level2Out124[19] , \Level4Out36[31] , 
        \Level2Out134[1] , \Level2Out172[18] , \Level4Out60[30] , 
        \Level1Out148[18] , \Level4Out36[28] , \ScanLink2[8] , 
        \Level1Out8[20] , \Level1Out9[8] , \ScanLink17[21] , \ScanLink18[5] , 
        \Level1Out20[4] , \ScanLink129[18] , \ScanLink222[6] , 
        \ScanLink142[3] , \Level8Out96[0] , \Level1Out23[7] , 
        \Level1Out28[13] , \Level1Out48[17] , \Level1Out85[13] , 
        \Level1Out90[27] , \ScanLink190[5] , \Level2Out110[7] , 
        \Level2Out120[28] , \Level1Out139[19] , \Level2Out120[31] , 
        \Level2Out176[30] , \Level4Out64[18] , \Level8Out128[16] , 
        \Level2Out176[29] , \Level4Out32[19] , \Level1Out161[8] , 
        \Level1Load206[0] , \Level2Out6[27] , \Level8Out216[14] , 
        \Level8Out240[15] , \ScanLink184[18] , \ScanLink193[6] , 
        \Level1Out194[19] , \Level16Out80[9] , \ScanLink221[5] , 
        \Level16Load80[0] , \Level16Out80[12] , \Level4Out124[4] , 
        \Level1Out85[20] , \ScanLink141[0] , \Level2Out74[18] , 
        \Level2Out98[1] , \Level8Out88[22] , \Level2Out22[19] , 
        \Level128Out128[14] , \Level4Out244[1] , \Level8Out128[25] , 
        \Level1Out90[14] , \Level1Out96[6] , \Level2Out174[3] , 
        \Level2Out214[6] , \Level4Out124[19] , \Level4Out172[18] , 
        \Level1Out28[20] , \Level1Out44[0] , \ScanLink246[2] , 
        \Level1Out47[3] , \ScanLink87[31] , \ScanLink87[28] , \ScanLink126[7] , 
        \Level1Out118[3] , \ScanLink217[30] , \ScanLink234[18] , 
        \ScanLink245[1] , \ScanLink125[4] , \ScanLink217[29] , 
        \ScanLink241[28] , \Level8Out88[11] , \Level4Out140[0] , 
        \ScanLink241[31] , \Level128Out128[27] , \Level4Out220[5] , 
        \Level1Out48[24] , \Level1Load65[0] , \Level4Out192[6] , 
        \Level16Out80[21] , \Level1Out95[5] , \Level1Out207[31] , 
        \Level8Out216[27] , \Level1Out224[19] , \Level1Out251[29] , 
        \Level2Out6[14] , \Level1Out207[28] , \ScanLink62[11] , 
        \ScanLink67[0] , \Level1Out104[23] , \Level1Out111[17] , 
        \Level1Out251[30] , \Level2Out248[18] , \Level8Out240[26] , 
        \Level1Out127[12] , \Level1Out132[26] , \Level1Out164[27] , 
        \Level1Out147[16] , \ScanLink224[8] , \Level2Out108[26] , 
        \Level16Out192[26] , \Level2Out168[22] , \Level1Out152[22] , 
        \Level2Out52[5] , \ScanLink137[13] , \Level1Out171[13] , 
        \Level32Out192[13] , \ScanLink99[10] , \ScanLink114[22] , 
        \ScanLink142[23] , \Level2Out116[9] , \ScanLink239[7] , 
        \Level2Out84[26] , \ScanLink161[12] , \Level1Out164[5] , 
        \ScanLink101[16] , \ScanLink122[27] , \ScanLink174[26] , 
        \Level2Out80[3] , \Level1Out204[0] , \ScanLink157[17] , 
        \ScanLink159[2] , \Level1Out167[6] , \ScanLink21[24] , 
        \ScanLink34[10] , \ScanLink41[20] , \ScanLink64[3] , \ScanLink54[14] , 
        \ScanLink195[8] , \Level1Out207[3] , \Level8Out96[30] , 
        \ScanLink209[11] , \ScanLink13[21] , \Level1Out15[30] , 
        \Level1Out15[29] , \Level1Out38[6] , \Level8Out96[29] , 
        \Level1Out43[31] , \ScanLink77[25] , \Level1Out219[10] , 
        \Level2Out108[5] , \Level2Out186[17] , \Level2Out200[21] , 
        \Level4Out64[8] , \Level4Out232[26] , \Level1Out60[19] , 
        \ScanLink188[7] , \Level4Out252[22] , \Level1Out25[9] , 
        \Level1Out43[28] , \Level2Out236[24] , \ScanLink17[12] , 
        \ScanLink21[17] , \Level1Out36[18] , \Level4Out204[23] , 
        \Level1Out90[8] , \Level1Out100[1] , \ScanLink101[25] , 
        \ScanLink174[15] , \ScanLink122[14] , \ScanLink157[24] , 
        \Level2Load108[0] , \ScanLink137[20] , \ScanLink142[10] , 
        \ScanLink161[21] , \ScanLink99[23] , \Level1Out104[10] , 
        \ScanLink114[11] , \Level2Out84[15] , \Level2Out212[8] , 
        \Level1Out127[21] , \Level1Out152[11] , \Level1Out171[20] , 
        \Level2Out168[11] , \Level32Out192[20] , \Level1Out111[24] , 
        \ScanLink120[9] , \Level1Out164[14] , \Level1Load119[0] , 
        \Level1Out132[15] , \Level1Out147[25] , \Level2Out36[1] , 
        \Level2Out108[15] , \Level16Out192[15] , \Level1Out219[23] , 
        \Level2Out186[24] , \Level2Out236[17] , \Level4Out204[10] , 
        \Level4Out252[11] , \Level2Out200[12] , \Level4Out232[15] , 
        \ScanLink54[27] , \ScanLink77[16] , \Level1Out103[2] , 
        \ScanLink209[22] , \ScanLink27[0] , \ScanLink34[23] , \ScanLink62[22] , 
        \ScanLink41[13] , \Level1Out100[23] , \Level1Out115[17] , 
        \Level1Out160[27] , \Level4Out168[20] , \Level8Out152[19] , 
        \Level1Out123[12] , \Level1Out136[26] , \Level1Out143[16] , 
        \Level1Out156[22] , \Level2Out12[5] , \Level4Out48[16] , 
        \Level8Out104[18] , \Level4Out28[12] , \Level1Out175[13] , 
        \Level4Out108[24] , \ScanLink133[13] , \ScanLink146[23] , 
        \Level2Out156[9] , \ScanLink88[24] , \ScanLink110[22] , 
        \ScanLink165[12] , \Level2Out80[26] , \Level1Out124[5] , 
        \ScanLink105[16] , \ScanLink170[26] , \ScanLink119[2] , 
        \ScanLink126[27] , \ScanLink153[17] , \Level1Out244[0] , 
        \ScanLink24[3] , \ScanLink30[10] , \ScanLink66[11] , \Level1Out127[6] , 
        \Level2Out58[16] , \ScanLink25[24] , \ScanLink45[20] , 
        \ScanLink218[25] , \ScanLink50[14] , \ScanLink73[25] , 
        \Level1Out247[3] , \Level2Out38[12] , \Level8Out8[15] , 
        \Level1Out78[6] , \Level2Out182[17] , \Level2Out252[20] , 
        \Level4Out24[8] , \Level1Out11[30] , \Level1Out11[29] , 
        \Level2Out148[5] , \Level2Out204[21] , \Level4Out236[26] , 
        \Level1Out32[18] , \Level1Out47[31] , \Level1Out64[19] , 
        \Level2Out228[0] , \Level4Out200[23] , \Level1Out47[28] , 
        \Level1Out65[9] , \Level2Out232[24] , \Level1Out208[24] , 
        \ScanLink4[6] , \Level1Out8[13] , \ScanLink43[4] , \ScanLink88[17] , 
        \ScanLink105[25] , \Level1Out140[1] , \ScanLink126[14] , 
        \ScanLink170[15] , \Level2Load148[0] , \ScanLink91[2] , 
        \Level1Out100[10] , \ScanLink110[11] , \ScanLink133[20] , 
        \ScanLink153[24] , \ScanLink146[10] , \Level1Out220[4] , 
        \Level2Out80[15] , \Level2Out252[8] , \Level1Out123[21] , 
        \ScanLink165[21] , \Level1Out156[11] , \Level1Out192[7] , 
        \Level4Out28[21] , \ScanLink92[1] , \Level1Out115[24] , 
        \Level1Out175[20] , \Level4Out108[17] , \Level4Out168[13] , 
        \Level1Out136[15] , \ScanLink160[9] , \Level1Out160[14] , 
        \Level1Out143[25] , \Level2Out76[1] , \Level4Out48[25] , 
        \Level1Load159[0] , \Level1Out191[4] , \Level1Out208[17] , 
        \Level2Out232[17] , \Level2Out252[13] , \Level4Out200[10] , 
        \Level2Out182[24] , \Level2Out204[12] , \ScanLink13[12] , 
        \ScanLink25[17] , \ScanLink50[27] , \Level4Out236[15] , 
        \Level2Out38[21] , \ScanLink40[7] , \ScanLink66[22] , \ScanLink73[16] , 
        \Level8Out8[26] , \Level1Out143[2] , \Level4Load8[0] , 
        \ScanLink30[23] , \ScanLink45[13] , \ScanLink218[16] , 
        \Level1Out223[7] , \Level2Out58[25] , \Level16Out0[3] , 
        \Level1Out39[27] , \Level1Out60[4] , \ScanLink102[3] , 
        \ScanLink158[31] , \ScanLink158[28] , \Level2Out182[1] , 
        \Level1Out81[13] , \Level1Out94[27] , \Level2Out150[7] , 
        \Level2Out172[30] , \Level4Out60[18] , \Level1Out121[8] , 
        \Level1Out148[30] , \Level2Out124[28] , \Level1Out148[29] , 
        \Level2Out124[31] , \Level2Out172[29] , \Level2Out230[2] , 
        \Level4Out36[19] , \Level1Load246[0] , \Level2Out2[27] , 
        \Level1Out59[23] , \Level4Out248[30] , \Level1Out63[7] , 
        \ScanLink180[18] , \Level1Out190[19] , \Level4Out248[29] , 
        \Level8Out224[11] , \Level4Out164[4] , \Level2Out70[18] , 
        \Level1Out81[20] , \ScanLink101[0] , \Level2Out26[19] , 
        \Level4Out204[1] , \Level2Out134[3] , \Level1Out1[2] , 
        \Level1Out6[24] , \ScanLink7[5] , \ScanLink58[5] , \Level1Out94[14] , 
        \Level1Out189[6] , \Level2Out254[6] , \Level4Out120[19] , 
        \Level4Out176[18] , \ScanLink78[30] , \ScanLink83[31] , 
        \ScanLink83[28] , \Level1Out194[9] , \ScanLink206[2] , 
        \Level1Out158[3] , \ScanLink166[7] , \ScanLink205[1] , 
        \ScanLink230[18] , \ScanLink245[28] , \Level4Out100[0] , 
        \ScanLink213[30] , \ScanLink213[29] , \ScanLink245[31] , 
        \ScanLink78[29] , \ScanLink165[4] , \Level1Out238[6] , \ScanLink15[2] , 
        \Level1Out15[18] , \ScanLink17[23] , \ScanLink18[7] , \Level1Out20[6] , 
        \Level1Out23[5] , \Level1Load25[0] , \Level1Out59[10] , 
        \Level64Out128[2] , \Level8Out224[22] , \Level1Out39[14] , 
        \ScanLink46[9] , \ScanLink89[0] , \Level1Out203[31] , 
        \Level1Out220[19] , \Level1Out225[9] , \Level1Out255[29] , 
        \Level2Out2[14] , \Level1Out203[28] , \Level1Out255[30] , 
        \ScanLink234[29] , \ScanLink241[19] , \Level2Out98[3] , 
        \Level8Out88[20] , \Level1Out28[11] , \ScanLink141[2] , 
        \ScanLink217[18] , \ScanLink234[30] , \Level4Out244[3] , 
        \ScanLink221[7] , \Level4Out124[6] , \Level128Out128[16] , 
        \Level1Out48[15] , \ScanLink193[4] , \Level8Out104[9] , 
        \Level16Out80[10] , \Level1Out224[28] , \Level8Out216[16] , 
        \Level1Out251[18] , \Level2Out248[30] , \Level2Out6[25] , 
        \Level1Out85[11] , \Level1Out207[19] , \Level1Out224[31] , 
        \Level2Out248[29] , \Level8Out128[14] , \Level8Out240[17] , 
        \Level1Out90[25] , \Level1Out162[9] , \ScanLink190[7] , 
        \Level4Out124[28] , \Level4Out172[30] , \Level2Out110[5] , 
        \Level4Out124[31] , \Level4Out172[29] , \ScanLink142[1] , 
        \Level8Out96[2] , \Level2Out54[9] , \Level1Out28[22] , 
        \Level1Out48[26] , \ScanLink87[19] , \ScanLink222[4] , 
        \Level1Out95[7] , \ScanLink138[9] , \Level2Out6[16] , 
        \Level4Load88[0] , \Level8Out216[25] , \Level8Out240[24] , 
        \Level4Out192[4] , \Level1Out44[2] , \Level1Out47[1] , 
        \Level1Out88[8] , \ScanLink125[6] , \Level1Out194[31] , 
        \Level8Out200[8] , \Level1Out194[28] , \Level4Out220[7] , 
        \Level16Out80[23] , \ScanLink184[30] , \Level1Out118[1] , 
        \ScanLink184[29] , \ScanLink245[3] , \Level2Out74[29] , 
        \Level4Out140[2] , \Level2Out22[31] , \Level8Out88[13] , 
        \Level2Out22[28] , \Level2Out74[30] , \Level128Out128[25] , 
        \Level2Load110[0] , \ScanLink126[5] , \ScanLink129[30] , 
        \ScanLink129[29] , \ScanLink21[26] , \Level1Out85[22] , 
        \Level1Out90[16] , \Level1Out96[4] , \Level1Load101[0] , 
        \ScanLink246[0] , \Level2Out214[4] , \Level2Out120[19] , 
        \Level4Out32[31] , \Level1Out139[31] , \Level2Out174[1] , 
        \Level4Out64[29] , \Level1Out139[28] , \Level2Out176[18] , 
        \Level4Out32[28] , \Level8Out128[27] , \Level4Out64[30] , 
        \ScanLink188[5] , \Level4Out252[20] , \Level1Out219[12] , 
        \Level2Out186[15] , \Level2Out236[26] , \Level4Out204[21] , 
        \ScanLink227[9] , \Level2Out108[7] , \Level2Out200[23] , 
        \Level4Out232[24] , \Level1Out38[4] , \ScanLink54[16] , 
        \ScanLink77[27] , \Level1Out207[1] , \ScanLink209[13] , 
        \ScanLink17[10] , \Level1Out26[8] , \ScanLink34[12] , \ScanLink62[13] , 
        \Level1Out167[4] , \Level8Load224[0] , \ScanLink41[22] , 
        \ScanLink64[1] , \ScanLink67[2] , \ScanLink101[14] , \ScanLink174[24] , 
        \Level2Out80[1] , \ScanLink122[25] , \ScanLink157[15] , 
        \ScanLink159[0] , \ScanLink196[9] , \Level1Out204[2] , 
        \ScanLink137[11] , \ScanLink142[21] , \ScanLink99[12] , 
        \ScanLink161[10] , \ScanLink114[20] , \Level1Out127[10] , 
        \Level1Out152[20] , \Level1Out164[7] , \ScanLink239[5] , 
        \Level2Out84[24] , \Level2Out52[7] , \ScanLink62[20] , 
        \Level1Out104[21] , \Level1Out171[11] , \Level2Out168[20] , 
        \Level32Out192[11] , \Level1Out111[15] , \Level1Out164[25] , 
        \Level1Out132[24] , \Level1Out147[14] , \Level2Out108[24] , 
        \Level16Out192[24] , \Level1Out179[8] , \Level1Out93[9] , 
        \ScanLink21[15] , \ScanLink34[21] , \ScanLink41[11] , \ScanLink54[25] , 
        \ScanLink209[20] , \Level1Out60[28] , \ScanLink77[14] , 
        \Level8Out96[18] , \Level1Out103[0] , \ScanLink123[8] , 
        \Level1Out219[21] , \Level2Out186[26] , \Level2Out200[10] , 
        \Level4Out232[17] , \Level4Out252[13] , \Level1Out36[30] , 
        \Level1Out36[29] , \Level1Out43[19] , \Level1Out60[31] , 
        \Level2Out236[15] , \Level1Out49[7] , \ScanLink99[21] , 
        \Level1Out104[12] , \Level1Out111[26] , \Level4Out204[12] , 
        \Level1Out127[23] , \Level1Out132[17] , \Level1Out164[16] , 
        \Level1Out147[27] , \Level2Out36[3] , \Level2Out108[17] , 
        \Level16Out192[17] , \Level2Out168[13] , \Level1Out152[13] , 
        \ScanLink114[13] , \ScanLink137[22] , \Level1Out171[22] , 
        \Level32Out192[22] , \ScanLink142[12] , \ScanLink161[23] , 
        \Level2Out84[17] , \Level1Out100[3] , \ScanLink101[27] , 
        \Level4Load148[0] , \ScanLink122[16] , \ScanLink174[17] , 
        \ScanLink157[26] , \Level1Out158[26] , \Level2Out0[5] , 
        \Level2Out134[27] , \Level1Out84[31] , \Level2Out102[22] , 
        \Level2Out162[26] , \Level1Out84[28] , \Level1Out116[7] , 
        \Level1Out138[22] , \Level2Out154[23] , \Level1Out29[31] , 
        \Level1Out54[8] , \ScanLink86[20] , \ScanLink128[23] , 
        \Level2Out20[7] , \ScanLink68[15] , \ScanLink93[14] , \Level1Out98[2] , 
        \ScanLink148[27] , \Level8Out72[18] , \ScanLink255[14] , 
        \Level2Out60[17] , \Level8Out24[19] , \ScanLink185[23] , 
        \ScanLink220[24] , \ScanLink190[17] , \ScanLink203[15] , 
        \Level2Out36[16] , \ScanLink216[21] , \Level2Out56[12] , 
        \ScanLink240[20] , \ScanLink235[10] , \ScanLink255[9] , 
        \Level32Out64[9] , \ScanLink128[3] , \Level1Out206[20] , 
        \Level1Out250[21] , \Level4Out188[11] , \Level16Out176[17] , 
        \Level1Out180[16] , \Level1Out225[11] , \Level1Out245[15] , 
        \ScanLink16[1] , \Level1Out195[22] , \Level1Out230[25] , 
        \Level1Out29[28] , \ScanLink93[27] , \Level1Out115[4] , 
        \Level1Out213[14] , \ScanLink248[6] , \Level2Out44[3] , 
        \Level1Out2[1] , \Level1Out6[17] , \ScanLink71[6] , \ScanLink86[13] , 
        \ScanLink128[10] , \ScanLink148[14] , \Level1Out138[11] , 
        \Level2Out96[5] , \Level1Out212[6] , \Level2Out102[11] , 
        \Level2Out154[10] , \Level1Out158[15] , \Level1Out172[3] , 
        \Level2Out134[14] , \Level2Out162[15] , \Level1Out195[11] , 
        \Level1Out230[16] , \Level1Out245[26] , \ScanLink72[5] , 
        \Level1Out171[0] , \Level1Out206[13] , \Level1Out211[5] , 
        \Level1Out213[27] , \Level16Out176[24] , \Level1Out180[25] , 
        \Level1Out225[22] , \ScanLink216[12] , \Level1Out250[12] , 
        \Level4Out188[22] , \ScanLink4[27] , \ScanLink4[14] , \Level1Out52[6] , 
        \ScanLink68[26] , \ScanLink151[8] , \ScanLink190[24] , 
        \Level2Out56[21] , \ScanLink235[23] , \Level1Out80[0] , 
        \ScanLink115[19] , \ScanLink136[31] , \ScanLink185[10] , 
        \ScanLink220[17] , \ScanLink240[13] , \Level2Out88[9] , 
        \ScanLink203[26] , \ScanLink255[27] , \Level2Out60[24] , 
        \Level2Out36[25] , \Level2Out202[0] , \ScanLink160[29] , 
        \Level1Out110[9] , \ScanLink136[28] , \ScanLink143[18] , 
        \ScanLink160[30] , \Level2Out90[30] , \Level2Out90[29] , 
        \Level2Out162[5] , \Level2Out26[9] , \Level1Out105[18] , 
        \Level1Out126[30] , \ScanLink130[1] , \Level8Out168[5] , 
        \Level1Out126[29] , \Level1Out170[28] , \Level16Out64[23] , 
        \Level128Out0[0] , \Level16Out32[22] , \Level1Out14[12] , 
        \Level1Out22[17] , \Level1Out57[27] , \Level1Out74[16] , 
        \Level1Out153[19] , \Level1Out170[31] , \ScanLink250[4] , 
        \Level4Out236[3] , \Level8Out208[0] , \ScanLink133[2] , 
        \Level4Out4[3] , \Level1Out37[23] , \Level1Out42[13] , 
        \Level1Out51[5] , \ScanLink253[7] , \Level4Out156[6] , 
        \Level1Out61[22] , \Level2Out192[18] , \Level4Out80[30] , 
        \Level1Out83[3] , \Level2Out38[5] , \Level4Out80[29] , 
        \Level8Out176[9] , \ScanLink154[5] , \Level1Out209[7] , 
        \Level2Out48[19] , \Level4Out184[0] , \Level16Out64[10] , 
        \Level8Out80[6] , \Level1Out9[19] , \Level1Out10[10] , 
        \ScanLink12[18] , \Level1Out14[21] , \ScanLink16[30] , 
        \ScanLink35[18] , \Level1Out36[2] , \Level16Out32[11] , 
        \ScanLink77[8] , \ScanLink98[18] , \Level1Out169[2] , \ScanLink234[0] , 
        \Level1Load173[0] , \ScanLink186[3] , \Level1Out214[8] , 
        \Level64Load64[0] , \Level2Out106[1] , \ScanLink185[0] , 
        \ScanLink208[19] , \ScanLink16[29] , \ScanLink40[28] , 
        \Level1Out35[1] , \Level1Out37[10] , \ScanLink40[31] , 
        \ScanLink63[19] , \Level1Out42[20] , \Level1Out22[24] , 
        \Level1Out61[11] , \ScanLink157[6] , \Level4Out252[7] , 
        \ScanLink69[4] , \Level4Out196[29] , \Level1Out74[25] , 
        \Level2Load162[0] , \Level4Out132[2] , \ScanLink31[29] , 
        \ScanLink44[19] , \Level1Out57[14] , \Level2Out222[18] , 
        \Level4Out196[30] , \Level1Out153[8] , \Level1Out218[18] , 
        \ScanLink237[3] , \Level1Load234[0] , \Level2Load194[0] , 
        \ScanLink67[31] , \ScanLink67[28] , \Level2Out78[7] , \ScanLink31[30] , 
        \Level1Out33[21] , \Level1Out46[11] , \Level4Out116[4] , 
        \ScanLink213[5] , \Level1Out65[20] , \Level2Out8[21] , 
        \Level1Out70[14] , \Level2Out226[30] , \Level4Out192[18] , 
        \Level1Out53[25] , \ScanLink173[0] , \ScanLink0[16] , \Level1Out11[7] , 
        \Level1Out26[15] , \Level2Out226[29] , \ScanLink81[8] , 
        \Level1Out12[4] , \Level1Load185[0] , \ScanLink210[6] , 
        \Level8Out248[2] , \Level1Out26[26] , \ScanLink29[6] , 
        \Level1Out70[27] , \ScanLink170[3] , \Level64Out128[20] , 
        \Level2Out122[7] , \Level8Out128[7] , \Level2Out242[2] , 
        \Level4Out108[8] , \Level4Out172[0] , \ScanLink0[25] , 
        \Level1Out10[23] , \Level1Out33[12] , \Level1Out53[16] , 
        \Level2Out196[29] , \Level1Out46[22] , \Level1Out75[3] , 
        \Level2Out196[30] , \Level4Out84[18] , \Level4Out212[5] , 
        \ScanLink34[9] , \Level1Load57[0] , \Level1Out65[13] , 
        \ScanLink117[4] , \Level2Out8[12] , \Level1Out101[29] , 
        \ScanLink109[8] , \ScanLink111[31] , \ScanLink111[28] , 
        \ScanLink147[30] , \ScanLink164[18] , \ScanLink147[29] , 
        \Level2Out146[3] , \ScanLink132[19] , \Level1Out129[0] , 
        \Level2Out94[18] , \Level2Out226[6] , \Level64Out128[13] , 
        \Level1Out157[31] , \Level2Out194[5] , \Level1Out174[19] , 
        \Level1Out249[5] , \ScanLink114[7] , \Level1Out2[26] , 
        \Level1Out76[0] , \Level1Out101[30] , \Level1Out157[28] , 
        \Level2Out118[18] , \Level8Out8[3] , \Level1Out122[18] , 
        \Level1Out2[15] , \ScanLink9[3] , \Level1Out17[9] , \ScanLink19[27] , 
        \ScanLink56[3] , \Level1Out191[20] , \Level1Out234[27] , 
        \Level1Out241[17] , \Level16Out144[10] , \Level32Out192[0] , 
        \ScanLink84[5] , \Level1Out155[6] , \ScanLink208[4] , 
        \Level2Out188[11] , \Level16Out112[11] , \Level1Out217[16] , 
        \ScanLink168[1] , \Level1Out202[22] , \Level2Out238[22] , 
        \Level1Out235[3] , \Level1Out254[23] , \Level1Out184[14] , 
        \ScanLink212[23] , \Level1Out221[13] , \Level2Out52[10] , 
        \ScanLink244[22] , \ScanLink79[23] , \Level1Out148[9] , 
        \Level1Out187[0] , \Level4Out56[8] , \ScanLink194[15] , 
        \ScanLink231[12] , \ScanLink251[16] , \Level2Out64[15] , 
        \ScanLink181[21] , \ScanLink224[26] , \ScanLink207[17] , 
        \Level2Out32[14] , \ScanLink19[14] , \ScanLink55[0] , \ScanLink82[22] , 
        \ScanLink87[6] , \ScanLink97[16] , \ScanLink139[15] , 
        \Level1Out184[3] , \ScanLink216[8] , \ScanLink159[11] , 
        \Level2Out60[5] , \Level1Out149[10] , \Level2Out106[20] , 
        \Level4Out48[4] , \Level1Out156[5] , \Level2Out124[9] , 
        \Level2Out150[21] , \ScanLink79[10] , \Level1Out129[14] , 
        \Level1Out236[0] , \Level2Out130[25] , \Level2Out166[24] , 
        \ScanLink181[12] , \ScanLink224[15] , \ScanLink194[26] , 
        \ScanLink207[24] , \ScanLink251[25] , \Level2Out64[26] , 
        \ScanLink212[10] , \Level2Out32[27] , \Level2Out52[23] , 
        \ScanLink231[21] , \ScanLink244[11] , \ScanLink32[7] , 
        \Level1Out131[2] , \Level1Out202[11] , \Level1Out184[27] , 
        \Level2Out238[11] , \Level1Out221[20] , \Level1Out58[30] , 
        \Level1Out254[10] , \Level1Out191[13] , \Level1Out234[14] , 
        \Level16Out144[23] , \Level1Out2[8] , \Level1Out4[6] , \Level1Out7[5] , 
        \ScanLink31[4] , \Level1Out58[29] , \Level1Out241[24] , 
        \Level1Out251[7] , \Level1Out217[25] , \Level2Out188[22] , 
        \Level16Out112[22] , \Level1Out80[19] , \Level1Out129[27] , 
        \Level2Out130[16] , \Level1Out132[1] , \Level2Out166[17] , 
        \Level1Out149[23] , \Level2Out220[8] , \Level2Out106[13] , 
        \Level2Out150[12] , \ScanLink82[11] , \ScanLink159[22] , 
        \Level1Out252[4] , \ScanLink97[25] , \Level1Out110[16] , 
        \ScanLink112[9] , \ScanLink139[26] , \Level1Out133[27] , 
        \Level1Out146[17] , \ScanLink234[9] , \Level1Out165[26] , 
        \Level1Out14[31] , \ScanLink16[20] , \ScanLink35[11] , \ScanLink77[1] , 
        \ScanLink98[11] , \Level1Out105[22] , \Level1Out170[12] , 
        \Level16Out64[19] , \Level1Out126[13] , \Level1Out153[23] , 
        \Level2Out42[4] , \Level16Out32[18] , \ScanLink160[13] , 
        \ScanLink115[23] , \ScanLink136[12] , \ScanLink143[22] , 
        \Level1Out174[4] , \ScanLink229[6] , \Level2Out106[8] , 
        \ScanLink100[17] , \ScanLink123[26] , \ScanLink149[3] , 
        \ScanLink156[16] , \Level1Out214[1] , \Level4Out4[25] , 
        \ScanLink175[27] , \Level2Out90[2] , \Level2Out90[13] , 
        \ScanLink40[21] , \ScanLink74[2] , \Level2Out28[27] , \ScanLink20[25] , 
        \Level1Out28[7] , \ScanLink63[10] , \Level1Out177[7] , 
        \ScanLink76[24] , \Level1Out37[19] , \ScanLink55[15] , 
        \Level2Out48[23] , \Level16Out96[6] , \Level8Out112[4] , 
        \ScanLink185[9] , \ScanLink208[10] , \Level1Out217[2] , 
        \Level1Out218[11] , \Level2Out118[4] , \Level4Out196[20] , 
        \Level2Out222[11] , \Level2Out192[22] , \Level1Out35[8] , 
        \Level1Out42[29] , \Level2Out242[15] , \Level2Out214[14] , 
        \Level4Out80[13] , \ScanLink10[6] , \ScanLink13[5] , \Level1Out14[28] , 
        \Level1Out42[30] , \Level1Out61[18] , \ScanLink198[6] , 
        \ScanLink123[15] , \Level4Out4[16] , \ScanLink20[16] , 
        \ScanLink55[26] , \ScanLink76[17] , \Level1Out80[9] , \ScanLink98[22] , 
        \ScanLink100[24] , \ScanLink156[25] , \Level4Out148[3] , 
        \Level1Out110[0] , \Level2Out90[20] , \ScanLink115[10] , 
        \ScanLink175[14] , \ScanLink160[20] , \Level2Out202[9] , 
        \Level1Out105[11] , \ScanLink136[21] , \ScanLink143[11] , 
        \Level4Out228[6] , \Level2Out6[2] , \Level1Out110[25] , 
        \Level1Out126[20] , \Level1Out170[21] , \Level128Out0[9] , 
        \Level1Out133[14] , \Level1Out153[10] , \Level8Out208[9] , 
        \Level1Out146[24] , \Level2Out26[0] , \ScanLink130[8] , 
        \Level1Out165[15] , \Level1Out218[22] , \Level2Out192[11] , 
        \Level2Out242[26] , \Level16Out192[7] , \Level2Out214[27] , 
        \Level4Out80[20] , \Level4Out196[13] , \Level2Out222[22] , 
        \Level4Out184[9] , \Level1Out113[3] , \Level8Out216[5] , 
        \ScanLink208[23] , \Level2Out48[10] , \ScanLink16[13] , 
        \ScanLink35[22] , \ScanLink40[12] , \Level2Out28[14] , 
        \ScanLink63[23] , \Level8Out176[0] , \Level1Out29[12] , 
        \Level1Out30[5] , \ScanLink128[19] , \ScanLink232[7] , 
        \Level1Out49[16] , \Level1Out84[12] , \Level1Out91[26] , 
        \ScanLink152[2] , \Level8Out24[23] , \Level8Out72[22] , 
        \Level2Out100[6] , \Level1Out138[18] , \Level2Out102[18] , 
        \Level2Out154[19] , \ScanLink180[4] , \Level1Out171[9] , 
        \ScanLink183[7] , \Level1Out195[18] , \Level8Out184[17] , 
        \ScanLink185[19] , \Level4Out72[7] , \ScanLink231[4] , 
        \Level4Load244[0] , \Level1Out9[23] , \Level1Out14[3] , 
        \ScanLink16[8] , \Level1Out33[6] , \ScanLink151[1] , \Level2Out56[28] , 
        \Level2Out56[31] , \Level2Out88[0] , \Level1Out54[1] , 
        \Level1Out84[21] , \ScanLink86[30] , \Level1Out86[7] , 
        \Level1Out91[15] , \Level2Out164[2] , \Level2Out204[7] , 
        \ScanLink256[3] , \Level8Out72[11] , \Level8Out24[10] , 
        \ScanLink86[29] , \ScanLink136[6] , \Level8Load128[0] , 
        \Level1Out57[2] , \Level1Out108[2] , \ScanLink216[31] , 
        \ScanLink216[28] , \ScanLink240[30] , \ScanLink235[19] , 
        \ScanLink240[29] , \ScanLink255[0] , \Level4Out16[3] , 
        \Level32Out64[0] , \ScanLink135[5] , \Level1Out17[0] , 
        \Level1Out29[21] , \Level1Out38[24] , \Level1Out49[25] , 
        \Level1Out85[4] , \Level1Load112[0] , \Level8Out184[24] , 
        \Level1Out250[31] , \Level1Out58[20] , \Level1Out73[4] , 
        \ScanLink111[3] , \Level1Out206[30] , \Level1Out206[29] , 
        \Level1Out225[18] , \Level1Out250[28] , \Level4Out188[18] , 
        \ScanLink212[19] , \ScanLink231[31] , \ScanLink231[28] , 
        \ScanLink244[18] , \ScanLink79[19] , \Level2Load244[0] , 
        \Level4Out32[5] , \Level1Out202[18] , \Level1Out221[30] , 
        \Level2Out238[18] , \Level1Out38[17] , \Level1Out70[7] , 
        \Level1Out80[10] , \Level1Out221[29] , \Level1Out254[19] , 
        \Level2Out220[1] , \Level32Out32[16] , \Level32Out64[17] , 
        \Level128Out0[25] , \Level1Out95[24] , \Level1Load255[0] , 
        \Level2Out140[4] , \Level1Out132[8] , \Level16Out48[15] , 
        \ScanLink82[18] , \ScanLink112[0] , \Level2Out192[2] , 
        \Level8Out16[24] , \Level8Out40[25] , \Level1Out58[13] , 
        \ScanLink99[3] , \ScanLink168[8] , \Level16Out144[19] , 
        \Level1Out191[29] , \Level2Out188[18] , \Level4Out84[7] , 
        \Level32Out192[9] , \Level16Out112[18] , \Level1Out191[30] , 
        \Level1Out148[0] , \ScanLink175[7] , \ScanLink181[28] , 
        \Level1Out228[5] , \ScanLink181[31] , \Level1Out187[9] , 
        \ScanLink215[2] , \Level2Out52[19] , \Level4Out56[1] , 
        \ScanLink159[18] , \Level8Out40[16] , \ScanLink176[4] , 
        \Level1Load36[0] , \ScanLink48[6] , \ScanLink216[1] , 
        \Level8Out16[17] , \Level1Out80[23] , \Level1Out95[17] , 
        \Level1Out149[19] , \Level1Out236[9] , \Level2Out244[5] , 
        \Level16Out48[26] , \Level1Out199[5] , \Level2Out106[29] , 
        \Level32Out64[24] , \Level2Out150[31] , \Level2Out106[30] , 
        \ScanLink55[9] , \Level2Out124[0] , \Level32Out32[25] , 
        \Level1Out209[27] , \Level2Out150[28] , \Level2Out196[20] , 
        \Level2Out238[3] , \Level128Out0[16] , \Level2Out246[17] , 
        \Level2Out210[16] , \Level4Out84[11] , \Level2Out158[6] , 
        \Level4Out192[22] , \Level2Out226[13] , \Level4Out172[9] , 
        \Level1Out9[10] , \ScanLink12[22] , \ScanLink24[27] , \Level1Out68[5] , 
        \ScanLink72[26] , \ScanLink31[13] , \ScanLink51[17] , 
        \Level8Out152[6] , \Level1Load98[0] , \ScanLink34[0] , 
        \ScanLink44[23] , \ScanLink219[26] , \ScanLink12[11] , 
        \ScanLink31[20] , \ScanLink37[3] , \ScanLink67[12] , \Level1Out137[5] , 
        \Level8Out232[3] , \ScanLink89[27] , \ScanLink109[1] , 
        \ScanLink127[24] , \ScanLink152[14] , \Level1Out254[3] , 
        \Level4Out0[27] , \ScanLink104[15] , \ScanLink171[25] , 
        \Level2Out94[11] , \ScanLink111[21] , \ScanLink164[11] , 
        \ScanLink132[10] , \Level1Out134[6] , \ScanLink147[20] , 
        \ScanLink44[10] , \Level1Out76[9] , \Level1Out101[20] , 
        \Level1Out174[10] , \Level1Out157[21] , \Level2Out118[11] , 
        \Level1Out114[14] , \Level1Out122[11] , \Level1Out129[9] , 
        \Level1Out137[25] , \Level1Out142[15] , \Level2Out178[15] , 
        \Level1Out161[24] , \ScanLink219[15] , \Level1Out233[4] , 
        \ScanLink67[21] , \Level8Out136[2] , \ScanLink24[14] , 
        \ScanLink51[24] , \ScanLink72[15] , \Level1Out153[1] , \ScanLink50[4] , 
        \Level1Out10[19] , \Level1Out33[28] , \Level1Out46[18] , 
        \ScanLink173[9] , \Level4Out192[11] , \Level2Out226[20] , 
        \Level1Out65[30] , \Level1Out209[14] , \Level2Out246[24] , 
        \Level1Out181[7] , \Level2Out8[31] , \Level2Out196[13] , 
        \Level1Out65[29] , \ScanLink82[2] , \Level1Out19[6] , 
        \Level1Out33[31] , \Level2Out8[28] , \Level4Out84[22] , 
        \ScanLink53[7] , \ScanLink81[1] , \Level1Out101[13] , 
        \Level1Out114[27] , \Level1Out137[16] , \Level2Out210[25] , 
        \Level1Out142[26] , \Level2Out66[2] , \Level2Out178[26] , 
        \Level64Out128[29] , \Level1Out161[17] , \Level64Out128[30] , 
        \ScanLink111[12] , \Level1Out122[22] , \Level1Out174[23] , 
        \Level1Out157[12] , \Level1Out182[4] , \Level2Out118[22] , 
        \ScanLink127[17] , \ScanLink132[23] , \ScanLink164[22] , 
        \ScanLink147[13] , \Level1Out230[7] , \Level4Out0[14] , 
        \ScanLink89[14] , \ScanLink104[26] , \ScanLink152[27] , 
        \Level2Out94[22] , \Level4Out108[1] , \Level1Out150[2] , 
        \ScanLink171[16] , \Level2Out112[17] , \Level4Out120[10] , 
        \ScanLink45[3] , \Level1Out81[29] , \Level1Out128[17] , 
        \Level1Out226[3] , \Level4Out56[27] , \Level4Out176[11] , 
        \Level32Out0[24] , \Level2Out144[16] , \Level2Out124[12] , 
        \Level4Out116[15] , \Level1Out81[30] , \Level4Out60[22] , 
        \Level1Out148[13] , \Level4Out36[23] , \ScanLink0[12] , 
        \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , \Level1Out3[25] , 
        \ScanLink18[24] , \ScanLink78[20] , \ScanLink83[21] , 
        \Level1Out146[6] , \Level2Out172[13] , \Level4Out140[14] , 
        \ScanLink96[15] , \ScanLink97[5] , \ScanLink138[16] , 
        \ScanLink158[12] , \Level2Out70[6] , \Level1Out194[0] , 
        \ScanLink206[14] , \Level2Out46[27] , \Level2Load86[0] , 
        \ScanLink250[15] , \ScanLink180[22] , \Level2Out10[26] , 
        \ScanLink225[25] , \ScanLink245[21] , \Level2Out70[22] , 
        \Level4Out100[9] , \Level1Out59[19] , \ScanLink94[6] , 
        \ScanLink195[16] , \Level1Out197[3] , \ScanLink205[8] , 
        \ScanLink230[11] , \ScanLink213[20] , \Level2Out26[23] , 
        \ScanLink178[2] , \Level1Out225[0] , \Level1Out255[20] , 
        \Level4Out228[17] , \Level1Out185[17] , \Level1Out220[10] , 
        \Level1Out203[21] , \Level8Out120[6] , \ScanLink218[7] , 
        \Level1Out145[5] , \Level1Out216[15] , \Level8Out240[3] , 
        \Level1Out3[16] , \ScanLink21[7] , \ScanLink46[0] , \ScanLink89[9] , 
        \Level1Out190[23] , \Level1Out240[14] , \Level1Out235[24] , 
        \Level4Out248[13] , \ScanLink83[12] , \ScanLink96[26] , 
        \ScanLink138[25] , \Level1Load138[0] , \Level2Out14[2] , 
        \Level1Out122[2] , \Level1Out128[24] , \Level1Out148[20] , 
        \ScanLink158[21] , \Level2Out182[8] , \Level1Out242[7] , 
        \Level2Out124[21] , \Level4Out60[11] , \Level2Out172[20] , 
        \Level4Out116[26] , \Level4Out140[27] , \Level4Out36[10] , 
        \Level2Out112[24] , \Level4Out56[14] , \Level4Out120[23] , 
        \Level2Out144[25] , \Level4Out176[22] , \Level32Out0[17] , 
        \Level1Out190[10] , \Level1Out216[26] , \Level8Out0[2] , 
        \Level8Out224[18] , \Level1Out235[17] , \Level4Out248[20] , 
        \ScanLink18[17] , \ScanLink22[4] , \Level1Out185[24] , 
        \Level1Out220[23] , \Level1Out240[27] , \Level8Out144[2] , 
        \Level1Out241[4] , \Level1Out121[1] , \Level1Out203[12] , 
        \Level1Out255[13] , \Level4Out228[24] , \ScanLink195[25] , 
        \ScanLink230[22] , \Level8Out224[7] , \ScanLink245[12] , 
        \Level2Out70[11] , \ScanLink78[13] , \ScanLink101[9] , 
        \ScanLink213[13] , \Level2Out26[10] , \Level4Out204[8] , 
        \ScanLink206[27] , \Level2Out46[14] , \ScanLink110[18] , 
        \ScanLink133[30] , \ScanLink133[29] , \ScanLink180[11] , 
        \Level2Out10[15] , \ScanLink225[16] , \ScanLink250[26] , 
        \ScanLink146[19] , \ScanLink165[31] , \ScanLink165[28] , 
        \Level2Out252[1] , \Level1Out123[28] , \Level1Out140[8] , 
        \ScanLink160[0] , \Level1Load227[0] , \Level2Out132[4] , 
        \Level2Out76[8] , \Level8Out152[23] , \Level8Out104[22] , 
        \ScanLink1[2] , \Level1Out11[13] , \Level1Out27[16] , 
        \Level1Out52[26] , \Level1Out100[19] , \Level1Out123[31] , 
        \Level1Out156[18] , \Level1Out175[30] , \ScanLink200[5] , 
        \Level4Out28[28] , \Level1Out175[29] , \Level4Out28[31] , 
        \Level1Load196[0] , \Level2Load236[0] , \Level1Out64[23] , 
        \Level1Out71[17] , \ScanLink163[3] , \ScanLink92[8] , 
        \Level1Out32[22] , \Level1Out47[12] , \Level4Out40[5] , 
        \ScanLink203[6] , \Level32Out32[6] , \Level2Out38[31] , 
        \Level2Out38[28] , \Level2Out68[4] , \Level4Out200[19] , 
        \Level4Out92[3] , \Level1Out2[22] , \ScanLink5[24] , \ScanLink5[17] , 
        \Level1Out8[30] , \Level1Out11[20] , \ScanLink13[31] , 
        \ScanLink13[28] , \ScanLink27[9] , \Level1Load44[0] , \Level1Out66[3] , 
        \ScanLink104[4] , \Level1Out139[3] , \Level2Out184[6] , 
        \Level4Out168[30] , \Level4Out168[29] , \Level8Out152[10] , 
        \Level8Out104[11] , \Level1Out244[9] , \Level2Out236[5] , 
        \Level2Out156[0] , \ScanLink30[19] , \ScanLink45[30] , 
        \ScanLink66[18] , \ScanLink45[29] , \Level1Out27[25] , 
        \Level1Out32[11] , \Level1Out64[10] , \ScanLink107[7] , 
        \Level2Out228[9] , \Level1Out47[21] , \Level1Out65[0] , 
        \Level2Out204[31] , \Level4Out24[1] , \Level1Out8[29] , 
        \Level1Out52[15] , \Level2Load28[0] , \Level2Out252[29] , 
        \Level2Out204[28] , \Level1Out15[11] , \ScanLink17[19] , 
        \ScanLink39[5] , \Level1Out71[24] , \Level2Out252[30] , 
        \ScanLink62[29] , \Level1Out103[9] , \ScanLink209[30] , 
        \ScanLink209[29] , \Level8Out96[11] , \Level2Out28[6] , 
        \Level1Out93[0] , \ScanLink34[31] , \ScanLink34[28] , \ScanLink41[18] , 
        \ScanLink62[30] , \Level1Out60[21] , \Level4Load236[0] , 
        \Level1Out23[14] , \Level1Out36[20] , \Level1Out43[10] , 
        \ScanLink243[4] , \Level1Out56[24] , \Level1Out219[28] , 
        \Level1Out41[6] , \Level1Out75[15] , \Level1Out219[31] , 
        \ScanLink123[1] , \Level2Out8[4] , \Level2Out200[19] , 
        \Level8Out208[27] , \Level1Out9[3] , \Level1Out15[22] , 
        \Level1Out23[27] , \Level1Out42[5] , \ScanLink120[2] , 
        \ScanLink240[7] , \Level8Out160[24] , \Level8Out136[25] , 
        \Level1Out90[3] , \ScanLink99[31] , \Level2Out172[6] , 
        \Level2Out212[3] , \ScanLink99[28] , \Level1Out56[17] , 
        \Level4Out64[3] , \Level1Out75[26] , \ScanLink79[7] , \ScanLink227[0] , 
        \Level8Out208[14] , \Level1Out25[2] , \Level1Out36[13] , 
        \Level1Out60[12] , \ScanLink147[5] , \Level4Out204[31] , 
        \Level4Out252[29] , \Level4Out204[28] , \Level1Out43[23] , 
        \ScanLink64[8] , \Level4Out252[30] , \ScanLink114[30] , 
        \ScanLink142[28] , \Level1Load160[0] , \ScanLink195[3] , 
        \Level1Out207[8] , \Level2Out116[2] , \Level8Out96[22] , 
        \ScanLink114[29] , \ScanLink137[18] , \ScanLink142[31] , 
        \ScanLink161[19] , \ScanLink159[9] , \ScanLink196[0] , 
        \Level2Out80[8] , \Level1Out179[1] , \ScanLink224[3] , 
        \Level8Out160[17] , \Level1Out7[27] , \Level1Out26[1] , 
        \Level1Out104[31] , \Level1Out152[29] , \Level2Out168[29] , 
        \Level1Out104[28] , \Level1Out127[19] , \Level1Out152[30] , 
        \Level1Out171[18] , \Level32Out192[18] , \Level1Out219[4] , 
        \Level8Out136[16] , \Level1Out105[7] , \ScanLink144[6] , 
        \Level2Out168[30] , \Level1Out212[17] , \Level2Out228[17] , 
        \Level8Out200[1] , \Level1Out244[16] , \Level1Out7[14] , 
        \Level1Out28[18] , \Level1Out47[8] , \ScanLink69[16] , 
        \ScanLink138[0] , \Level1Out194[21] , \Level1Out231[26] , 
        \Level1Out251[22] , \Level1Out181[15] , \Level1Out224[12] , 
        \ScanLink191[14] , \Level1Out207[23] , \Level2Out198[24] , 
        \Level8Out160[4] , \ScanLink234[13] , \ScanLink241[23] , 
        \Level2Out74[20] , \Level2Out248[13] , \Level1Out88[1] , 
        \Level1Out118[8] , \ScanLink202[16] , \ScanLink217[22] , 
        \Level2Out22[21] , \Level2Out42[25] , \ScanLink254[17] , 
        \ScanLink184[20] , \ScanLink221[27] , \Level2Out14[24] , 
        \Level1Out59[4] , \ScanLink87[23] , \ScanLink92[17] , 
        \ScanLink149[24] , \ScanLink246[9] , \Level1Out106[4] , 
        \ScanLink129[20] , \Level2Out30[4] , \Level1Out139[21] , 
        \Level2Out120[10] , \Level4Out112[17] , \Level2Out174[8] , 
        \Level4Out32[21] , \Level4Out64[20] , \Level4Out144[16] , 
        \Level1Out159[25] , \Level2Out176[11] , \Level2Out116[15] , 
        \Level4Out124[12] , \ScanLink62[6] , \ScanLink69[25] , 
        \ScanLink184[13] , \ScanLink202[25] , \Level2Out140[14] , 
        \Level4Out52[25] , \Level4Out172[13] , \Level2Out42[16] , 
        \ScanLink191[27] , \ScanLink221[14] , \ScanLink234[20] , 
        \ScanLink254[24] , \Level2Out14[17] , \Level8Out88[29] , 
        \Level1Out181[26] , \ScanLink217[11] , \ScanLink241[10] , 
        \Level2Out74[13] , \Level2Load2[0] , \Level2Out22[12] , 
        \Level1Out224[21] , \Level8Out88[30] , \Level1Out161[3] , 
        \Level1Out207[10] , \Level1Out251[11] , \Level2Out248[20] , 
        \Level1Out212[24] , \Level2Out198[17] , \Level2Out228[24] , 
        \Level1Out194[12] , \Level16Out80[2] , \Level1Out231[15] , 
        \Level1Out244[25] , \Level16Out80[19] , \Level8Out104[0] , 
        \ScanLink9[7] , \ScanLink55[4] , \ScanLink61[5] , \Level1Out159[16] , 
        \Level1Out162[0] , \Level1Out201[6] , \Level8Out88[7] , 
        \Level2Load70[0] , \Level4Out52[16] , \Level2Out116[26] , 
        \Level2Out140[27] , \Level4Out124[21] , \Level4Out172[20] , 
        \Level1Out85[18] , \Level1Out202[5] , \Level2Out120[23] , 
        \Level4Out64[13] , \Level4Out112[24] , \ScanLink87[10] , 
        \Level1Out139[12] , \Level2Out86[6] , \Level2Out176[22] , 
        \Level4Out32[12] , \Level4Out144[25] , \ScanLink92[24] , 
        \ScanLink129[13] , \ScanLink142[8] , \ScanLink149[17] , 
        \Level2Out54[0] , \Level1Out129[10] , \Level2Out166[20] , 
        \Level2Out244[8] , \Level1Out236[4] , \Level2Out130[21] , 
        \Level2Out150[25] , \Level32Out64[30] , \ScanLink82[26] , 
        \Level1Out149[14] , \Level2Out106[24] , \Level4Out48[0] , 
        \Level32Out32[28] , \Level32Out64[29] , \Level1Out156[1] , 
        \Level1Out199[8] , \Level32Out32[31] , \ScanLink87[2] , 
        \ScanLink139[11] , \ScanLink159[15] , \Level2Out60[1] , 
        \ScanLink176[9] , \ScanLink19[23] , \ScanLink79[27] , \ScanLink97[12] , 
        \Level1Out184[7] , \ScanLink207[13] , \Level1Out228[8] , 
        \Level2Out32[10] , \ScanLink251[12] , \Level2Out64[11] , 
        \ScanLink181[25] , \ScanLink224[22] , \ScanLink244[26] , 
        \ScanLink84[1] , \Level1Out187[4] , \ScanLink194[11] , 
        \ScanLink212[27] , \ScanLink231[16] , \Level2Out52[14] , 
        \Level1Out155[2] , \ScanLink168[5] , \Level1Out235[7] , 
        \Level1Out254[27] , \Level1Out184[10] , \Level1Out202[26] , 
        \Level1Out221[17] , \Level2Out238[26] , \ScanLink208[0] , 
        \Level2Out188[15] , \Level16Out112[15] , \Level1Out217[12] , 
        \Level1Out241[13] , \Level1Out2[11] , \ScanLink31[0] , \ScanLink56[7] , 
        \Level1Out191[24] , \Level1Out234[23] , \Level32Out192[4] , 
        \Level16Out144[14] , \ScanLink82[15] , \ScanLink97[21] , 
        \ScanLink139[22] , \Level8Out16[29] , \Level8Out40[31] , 
        \Level1Out95[30] , \Level1Out129[23] , \Level1Out149[27] , 
        \ScanLink159[26] , \Level8Out16[30] , \Level8Out40[28] , 
        \Level1Out252[0] , \Level2Out150[16] , \Level128Out0[28] , 
        \Level128Out0[31] , \Level2Out106[17] , \Level2Out166[13] , 
        \Level16Out48[18] , \Level1Out132[5] , \Level2Out140[9] , 
        \Level1Out95[29] , \Level1Out191[17] , \Level1Out217[21] , 
        \Level2Out130[12] , \Level1Out234[10] , \Level2Out188[26] , 
        \Level16Out112[26] , \Level16Out144[27] , \Level1Out241[20] , 
        \Level1Out12[0] , \ScanLink19[10] , \ScanLink32[3] , 
        \Level1Out184[23] , \Level1Out251[3] , \Level1Out221[24] , 
        \Level1Out38[30] , \Level1Out38[29] , \Level1Out131[6] , 
        \Level1Out202[15] , \Level1Out254[14] , \Level1Out73[9] , 
        \ScanLink194[22] , \Level2Out238[15] , \ScanLink231[25] , 
        \ScanLink244[15] , \ScanLink79[14] , \ScanLink207[20] , 
        \ScanLink212[14] , \Level2Out32[23] , \Level2Out52[27] , 
        \ScanLink89[19] , \ScanLink181[16] , \ScanLink224[11] , 
        \Level4Out32[8] , \ScanLink251[21] , \Level2Out64[22] , 
        \Level2Out242[6] , \ScanLink170[7] , \Level2Out122[3] , 
        \Level4Out0[19] , \Level4Load68[0] , \Level8Out128[3] , 
        \Level64Out128[24] , \Level1Out53[21] , \Level1Out182[9] , 
        \ScanLink210[2] , \Level8Out248[6] , \ScanLink0[21] , 
        \Level1Out10[14] , \Level1Out11[3] , \Level1Out26[11] , 
        \Level1Out65[24] , \Level1Out70[10] , \ScanLink173[4] , 
        \Level2Out8[25] , \Level2Out246[30] , \Level2Out210[28] , 
        \ScanLink24[19] , \Level1Load33[0] , \Level1Out33[25] , 
        \Level1Out46[15] , \Level2Out246[29] , \Level1Out209[19] , 
        \ScanLink213[1] , \Level4Out116[0] , \Level2Out210[31] , 
        \ScanLink219[18] , \Level2Out78[3] , \Level1Out233[9] , 
        \ScanLink51[29] , \ScanLink50[9] , \ScanLink51[30] , \ScanLink72[18] , 
        \Level1Out10[27] , \Level1Out68[8] , \Level1Out76[4] , \Level8Out8[7] , 
        \ScanLink104[18] , \ScanLink114[3] , \Level1Out249[1] , 
        \Level1Out114[19] , \Level1Out137[31] , \Level1Out161[29] , 
        \Level2Out194[1] , \ScanLink127[30] , \Level1Out129[4] , 
        \Level1Out137[28] , \Level1Out142[18] , \Level1Out161[30] , 
        \Level64Out128[17] , \Level2Out178[18] , \ScanLink171[28] , 
        \Level2Out226[2] , \ScanLink127[29] , \ScanLink152[19] , 
        \ScanLink171[31] , \Level2Out146[7] , \Level1Out137[8] , 
        \Level1Load250[0] , \Level1Out26[22] , \Level1Out33[16] , 
        \Level1Out65[17] , \ScanLink117[0] , \Level2Out8[16] , 
        \Level4Out212[1] , \Level1Out46[26] , \Level1Out75[7] , 
        \Level4Out172[4] , \Level1Out1[6] , \Level1Out2[5] , \ScanLink4[23] , 
        \ScanLink4[10] , \Level1Out14[16] , \ScanLink29[2] , \Level1Out53[12] , 
        \Level1Out61[26] , \Level1Out70[23] , \Level1Out83[7] , 
        \Level2Out38[1] , \Level4Out184[4] , \Level8Out216[8] , 
        \Level2Out28[19] , \Level2Load106[0] , \Level1Out22[13] , 
        \Level1Out37[27] , \Level1Out42[17] , \Level4Out156[2] , 
        \ScanLink253[3] , \Level1Out57[23] , \Level4Out4[7] , \Level1Out51[1] , 
        \Level1Out74[12] , \ScanLink133[6] , \Level4Out236[7] , 
        \Level16Out32[26] , \ScanLink13[8] , \Level1Out52[2] , 
        \Level1Out110[31] , \Level1Out110[28] , \ScanLink250[0] , 
        \Level8Out208[4] , \Level16Out64[27] , \Level128Out0[4] , 
        \ScanLink130[5] , \Level1Out146[30] , \Level1Out165[18] , 
        \Level8Out168[1] , \Level1Out133[19] , \ScanLink100[30] , 
        \ScanLink100[29] , \Level1Out146[29] , \ScanLink156[31] , 
        \ScanLink175[19] , \ScanLink123[18] , \Level2Out162[1] , 
        \Level1Out14[25] , \Level1Out22[20] , \Level1Out80[4] , 
        \Level1Load117[0] , \ScanLink156[28] , \Level2Out202[4] , 
        \Level1Out57[10] , \Level4Out132[6] , \ScanLink69[0] , 
        \Level1Out74[21] , \ScanLink237[7] , \Level2Out118[9] , 
        \Level4Out252[3] , \ScanLink20[31] , \ScanLink20[28] , 
        \Level1Out35[5] , \Level1Out37[14] , \Level1Out61[15] , 
        \ScanLink157[2] , \Level2Out214[19] , \Level1Out42[24] , 
        \Level2Out242[18] , \ScanLink55[18] , \ScanLink76[30] , 
        \Level8Out112[9] , \ScanLink185[4] , \ScanLink76[29] , 
        \Level1Out169[6] , \Level1Out174[9] , \Level2Out106[5] , 
        \ScanLink186[7] , \Level4Out4[31] , \Level4Out4[28] , \ScanLink234[4] , 
        \Level1Out6[20] , \Level1Out7[8] , \Level1Out36[6] , \Level2Out42[9] , 
        \Level16Out32[15] , \Level1Out115[0] , \ScanLink154[1] , 
        \Level1Out209[3] , \Level16Out64[14] , \Level1Out213[10] , 
        \ScanLink248[2] , \Level8Out80[2] , \Level8Out184[29] , 
        \ScanLink15[6] , \ScanLink16[5] , \Level1Out195[26] , 
        \Level1Out230[21] , \Level1Out245[11] , \Level8Out184[30] , 
        \Level1Out49[31] , \Level1Out250[25] , \Level4Out188[15] , 
        \Level1Out49[28] , \Level1Out85[9] , \ScanLink128[7] , 
        \Level1Out180[12] , \Level1Out225[15] , \ScanLink68[11] , 
        \ScanLink190[13] , \Level1Out206[24] , \ScanLink240[24] , 
        \Level16Out176[13] , \ScanLink235[14] , \ScanLink86[24] , 
        \ScanLink93[10] , \Level1Out98[6] , \ScanLink135[8] , 
        \ScanLink203[11] , \ScanLink216[25] , \Level2Out56[16] , 
        \Level2Out36[12] , \ScanLink255[10] , \Level2Out60[13] , 
        \ScanLink148[23] , \ScanLink185[27] , \ScanLink220[20] , 
        \ScanLink128[27] , \Level2Out20[3] , \Level2Out154[27] , 
        \Level1Out49[3] , \Level1Out116[3] , \Level2Out102[26] , 
        \Level1Out138[26] , \Level1Out158[22] , \ScanLink68[22] , 
        \Level1Out91[18] , \Level2Out134[23] , \Level2Out162[22] , 
        \ScanLink185[14] , \ScanLink203[22] , \Level2Out0[1] , 
        \ScanLink220[13] , \Level2Out36[21] , \ScanLink190[20] , 
        \ScanLink231[9] , \ScanLink255[23] , \Level2Out60[20] , 
        \ScanLink235[27] , \ScanLink216[16] , \ScanLink240[17] , 
        \Level1Out6[13] , \ScanLink72[1] , \Level1Out180[21] , 
        \Level2Out56[25] , \Level1Out225[26] , \Level1Out171[4] , 
        \Level1Out206[17] , \Level1Out250[16] , \Level4Out188[26] , 
        \Level16Out176[20] , \Level8Load232[0] , \Level1Out195[15] , 
        \Level1Out213[23] , \Level1Out230[12] , \ScanLink71[2] , 
        \Level1Out158[11] , \Level1Out211[1] , \Level1Out245[22] , 
        \Level2Out162[11] , \Level1Out172[7] , \ScanLink86[17] , 
        \Level1Out138[15] , \ScanLink180[9] , \Level2Out134[10] , 
        \Level2Out154[14] , \Level1Out212[2] , \Level2Out96[1] , 
        \Level2Out102[15] , \ScanLink128[14] , \Level1Load208[0] , 
        \Level1Out3[31] , \Level1Out3[28] , \ScanLink5[30] , \Level1Load19[0] , 
        \Level1Out30[8] , \ScanLink148[10] , \Level2Out44[7] , 
        \ScanLink93[23] , \Level1Out132[20] , \Level1Out147[10] , 
        \Level2Out108[20] , \Level16Out192[20] , \Level1Out111[11] , 
        \Level1Out164[21] , \ScanLink5[29] , \Level1Out104[25] , 
        \Level1Out171[15] , \Level1Out219[9] , \Level32Out192[15] , 
        \Level1Out7[19] , \ScanLink17[27] , \ScanLink34[16] , \ScanLink67[6] , 
        \ScanLink99[16] , \Level1Out127[14] , \Level1Out152[24] , 
        \Level2Out52[3] , \ScanLink161[14] , \Level2Out168[24] , 
        \ScanLink114[24] , \ScanLink239[1] , \Level2Out84[20] , 
        \ScanLink137[15] , \ScanLink142[25] , \Level1Out164[3] , 
        \ScanLink101[10] , \ScanLink122[21] , \ScanLink157[11] , 
        \Level1Out204[6] , \ScanLink159[4] , \ScanLink174[20] , 
        \Level2Out80[5] , \ScanLink41[26] , \ScanLink64[5] , \ScanLink17[14] , 
        \ScanLink21[22] , \Level1Out38[0] , \ScanLink62[17] , 
        \Level1Out167[0] , \ScanLink77[23] , \ScanLink21[11] , 
        \Level1Out23[19] , \Level1Out42[8] , \ScanLink54[12] , 
        \ScanLink99[25] , \Level1Out100[7] , \ScanLink101[23] , 
        \ScanLink122[12] , \ScanLink147[8] , \Level1Out207[5] , 
        \ScanLink209[17] , \Level1Out219[16] , \Level2Out108[3] , 
        \Level2Out200[27] , \Level4Out232[20] , \Level2Out186[11] , 
        \Level8Out208[19] , \Level2Out236[22] , \Level4Out204[25] , 
        \ScanLink188[1] , \Level4Out252[24] , \ScanLink157[22] , 
        \ScanLink114[17] , \ScanLink174[13] , \Level2Out84[13] , 
        \ScanLink161[27] , \Level1Out104[16] , \ScanLink137[26] , 
        \ScanLink142[16] , \Level8Out136[28] , \Level1Out127[27] , 
        \Level1Out171[26] , \Level8Out160[30] , \Level2Out168[17] , 
        \Level8Out136[31] , \Level32Out192[26] , \Level1Out132[13] , 
        \Level1Out152[17] , \Level8Out160[29] , \Level1Out147[23] , 
        \Level2Out36[7] , \Level2Out108[13] , \Level16Out192[13] , 
        \Level1Out56[30] , \Level1Out75[18] , \Level1Out111[22] , 
        \Level1Out164[12] , \ScanLink243[9] , \Level2Out236[11] , 
        \Level4Out204[16] , \Level4Out252[17] , \Level1Out56[29] , 
        \Level2Out8[9] , \Level2Out200[14] , \Level4Out232[13] , 
        \Level1Out219[25] , \ScanLink54[21] , \ScanLink77[10] , 
        \Level2Out186[22] , \Level1Out103[4] , \Level8Load240[0] , 
        \ScanLink209[24] , \ScanLink34[25] , \ScanLink41[15] , 
        \ScanLink62[24] , \Level1Out20[2] , \ScanLink92[29] , \ScanLink222[0] , 
        \Level1Out48[11] , \ScanLink61[8] , \ScanLink92[30] , \ScanLink142[5] , 
        \Level2Out110[1] , \Level8Out96[6] , \Level1Out85[15] , 
        \Level1Out90[21] , \Level1Load165[0] , \Level4Out144[28] , 
        \Level4Out112[30] , \Level4Out112[29] , \Level4Out144[31] , 
        \Level8Out128[10] , \ScanLink190[3] , \Level1Out202[8] , 
        \Level1Out212[30] , \Level1Out231[18] , \Level2Out6[21] , 
        \Level8Out216[12] , \Level8Out240[13] , \Level1Out244[28] , 
        \Level16Out80[14] , \ScanLink18[3] , \Level1Out23[1] , 
        \Level1Out28[15] , \ScanLink193[0] , \Level2Out228[30] , 
        \Level1Out212[29] , \ScanLink69[31] , \ScanLink202[31] , 
        \ScanLink221[19] , \Level1Out244[31] , \Level2Out228[29] , 
        \Level4Out124[2] , \ScanLink202[28] , \ScanLink221[3] , 
        \ScanLink254[29] , \ScanLink254[30] , \Level2Load174[0] , 
        \Level4Out244[7] , \ScanLink69[28] , \ScanLink141[6] , 
        \Level128Out128[12] , \Level2Out98[7] , \Level8Out88[24] , 
        \Level1Out59[9] , \Level1Out85[26] , \Level1Out106[9] , 
        \Level1Out90[12] , \Level2Out174[5] , \Level8Out128[23] , 
        \Level1Out159[31] , \Level1Out159[28] , \Level2Out116[18] , 
        \Level2Out140[19] , \Level4Out52[31] , \Level2Out214[0] , 
        \Level1Out96[0] , \Level4Out52[28] , \ScanLink149[30] , 
        \ScanLink149[29] , \ScanLink246[4] , \ScanLink22[9] , 
        \Level1Out28[26] , \Level1Out44[6] , \ScanLink126[1] , 
        \Level2Out30[9] , \Level1Out47[5] , \Level1Out118[5] , 
        \ScanLink191[19] , \Level4Out140[6] , \Level128Out128[21] , 
        \ScanLink245[7] , \Level2Out42[31] , \Level8Out88[17] , 
        \ScanLink125[2] , \Level2Out14[29] , \Level2Out42[28] , 
        \Level4Out220[3] , \Level2Out14[30] , \Level16Out80[27] , 
        \Level1Out39[23] , \Level1Out48[22] , \Level1Out95[3] , 
        \Level2Out198[29] , \Level4Out192[0] , \Level8Out240[20] , 
        \Level1Out59[27] , \Level1Out63[3] , \ScanLink101[4] , 
        \Level1Out181[18] , \Level2Out6[12] , \Level2Out198[30] , 
        \Level8Out160[9] , \Level8Out216[21] , \ScanLink195[31] , 
        \Level4Out204[5] , \ScanLink195[28] , \Level1Out241[9] , 
        \Level2Out10[18] , \Level4Out164[0] , \Level2Out46[19] , 
        \Level1Out185[30] , \Level8Out224[15] , \Level4Out228[30] , 
        \Level1Load41[0] , \Level1Out185[29] , \Level1Out39[10] , 
        \Level1Out60[0] , \Level1Out81[17] , \Level2Out2[23] , 
        \Level4Out228[29] , \Level2Out230[6] , \Level1Out94[23] , 
        \Level1Out128[30] , \Level2Out144[28] , \Level2Out150[3] , 
        \Level2Out112[30] , \Level1Out128[29] , \Level2Out144[31] , 
        \Level4Out56[19] , \ScanLink138[31] , \Level2Out112[29] , 
        \ScanLink102[7] , \ScanLink138[28] , \Level2Out182[5] , 
        \Level1Load222[0] , \Level2Out2[10] , \ScanLink89[4] , 
        \Level1Out240[19] , \Level2Load182[0] , \Level1Out235[29] , 
        \ScanLink4[2] , \ScanLink7[1] , \Level64Out128[6] , \ScanLink18[30] , 
        \Level1Out59[14] , \Level1Out145[8] , \Level1Out216[18] , 
        \Level1Out235[30] , \Level8Out224[26] , \ScanLink165[0] , 
        \ScanLink206[19] , \ScanLink225[28] , \ScanLink250[18] , 
        \Level1Out238[2] , \ScanLink225[31] , \ScanLink18[29] , 
        \ScanLink58[1] , \ScanLink96[18] , \Level1Out158[7] , \ScanLink205[5] , 
        \Level4Out100[4] , \ScanLink166[3] , \Level1Load193[0] , 
        \ScanLink206[6] , \Level1Out94[10] , \ScanLink97[8] , 
        \Level32Out0[29] , \Level2Out254[2] , \Level32Out0[30] , 
        \ScanLink0[31] , \ScanLink0[28] , \ScanLink1[22] , \ScanLink1[18] , 
        \Level1Out8[24] , \Level1Out81[24] , \Level1Out189[2] , 
        \Level4Out140[19] , \Level1Out208[20] , \Level2Out134[7] , 
        \Level4Out116[18] , \Level2Out228[4] , \Level2Out232[20] , 
        \Level4Out200[27] , \Level4Out236[22] , \Level1Out8[17] , 
        \ScanLink13[25] , \ScanLink24[7] , \ScanLink25[20] , \Level1Out27[31] , 
        \Level1Out27[28] , \ScanLink39[8] , \Level1Out71[29] , 
        \Level2Out148[1] , \Level2Out204[25] , \Level2Out182[13] , 
        \Level1Out52[18] , \Level1Out71[30] , \Level2Out252[24] , 
        \ScanLink73[21] , \Level1Out78[2] , \Level8Out8[11] , \ScanLink30[14] , 
        \ScanLink50[10] , \Level1Out247[7] , \Level2Out38[16] , 
        \Level2Out58[12] , \ScanLink45[24] , \ScanLink218[21] , 
        \ScanLink13[16] , \ScanLink27[4] , \ScanLink66[15] , \Level1Out127[2] , 
        \ScanLink88[20] , \ScanLink119[6] , \ScanLink153[13] , 
        \Level1Out244[4] , \ScanLink126[23] , \ScanLink105[12] , 
        \ScanLink170[22] , \Level2Out236[8] , \ScanLink110[26] , 
        \ScanLink165[16] , \Level1Out124[1] , \Level2Out80[22] , 
        \ScanLink133[17] , \ScanLink146[27] , \ScanLink30[27] , 
        \ScanLink45[17] , \Level1Out100[27] , \ScanLink104[9] , 
        \Level1Out175[17] , \Level4Out108[20] , \Level1Out115[13] , 
        \Level1Out123[16] , \Level1Out156[26] , \Level2Out12[1] , 
        \Level4Out28[16] , \Level1Out136[22] , \Level1Out143[12] , 
        \Level1Out160[23] , \Level4Out48[12] , \Level4Out168[24] , 
        \ScanLink218[12] , \Level1Out223[3] , \Level2Out58[21] , 
        \ScanLink66[26] , \Level16Out0[7] , \Level2Out68[9] , \ScanLink25[13] , 
        \ScanLink50[23] , \ScanLink73[12] , \Level1Out143[6] , 
        \Level8Out8[22] , \Level2Out38[25] , \ScanLink40[3] , 
        \Level2Out204[16] , \Level4Out236[11] , \ScanLink91[6] , 
        \ScanLink92[5] , \Level1Out191[0] , \Level1Out208[13] , 
        \Level2Out182[20] , \Level2Out252[17] , \Level4Out40[8] , 
        \Level2Out232[13] , \Level4Out200[14] , \Level1Out100[14] , 
        \Level1Out115[20] , \Level1Out136[11] , \Level1Out143[21] , 
        \Level2Out76[5] , \Level4Out48[21] , \Level4Out168[17] , 
        \Level1Out160[10] , \Level4Out108[13] , \Level1Out123[25] , 
        \Level1Out175[24] , \ScanLink1[11] , \ScanLink1[6] , \ScanLink5[20] , 
        \ScanLink5[13] , \Level1Out7[23] , \ScanLink43[0] , \ScanLink110[15] , 
        \Level1Out156[15] , \Level1Out192[3] , \ScanLink200[8] , 
        \Level4Out28[25] , \ScanLink126[10] , \ScanLink133[24] , 
        \ScanLink165[25] , \Level2Out80[11] , \ScanLink146[14] , 
        \Level1Out220[0] , \Level2Out132[9] , \Level1Out59[0] , 
        \ScanLink88[13] , \ScanLink105[21] , \ScanLink153[20] , 
        \Level1Out140[5] , \Level1Out159[21] , \ScanLink170[11] , 
        \Level2Out140[10] , \Level4Out172[17] , \Level2Out214[9] , 
        \Level2Out116[11] , \Level4Out124[16] , \ScanLink69[12] , 
        \Level1Load78[0] , \ScanLink87[27] , \Level1Out96[9] , 
        \Level1Out106[0] , \Level4Out32[25] , \Level4Out52[21] , 
        \ScanLink126[8] , \Level1Out139[25] , \Level2Load14[0] , 
        \Level4Out144[12] , \Level2Out120[14] , \Level2Out176[15] , 
        \Level4Out112[13] , \Level4Out64[24] , \ScanLink129[24] , 
        \Level2Out30[0] , \Level1Out88[5] , \ScanLink92[13] , 
        \ScanLink149[20] , \ScanLink254[13] , \ScanLink184[24] , 
        \Level2Out14[20] , \ScanLink202[12] , \ScanLink221[23] , 
        \Level2Out42[21] , \ScanLink191[10] , \ScanLink217[26] , 
        \Level128Out128[28] , \ScanLink234[17] , \ScanLink241[27] , 
        \Level2Out22[25] , \Level2Out74[24] , \Level128Out128[31] , 
        \ScanLink138[4] , \Level1Out207[27] , \Level2Out198[20] , 
        \Level8Out240[29] , \Level8Out216[31] , \Level1Out251[26] , 
        \Level2Out248[17] , \Level8Out240[30] , \Level8Out216[28] , 
        \Level1Out181[11] , \Level1Out224[16] , \Level8Out160[0] , 
        \Level1Out7[10] , \ScanLink61[1] , \ScanLink87[14] , \ScanLink92[20] , 
        \Level1Out105[3] , \Level1Out194[25] , \Level1Out244[12] , 
        \Level1Out212[13] , \Level1Out231[22] , \Level2Out228[13] , 
        \Level4Out192[9] , \Level8Out200[5] , \Level2Out54[4] , 
        \ScanLink129[17] , \ScanLink149[13] , \Level1Out90[28] , 
        \Level1Out139[16] , \ScanLink222[9] , \Level2Out86[2] , 
        \Level2Out176[26] , \Level1Out202[1] , \Level2Out120[27] , 
        \Level4Out32[16] , \Level4Out144[21] , \Level4Out64[17] , 
        \Level8Out128[19] , \Level2Out110[8] , \Level4Out112[20] , 
        \Level2Out140[23] , \Level4Out172[24] , \Level1Out90[31] , 
        \Level2Out116[22] , \Level4Out52[12] , \Level1Out159[12] , 
        \Level1Out162[4] , \Level4Out124[25] , \Level1Out194[16] , 
        \Level1Out231[11] , \Level16Out80[6] , \Level1Out23[8] , 
        \Level1Out48[18] , \ScanLink193[9] , \Level1Out244[21] , 
        \Level8Out88[3] , \Level8Out104[4] , \Level1Out201[2] , 
        \Level1Out212[20] , \Level2Out228[20] , \Level2Out248[24] , 
        \ScanLink62[2] , \Level1Out161[7] , \Level1Out207[14] , 
        \Level1Out181[22] , \Level1Out224[25] , \Level2Out6[31] , 
        \Level2Out198[13] , \ScanLink69[21] , \ScanLink191[23] , 
        \ScanLink217[15] , \Level1Out251[15] , \Level2Out6[28] , 
        \ScanLink234[24] , \Level2Out22[16] , \Level1Out42[1] , 
        \Level1Out90[7] , \ScanLink184[17] , \ScanLink241[14] , 
        \Level2Out14[13] , \Level2Out74[17] , \ScanLink202[21] , 
        \ScanLink221[10] , \ScanLink254[20] , \Level2Out42[12] , 
        \Level2Out212[7] , \Level2Out172[2] , \ScanLink120[6] , 
        \Level8Out136[21] , \Level1Out15[15] , \Level1Out23[10] , 
        \Level1Out56[20] , \Level1Out75[11] , \ScanLink240[3] , 
        \Level8Out160[20] , \ScanLink123[5] , \Level8Out208[23] , 
        \Level2Out8[0] , \Level1Out36[24] , \Level1Out41[2] , 
        \Level1Out43[14] , \ScanLink243[0] , \Level1Out60[25] , 
        \Level2Out236[18] , \ScanLink21[18] , \ScanLink54[31] , 
        \ScanLink77[19] , \Level1Out93[4] , \Level1Load104[0] , 
        \Level2Out28[2] , \ScanLink54[28] , \Level8Out96[15] , 
        \ScanLink144[2] , \Level1Out219[0] , \Level8Out136[12] , 
        \Level8Out160[13] , \Level1Out9[7] , \Level1Out26[5] , 
        \Level1Out38[9] , \ScanLink101[19] , \Level1Out111[18] , 
        \Level1Out132[30] , \Level1Out132[29] , \Level1Out147[19] , 
        \Level1Out164[31] , \Level2Out108[29] , \Level16Out192[29] , 
        \Level1Out164[28] , \Level1Out179[5] , \ScanLink224[7] , 
        \Level2Out108[30] , \Level16Out192[30] , \ScanLink122[31] , 
        \ScanLink122[28] , \ScanLink157[18] , \ScanLink174[30] , 
        \ScanLink196[4] , \ScanLink174[29] , \ScanLink239[8] , 
        \Level2Out84[29] , \Level2Out84[30] , \Level2Out116[6] , 
        \Level8Out96[26] , \Level1Out15[26] , \Level1Out25[6] , 
        \Level1Out36[17] , \Level1Out167[9] , \ScanLink195[7] , 
        \Level1Out43[27] , \Level1Out23[23] , \Level1Out60[16] , 
        \ScanLink147[1] , \ScanLink188[8] , \Level1Out75[22] , 
        \Level4Out232[29] , \ScanLink79[3] , \Level4Load252[0] , 
        \Level8Out208[10] , \Level1Out56[13] , \Level2Out186[18] , 
        \Level4Out64[7] , \Level4Out232[30] , \ScanLink227[4] , 
        \Level4Out92[7] , \Level1Out11[17] , \Level1Out32[26] , 
        \Level1Out47[16] , \Level2Out58[31] , \Level2Out58[28] , 
        \Level2Out68[0] , \Level4Out40[1] , \Level1Out191[9] , 
        \ScanLink203[2] , \Level32Out32[2] , \Level1Out64[27] , 
        \Level1Out27[12] , \Level1Out52[22] , \Level1Out71[13] , 
        \ScanLink163[7] , \Level2Out182[30] , \Level4Out236[18] , 
        \Level2Out182[29] , \ScanLink2[5] , \Level1Load20[0] , 
        \ScanLink105[31] , \Level1Out115[30] , \ScanLink200[1] , 
        \Level1Out115[29] , \Level1Out136[18] , \Level4Out48[28] , 
        \Level1Out143[28] , \Level8Out104[26] , \Level1Out143[31] , 
        \Level4Out48[31] , \ScanLink160[4] , \Level1Out160[19] , 
        \Level8Out152[27] , \ScanLink43[9] , \ScanLink126[19] , 
        \Level2Out132[0] , \ScanLink153[29] , \Level1Out11[24] , 
        \Level1Out27[21] , \ScanLink39[1] , \ScanLink105[28] , 
        \ScanLink153[30] , \ScanLink170[18] , \Level1Out220[9] , 
        \Level2Out80[18] , \Level2Out252[5] , \Level2Out148[8] , 
        \Level1Out71[20] , \Level1Out32[15] , \Level1Out52[11] , 
        \Level4Out24[5] , \Level2Out232[29] , \Level1Out47[25] , 
        \Level1Out65[4] , \Level1Out208[29] , \Level2Out232[30] , 
        \Level2Load252[0] , \ScanLink25[30] , \Level1Out64[14] , 
        \ScanLink107[3] , \Level1Out208[30] , \ScanLink218[31] , 
        \ScanLink218[28] , \ScanLink25[29] , \ScanLink73[28] , 
        \Level8Out8[18] , \ScanLink50[19] , \ScanLink73[31] , \ScanLink88[30] , 
        \Level1Out124[8] , \Level1Load243[0] , \Level2Out156[4] , 
        \ScanLink88[29] , \ScanLink104[0] , \Level1Out139[7] , 
        \Level2Out236[1] , \Level8Out104[15] , \Level2Out184[2] , 
        \Level8Out152[14] , \Level4Out108[29] , \Level1Out3[21] , 
        \Level1Out66[7] , \Level2Out12[8] , \Level4Out108[30] , 
        \Level1Out240[10] , \Level1Out3[12] , \ScanLink7[8] , \ScanLink46[4] , 
        \Level1Out190[27] , \Level1Out235[20] , \Level4Out248[17] , 
        \ScanLink18[20] , \Level1Out39[19] , \Level1Out145[1] , 
        \Level1Out216[11] , \ScanLink218[3] , \Level8Out240[7] , 
        \ScanLink94[2] , \ScanLink178[6] , \Level1Out203[25] , 
        \Level1Out225[4] , \Level1Out255[24] , \Level2Out2[19] , 
        \Level4Out228[13] , \Level1Out185[13] , \Level1Out220[14] , 
        \Level8Out120[2] , \ScanLink213[24] , \Level2Out26[27] , 
        \ScanLink245[25] , \Level2Out70[26] , \ScanLink18[13] , 
        \Level1Out19[2] , \ScanLink45[7] , \ScanLink58[8] , \ScanLink78[24] , 
        \ScanLink195[12] , \Level1Out197[7] , \ScanLink230[15] , 
        \ScanLink250[11] , \ScanLink96[11] , \ScanLink165[9] , 
        \ScanLink180[26] , \ScanLink225[21] , \Level2Out10[22] , 
        \Level2Out46[23] , \ScanLink206[10] , \Level1Out194[4] , 
        \ScanLink83[25] , \ScanLink97[1] , \ScanLink138[12] , 
        \ScanLink158[16] , \Level2Out70[2] , \Level1Out146[2] , 
        \Level1Out148[17] , \Level4Out36[27] , \Level4Out140[10] , 
        \Level2Out124[16] , \Level2Out172[17] , \Level4Out116[11] , 
        \Level1Out94[19] , \Level4Out60[26] , \Level32Out0[20] , 
        \Level1Out226[7] , \Level2Out112[13] , \Level2Out144[12] , 
        \Level4Out176[15] , \Level4Out120[14] , \ScanLink78[17] , 
        \Level1Out128[13] , \Level4Out56[23] , \ScanLink180[15] , 
        \Level4Out164[9] , \ScanLink195[21] , \ScanLink206[23] , 
        \ScanLink225[12] , \ScanLink250[22] , \Level2Out10[11] , 
        \ScanLink213[17] , \Level2Out26[14] , \Level2Out46[10] , 
        \ScanLink230[26] , \ScanLink245[16] , \Level2Out70[15] , 
        \ScanLink22[0] , \Level1Out121[5] , \Level1Out203[16] , 
        \Level1Out185[20] , \Level1Out220[27] , \Level8Out224[3] , 
        \Level1Out190[14] , \Level1Out255[17] , \Level4Out228[20] , 
        \Level1Out235[13] , \Level1Out240[23] , \Level4Out248[24] , 
        \Level8Out144[6] , \ScanLink21[3] , \Level1Out216[22] , 
        \Level1Out241[0] , \Level2Out144[21] , \Level8Out0[6] , 
        \Level4Out176[26] , \Level32Out0[13] , \Level1Out60[9] , 
        \ScanLink83[16] , \Level1Out122[6] , \Level1Out128[20] , 
        \Level2Out112[20] , \Level4Out56[10] , \Level1Out148[24] , 
        \Level2Out172[24] , \Level4Out120[27] , \Level4Out140[23] , 
        \ScanLink158[25] , \Level1Out242[3] , \Level2Out124[25] , 
        \Level4Out36[14] , \Level4Out60[15] , \Level4Out116[22] , 
        \Level2Out14[6] , \ScanLink96[22] , \Level1Out114[10] , 
        \ScanLink138[21] , \Level1Out161[20] , \Level2Out194[8] , 
        \Level1Out137[21] , \Level1Out142[11] , \Level2Out178[11] , 
        \Level1Out122[15] , \Level1Out157[25] , \Level2Out118[15] , 
        \Level1Out2[18] , \Level1Out9[27] , \ScanLink12[26] , \ScanLink37[7] , 
        \Level1Out101[24] , \Level1Out174[14] , \Level1Out249[8] , 
        \ScanLink132[14] , \ScanLink147[24] , \ScanLink89[23] , 
        \ScanLink111[25] , \ScanLink164[15] , \Level1Out134[2] , 
        \ScanLink104[11] , \ScanLink171[21] , \ScanLink109[5] , 
        \ScanLink152[10] , \Level2Out94[15] , \Level1Out254[7] , 
        \Level4Out0[23] , \ScanLink127[20] , \ScanLink24[23] , 
        \ScanLink31[17] , \ScanLink67[16] , \Level1Out137[1] , 
        \Level8Out232[7] , \ScanLink34[4] , \ScanLink44[27] , 
        \ScanLink219[22] , \ScanLink51[13] , \Level8Out152[2] , 
        \Level1Out68[1] , \ScanLink72[22] , \Level2Out226[17] , 
        \Level4Out192[26] , \Level1Out9[14] , \Level1Out12[9] , 
        \ScanLink53[3] , \ScanLink89[10] , \ScanLink104[22] , \ScanLink117[9] , 
        \Level2Out158[2] , \Level2Out210[12] , \Level4Out84[15] , 
        \Level4Out212[8] , \Level1Out209[23] , \Level2Out196[24] , 
        \Level2Out238[7] , \Level2Out246[13] , \Level4Out108[5] , 
        \Level1Out150[6] , \Level2Out94[26] , \ScanLink127[13] , 
        \ScanLink171[12] , \Level4Out0[10] , \ScanLink81[5] , 
        \Level1Out101[17] , \ScanLink111[16] , \ScanLink132[27] , 
        \ScanLink152[23] , \ScanLink147[17] , \Level1Out230[3] , 
        \Level1Out122[26] , \ScanLink164[26] , \Level1Out157[16] , 
        \Level1Out182[0] , \Level2Load90[0] , \Level2Out118[26] , 
        \Level1Out114[23] , \Level1Out174[27] , \Level1Out137[12] , 
        \Level1Out161[13] , \Level2Out66[6] , \Level2Out178[22] , 
        \Level1Out26[18] , \Level1Out53[28] , \ScanLink82[6] , 
        \Level1Out142[22] , \Level1Out181[3] , \Level1Out209[10] , 
        \Level2Out210[21] , \Level4Out84[26] , \Level2Out246[20] , 
        \Level4Out116[9] , \ScanLink213[8] , \Level2Out196[17] , 
        \Level1Out53[31] , \Level1Out70[19] , \Level2Out226[24] , 
        \Level4Out192[15] , \ScanLink12[15] , \ScanLink24[10] , 
        \ScanLink51[20] , \ScanLink50[0] , \ScanLink67[25] , \ScanLink72[11] , 
        \Level1Out153[5] , \ScanLink31[24] , \ScanLink44[14] , 
        \ScanLink219[11] , \Level1Out233[0] , \ScanLink31[9] , 
        \Level1Load52[0] , \Level1Out70[3] , \ScanLink97[31] , 
        \Level2Out192[6] , \Level8Out16[20] , \Level8Out136[6] , 
        \Level8Out40[21] , \ScanLink97[28] , \ScanLink112[4] , 
        \Level2Out140[0] , \Level16Out48[11] , \Level1Out95[20] , 
        \Level1Out38[20] , \Level1Out80[14] , \Level1Out252[9] , 
        \Level32Out32[12] , \Level128Out0[21] , \Level2Out220[5] , 
        \Level32Out64[13] , \Level1Out58[24] , \Level1Out217[31] , 
        \Level1Out217[28] , \Level1Out234[19] , \Level1Out241[30] , 
        \ScanLink4[19] , \Level1Out4[2] , \Level1Out6[30] , \Level1Out14[7] , 
        \ScanLink19[19] , \Level1Out73[0] , \ScanLink207[30] , 
        \ScanLink207[29] , \Level1Out241[29] , \ScanLink224[18] , 
        \ScanLink251[31] , \Level4Out32[1] , \ScanLink251[28] , 
        \ScanLink48[2] , \Level1Out80[27] , \ScanLink111[7] , 
        \Level1Out95[13] , \Level1Out129[19] , \Level1Out156[8] , 
        \Level1Load231[0] , \Level2Out124[4] , \Level4Out48[9] , 
        \Level32Out32[21] , \Level32Out64[20] , \Level128Out0[12] , 
        \Level1Out199[1] , \Level2Out130[31] , \Level2Out244[1] , 
        \Level16Out48[22] , \Level2Out166[29] , \ScanLink139[18] , 
        \Level2Out130[28] , \Level2Out166[30] , \ScanLink216[5] , 
        \Level2Out60[8] , \Level8Out16[13] , \Level1Out17[4] , \ScanLink84[8] , 
        \Level1Out148[4] , \ScanLink176[0] , \Level8Out40[12] , 
        \ScanLink194[18] , \ScanLink215[6] , \Level4Out56[5] , 
        \ScanLink175[3] , \Level1Out228[1] , \Level2Out32[19] , 
        \Level1Load180[0] , \Level2Out64[18] , \Level2Load220[0] , 
        \Level1Out29[16] , \Level1Out33[2] , \Level1Out38[13] , 
        \Level1Out58[17] , \Level4Out84[3] , \ScanLink99[7] , \ScanLink208[9] , 
        \Level1Out184[19] , \ScanLink190[29] , \Level2Out88[4] , 
        \ScanLink151[5] , \ScanLink190[30] , \Level1Load176[0] , 
        \ScanLink231[0] , \Level2Out36[31] , \Level2Out36[28] , 
        \Level2Out60[30] , \Level4Out72[3] , \Level2Out60[29] , 
        \Level8Out184[13] , \Level1Out30[1] , \Level1Out49[12] , 
        \ScanLink72[8] , \Level1Out180[28] , \ScanLink183[3] , 
        \Level1Out211[8] , \Level16Out176[30] , \Level1Out84[16] , 
        \Level1Out180[31] , \Level16Out176[29] , \Level1Out91[22] , 
        \Level1Out158[18] , \ScanLink180[0] , \Level2Out96[8] , 
        \Level2Out162[18] , \Level2Out100[2] , \Level2Out134[19] , 
        \ScanLink148[19] , \Level8Out24[27] , \ScanLink152[6] , 
        \Level8Out72[26] , \Level1Out49[21] , \Level1Out85[0] , 
        \ScanLink232[3] , \Level1Out6[29] , \Level1Out29[25] , 
        \Level1Out115[9] , \Level1Out213[19] , \Level1Out230[31] , 
        \Level8Out184[20] , \Level1Out245[18] , \Level1Out54[5] , 
        \Level1Out57[6] , \ScanLink135[1] , \Level1Out230[28] , 
        \ScanLink203[18] , \ScanLink220[30] , \ScanLink255[19] , 
        \ScanLink68[18] , \Level1Out108[6] , \ScanLink220[29] , 
        \ScanLink255[4] , \Level4Out16[7] , \Level32Out64[4] , 
        \Level4Load220[0] , \Level1Out84[25] , \Level1Out86[3] , 
        \ScanLink93[19] , \ScanLink136[2] , \Level8Out24[14] , 
        \Level8Out72[15] , \ScanLink256[7] , \Level2Out204[3] , 
        \Level1Out91[11] , \Level2Out0[8] , \Level2Out164[6] , 
        \Level2Out214[10] , \Level1Out7[1] , \ScanLink16[24] , 
        \ScanLink20[21] , \Level1Out22[30] , \Level1Out22[29] , 
        \ScanLink198[2] , \Level4Out80[17] , \Level2Out192[26] , 
        \Level2Out222[15] , \Level2Out242[11] , \Level1Out57[19] , 
        \Level1Out74[31] , \Level1Out218[15] , \Level4Out196[24] , 
        \ScanLink69[9] , \Level2Out118[0] , \Level1Out74[28] , 
        \Level1Out28[3] , \ScanLink55[11] , \Level2Out48[27] , 
        \Level16Out96[2] , \Level8Out112[0] , \ScanLink76[20] , 
        \ScanLink208[14] , \Level1Out217[6] , \ScanLink35[15] , 
        \ScanLink63[14] , \Level1Out177[3] , \ScanLink40[25] , \ScanLink74[6] , 
        \Level2Out28[23] , \ScanLink77[5] , \ScanLink100[13] , 
        \ScanLink175[23] , \Level2Out90[6] , \Level2Out90[17] , 
        \ScanLink123[22] , \ScanLink156[12] , \Level1Out214[5] , 
        \Level4Out4[21] , \ScanLink136[16] , \ScanLink143[26] , 
        \ScanLink149[7] , \ScanLink98[15] , \ScanLink160[17] , 
        \ScanLink115[27] , \ScanLink229[2] , \Level1Out126[17] , 
        \Level1Out153[27] , \Level1Out174[0] , \Level2Load66[0] , 
        \Level2Out42[0] , \ScanLink10[2] , \ScanLink16[17] , \ScanLink63[27] , 
        \Level1Out105[26] , \ScanLink154[8] , \Level1Out170[16] , 
        \Level1Out110[12] , \Level1Out165[22] , \Level1Out133[23] , 
        \Level1Out146[13] , \Level2Out38[8] , \ScanLink20[12] , 
        \ScanLink35[26] , \ScanLink40[16] , \Level2Out28[10] , 
        \ScanLink55[22] , \Level8Out176[4] , \ScanLink208[27] , 
        \Level2Out48[14] , \Level1Out51[8] , \ScanLink76[13] , 
        \Level1Out113[7] , \Level8Out216[1] , \Level1Out218[26] , 
        \Level2Out222[26] , \Level1Out110[21] , \Level2Out192[15] , 
        \Level2Out214[23] , \Level4Out80[24] , \Level4Out196[17] , 
        \Level2Out242[22] , \Level16Out192[3] , \Level1Out126[24] , 
        \Level1Out133[10] , \Level1Out165[11] , \Level8Out168[8] , 
        \Level1Out146[20] , \Level2Out26[4] , \ScanLink98[26] , 
        \Level1Out105[15] , \Level1Out153[14] , \ScanLink250[9] , 
        \ScanLink115[14] , \ScanLink136[25] , \Level1Out170[25] , 
        \ScanLink143[15] , \Level2Out6[6] , \Level4Out228[2] , 
        \ScanLink160[24] , \ScanLink100[20] , \Level2Out90[24] , 
        \Level4Out148[7] , \Level1Out110[4] , \ScanLink123[11] , 
        \ScanLink175[10] , \Level4Out4[12] , \Level2Out162[8] , 
        \ScanLink13[1] , \ScanLink156[21] ;
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanOut({\ScanLink2[31] , 
        \ScanLink2[30] , \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , 
        \ScanLink2[26] , \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , 
        \ScanLink2[22] , \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , 
        \ScanLink2[18] , \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , 
        \ScanLink2[14] , \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , 
        \ScanLink2[10] , \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , 
        \ScanLink2[6] , \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , 
        \ScanLink2[2] , \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load1[0] ), .Out({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_21 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanOut({\ScanLink22[31] , 
        \ScanLink22[30] , \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , 
        \ScanLink22[26] , \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , 
        \ScanLink22[22] , \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , 
        \ScanLink22[18] , \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , 
        \ScanLink22[14] , \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , 
        \ScanLink22[10] , \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , 
        \ScanLink22[6] , \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , 
        \ScanLink22[2] , \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load21[0] ), .Out({
        \Level1Out21[31] , \Level1Out21[30] , \Level1Out21[29] , 
        \Level1Out21[28] , \Level1Out21[27] , \Level1Out21[26] , 
        \Level1Out21[25] , \Level1Out21[24] , \Level1Out21[23] , 
        \Level1Out21[22] , \Level1Out21[21] , \Level1Out21[20] , 
        \Level1Out21[19] , \Level1Out21[18] , \Level1Out21[17] , 
        \Level1Out21[16] , \Level1Out21[15] , \Level1Out21[14] , 
        \Level1Out21[13] , \Level1Out21[12] , \Level1Out21[11] , 
        \Level1Out21[10] , \Level1Out21[9] , \Level1Out21[8] , 
        \Level1Out21[7] , \Level1Out21[6] , \Level1Out21[5] , \Level1Out21[4] , 
        \Level1Out21[3] , \Level1Out21[2] , \Level1Out21[1] , \Level1Out21[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_103 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink103[31] , \ScanLink103[30] , 
        \ScanLink103[29] , \ScanLink103[28] , \ScanLink103[27] , 
        \ScanLink103[26] , \ScanLink103[25] , \ScanLink103[24] , 
        \ScanLink103[23] , \ScanLink103[22] , \ScanLink103[21] , 
        \ScanLink103[20] , \ScanLink103[19] , \ScanLink103[18] , 
        \ScanLink103[17] , \ScanLink103[16] , \ScanLink103[15] , 
        \ScanLink103[14] , \ScanLink103[13] , \ScanLink103[12] , 
        \ScanLink103[11] , \ScanLink103[10] , \ScanLink103[9] , 
        \ScanLink103[8] , \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , 
        \ScanLink103[4] , \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , 
        \ScanLink103[0] }), .ScanOut({\ScanLink104[31] , \ScanLink104[30] , 
        \ScanLink104[29] , \ScanLink104[28] , \ScanLink104[27] , 
        \ScanLink104[26] , \ScanLink104[25] , \ScanLink104[24] , 
        \ScanLink104[23] , \ScanLink104[22] , \ScanLink104[21] , 
        \ScanLink104[20] , \ScanLink104[19] , \ScanLink104[18] , 
        \ScanLink104[17] , \ScanLink104[16] , \ScanLink104[15] , 
        \ScanLink104[14] , \ScanLink104[13] , \ScanLink104[12] , 
        \ScanLink104[11] , \ScanLink104[10] , \ScanLink104[9] , 
        \ScanLink104[8] , \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , 
        \ScanLink104[4] , \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , 
        \ScanLink104[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load103[0] ), .Out({\Level1Out103[31] , \Level1Out103[30] , 
        \Level1Out103[29] , \Level1Out103[28] , \Level1Out103[27] , 
        \Level1Out103[26] , \Level1Out103[25] , \Level1Out103[24] , 
        \Level1Out103[23] , \Level1Out103[22] , \Level1Out103[21] , 
        \Level1Out103[20] , \Level1Out103[19] , \Level1Out103[18] , 
        \Level1Out103[17] , \Level1Out103[16] , \Level1Out103[15] , 
        \Level1Out103[14] , \Level1Out103[13] , \Level1Out103[12] , 
        \Level1Out103[11] , \Level1Out103[10] , \Level1Out103[9] , 
        \Level1Out103[8] , \Level1Out103[7] , \Level1Out103[6] , 
        \Level1Out103[5] , \Level1Out103[4] , \Level1Out103[3] , 
        \Level1Out103[2] , \Level1Out103[1] , \Level1Out103[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_124 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink124[31] , \ScanLink124[30] , 
        \ScanLink124[29] , \ScanLink124[28] , \ScanLink124[27] , 
        \ScanLink124[26] , \ScanLink124[25] , \ScanLink124[24] , 
        \ScanLink124[23] , \ScanLink124[22] , \ScanLink124[21] , 
        \ScanLink124[20] , \ScanLink124[19] , \ScanLink124[18] , 
        \ScanLink124[17] , \ScanLink124[16] , \ScanLink124[15] , 
        \ScanLink124[14] , \ScanLink124[13] , \ScanLink124[12] , 
        \ScanLink124[11] , \ScanLink124[10] , \ScanLink124[9] , 
        \ScanLink124[8] , \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , 
        \ScanLink124[4] , \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , 
        \ScanLink124[0] }), .ScanOut({\ScanLink125[31] , \ScanLink125[30] , 
        \ScanLink125[29] , \ScanLink125[28] , \ScanLink125[27] , 
        \ScanLink125[26] , \ScanLink125[25] , \ScanLink125[24] , 
        \ScanLink125[23] , \ScanLink125[22] , \ScanLink125[21] , 
        \ScanLink125[20] , \ScanLink125[19] , \ScanLink125[18] , 
        \ScanLink125[17] , \ScanLink125[16] , \ScanLink125[15] , 
        \ScanLink125[14] , \ScanLink125[13] , \ScanLink125[12] , 
        \ScanLink125[11] , \ScanLink125[10] , \ScanLink125[9] , 
        \ScanLink125[8] , \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , 
        \ScanLink125[4] , \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , 
        \ScanLink125[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load124[0] ), .Out({\Level1Out124[31] , \Level1Out124[30] , 
        \Level1Out124[29] , \Level1Out124[28] , \Level1Out124[27] , 
        \Level1Out124[26] , \Level1Out124[25] , \Level1Out124[24] , 
        \Level1Out124[23] , \Level1Out124[22] , \Level1Out124[21] , 
        \Level1Out124[20] , \Level1Out124[19] , \Level1Out124[18] , 
        \Level1Out124[17] , \Level1Out124[16] , \Level1Out124[15] , 
        \Level1Out124[14] , \Level1Out124[13] , \Level1Out124[12] , 
        \Level1Out124[11] , \Level1Out124[10] , \Level1Out124[9] , 
        \Level1Out124[8] , \Level1Out124[7] , \Level1Out124[6] , 
        \Level1Out124[5] , \Level1Out124[4] , \Level1Out124[3] , 
        \Level1Out124[2] , \Level1Out124[1] , \Level1Out124[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_214 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink214[31] , \ScanLink214[30] , 
        \ScanLink214[29] , \ScanLink214[28] , \ScanLink214[27] , 
        \ScanLink214[26] , \ScanLink214[25] , \ScanLink214[24] , 
        \ScanLink214[23] , \ScanLink214[22] , \ScanLink214[21] , 
        \ScanLink214[20] , \ScanLink214[19] , \ScanLink214[18] , 
        \ScanLink214[17] , \ScanLink214[16] , \ScanLink214[15] , 
        \ScanLink214[14] , \ScanLink214[13] , \ScanLink214[12] , 
        \ScanLink214[11] , \ScanLink214[10] , \ScanLink214[9] , 
        \ScanLink214[8] , \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , 
        \ScanLink214[4] , \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , 
        \ScanLink214[0] }), .ScanOut({\ScanLink215[31] , \ScanLink215[30] , 
        \ScanLink215[29] , \ScanLink215[28] , \ScanLink215[27] , 
        \ScanLink215[26] , \ScanLink215[25] , \ScanLink215[24] , 
        \ScanLink215[23] , \ScanLink215[22] , \ScanLink215[21] , 
        \ScanLink215[20] , \ScanLink215[19] , \ScanLink215[18] , 
        \ScanLink215[17] , \ScanLink215[16] , \ScanLink215[15] , 
        \ScanLink215[14] , \ScanLink215[13] , \ScanLink215[12] , 
        \ScanLink215[11] , \ScanLink215[10] , \ScanLink215[9] , 
        \ScanLink215[8] , \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , 
        \ScanLink215[4] , \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , 
        \ScanLink215[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load214[0] ), .Out({\Level1Out214[31] , \Level1Out214[30] , 
        \Level1Out214[29] , \Level1Out214[28] , \Level1Out214[27] , 
        \Level1Out214[26] , \Level1Out214[25] , \Level1Out214[24] , 
        \Level1Out214[23] , \Level1Out214[22] , \Level1Out214[21] , 
        \Level1Out214[20] , \Level1Out214[19] , \Level1Out214[18] , 
        \Level1Out214[17] , \Level1Out214[16] , \Level1Out214[15] , 
        \Level1Out214[14] , \Level1Out214[13] , \Level1Out214[12] , 
        \Level1Out214[11] , \Level1Out214[10] , \Level1Out214[9] , 
        \Level1Out214[8] , \Level1Out214[7] , \Level1Out214[6] , 
        \Level1Out214[5] , \Level1Out214[4] , \Level1Out214[3] , 
        \Level1Out214[2] , \Level1Out214[1] , \Level1Out214[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_233 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink233[31] , \ScanLink233[30] , 
        \ScanLink233[29] , \ScanLink233[28] , \ScanLink233[27] , 
        \ScanLink233[26] , \ScanLink233[25] , \ScanLink233[24] , 
        \ScanLink233[23] , \ScanLink233[22] , \ScanLink233[21] , 
        \ScanLink233[20] , \ScanLink233[19] , \ScanLink233[18] , 
        \ScanLink233[17] , \ScanLink233[16] , \ScanLink233[15] , 
        \ScanLink233[14] , \ScanLink233[13] , \ScanLink233[12] , 
        \ScanLink233[11] , \ScanLink233[10] , \ScanLink233[9] , 
        \ScanLink233[8] , \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , 
        \ScanLink233[4] , \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , 
        \ScanLink233[0] }), .ScanOut({\ScanLink234[31] , \ScanLink234[30] , 
        \ScanLink234[29] , \ScanLink234[28] , \ScanLink234[27] , 
        \ScanLink234[26] , \ScanLink234[25] , \ScanLink234[24] , 
        \ScanLink234[23] , \ScanLink234[22] , \ScanLink234[21] , 
        \ScanLink234[20] , \ScanLink234[19] , \ScanLink234[18] , 
        \ScanLink234[17] , \ScanLink234[16] , \ScanLink234[15] , 
        \ScanLink234[14] , \ScanLink234[13] , \ScanLink234[12] , 
        \ScanLink234[11] , \ScanLink234[10] , \ScanLink234[9] , 
        \ScanLink234[8] , \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , 
        \ScanLink234[4] , \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , 
        \ScanLink234[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load233[0] ), .Out({\Level1Out233[31] , \Level1Out233[30] , 
        \Level1Out233[29] , \Level1Out233[28] , \Level1Out233[27] , 
        \Level1Out233[26] , \Level1Out233[25] , \Level1Out233[24] , 
        \Level1Out233[23] , \Level1Out233[22] , \Level1Out233[21] , 
        \Level1Out233[20] , \Level1Out233[19] , \Level1Out233[18] , 
        \Level1Out233[17] , \Level1Out233[16] , \Level1Out233[15] , 
        \Level1Out233[14] , \Level1Out233[13] , \Level1Out233[12] , 
        \Level1Out233[11] , \Level1Out233[10] , \Level1Out233[9] , 
        \Level1Out233[8] , \Level1Out233[7] , \Level1Out233[6] , 
        \Level1Out233[5] , \Level1Out233[4] , \Level1Out233[3] , 
        \Level1Out233[2] , \Level1Out233[1] , \Level1Out233[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_188 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink188[31] , \ScanLink188[30] , 
        \ScanLink188[29] , \ScanLink188[28] , \ScanLink188[27] , 
        \ScanLink188[26] , \ScanLink188[25] , \ScanLink188[24] , 
        \ScanLink188[23] , \ScanLink188[22] , \ScanLink188[21] , 
        \ScanLink188[20] , \ScanLink188[19] , \ScanLink188[18] , 
        \ScanLink188[17] , \ScanLink188[16] , \ScanLink188[15] , 
        \ScanLink188[14] , \ScanLink188[13] , \ScanLink188[12] , 
        \ScanLink188[11] , \ScanLink188[10] , \ScanLink188[9] , 
        \ScanLink188[8] , \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , 
        \ScanLink188[4] , \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , 
        \ScanLink188[0] }), .ScanOut({\ScanLink189[31] , \ScanLink189[30] , 
        \ScanLink189[29] , \ScanLink189[28] , \ScanLink189[27] , 
        \ScanLink189[26] , \ScanLink189[25] , \ScanLink189[24] , 
        \ScanLink189[23] , \ScanLink189[22] , \ScanLink189[21] , 
        \ScanLink189[20] , \ScanLink189[19] , \ScanLink189[18] , 
        \ScanLink189[17] , \ScanLink189[16] , \ScanLink189[15] , 
        \ScanLink189[14] , \ScanLink189[13] , \ScanLink189[12] , 
        \ScanLink189[11] , \ScanLink189[10] , \ScanLink189[9] , 
        \ScanLink189[8] , \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , 
        \ScanLink189[4] , \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , 
        \ScanLink189[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load188[0] ), .Out({\Level1Out188[31] , \Level1Out188[30] , 
        \Level1Out188[29] , \Level1Out188[28] , \Level1Out188[27] , 
        \Level1Out188[26] , \Level1Out188[25] , \Level1Out188[24] , 
        \Level1Out188[23] , \Level1Out188[22] , \Level1Out188[21] , 
        \Level1Out188[20] , \Level1Out188[19] , \Level1Out188[18] , 
        \Level1Out188[17] , \Level1Out188[16] , \Level1Out188[15] , 
        \Level1Out188[14] , \Level1Out188[13] , \Level1Out188[12] , 
        \Level1Out188[11] , \Level1Out188[10] , \Level1Out188[9] , 
        \Level1Out188[8] , \Level1Out188[7] , \Level1Out188[6] , 
        \Level1Out188[5] , \Level1Out188[4] , \Level1Out188[3] , 
        \Level1Out188[2] , \Level1Out188[1] , \Level1Out188[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_68 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink68[31] , \ScanLink68[30] , 
        \ScanLink68[29] , \ScanLink68[28] , \ScanLink68[27] , \ScanLink68[26] , 
        \ScanLink68[25] , \ScanLink68[24] , \ScanLink68[23] , \ScanLink68[22] , 
        \ScanLink68[21] , \ScanLink68[20] , \ScanLink68[19] , \ScanLink68[18] , 
        \ScanLink68[17] , \ScanLink68[16] , \ScanLink68[15] , \ScanLink68[14] , 
        \ScanLink68[13] , \ScanLink68[12] , \ScanLink68[11] , \ScanLink68[10] , 
        \ScanLink68[9] , \ScanLink68[8] , \ScanLink68[7] , \ScanLink68[6] , 
        \ScanLink68[5] , \ScanLink68[4] , \ScanLink68[3] , \ScanLink68[2] , 
        \ScanLink68[1] , \ScanLink68[0] }), .ScanOut({\ScanLink69[31] , 
        \ScanLink69[30] , \ScanLink69[29] , \ScanLink69[28] , \ScanLink69[27] , 
        \ScanLink69[26] , \ScanLink69[25] , \ScanLink69[24] , \ScanLink69[23] , 
        \ScanLink69[22] , \ScanLink69[21] , \ScanLink69[20] , \ScanLink69[19] , 
        \ScanLink69[18] , \ScanLink69[17] , \ScanLink69[16] , \ScanLink69[15] , 
        \ScanLink69[14] , \ScanLink69[13] , \ScanLink69[12] , \ScanLink69[11] , 
        \ScanLink69[10] , \ScanLink69[9] , \ScanLink69[8] , \ScanLink69[7] , 
        \ScanLink69[6] , \ScanLink69[5] , \ScanLink69[4] , \ScanLink69[3] , 
        \ScanLink69[2] , \ScanLink69[1] , \ScanLink69[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load68[0] ), .Out({
        \Level1Out68[31] , \Level1Out68[30] , \Level1Out68[29] , 
        \Level1Out68[28] , \Level1Out68[27] , \Level1Out68[26] , 
        \Level1Out68[25] , \Level1Out68[24] , \Level1Out68[23] , 
        \Level1Out68[22] , \Level1Out68[21] , \Level1Out68[20] , 
        \Level1Out68[19] , \Level1Out68[18] , \Level1Out68[17] , 
        \Level1Out68[16] , \Level1Out68[15] , \Level1Out68[14] , 
        \Level1Out68[13] , \Level1Out68[12] , \Level1Out68[11] , 
        \Level1Out68[10] , \Level1Out68[9] , \Level1Out68[8] , 
        \Level1Out68[7] , \Level1Out68[6] , \Level1Out68[5] , \Level1Out68[4] , 
        \Level1Out68[3] , \Level1Out68[2] , \Level1Out68[1] , \Level1Out68[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_36_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load36[0] ), .Out({\Level2Out36[31] , \Level2Out36[30] , 
        \Level2Out36[29] , \Level2Out36[28] , \Level2Out36[27] , 
        \Level2Out36[26] , \Level2Out36[25] , \Level2Out36[24] , 
        \Level2Out36[23] , \Level2Out36[22] , \Level2Out36[21] , 
        \Level2Out36[20] , \Level2Out36[19] , \Level2Out36[18] , 
        \Level2Out36[17] , \Level2Out36[16] , \Level2Out36[15] , 
        \Level2Out36[14] , \Level2Out36[13] , \Level2Out36[12] , 
        \Level2Out36[11] , \Level2Out36[10] , \Level2Out36[9] , 
        \Level2Out36[8] , \Level2Out36[7] , \Level2Out36[6] , \Level2Out36[5] , 
        \Level2Out36[4] , \Level2Out36[3] , \Level2Out36[2] , \Level2Out36[1] , 
        \Level2Out36[0] }), .In1({\Level1Out36[31] , \Level1Out36[30] , 
        \Level1Out36[29] , \Level1Out36[28] , \Level1Out36[27] , 
        \Level1Out36[26] , \Level1Out36[25] , \Level1Out36[24] , 
        \Level1Out36[23] , \Level1Out36[22] , \Level1Out36[21] , 
        \Level1Out36[20] , \Level1Out36[19] , \Level1Out36[18] , 
        \Level1Out36[17] , \Level1Out36[16] , \Level1Out36[15] , 
        \Level1Out36[14] , \Level1Out36[13] , \Level1Out36[12] , 
        \Level1Out36[11] , \Level1Out36[10] , \Level1Out36[9] , 
        \Level1Out36[8] , \Level1Out36[7] , \Level1Out36[6] , \Level1Out36[5] , 
        \Level1Out36[4] , \Level1Out36[3] , \Level1Out36[2] , \Level1Out36[1] , 
        \Level1Out36[0] }), .In2({\Level1Out37[31] , \Level1Out37[30] , 
        \Level1Out37[29] , \Level1Out37[28] , \Level1Out37[27] , 
        \Level1Out37[26] , \Level1Out37[25] , \Level1Out37[24] , 
        \Level1Out37[23] , \Level1Out37[22] , \Level1Out37[21] , 
        \Level1Out37[20] , \Level1Out37[19] , \Level1Out37[18] , 
        \Level1Out37[17] , \Level1Out37[16] , \Level1Out37[15] , 
        \Level1Out37[14] , \Level1Out37[13] , \Level1Out37[12] , 
        \Level1Out37[11] , \Level1Out37[10] , \Level1Out37[9] , 
        \Level1Out37[8] , \Level1Out37[7] , \Level1Out37[6] , \Level1Out37[5] , 
        \Level1Out37[4] , \Level1Out37[3] , \Level1Out37[2] , \Level1Out37[1] , 
        \Level1Out37[0] }), .Read1(\Level1Load36[0] ), .Read2(
        \Level1Load37[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_244_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load244[0] ), .Out({\Level2Out244[31] , \Level2Out244[30] , 
        \Level2Out244[29] , \Level2Out244[28] , \Level2Out244[27] , 
        \Level2Out244[26] , \Level2Out244[25] , \Level2Out244[24] , 
        \Level2Out244[23] , \Level2Out244[22] , \Level2Out244[21] , 
        \Level2Out244[20] , \Level2Out244[19] , \Level2Out244[18] , 
        \Level2Out244[17] , \Level2Out244[16] , \Level2Out244[15] , 
        \Level2Out244[14] , \Level2Out244[13] , \Level2Out244[12] , 
        \Level2Out244[11] , \Level2Out244[10] , \Level2Out244[9] , 
        \Level2Out244[8] , \Level2Out244[7] , \Level2Out244[6] , 
        \Level2Out244[5] , \Level2Out244[4] , \Level2Out244[3] , 
        \Level2Out244[2] , \Level2Out244[1] , \Level2Out244[0] }), .In1({
        \Level1Out244[31] , \Level1Out244[30] , \Level1Out244[29] , 
        \Level1Out244[28] , \Level1Out244[27] , \Level1Out244[26] , 
        \Level1Out244[25] , \Level1Out244[24] , \Level1Out244[23] , 
        \Level1Out244[22] , \Level1Out244[21] , \Level1Out244[20] , 
        \Level1Out244[19] , \Level1Out244[18] , \Level1Out244[17] , 
        \Level1Out244[16] , \Level1Out244[15] , \Level1Out244[14] , 
        \Level1Out244[13] , \Level1Out244[12] , \Level1Out244[11] , 
        \Level1Out244[10] , \Level1Out244[9] , \Level1Out244[8] , 
        \Level1Out244[7] , \Level1Out244[6] , \Level1Out244[5] , 
        \Level1Out244[4] , \Level1Out244[3] , \Level1Out244[2] , 
        \Level1Out244[1] , \Level1Out244[0] }), .In2({\Level1Out245[31] , 
        \Level1Out245[30] , \Level1Out245[29] , \Level1Out245[28] , 
        \Level1Out245[27] , \Level1Out245[26] , \Level1Out245[25] , 
        \Level1Out245[24] , \Level1Out245[23] , \Level1Out245[22] , 
        \Level1Out245[21] , \Level1Out245[20] , \Level1Out245[19] , 
        \Level1Out245[18] , \Level1Out245[17] , \Level1Out245[16] , 
        \Level1Out245[15] , \Level1Out245[14] , \Level1Out245[13] , 
        \Level1Out245[12] , \Level1Out245[11] , \Level1Out245[10] , 
        \Level1Out245[9] , \Level1Out245[8] , \Level1Out245[7] , 
        \Level1Out245[6] , \Level1Out245[5] , \Level1Out245[4] , 
        \Level1Out245[3] , \Level1Out245[2] , \Level1Out245[1] , 
        \Level1Out245[0] }), .Read1(\Level1Load244[0] ), .Read2(
        \Level1Load245[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_170_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load170[0] ), .Out({\Level2Out170[31] , \Level2Out170[30] , 
        \Level2Out170[29] , \Level2Out170[28] , \Level2Out170[27] , 
        \Level2Out170[26] , \Level2Out170[25] , \Level2Out170[24] , 
        \Level2Out170[23] , \Level2Out170[22] , \Level2Out170[21] , 
        \Level2Out170[20] , \Level2Out170[19] , \Level2Out170[18] , 
        \Level2Out170[17] , \Level2Out170[16] , \Level2Out170[15] , 
        \Level2Out170[14] , \Level2Out170[13] , \Level2Out170[12] , 
        \Level2Out170[11] , \Level2Out170[10] , \Level2Out170[9] , 
        \Level2Out170[8] , \Level2Out170[7] , \Level2Out170[6] , 
        \Level2Out170[5] , \Level2Out170[4] , \Level2Out170[3] , 
        \Level2Out170[2] , \Level2Out170[1] , \Level2Out170[0] }), .In1({
        \Level1Out170[31] , \Level1Out170[30] , \Level1Out170[29] , 
        \Level1Out170[28] , \Level1Out170[27] , \Level1Out170[26] , 
        \Level1Out170[25] , \Level1Out170[24] , \Level1Out170[23] , 
        \Level1Out170[22] , \Level1Out170[21] , \Level1Out170[20] , 
        \Level1Out170[19] , \Level1Out170[18] , \Level1Out170[17] , 
        \Level1Out170[16] , \Level1Out170[15] , \Level1Out170[14] , 
        \Level1Out170[13] , \Level1Out170[12] , \Level1Out170[11] , 
        \Level1Out170[10] , \Level1Out170[9] , \Level1Out170[8] , 
        \Level1Out170[7] , \Level1Out170[6] , \Level1Out170[5] , 
        \Level1Out170[4] , \Level1Out170[3] , \Level1Out170[2] , 
        \Level1Out170[1] , \Level1Out170[0] }), .In2({\Level1Out171[31] , 
        \Level1Out171[30] , \Level1Out171[29] , \Level1Out171[28] , 
        \Level1Out171[27] , \Level1Out171[26] , \Level1Out171[25] , 
        \Level1Out171[24] , \Level1Out171[23] , \Level1Out171[22] , 
        \Level1Out171[21] , \Level1Out171[20] , \Level1Out171[19] , 
        \Level1Out171[18] , \Level1Out171[17] , \Level1Out171[16] , 
        \Level1Out171[15] , \Level1Out171[14] , \Level1Out171[13] , 
        \Level1Out171[12] , \Level1Out171[11] , \Level1Out171[10] , 
        \Level1Out171[9] , \Level1Out171[8] , \Level1Out171[7] , 
        \Level1Out171[6] , \Level1Out171[5] , \Level1Out171[4] , 
        \Level1Out171[3] , \Level1Out171[2] , \Level1Out171[1] , 
        \Level1Out171[0] }), .Read1(\Level1Load170[0] ), .Read2(
        \Level1Load171[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_54 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanOut({\ScanLink55[31] , 
        \ScanLink55[30] , \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , 
        \ScanLink55[26] , \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , 
        \ScanLink55[22] , \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , 
        \ScanLink55[18] , \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , 
        \ScanLink55[14] , \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , 
        \ScanLink55[10] , \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , 
        \ScanLink55[6] , \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , 
        \ScanLink55[2] , \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load54[0] ), .Out({
        \Level1Out54[31] , \Level1Out54[30] , \Level1Out54[29] , 
        \Level1Out54[28] , \Level1Out54[27] , \Level1Out54[26] , 
        \Level1Out54[25] , \Level1Out54[24] , \Level1Out54[23] , 
        \Level1Out54[22] , \Level1Out54[21] , \Level1Out54[20] , 
        \Level1Out54[19] , \Level1Out54[18] , \Level1Out54[17] , 
        \Level1Out54[16] , \Level1Out54[15] , \Level1Out54[14] , 
        \Level1Out54[13] , \Level1Out54[12] , \Level1Out54[11] , 
        \Level1Out54[10] , \Level1Out54[9] , \Level1Out54[8] , 
        \Level1Out54[7] , \Level1Out54[6] , \Level1Out54[5] , \Level1Out54[4] , 
        \Level1Out54[3] , \Level1Out54[2] , \Level1Out54[1] , \Level1Out54[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_73 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink73[31] , \ScanLink73[30] , 
        \ScanLink73[29] , \ScanLink73[28] , \ScanLink73[27] , \ScanLink73[26] , 
        \ScanLink73[25] , \ScanLink73[24] , \ScanLink73[23] , \ScanLink73[22] , 
        \ScanLink73[21] , \ScanLink73[20] , \ScanLink73[19] , \ScanLink73[18] , 
        \ScanLink73[17] , \ScanLink73[16] , \ScanLink73[15] , \ScanLink73[14] , 
        \ScanLink73[13] , \ScanLink73[12] , \ScanLink73[11] , \ScanLink73[10] , 
        \ScanLink73[9] , \ScanLink73[8] , \ScanLink73[7] , \ScanLink73[6] , 
        \ScanLink73[5] , \ScanLink73[4] , \ScanLink73[3] , \ScanLink73[2] , 
        \ScanLink73[1] , \ScanLink73[0] }), .ScanOut({\ScanLink74[31] , 
        \ScanLink74[30] , \ScanLink74[29] , \ScanLink74[28] , \ScanLink74[27] , 
        \ScanLink74[26] , \ScanLink74[25] , \ScanLink74[24] , \ScanLink74[23] , 
        \ScanLink74[22] , \ScanLink74[21] , \ScanLink74[20] , \ScanLink74[19] , 
        \ScanLink74[18] , \ScanLink74[17] , \ScanLink74[16] , \ScanLink74[15] , 
        \ScanLink74[14] , \ScanLink74[13] , \ScanLink74[12] , \ScanLink74[11] , 
        \ScanLink74[10] , \ScanLink74[9] , \ScanLink74[8] , \ScanLink74[7] , 
        \ScanLink74[6] , \ScanLink74[5] , \ScanLink74[4] , \ScanLink74[3] , 
        \ScanLink74[2] , \ScanLink74[1] , \ScanLink74[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load73[0] ), .Out({
        \Level1Out73[31] , \Level1Out73[30] , \Level1Out73[29] , 
        \Level1Out73[28] , \Level1Out73[27] , \Level1Out73[26] , 
        \Level1Out73[25] , \Level1Out73[24] , \Level1Out73[23] , 
        \Level1Out73[22] , \Level1Out73[21] , \Level1Out73[20] , 
        \Level1Out73[19] , \Level1Out73[18] , \Level1Out73[17] , 
        \Level1Out73[16] , \Level1Out73[15] , \Level1Out73[14] , 
        \Level1Out73[13] , \Level1Out73[12] , \Level1Out73[11] , 
        \Level1Out73[10] , \Level1Out73[9] , \Level1Out73[8] , 
        \Level1Out73[7] , \Level1Out73[6] , \Level1Out73[5] , \Level1Out73[4] , 
        \Level1Out73[3] , \Level1Out73[2] , \Level1Out73[1] , \Level1Out73[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_151 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink151[31] , \ScanLink151[30] , 
        \ScanLink151[29] , \ScanLink151[28] , \ScanLink151[27] , 
        \ScanLink151[26] , \ScanLink151[25] , \ScanLink151[24] , 
        \ScanLink151[23] , \ScanLink151[22] , \ScanLink151[21] , 
        \ScanLink151[20] , \ScanLink151[19] , \ScanLink151[18] , 
        \ScanLink151[17] , \ScanLink151[16] , \ScanLink151[15] , 
        \ScanLink151[14] , \ScanLink151[13] , \ScanLink151[12] , 
        \ScanLink151[11] , \ScanLink151[10] , \ScanLink151[9] , 
        \ScanLink151[8] , \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , 
        \ScanLink151[4] , \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , 
        \ScanLink151[0] }), .ScanOut({\ScanLink152[31] , \ScanLink152[30] , 
        \ScanLink152[29] , \ScanLink152[28] , \ScanLink152[27] , 
        \ScanLink152[26] , \ScanLink152[25] , \ScanLink152[24] , 
        \ScanLink152[23] , \ScanLink152[22] , \ScanLink152[21] , 
        \ScanLink152[20] , \ScanLink152[19] , \ScanLink152[18] , 
        \ScanLink152[17] , \ScanLink152[16] , \ScanLink152[15] , 
        \ScanLink152[14] , \ScanLink152[13] , \ScanLink152[12] , 
        \ScanLink152[11] , \ScanLink152[10] , \ScanLink152[9] , 
        \ScanLink152[8] , \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , 
        \ScanLink152[4] , \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , 
        \ScanLink152[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load151[0] ), .Out({\Level1Out151[31] , \Level1Out151[30] , 
        \Level1Out151[29] , \Level1Out151[28] , \Level1Out151[27] , 
        \Level1Out151[26] , \Level1Out151[25] , \Level1Out151[24] , 
        \Level1Out151[23] , \Level1Out151[22] , \Level1Out151[21] , 
        \Level1Out151[20] , \Level1Out151[19] , \Level1Out151[18] , 
        \Level1Out151[17] , \Level1Out151[16] , \Level1Out151[15] , 
        \Level1Out151[14] , \Level1Out151[13] , \Level1Out151[12] , 
        \Level1Out151[11] , \Level1Out151[10] , \Level1Out151[9] , 
        \Level1Out151[8] , \Level1Out151[7] , \Level1Out151[6] , 
        \Level1Out151[5] , \Level1Out151[4] , \Level1Out151[3] , 
        \Level1Out151[2] , \Level1Out151[1] , \Level1Out151[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_176 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink176[31] , \ScanLink176[30] , 
        \ScanLink176[29] , \ScanLink176[28] , \ScanLink176[27] , 
        \ScanLink176[26] , \ScanLink176[25] , \ScanLink176[24] , 
        \ScanLink176[23] , \ScanLink176[22] , \ScanLink176[21] , 
        \ScanLink176[20] , \ScanLink176[19] , \ScanLink176[18] , 
        \ScanLink176[17] , \ScanLink176[16] , \ScanLink176[15] , 
        \ScanLink176[14] , \ScanLink176[13] , \ScanLink176[12] , 
        \ScanLink176[11] , \ScanLink176[10] , \ScanLink176[9] , 
        \ScanLink176[8] , \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , 
        \ScanLink176[4] , \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , 
        \ScanLink176[0] }), .ScanOut({\ScanLink177[31] , \ScanLink177[30] , 
        \ScanLink177[29] , \ScanLink177[28] , \ScanLink177[27] , 
        \ScanLink177[26] , \ScanLink177[25] , \ScanLink177[24] , 
        \ScanLink177[23] , \ScanLink177[22] , \ScanLink177[21] , 
        \ScanLink177[20] , \ScanLink177[19] , \ScanLink177[18] , 
        \ScanLink177[17] , \ScanLink177[16] , \ScanLink177[15] , 
        \ScanLink177[14] , \ScanLink177[13] , \ScanLink177[12] , 
        \ScanLink177[11] , \ScanLink177[10] , \ScanLink177[9] , 
        \ScanLink177[8] , \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , 
        \ScanLink177[4] , \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , 
        \ScanLink177[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load176[0] ), .Out({\Level1Out176[31] , \Level1Out176[30] , 
        \Level1Out176[29] , \Level1Out176[28] , \Level1Out176[27] , 
        \Level1Out176[26] , \Level1Out176[25] , \Level1Out176[24] , 
        \Level1Out176[23] , \Level1Out176[22] , \Level1Out176[21] , 
        \Level1Out176[20] , \Level1Out176[19] , \Level1Out176[18] , 
        \Level1Out176[17] , \Level1Out176[16] , \Level1Out176[15] , 
        \Level1Out176[14] , \Level1Out176[13] , \Level1Out176[12] , 
        \Level1Out176[11] , \Level1Out176[10] , \Level1Out176[9] , 
        \Level1Out176[8] , \Level1Out176[7] , \Level1Out176[6] , 
        \Level1Out176[5] , \Level1Out176[4] , \Level1Out176[3] , 
        \Level1Out176[2] , \Level1Out176[1] , \Level1Out176[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_246 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink246[31] , \ScanLink246[30] , 
        \ScanLink246[29] , \ScanLink246[28] , \ScanLink246[27] , 
        \ScanLink246[26] , \ScanLink246[25] , \ScanLink246[24] , 
        \ScanLink246[23] , \ScanLink246[22] , \ScanLink246[21] , 
        \ScanLink246[20] , \ScanLink246[19] , \ScanLink246[18] , 
        \ScanLink246[17] , \ScanLink246[16] , \ScanLink246[15] , 
        \ScanLink246[14] , \ScanLink246[13] , \ScanLink246[12] , 
        \ScanLink246[11] , \ScanLink246[10] , \ScanLink246[9] , 
        \ScanLink246[8] , \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , 
        \ScanLink246[4] , \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , 
        \ScanLink246[0] }), .ScanOut({\ScanLink247[31] , \ScanLink247[30] , 
        \ScanLink247[29] , \ScanLink247[28] , \ScanLink247[27] , 
        \ScanLink247[26] , \ScanLink247[25] , \ScanLink247[24] , 
        \ScanLink247[23] , \ScanLink247[22] , \ScanLink247[21] , 
        \ScanLink247[20] , \ScanLink247[19] , \ScanLink247[18] , 
        \ScanLink247[17] , \ScanLink247[16] , \ScanLink247[15] , 
        \ScanLink247[14] , \ScanLink247[13] , \ScanLink247[12] , 
        \ScanLink247[11] , \ScanLink247[10] , \ScanLink247[9] , 
        \ScanLink247[8] , \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , 
        \ScanLink247[4] , \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , 
        \ScanLink247[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load246[0] ), .Out({\Level1Out246[31] , \Level1Out246[30] , 
        \Level1Out246[29] , \Level1Out246[28] , \Level1Out246[27] , 
        \Level1Out246[26] , \Level1Out246[25] , \Level1Out246[24] , 
        \Level1Out246[23] , \Level1Out246[22] , \Level1Out246[21] , 
        \Level1Out246[20] , \Level1Out246[19] , \Level1Out246[18] , 
        \Level1Out246[17] , \Level1Out246[16] , \Level1Out246[15] , 
        \Level1Out246[14] , \Level1Out246[13] , \Level1Out246[12] , 
        \Level1Out246[11] , \Level1Out246[10] , \Level1Out246[9] , 
        \Level1Out246[8] , \Level1Out246[7] , \Level1Out246[6] , 
        \Level1Out246[5] , \Level1Out246[4] , \Level1Out246[3] , 
        \Level1Out246[2] , \Level1Out246[1] , \Level1Out246[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load32[0] ), .Out({\Level4Out32[31] , \Level4Out32[30] , 
        \Level4Out32[29] , \Level4Out32[28] , \Level4Out32[27] , 
        \Level4Out32[26] , \Level4Out32[25] , \Level4Out32[24] , 
        \Level4Out32[23] , \Level4Out32[22] , \Level4Out32[21] , 
        \Level4Out32[20] , \Level4Out32[19] , \Level4Out32[18] , 
        \Level4Out32[17] , \Level4Out32[16] , \Level4Out32[15] , 
        \Level4Out32[14] , \Level4Out32[13] , \Level4Out32[12] , 
        \Level4Out32[11] , \Level4Out32[10] , \Level4Out32[9] , 
        \Level4Out32[8] , \Level4Out32[7] , \Level4Out32[6] , \Level4Out32[5] , 
        \Level4Out32[4] , \Level4Out32[3] , \Level4Out32[2] , \Level4Out32[1] , 
        \Level4Out32[0] }), .In1({\Level2Out32[31] , \Level2Out32[30] , 
        \Level2Out32[29] , \Level2Out32[28] , \Level2Out32[27] , 
        \Level2Out32[26] , \Level2Out32[25] , \Level2Out32[24] , 
        \Level2Out32[23] , \Level2Out32[22] , \Level2Out32[21] , 
        \Level2Out32[20] , \Level2Out32[19] , \Level2Out32[18] , 
        \Level2Out32[17] , \Level2Out32[16] , \Level2Out32[15] , 
        \Level2Out32[14] , \Level2Out32[13] , \Level2Out32[12] , 
        \Level2Out32[11] , \Level2Out32[10] , \Level2Out32[9] , 
        \Level2Out32[8] , \Level2Out32[7] , \Level2Out32[6] , \Level2Out32[5] , 
        \Level2Out32[4] , \Level2Out32[3] , \Level2Out32[2] , \Level2Out32[1] , 
        \Level2Out32[0] }), .In2({\Level2Out34[31] , \Level2Out34[30] , 
        \Level2Out34[29] , \Level2Out34[28] , \Level2Out34[27] , 
        \Level2Out34[26] , \Level2Out34[25] , \Level2Out34[24] , 
        \Level2Out34[23] , \Level2Out34[22] , \Level2Out34[21] , 
        \Level2Out34[20] , \Level2Out34[19] , \Level2Out34[18] , 
        \Level2Out34[17] , \Level2Out34[16] , \Level2Out34[15] , 
        \Level2Out34[14] , \Level2Out34[13] , \Level2Out34[12] , 
        \Level2Out34[11] , \Level2Out34[10] , \Level2Out34[9] , 
        \Level2Out34[8] , \Level2Out34[7] , \Level2Out34[6] , \Level2Out34[5] , 
        \Level2Out34[4] , \Level2Out34[3] , \Level2Out34[2] , \Level2Out34[1] , 
        \Level2Out34[0] }), .Read1(\Level2Load32[0] ), .Read2(
        \Level2Load34[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_96_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load96[0] ), .Out({\Level4Out96[31] , \Level4Out96[30] , 
        \Level4Out96[29] , \Level4Out96[28] , \Level4Out96[27] , 
        \Level4Out96[26] , \Level4Out96[25] , \Level4Out96[24] , 
        \Level4Out96[23] , \Level4Out96[22] , \Level4Out96[21] , 
        \Level4Out96[20] , \Level4Out96[19] , \Level4Out96[18] , 
        \Level4Out96[17] , \Level4Out96[16] , \Level4Out96[15] , 
        \Level4Out96[14] , \Level4Out96[13] , \Level4Out96[12] , 
        \Level4Out96[11] , \Level4Out96[10] , \Level4Out96[9] , 
        \Level4Out96[8] , \Level4Out96[7] , \Level4Out96[6] , \Level4Out96[5] , 
        \Level4Out96[4] , \Level4Out96[3] , \Level4Out96[2] , \Level4Out96[1] , 
        \Level4Out96[0] }), .In1({\Level2Out96[31] , \Level2Out96[30] , 
        \Level2Out96[29] , \Level2Out96[28] , \Level2Out96[27] , 
        \Level2Out96[26] , \Level2Out96[25] , \Level2Out96[24] , 
        \Level2Out96[23] , \Level2Out96[22] , \Level2Out96[21] , 
        \Level2Out96[20] , \Level2Out96[19] , \Level2Out96[18] , 
        \Level2Out96[17] , \Level2Out96[16] , \Level2Out96[15] , 
        \Level2Out96[14] , \Level2Out96[13] , \Level2Out96[12] , 
        \Level2Out96[11] , \Level2Out96[10] , \Level2Out96[9] , 
        \Level2Out96[8] , \Level2Out96[7] , \Level2Out96[6] , \Level2Out96[5] , 
        \Level2Out96[4] , \Level2Out96[3] , \Level2Out96[2] , \Level2Out96[1] , 
        \Level2Out96[0] }), .In2({\Level2Out98[31] , \Level2Out98[30] , 
        \Level2Out98[29] , \Level2Out98[28] , \Level2Out98[27] , 
        \Level2Out98[26] , \Level2Out98[25] , \Level2Out98[24] , 
        \Level2Out98[23] , \Level2Out98[22] , \Level2Out98[21] , 
        \Level2Out98[20] , \Level2Out98[19] , \Level2Out98[18] , 
        \Level2Out98[17] , \Level2Out98[16] , \Level2Out98[15] , 
        \Level2Out98[14] , \Level2Out98[13] , \Level2Out98[12] , 
        \Level2Out98[11] , \Level2Out98[10] , \Level2Out98[9] , 
        \Level2Out98[8] , \Level2Out98[7] , \Level2Out98[6] , \Level2Out98[5] , 
        \Level2Out98[4] , \Level2Out98[3] , \Level2Out98[2] , \Level2Out98[1] , 
        \Level2Out98[0] }), .Read1(\Level2Load96[0] ), .Read2(
        \Level2Load98[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_144_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load144[0] ), .Out({\Level8Out144[31] , \Level8Out144[30] , 
        \Level8Out144[29] , \Level8Out144[28] , \Level8Out144[27] , 
        \Level8Out144[26] , \Level8Out144[25] , \Level8Out144[24] , 
        \Level8Out144[23] , \Level8Out144[22] , \Level8Out144[21] , 
        \Level8Out144[20] , \Level8Out144[19] , \Level8Out144[18] , 
        \Level8Out144[17] , \Level8Out144[16] , \Level8Out144[15] , 
        \Level8Out144[14] , \Level8Out144[13] , \Level8Out144[12] , 
        \Level8Out144[11] , \Level8Out144[10] , \Level8Out144[9] , 
        \Level8Out144[8] , \Level8Out144[7] , \Level8Out144[6] , 
        \Level8Out144[5] , \Level8Out144[4] , \Level8Out144[3] , 
        \Level8Out144[2] , \Level8Out144[1] , \Level8Out144[0] }), .In1({
        \Level4Out144[31] , \Level4Out144[30] , \Level4Out144[29] , 
        \Level4Out144[28] , \Level4Out144[27] , \Level4Out144[26] , 
        \Level4Out144[25] , \Level4Out144[24] , \Level4Out144[23] , 
        \Level4Out144[22] , \Level4Out144[21] , \Level4Out144[20] , 
        \Level4Out144[19] , \Level4Out144[18] , \Level4Out144[17] , 
        \Level4Out144[16] , \Level4Out144[15] , \Level4Out144[14] , 
        \Level4Out144[13] , \Level4Out144[12] , \Level4Out144[11] , 
        \Level4Out144[10] , \Level4Out144[9] , \Level4Out144[8] , 
        \Level4Out144[7] , \Level4Out144[6] , \Level4Out144[5] , 
        \Level4Out144[4] , \Level4Out144[3] , \Level4Out144[2] , 
        \Level4Out144[1] , \Level4Out144[0] }), .In2({\Level4Out148[31] , 
        \Level4Out148[30] , \Level4Out148[29] , \Level4Out148[28] , 
        \Level4Out148[27] , \Level4Out148[26] , \Level4Out148[25] , 
        \Level4Out148[24] , \Level4Out148[23] , \Level4Out148[22] , 
        \Level4Out148[21] , \Level4Out148[20] , \Level4Out148[19] , 
        \Level4Out148[18] , \Level4Out148[17] , \Level4Out148[16] , 
        \Level4Out148[15] , \Level4Out148[14] , \Level4Out148[13] , 
        \Level4Out148[12] , \Level4Out148[11] , \Level4Out148[10] , 
        \Level4Out148[9] , \Level4Out148[8] , \Level4Out148[7] , 
        \Level4Out148[6] , \Level4Out148[5] , \Level4Out148[4] , 
        \Level4Out148[3] , \Level4Out148[2] , \Level4Out148[1] , 
        \Level4Out148[0] }), .Read1(\Level4Load144[0] ), .Read2(
        \Level4Load148[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_142_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load142[0] ), .Out({\Level2Out142[31] , \Level2Out142[30] , 
        \Level2Out142[29] , \Level2Out142[28] , \Level2Out142[27] , 
        \Level2Out142[26] , \Level2Out142[25] , \Level2Out142[24] , 
        \Level2Out142[23] , \Level2Out142[22] , \Level2Out142[21] , 
        \Level2Out142[20] , \Level2Out142[19] , \Level2Out142[18] , 
        \Level2Out142[17] , \Level2Out142[16] , \Level2Out142[15] , 
        \Level2Out142[14] , \Level2Out142[13] , \Level2Out142[12] , 
        \Level2Out142[11] , \Level2Out142[10] , \Level2Out142[9] , 
        \Level2Out142[8] , \Level2Out142[7] , \Level2Out142[6] , 
        \Level2Out142[5] , \Level2Out142[4] , \Level2Out142[3] , 
        \Level2Out142[2] , \Level2Out142[1] , \Level2Out142[0] }), .In1({
        \Level1Out142[31] , \Level1Out142[30] , \Level1Out142[29] , 
        \Level1Out142[28] , \Level1Out142[27] , \Level1Out142[26] , 
        \Level1Out142[25] , \Level1Out142[24] , \Level1Out142[23] , 
        \Level1Out142[22] , \Level1Out142[21] , \Level1Out142[20] , 
        \Level1Out142[19] , \Level1Out142[18] , \Level1Out142[17] , 
        \Level1Out142[16] , \Level1Out142[15] , \Level1Out142[14] , 
        \Level1Out142[13] , \Level1Out142[12] , \Level1Out142[11] , 
        \Level1Out142[10] , \Level1Out142[9] , \Level1Out142[8] , 
        \Level1Out142[7] , \Level1Out142[6] , \Level1Out142[5] , 
        \Level1Out142[4] , \Level1Out142[3] , \Level1Out142[2] , 
        \Level1Out142[1] , \Level1Out142[0] }), .In2({\Level1Out143[31] , 
        \Level1Out143[30] , \Level1Out143[29] , \Level1Out143[28] , 
        \Level1Out143[27] , \Level1Out143[26] , \Level1Out143[25] , 
        \Level1Out143[24] , \Level1Out143[23] , \Level1Out143[22] , 
        \Level1Out143[21] , \Level1Out143[20] , \Level1Out143[19] , 
        \Level1Out143[18] , \Level1Out143[17] , \Level1Out143[16] , 
        \Level1Out143[15] , \Level1Out143[14] , \Level1Out143[13] , 
        \Level1Out143[12] , \Level1Out143[11] , \Level1Out143[10] , 
        \Level1Out143[9] , \Level1Out143[8] , \Level1Out143[7] , 
        \Level1Out143[6] , \Level1Out143[5] , \Level1Out143[4] , 
        \Level1Out143[3] , \Level1Out143[2] , \Level1Out143[1] , 
        \Level1Out143[0] }), .Read1(\Level1Load142[0] ), .Read2(
        \Level1Load143[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_168_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load168[0] ), .Out({\Level2Out168[31] , \Level2Out168[30] , 
        \Level2Out168[29] , \Level2Out168[28] , \Level2Out168[27] , 
        \Level2Out168[26] , \Level2Out168[25] , \Level2Out168[24] , 
        \Level2Out168[23] , \Level2Out168[22] , \Level2Out168[21] , 
        \Level2Out168[20] , \Level2Out168[19] , \Level2Out168[18] , 
        \Level2Out168[17] , \Level2Out168[16] , \Level2Out168[15] , 
        \Level2Out168[14] , \Level2Out168[13] , \Level2Out168[12] , 
        \Level2Out168[11] , \Level2Out168[10] , \Level2Out168[9] , 
        \Level2Out168[8] , \Level2Out168[7] , \Level2Out168[6] , 
        \Level2Out168[5] , \Level2Out168[4] , \Level2Out168[3] , 
        \Level2Out168[2] , \Level2Out168[1] , \Level2Out168[0] }), .In1({
        \Level1Out168[31] , \Level1Out168[30] , \Level1Out168[29] , 
        \Level1Out168[28] , \Level1Out168[27] , \Level1Out168[26] , 
        \Level1Out168[25] , \Level1Out168[24] , \Level1Out168[23] , 
        \Level1Out168[22] , \Level1Out168[21] , \Level1Out168[20] , 
        \Level1Out168[19] , \Level1Out168[18] , \Level1Out168[17] , 
        \Level1Out168[16] , \Level1Out168[15] , \Level1Out168[14] , 
        \Level1Out168[13] , \Level1Out168[12] , \Level1Out168[11] , 
        \Level1Out168[10] , \Level1Out168[9] , \Level1Out168[8] , 
        \Level1Out168[7] , \Level1Out168[6] , \Level1Out168[5] , 
        \Level1Out168[4] , \Level1Out168[3] , \Level1Out168[2] , 
        \Level1Out168[1] , \Level1Out168[0] }), .In2({\Level1Out169[31] , 
        \Level1Out169[30] , \Level1Out169[29] , \Level1Out169[28] , 
        \Level1Out169[27] , \Level1Out169[26] , \Level1Out169[25] , 
        \Level1Out169[24] , \Level1Out169[23] , \Level1Out169[22] , 
        \Level1Out169[21] , \Level1Out169[20] , \Level1Out169[19] , 
        \Level1Out169[18] , \Level1Out169[17] , \Level1Out169[16] , 
        \Level1Out169[15] , \Level1Out169[14] , \Level1Out169[13] , 
        \Level1Out169[12] , \Level1Out169[11] , \Level1Out169[10] , 
        \Level1Out169[9] , \Level1Out169[8] , \Level1Out169[7] , 
        \Level1Out169[6] , \Level1Out169[5] , \Level1Out169[4] , 
        \Level1Out169[3] , \Level1Out169[2] , \Level1Out169[1] , 
        \Level1Out169[0] }), .Read1(\Level1Load168[0] ), .Read2(
        \Level1Load169[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_240_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load240[0] ), .Out({\Level4Out240[31] , \Level4Out240[30] , 
        \Level4Out240[29] , \Level4Out240[28] , \Level4Out240[27] , 
        \Level4Out240[26] , \Level4Out240[25] , \Level4Out240[24] , 
        \Level4Out240[23] , \Level4Out240[22] , \Level4Out240[21] , 
        \Level4Out240[20] , \Level4Out240[19] , \Level4Out240[18] , 
        \Level4Out240[17] , \Level4Out240[16] , \Level4Out240[15] , 
        \Level4Out240[14] , \Level4Out240[13] , \Level4Out240[12] , 
        \Level4Out240[11] , \Level4Out240[10] , \Level4Out240[9] , 
        \Level4Out240[8] , \Level4Out240[7] , \Level4Out240[6] , 
        \Level4Out240[5] , \Level4Out240[4] , \Level4Out240[3] , 
        \Level4Out240[2] , \Level4Out240[1] , \Level4Out240[0] }), .In1({
        \Level2Out240[31] , \Level2Out240[30] , \Level2Out240[29] , 
        \Level2Out240[28] , \Level2Out240[27] , \Level2Out240[26] , 
        \Level2Out240[25] , \Level2Out240[24] , \Level2Out240[23] , 
        \Level2Out240[22] , \Level2Out240[21] , \Level2Out240[20] , 
        \Level2Out240[19] , \Level2Out240[18] , \Level2Out240[17] , 
        \Level2Out240[16] , \Level2Out240[15] , \Level2Out240[14] , 
        \Level2Out240[13] , \Level2Out240[12] , \Level2Out240[11] , 
        \Level2Out240[10] , \Level2Out240[9] , \Level2Out240[8] , 
        \Level2Out240[7] , \Level2Out240[6] , \Level2Out240[5] , 
        \Level2Out240[4] , \Level2Out240[3] , \Level2Out240[2] , 
        \Level2Out240[1] , \Level2Out240[0] }), .In2({\Level2Out242[31] , 
        \Level2Out242[30] , \Level2Out242[29] , \Level2Out242[28] , 
        \Level2Out242[27] , \Level2Out242[26] , \Level2Out242[25] , 
        \Level2Out242[24] , \Level2Out242[23] , \Level2Out242[22] , 
        \Level2Out242[21] , \Level2Out242[20] , \Level2Out242[19] , 
        \Level2Out242[18] , \Level2Out242[17] , \Level2Out242[16] , 
        \Level2Out242[15] , \Level2Out242[14] , \Level2Out242[13] , 
        \Level2Out242[12] , \Level2Out242[11] , \Level2Out242[10] , 
        \Level2Out242[9] , \Level2Out242[8] , \Level2Out242[7] , 
        \Level2Out242[6] , \Level2Out242[5] , \Level2Out242[4] , 
        \Level2Out242[3] , \Level2Out242[2] , \Level2Out242[1] , 
        \Level2Out242[0] }), .Read1(\Level2Load240[0] ), .Read2(
        \Level2Load242[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_176_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load176[0] ), .Out({\Level8Out176[31] , \Level8Out176[30] , 
        \Level8Out176[29] , \Level8Out176[28] , \Level8Out176[27] , 
        \Level8Out176[26] , \Level8Out176[25] , \Level8Out176[24] , 
        \Level8Out176[23] , \Level8Out176[22] , \Level8Out176[21] , 
        \Level8Out176[20] , \Level8Out176[19] , \Level8Out176[18] , 
        \Level8Out176[17] , \Level8Out176[16] , \Level8Out176[15] , 
        \Level8Out176[14] , \Level8Out176[13] , \Level8Out176[12] , 
        \Level8Out176[11] , \Level8Out176[10] , \Level8Out176[9] , 
        \Level8Out176[8] , \Level8Out176[7] , \Level8Out176[6] , 
        \Level8Out176[5] , \Level8Out176[4] , \Level8Out176[3] , 
        \Level8Out176[2] , \Level8Out176[1] , \Level8Out176[0] }), .In1({
        \Level4Out176[31] , \Level4Out176[30] , \Level4Out176[29] , 
        \Level4Out176[28] , \Level4Out176[27] , \Level4Out176[26] , 
        \Level4Out176[25] , \Level4Out176[24] , \Level4Out176[23] , 
        \Level4Out176[22] , \Level4Out176[21] , \Level4Out176[20] , 
        \Level4Out176[19] , \Level4Out176[18] , \Level4Out176[17] , 
        \Level4Out176[16] , \Level4Out176[15] , \Level4Out176[14] , 
        \Level4Out176[13] , \Level4Out176[12] , \Level4Out176[11] , 
        \Level4Out176[10] , \Level4Out176[9] , \Level4Out176[8] , 
        \Level4Out176[7] , \Level4Out176[6] , \Level4Out176[5] , 
        \Level4Out176[4] , \Level4Out176[3] , \Level4Out176[2] , 
        \Level4Out176[1] , \Level4Out176[0] }), .In2({\Level4Out180[31] , 
        \Level4Out180[30] , \Level4Out180[29] , \Level4Out180[28] , 
        \Level4Out180[27] , \Level4Out180[26] , \Level4Out180[25] , 
        \Level4Out180[24] , \Level4Out180[23] , \Level4Out180[22] , 
        \Level4Out180[21] , \Level4Out180[20] , \Level4Out180[19] , 
        \Level4Out180[18] , \Level4Out180[17] , \Level4Out180[16] , 
        \Level4Out180[15] , \Level4Out180[14] , \Level4Out180[13] , 
        \Level4Out180[12] , \Level4Out180[11] , \Level4Out180[10] , 
        \Level4Out180[9] , \Level4Out180[8] , \Level4Out180[7] , 
        \Level4Out180[6] , \Level4Out180[5] , \Level4Out180[4] , 
        \Level4Out180[3] , \Level4Out180[2] , \Level4Out180[1] , 
        \Level4Out180[0] }), .Read1(\Level4Load176[0] ), .Read2(
        \Level4Load180[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_96 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink96[31] , \ScanLink96[30] , 
        \ScanLink96[29] , \ScanLink96[28] , \ScanLink96[27] , \ScanLink96[26] , 
        \ScanLink96[25] , \ScanLink96[24] , \ScanLink96[23] , \ScanLink96[22] , 
        \ScanLink96[21] , \ScanLink96[20] , \ScanLink96[19] , \ScanLink96[18] , 
        \ScanLink96[17] , \ScanLink96[16] , \ScanLink96[15] , \ScanLink96[14] , 
        \ScanLink96[13] , \ScanLink96[12] , \ScanLink96[11] , \ScanLink96[10] , 
        \ScanLink96[9] , \ScanLink96[8] , \ScanLink96[7] , \ScanLink96[6] , 
        \ScanLink96[5] , \ScanLink96[4] , \ScanLink96[3] , \ScanLink96[2] , 
        \ScanLink96[1] , \ScanLink96[0] }), .ScanOut({\ScanLink97[31] , 
        \ScanLink97[30] , \ScanLink97[29] , \ScanLink97[28] , \ScanLink97[27] , 
        \ScanLink97[26] , \ScanLink97[25] , \ScanLink97[24] , \ScanLink97[23] , 
        \ScanLink97[22] , \ScanLink97[21] , \ScanLink97[20] , \ScanLink97[19] , 
        \ScanLink97[18] , \ScanLink97[17] , \ScanLink97[16] , \ScanLink97[15] , 
        \ScanLink97[14] , \ScanLink97[13] , \ScanLink97[12] , \ScanLink97[11] , 
        \ScanLink97[10] , \ScanLink97[9] , \ScanLink97[8] , \ScanLink97[7] , 
        \ScanLink97[6] , \ScanLink97[5] , \ScanLink97[4] , \ScanLink97[3] , 
        \ScanLink97[2] , \ScanLink97[1] , \ScanLink97[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load96[0] ), .Out({
        \Level1Out96[31] , \Level1Out96[30] , \Level1Out96[29] , 
        \Level1Out96[28] , \Level1Out96[27] , \Level1Out96[26] , 
        \Level1Out96[25] , \Level1Out96[24] , \Level1Out96[23] , 
        \Level1Out96[22] , \Level1Out96[21] , \Level1Out96[20] , 
        \Level1Out96[19] , \Level1Out96[18] , \Level1Out96[17] , 
        \Level1Out96[16] , \Level1Out96[15] , \Level1Out96[14] , 
        \Level1Out96[13] , \Level1Out96[12] , \Level1Out96[11] , 
        \Level1Out96[10] , \Level1Out96[9] , \Level1Out96[8] , 
        \Level1Out96[7] , \Level1Out96[6] , \Level1Out96[5] , \Level1Out96[4] , 
        \Level1Out96[3] , \Level1Out96[2] , \Level1Out96[1] , \Level1Out96[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_118 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink118[31] , \ScanLink118[30] , 
        \ScanLink118[29] , \ScanLink118[28] , \ScanLink118[27] , 
        \ScanLink118[26] , \ScanLink118[25] , \ScanLink118[24] , 
        \ScanLink118[23] , \ScanLink118[22] , \ScanLink118[21] , 
        \ScanLink118[20] , \ScanLink118[19] , \ScanLink118[18] , 
        \ScanLink118[17] , \ScanLink118[16] , \ScanLink118[15] , 
        \ScanLink118[14] , \ScanLink118[13] , \ScanLink118[12] , 
        \ScanLink118[11] , \ScanLink118[10] , \ScanLink118[9] , 
        \ScanLink118[8] , \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , 
        \ScanLink118[4] , \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , 
        \ScanLink118[0] }), .ScanOut({\ScanLink119[31] , \ScanLink119[30] , 
        \ScanLink119[29] , \ScanLink119[28] , \ScanLink119[27] , 
        \ScanLink119[26] , \ScanLink119[25] , \ScanLink119[24] , 
        \ScanLink119[23] , \ScanLink119[22] , \ScanLink119[21] , 
        \ScanLink119[20] , \ScanLink119[19] , \ScanLink119[18] , 
        \ScanLink119[17] , \ScanLink119[16] , \ScanLink119[15] , 
        \ScanLink119[14] , \ScanLink119[13] , \ScanLink119[12] , 
        \ScanLink119[11] , \ScanLink119[10] , \ScanLink119[9] , 
        \ScanLink119[8] , \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , 
        \ScanLink119[4] , \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , 
        \ScanLink119[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load118[0] ), .Out({\Level1Out118[31] , \Level1Out118[30] , 
        \Level1Out118[29] , \Level1Out118[28] , \Level1Out118[27] , 
        \Level1Out118[26] , \Level1Out118[25] , \Level1Out118[24] , 
        \Level1Out118[23] , \Level1Out118[22] , \Level1Out118[21] , 
        \Level1Out118[20] , \Level1Out118[19] , \Level1Out118[18] , 
        \Level1Out118[17] , \Level1Out118[16] , \Level1Out118[15] , 
        \Level1Out118[14] , \Level1Out118[13] , \Level1Out118[12] , 
        \Level1Out118[11] , \Level1Out118[10] , \Level1Out118[9] , 
        \Level1Out118[8] , \Level1Out118[7] , \Level1Out118[6] , 
        \Level1Out118[5] , \Level1Out118[4] , \Level1Out118[3] , 
        \Level1Out118[2] , \Level1Out118[1] , \Level1Out118[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_193 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink193[31] , \ScanLink193[30] , 
        \ScanLink193[29] , \ScanLink193[28] , \ScanLink193[27] , 
        \ScanLink193[26] , \ScanLink193[25] , \ScanLink193[24] , 
        \ScanLink193[23] , \ScanLink193[22] , \ScanLink193[21] , 
        \ScanLink193[20] , \ScanLink193[19] , \ScanLink193[18] , 
        \ScanLink193[17] , \ScanLink193[16] , \ScanLink193[15] , 
        \ScanLink193[14] , \ScanLink193[13] , \ScanLink193[12] , 
        \ScanLink193[11] , \ScanLink193[10] , \ScanLink193[9] , 
        \ScanLink193[8] , \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , 
        \ScanLink193[4] , \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , 
        \ScanLink193[0] }), .ScanOut({\ScanLink194[31] , \ScanLink194[30] , 
        \ScanLink194[29] , \ScanLink194[28] , \ScanLink194[27] , 
        \ScanLink194[26] , \ScanLink194[25] , \ScanLink194[24] , 
        \ScanLink194[23] , \ScanLink194[22] , \ScanLink194[21] , 
        \ScanLink194[20] , \ScanLink194[19] , \ScanLink194[18] , 
        \ScanLink194[17] , \ScanLink194[16] , \ScanLink194[15] , 
        \ScanLink194[14] , \ScanLink194[13] , \ScanLink194[12] , 
        \ScanLink194[11] , \ScanLink194[10] , \ScanLink194[9] , 
        \ScanLink194[8] , \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , 
        \ScanLink194[4] , \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , 
        \ScanLink194[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load193[0] ), .Out({\Level1Out193[31] , \Level1Out193[30] , 
        \Level1Out193[29] , \Level1Out193[28] , \Level1Out193[27] , 
        \Level1Out193[26] , \Level1Out193[25] , \Level1Out193[24] , 
        \Level1Out193[23] , \Level1Out193[22] , \Level1Out193[21] , 
        \Level1Out193[20] , \Level1Out193[19] , \Level1Out193[18] , 
        \Level1Out193[17] , \Level1Out193[16] , \Level1Out193[15] , 
        \Level1Out193[14] , \Level1Out193[13] , \Level1Out193[12] , 
        \Level1Out193[11] , \Level1Out193[10] , \Level1Out193[9] , 
        \Level1Out193[8] , \Level1Out193[7] , \Level1Out193[6] , 
        \Level1Out193[5] , \Level1Out193[4] , \Level1Out193[3] , 
        \Level1Out193[2] , \Level1Out193[1] , \Level1Out193[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_92_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load92[0] ), .Out({\Level2Out92[31] , \Level2Out92[30] , 
        \Level2Out92[29] , \Level2Out92[28] , \Level2Out92[27] , 
        \Level2Out92[26] , \Level2Out92[25] , \Level2Out92[24] , 
        \Level2Out92[23] , \Level2Out92[22] , \Level2Out92[21] , 
        \Level2Out92[20] , \Level2Out92[19] , \Level2Out92[18] , 
        \Level2Out92[17] , \Level2Out92[16] , \Level2Out92[15] , 
        \Level2Out92[14] , \Level2Out92[13] , \Level2Out92[12] , 
        \Level2Out92[11] , \Level2Out92[10] , \Level2Out92[9] , 
        \Level2Out92[8] , \Level2Out92[7] , \Level2Out92[6] , \Level2Out92[5] , 
        \Level2Out92[4] , \Level2Out92[3] , \Level2Out92[2] , \Level2Out92[1] , 
        \Level2Out92[0] }), .In1({\Level1Out92[31] , \Level1Out92[30] , 
        \Level1Out92[29] , \Level1Out92[28] , \Level1Out92[27] , 
        \Level1Out92[26] , \Level1Out92[25] , \Level1Out92[24] , 
        \Level1Out92[23] , \Level1Out92[22] , \Level1Out92[21] , 
        \Level1Out92[20] , \Level1Out92[19] , \Level1Out92[18] , 
        \Level1Out92[17] , \Level1Out92[16] , \Level1Out92[15] , 
        \Level1Out92[14] , \Level1Out92[13] , \Level1Out92[12] , 
        \Level1Out92[11] , \Level1Out92[10] , \Level1Out92[9] , 
        \Level1Out92[8] , \Level1Out92[7] , \Level1Out92[6] , \Level1Out92[5] , 
        \Level1Out92[4] , \Level1Out92[3] , \Level1Out92[2] , \Level1Out92[1] , 
        \Level1Out92[0] }), .In2({\Level1Out93[31] , \Level1Out93[30] , 
        \Level1Out93[29] , \Level1Out93[28] , \Level1Out93[27] , 
        \Level1Out93[26] , \Level1Out93[25] , \Level1Out93[24] , 
        \Level1Out93[23] , \Level1Out93[22] , \Level1Out93[21] , 
        \Level1Out93[20] , \Level1Out93[19] , \Level1Out93[18] , 
        \Level1Out93[17] , \Level1Out93[16] , \Level1Out93[15] , 
        \Level1Out93[14] , \Level1Out93[13] , \Level1Out93[12] , 
        \Level1Out93[11] , \Level1Out93[10] , \Level1Out93[9] , 
        \Level1Out93[8] , \Level1Out93[7] , \Level1Out93[6] , \Level1Out93[5] , 
        \Level1Out93[4] , \Level1Out93[3] , \Level1Out93[2] , \Level1Out93[1] , 
        \Level1Out93[0] }), .Read1(\Level1Load92[0] ), .Read2(
        \Level1Load93[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_228 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink228[31] , \ScanLink228[30] , 
        \ScanLink228[29] , \ScanLink228[28] , \ScanLink228[27] , 
        \ScanLink228[26] , \ScanLink228[25] , \ScanLink228[24] , 
        \ScanLink228[23] , \ScanLink228[22] , \ScanLink228[21] , 
        \ScanLink228[20] , \ScanLink228[19] , \ScanLink228[18] , 
        \ScanLink228[17] , \ScanLink228[16] , \ScanLink228[15] , 
        \ScanLink228[14] , \ScanLink228[13] , \ScanLink228[12] , 
        \ScanLink228[11] , \ScanLink228[10] , \ScanLink228[9] , 
        \ScanLink228[8] , \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , 
        \ScanLink228[4] , \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , 
        \ScanLink228[0] }), .ScanOut({\ScanLink229[31] , \ScanLink229[30] , 
        \ScanLink229[29] , \ScanLink229[28] , \ScanLink229[27] , 
        \ScanLink229[26] , \ScanLink229[25] , \ScanLink229[24] , 
        \ScanLink229[23] , \ScanLink229[22] , \ScanLink229[21] , 
        \ScanLink229[20] , \ScanLink229[19] , \ScanLink229[18] , 
        \ScanLink229[17] , \ScanLink229[16] , \ScanLink229[15] , 
        \ScanLink229[14] , \ScanLink229[13] , \ScanLink229[12] , 
        \ScanLink229[11] , \ScanLink229[10] , \ScanLink229[9] , 
        \ScanLink229[8] , \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , 
        \ScanLink229[4] , \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , 
        \ScanLink229[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load228[0] ), .Out({\Level1Out228[31] , \Level1Out228[30] , 
        \Level1Out228[29] , \Level1Out228[28] , \Level1Out228[27] , 
        \Level1Out228[26] , \Level1Out228[25] , \Level1Out228[24] , 
        \Level1Out228[23] , \Level1Out228[22] , \Level1Out228[21] , 
        \Level1Out228[20] , \Level1Out228[19] , \Level1Out228[18] , 
        \Level1Out228[17] , \Level1Out228[16] , \Level1Out228[15] , 
        \Level1Out228[14] , \Level1Out228[13] , \Level1Out228[12] , 
        \Level1Out228[11] , \Level1Out228[10] , \Level1Out228[9] , 
        \Level1Out228[8] , \Level1Out228[7] , \Level1Out228[6] , 
        \Level1Out228[5] , \Level1Out228[4] , \Level1Out228[3] , 
        \Level1Out228[2] , \Level1Out228[1] , \Level1Out228[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink1[31] , 
        \ScanLink1[30] , \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , 
        \ScanLink1[26] , \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , 
        \ScanLink1[22] , \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , 
        \ScanLink1[18] , \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , 
        \ScanLink1[14] , \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , 
        \ScanLink1[10] , \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , 
        \ScanLink1[6] , \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , 
        \ScanLink1[2] , \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load0[0] ), .Out({
        \Level1Out0[31] , \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , 
        \Level1Out0[27] , \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , 
        \Level1Out0[23] , \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , 
        \Level1Out0[19] , \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , 
        \Level1Out0[15] , \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , 
        \Level1Out0[11] , \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , 
        \Level1Out0[7] , \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , 
        \Level1Out0[3] , \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanOut({\ScanLink7[31] , 
        \ScanLink7[30] , \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , 
        \ScanLink7[26] , \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , 
        \ScanLink7[22] , \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , 
        \ScanLink7[18] , \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , 
        \ScanLink7[14] , \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , 
        \ScanLink7[10] , \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , 
        \ScanLink7[6] , \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , 
        \ScanLink7[2] , \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load6[0] ), .Out({
        \Level1Out6[31] , \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , 
        \Level1Out6[27] , \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , 
        \Level1Out6[23] , \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , 
        \Level1Out6[19] , \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , 
        \Level1Out6[15] , \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , 
        \Level1Out6[11] , \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , 
        \Level1Out6[7] , \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , 
        \Level1Out6[3] , \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanOut({\ScanLink9[31] , 
        \ScanLink9[30] , \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , 
        \ScanLink9[26] , \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , 
        \ScanLink9[22] , \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , 
        \ScanLink9[18] , \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , 
        \ScanLink9[14] , \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , 
        \ScanLink9[10] , \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , 
        \ScanLink9[6] , \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , 
        \ScanLink9[2] , \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load8[0] ), .Out({
        \Level1Out8[31] , \Level1Out8[30] , \Level1Out8[29] , \Level1Out8[28] , 
        \Level1Out8[27] , \Level1Out8[26] , \Level1Out8[25] , \Level1Out8[24] , 
        \Level1Out8[23] , \Level1Out8[22] , \Level1Out8[21] , \Level1Out8[20] , 
        \Level1Out8[19] , \Level1Out8[18] , \Level1Out8[17] , \Level1Out8[16] , 
        \Level1Out8[15] , \Level1Out8[14] , \Level1Out8[13] , \Level1Out8[12] , 
        \Level1Out8[11] , \Level1Out8[10] , \Level1Out8[9] , \Level1Out8[8] , 
        \Level1Out8[7] , \Level1Out8[6] , \Level1Out8[5] , \Level1Out8[4] , 
        \Level1Out8[3] , \Level1Out8[2] , \Level1Out8[1] , \Level1Out8[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_28 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanOut({\ScanLink29[31] , 
        \ScanLink29[30] , \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , 
        \ScanLink29[26] , \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , 
        \ScanLink29[22] , \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , 
        \ScanLink29[18] , \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , 
        \ScanLink29[14] , \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , 
        \ScanLink29[10] , \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , 
        \ScanLink29[6] , \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , 
        \ScanLink29[2] , \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load28[0] ), .Out({
        \Level1Out28[31] , \Level1Out28[30] , \Level1Out28[29] , 
        \Level1Out28[28] , \Level1Out28[27] , \Level1Out28[26] , 
        \Level1Out28[25] , \Level1Out28[24] , \Level1Out28[23] , 
        \Level1Out28[22] , \Level1Out28[21] , \Level1Out28[20] , 
        \Level1Out28[19] , \Level1Out28[18] , \Level1Out28[17] , 
        \Level1Out28[16] , \Level1Out28[15] , \Level1Out28[14] , 
        \Level1Out28[13] , \Level1Out28[12] , \Level1Out28[11] , 
        \Level1Out28[10] , \Level1Out28[9] , \Level1Out28[8] , 
        \Level1Out28[7] , \Level1Out28[6] , \Level1Out28[5] , \Level1Out28[4] , 
        \Level1Out28[3] , \Level1Out28[2] , \Level1Out28[1] , \Level1Out28[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_84 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink84[31] , \ScanLink84[30] , 
        \ScanLink84[29] , \ScanLink84[28] , \ScanLink84[27] , \ScanLink84[26] , 
        \ScanLink84[25] , \ScanLink84[24] , \ScanLink84[23] , \ScanLink84[22] , 
        \ScanLink84[21] , \ScanLink84[20] , \ScanLink84[19] , \ScanLink84[18] , 
        \ScanLink84[17] , \ScanLink84[16] , \ScanLink84[15] , \ScanLink84[14] , 
        \ScanLink84[13] , \ScanLink84[12] , \ScanLink84[11] , \ScanLink84[10] , 
        \ScanLink84[9] , \ScanLink84[8] , \ScanLink84[7] , \ScanLink84[6] , 
        \ScanLink84[5] , \ScanLink84[4] , \ScanLink84[3] , \ScanLink84[2] , 
        \ScanLink84[1] , \ScanLink84[0] }), .ScanOut({\ScanLink85[31] , 
        \ScanLink85[30] , \ScanLink85[29] , \ScanLink85[28] , \ScanLink85[27] , 
        \ScanLink85[26] , \ScanLink85[25] , \ScanLink85[24] , \ScanLink85[23] , 
        \ScanLink85[22] , \ScanLink85[21] , \ScanLink85[20] , \ScanLink85[19] , 
        \ScanLink85[18] , \ScanLink85[17] , \ScanLink85[16] , \ScanLink85[15] , 
        \ScanLink85[14] , \ScanLink85[13] , \ScanLink85[12] , \ScanLink85[11] , 
        \ScanLink85[10] , \ScanLink85[9] , \ScanLink85[8] , \ScanLink85[7] , 
        \ScanLink85[6] , \ScanLink85[5] , \ScanLink85[4] , \ScanLink85[3] , 
        \ScanLink85[2] , \ScanLink85[1] , \ScanLink85[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load84[0] ), .Out({
        \Level1Out84[31] , \Level1Out84[30] , \Level1Out84[29] , 
        \Level1Out84[28] , \Level1Out84[27] , \Level1Out84[26] , 
        \Level1Out84[25] , \Level1Out84[24] , \Level1Out84[23] , 
        \Level1Out84[22] , \Level1Out84[21] , \Level1Out84[20] , 
        \Level1Out84[19] , \Level1Out84[18] , \Level1Out84[17] , 
        \Level1Out84[16] , \Level1Out84[15] , \Level1Out84[14] , 
        \Level1Out84[13] , \Level1Out84[12] , \Level1Out84[11] , 
        \Level1Out84[10] , \Level1Out84[9] , \Level1Out84[8] , 
        \Level1Out84[7] , \Level1Out84[6] , \Level1Out84[5] , \Level1Out84[4] , 
        \Level1Out84[3] , \Level1Out84[2] , \Level1Out84[1] , \Level1Out84[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_184_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load184[0] ), .Out({\Level2Out184[31] , \Level2Out184[30] , 
        \Level2Out184[29] , \Level2Out184[28] , \Level2Out184[27] , 
        \Level2Out184[26] , \Level2Out184[25] , \Level2Out184[24] , 
        \Level2Out184[23] , \Level2Out184[22] , \Level2Out184[21] , 
        \Level2Out184[20] , \Level2Out184[19] , \Level2Out184[18] , 
        \Level2Out184[17] , \Level2Out184[16] , \Level2Out184[15] , 
        \Level2Out184[14] , \Level2Out184[13] , \Level2Out184[12] , 
        \Level2Out184[11] , \Level2Out184[10] , \Level2Out184[9] , 
        \Level2Out184[8] , \Level2Out184[7] , \Level2Out184[6] , 
        \Level2Out184[5] , \Level2Out184[4] , \Level2Out184[3] , 
        \Level2Out184[2] , \Level2Out184[1] , \Level2Out184[0] }), .In1({
        \Level1Out184[31] , \Level1Out184[30] , \Level1Out184[29] , 
        \Level1Out184[28] , \Level1Out184[27] , \Level1Out184[26] , 
        \Level1Out184[25] , \Level1Out184[24] , \Level1Out184[23] , 
        \Level1Out184[22] , \Level1Out184[21] , \Level1Out184[20] , 
        \Level1Out184[19] , \Level1Out184[18] , \Level1Out184[17] , 
        \Level1Out184[16] , \Level1Out184[15] , \Level1Out184[14] , 
        \Level1Out184[13] , \Level1Out184[12] , \Level1Out184[11] , 
        \Level1Out184[10] , \Level1Out184[9] , \Level1Out184[8] , 
        \Level1Out184[7] , \Level1Out184[6] , \Level1Out184[5] , 
        \Level1Out184[4] , \Level1Out184[3] , \Level1Out184[2] , 
        \Level1Out184[1] , \Level1Out184[0] }), .In2({\Level1Out185[31] , 
        \Level1Out185[30] , \Level1Out185[29] , \Level1Out185[28] , 
        \Level1Out185[27] , \Level1Out185[26] , \Level1Out185[25] , 
        \Level1Out185[24] , \Level1Out185[23] , \Level1Out185[22] , 
        \Level1Out185[21] , \Level1Out185[20] , \Level1Out185[19] , 
        \Level1Out185[18] , \Level1Out185[17] , \Level1Out185[16] , 
        \Level1Out185[15] , \Level1Out185[14] , \Level1Out185[13] , 
        \Level1Out185[12] , \Level1Out185[11] , \Level1Out185[10] , 
        \Level1Out185[9] , \Level1Out185[8] , \Level1Out185[7] , 
        \Level1Out185[6] , \Level1Out185[5] , \Level1Out185[4] , 
        \Level1Out185[3] , \Level1Out185[2] , \Level1Out185[1] , 
        \Level1Out185[0] }), .Read1(\Level1Load184[0] ), .Read2(
        \Level1Load185[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load48[0] ), .Out({\Level4Out48[31] , \Level4Out48[30] , 
        \Level4Out48[29] , \Level4Out48[28] , \Level4Out48[27] , 
        \Level4Out48[26] , \Level4Out48[25] , \Level4Out48[24] , 
        \Level4Out48[23] , \Level4Out48[22] , \Level4Out48[21] , 
        \Level4Out48[20] , \Level4Out48[19] , \Level4Out48[18] , 
        \Level4Out48[17] , \Level4Out48[16] , \Level4Out48[15] , 
        \Level4Out48[14] , \Level4Out48[13] , \Level4Out48[12] , 
        \Level4Out48[11] , \Level4Out48[10] , \Level4Out48[9] , 
        \Level4Out48[8] , \Level4Out48[7] , \Level4Out48[6] , \Level4Out48[5] , 
        \Level4Out48[4] , \Level4Out48[3] , \Level4Out48[2] , \Level4Out48[1] , 
        \Level4Out48[0] }), .In1({\Level2Out48[31] , \Level2Out48[30] , 
        \Level2Out48[29] , \Level2Out48[28] , \Level2Out48[27] , 
        \Level2Out48[26] , \Level2Out48[25] , \Level2Out48[24] , 
        \Level2Out48[23] , \Level2Out48[22] , \Level2Out48[21] , 
        \Level2Out48[20] , \Level2Out48[19] , \Level2Out48[18] , 
        \Level2Out48[17] , \Level2Out48[16] , \Level2Out48[15] , 
        \Level2Out48[14] , \Level2Out48[13] , \Level2Out48[12] , 
        \Level2Out48[11] , \Level2Out48[10] , \Level2Out48[9] , 
        \Level2Out48[8] , \Level2Out48[7] , \Level2Out48[6] , \Level2Out48[5] , 
        \Level2Out48[4] , \Level2Out48[3] , \Level2Out48[2] , \Level2Out48[1] , 
        \Level2Out48[0] }), .In2({\Level2Out50[31] , \Level2Out50[30] , 
        \Level2Out50[29] , \Level2Out50[28] , \Level2Out50[27] , 
        \Level2Out50[26] , \Level2Out50[25] , \Level2Out50[24] , 
        \Level2Out50[23] , \Level2Out50[22] , \Level2Out50[21] , 
        \Level2Out50[20] , \Level2Out50[19] , \Level2Out50[18] , 
        \Level2Out50[17] , \Level2Out50[16] , \Level2Out50[15] , 
        \Level2Out50[14] , \Level2Out50[13] , \Level2Out50[12] , 
        \Level2Out50[11] , \Level2Out50[10] , \Level2Out50[9] , 
        \Level2Out50[8] , \Level2Out50[7] , \Level2Out50[6] , \Level2Out50[5] , 
        \Level2Out50[4] , \Level2Out50[3] , \Level2Out50[2] , \Level2Out50[1] , 
        \Level2Out50[0] }), .Read1(\Level2Load48[0] ), .Read2(
        \Level2Load50[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_46 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanOut({\ScanLink47[31] , 
        \ScanLink47[30] , \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , 
        \ScanLink47[26] , \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , 
        \ScanLink47[22] , \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , 
        \ScanLink47[18] , \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , 
        \ScanLink47[14] , \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , 
        \ScanLink47[10] , \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , 
        \ScanLink47[6] , \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , 
        \ScanLink47[2] , \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load46[0] ), .Out({
        \Level1Out46[31] , \Level1Out46[30] , \Level1Out46[29] , 
        \Level1Out46[28] , \Level1Out46[27] , \Level1Out46[26] , 
        \Level1Out46[25] , \Level1Out46[24] , \Level1Out46[23] , 
        \Level1Out46[22] , \Level1Out46[21] , \Level1Out46[20] , 
        \Level1Out46[19] , \Level1Out46[18] , \Level1Out46[17] , 
        \Level1Out46[16] , \Level1Out46[15] , \Level1Out46[14] , 
        \Level1Out46[13] , \Level1Out46[12] , \Level1Out46[11] , 
        \Level1Out46[10] , \Level1Out46[9] , \Level1Out46[8] , 
        \Level1Out46[7] , \Level1Out46[6] , \Level1Out46[5] , \Level1Out46[4] , 
        \Level1Out46[3] , \Level1Out46[2] , \Level1Out46[1] , \Level1Out46[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_61 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanOut({\ScanLink62[31] , 
        \ScanLink62[30] , \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , 
        \ScanLink62[26] , \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , 
        \ScanLink62[22] , \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , 
        \ScanLink62[18] , \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , 
        \ScanLink62[14] , \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , 
        \ScanLink62[10] , \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , 
        \ScanLink62[6] , \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , 
        \ScanLink62[2] , \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load61[0] ), .Out({
        \Level1Out61[31] , \Level1Out61[30] , \Level1Out61[29] , 
        \Level1Out61[28] , \Level1Out61[27] , \Level1Out61[26] , 
        \Level1Out61[25] , \Level1Out61[24] , \Level1Out61[23] , 
        \Level1Out61[22] , \Level1Out61[21] , \Level1Out61[20] , 
        \Level1Out61[19] , \Level1Out61[18] , \Level1Out61[17] , 
        \Level1Out61[16] , \Level1Out61[15] , \Level1Out61[14] , 
        \Level1Out61[13] , \Level1Out61[12] , \Level1Out61[11] , 
        \Level1Out61[10] , \Level1Out61[9] , \Level1Out61[8] , 
        \Level1Out61[7] , \Level1Out61[6] , \Level1Out61[5] , \Level1Out61[4] , 
        \Level1Out61[3] , \Level1Out61[2] , \Level1Out61[1] , \Level1Out61[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_181 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink181[31] , \ScanLink181[30] , 
        \ScanLink181[29] , \ScanLink181[28] , \ScanLink181[27] , 
        \ScanLink181[26] , \ScanLink181[25] , \ScanLink181[24] , 
        \ScanLink181[23] , \ScanLink181[22] , \ScanLink181[21] , 
        \ScanLink181[20] , \ScanLink181[19] , \ScanLink181[18] , 
        \ScanLink181[17] , \ScanLink181[16] , \ScanLink181[15] , 
        \ScanLink181[14] , \ScanLink181[13] , \ScanLink181[12] , 
        \ScanLink181[11] , \ScanLink181[10] , \ScanLink181[9] , 
        \ScanLink181[8] , \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , 
        \ScanLink181[4] , \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , 
        \ScanLink181[0] }), .ScanOut({\ScanLink182[31] , \ScanLink182[30] , 
        \ScanLink182[29] , \ScanLink182[28] , \ScanLink182[27] , 
        \ScanLink182[26] , \ScanLink182[25] , \ScanLink182[24] , 
        \ScanLink182[23] , \ScanLink182[22] , \ScanLink182[21] , 
        \ScanLink182[20] , \ScanLink182[19] , \ScanLink182[18] , 
        \ScanLink182[17] , \ScanLink182[16] , \ScanLink182[15] , 
        \ScanLink182[14] , \ScanLink182[13] , \ScanLink182[12] , 
        \ScanLink182[11] , \ScanLink182[10] , \ScanLink182[9] , 
        \ScanLink182[8] , \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , 
        \ScanLink182[4] , \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , 
        \ScanLink182[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load181[0] ), .Out({\Level1Out181[31] , \Level1Out181[30] , 
        \Level1Out181[29] , \Level1Out181[28] , \Level1Out181[27] , 
        \Level1Out181[26] , \Level1Out181[25] , \Level1Out181[24] , 
        \Level1Out181[23] , \Level1Out181[22] , \Level1Out181[21] , 
        \Level1Out181[20] , \Level1Out181[19] , \Level1Out181[18] , 
        \Level1Out181[17] , \Level1Out181[16] , \Level1Out181[15] , 
        \Level1Out181[14] , \Level1Out181[13] , \Level1Out181[12] , 
        \Level1Out181[11] , \Level1Out181[10] , \Level1Out181[9] , 
        \Level1Out181[8] , \Level1Out181[7] , \Level1Out181[6] , 
        \Level1Out181[5] , \Level1Out181[4] , \Level1Out181[3] , 
        \Level1Out181[2] , \Level1Out181[1] , \Level1Out181[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_54_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load54[0] ), .Out({\Level2Out54[31] , \Level2Out54[30] , 
        \Level2Out54[29] , \Level2Out54[28] , \Level2Out54[27] , 
        \Level2Out54[26] , \Level2Out54[25] , \Level2Out54[24] , 
        \Level2Out54[23] , \Level2Out54[22] , \Level2Out54[21] , 
        \Level2Out54[20] , \Level2Out54[19] , \Level2Out54[18] , 
        \Level2Out54[17] , \Level2Out54[16] , \Level2Out54[15] , 
        \Level2Out54[14] , \Level2Out54[13] , \Level2Out54[12] , 
        \Level2Out54[11] , \Level2Out54[10] , \Level2Out54[9] , 
        \Level2Out54[8] , \Level2Out54[7] , \Level2Out54[6] , \Level2Out54[5] , 
        \Level2Out54[4] , \Level2Out54[3] , \Level2Out54[2] , \Level2Out54[1] , 
        \Level2Out54[0] }), .In1({\Level1Out54[31] , \Level1Out54[30] , 
        \Level1Out54[29] , \Level1Out54[28] , \Level1Out54[27] , 
        \Level1Out54[26] , \Level1Out54[25] , \Level1Out54[24] , 
        \Level1Out54[23] , \Level1Out54[22] , \Level1Out54[21] , 
        \Level1Out54[20] , \Level1Out54[19] , \Level1Out54[18] , 
        \Level1Out54[17] , \Level1Out54[16] , \Level1Out54[15] , 
        \Level1Out54[14] , \Level1Out54[13] , \Level1Out54[12] , 
        \Level1Out54[11] , \Level1Out54[10] , \Level1Out54[9] , 
        \Level1Out54[8] , \Level1Out54[7] , \Level1Out54[6] , \Level1Out54[5] , 
        \Level1Out54[4] , \Level1Out54[3] , \Level1Out54[2] , \Level1Out54[1] , 
        \Level1Out54[0] }), .In2({\Level1Out55[31] , \Level1Out55[30] , 
        \Level1Out55[29] , \Level1Out55[28] , \Level1Out55[27] , 
        \Level1Out55[26] , \Level1Out55[25] , \Level1Out55[24] , 
        \Level1Out55[23] , \Level1Out55[22] , \Level1Out55[21] , 
        \Level1Out55[20] , \Level1Out55[19] , \Level1Out55[18] , 
        \Level1Out55[17] , \Level1Out55[16] , \Level1Out55[15] , 
        \Level1Out55[14] , \Level1Out55[13] , \Level1Out55[12] , 
        \Level1Out55[11] , \Level1Out55[10] , \Level1Out55[9] , 
        \Level1Out55[8] , \Level1Out55[7] , \Level1Out55[6] , \Level1Out55[5] , 
        \Level1Out55[4] , \Level1Out55[3] , \Level1Out55[2] , \Level1Out55[1] , 
        \Level1Out55[0] }), .Read1(\Level1Load54[0] ), .Read2(
        \Level1Load55[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_112_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load112[0] ), .Out({\Level2Out112[31] , \Level2Out112[30] , 
        \Level2Out112[29] , \Level2Out112[28] , \Level2Out112[27] , 
        \Level2Out112[26] , \Level2Out112[25] , \Level2Out112[24] , 
        \Level2Out112[23] , \Level2Out112[22] , \Level2Out112[21] , 
        \Level2Out112[20] , \Level2Out112[19] , \Level2Out112[18] , 
        \Level2Out112[17] , \Level2Out112[16] , \Level2Out112[15] , 
        \Level2Out112[14] , \Level2Out112[13] , \Level2Out112[12] , 
        \Level2Out112[11] , \Level2Out112[10] , \Level2Out112[9] , 
        \Level2Out112[8] , \Level2Out112[7] , \Level2Out112[6] , 
        \Level2Out112[5] , \Level2Out112[4] , \Level2Out112[3] , 
        \Level2Out112[2] , \Level2Out112[1] , \Level2Out112[0] }), .In1({
        \Level1Out112[31] , \Level1Out112[30] , \Level1Out112[29] , 
        \Level1Out112[28] , \Level1Out112[27] , \Level1Out112[26] , 
        \Level1Out112[25] , \Level1Out112[24] , \Level1Out112[23] , 
        \Level1Out112[22] , \Level1Out112[21] , \Level1Out112[20] , 
        \Level1Out112[19] , \Level1Out112[18] , \Level1Out112[17] , 
        \Level1Out112[16] , \Level1Out112[15] , \Level1Out112[14] , 
        \Level1Out112[13] , \Level1Out112[12] , \Level1Out112[11] , 
        \Level1Out112[10] , \Level1Out112[9] , \Level1Out112[8] , 
        \Level1Out112[7] , \Level1Out112[6] , \Level1Out112[5] , 
        \Level1Out112[4] , \Level1Out112[3] , \Level1Out112[2] , 
        \Level1Out112[1] , \Level1Out112[0] }), .In2({\Level1Out113[31] , 
        \Level1Out113[30] , \Level1Out113[29] , \Level1Out113[28] , 
        \Level1Out113[27] , \Level1Out113[26] , \Level1Out113[25] , 
        \Level1Out113[24] , \Level1Out113[23] , \Level1Out113[22] , 
        \Level1Out113[21] , \Level1Out113[20] , \Level1Out113[19] , 
        \Level1Out113[18] , \Level1Out113[17] , \Level1Out113[16] , 
        \Level1Out113[15] , \Level1Out113[14] , \Level1Out113[13] , 
        \Level1Out113[12] , \Level1Out113[11] , \Level1Out113[10] , 
        \Level1Out113[9] , \Level1Out113[8] , \Level1Out113[7] , 
        \Level1Out113[6] , \Level1Out113[5] , \Level1Out113[4] , 
        \Level1Out113[3] , \Level1Out113[2] , \Level1Out113[1] , 
        \Level1Out113[0] }), .Read1(\Level1Load112[0] ), .Read2(
        \Level1Load113[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_138_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load138[0] ), .Out({\Level2Out138[31] , \Level2Out138[30] , 
        \Level2Out138[29] , \Level2Out138[28] , \Level2Out138[27] , 
        \Level2Out138[26] , \Level2Out138[25] , \Level2Out138[24] , 
        \Level2Out138[23] , \Level2Out138[22] , \Level2Out138[21] , 
        \Level2Out138[20] , \Level2Out138[19] , \Level2Out138[18] , 
        \Level2Out138[17] , \Level2Out138[16] , \Level2Out138[15] , 
        \Level2Out138[14] , \Level2Out138[13] , \Level2Out138[12] , 
        \Level2Out138[11] , \Level2Out138[10] , \Level2Out138[9] , 
        \Level2Out138[8] , \Level2Out138[7] , \Level2Out138[6] , 
        \Level2Out138[5] , \Level2Out138[4] , \Level2Out138[3] , 
        \Level2Out138[2] , \Level2Out138[1] , \Level2Out138[0] }), .In1({
        \Level1Out138[31] , \Level1Out138[30] , \Level1Out138[29] , 
        \Level1Out138[28] , \Level1Out138[27] , \Level1Out138[26] , 
        \Level1Out138[25] , \Level1Out138[24] , \Level1Out138[23] , 
        \Level1Out138[22] , \Level1Out138[21] , \Level1Out138[20] , 
        \Level1Out138[19] , \Level1Out138[18] , \Level1Out138[17] , 
        \Level1Out138[16] , \Level1Out138[15] , \Level1Out138[14] , 
        \Level1Out138[13] , \Level1Out138[12] , \Level1Out138[11] , 
        \Level1Out138[10] , \Level1Out138[9] , \Level1Out138[8] , 
        \Level1Out138[7] , \Level1Out138[6] , \Level1Out138[5] , 
        \Level1Out138[4] , \Level1Out138[3] , \Level1Out138[2] , 
        \Level1Out138[1] , \Level1Out138[0] }), .In2({\Level1Out139[31] , 
        \Level1Out139[30] , \Level1Out139[29] , \Level1Out139[28] , 
        \Level1Out139[27] , \Level1Out139[26] , \Level1Out139[25] , 
        \Level1Out139[24] , \Level1Out139[23] , \Level1Out139[22] , 
        \Level1Out139[21] , \Level1Out139[20] , \Level1Out139[19] , 
        \Level1Out139[18] , \Level1Out139[17] , \Level1Out139[16] , 
        \Level1Out139[15] , \Level1Out139[14] , \Level1Out139[13] , 
        \Level1Out139[12] , \Level1Out139[11] , \Level1Out139[10] , 
        \Level1Out139[9] , \Level1Out139[8] , \Level1Out139[7] , 
        \Level1Out139[6] , \Level1Out139[5] , \Level1Out139[4] , 
        \Level1Out139[3] , \Level1Out139[2] , \Level1Out139[1] , 
        \Level1Out139[0] }), .Read1(\Level1Load138[0] ), .Read2(
        \Level1Load139[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_226_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load226[0] ), .Out({\Level2Out226[31] , \Level2Out226[30] , 
        \Level2Out226[29] , \Level2Out226[28] , \Level2Out226[27] , 
        \Level2Out226[26] , \Level2Out226[25] , \Level2Out226[24] , 
        \Level2Out226[23] , \Level2Out226[22] , \Level2Out226[21] , 
        \Level2Out226[20] , \Level2Out226[19] , \Level2Out226[18] , 
        \Level2Out226[17] , \Level2Out226[16] , \Level2Out226[15] , 
        \Level2Out226[14] , \Level2Out226[13] , \Level2Out226[12] , 
        \Level2Out226[11] , \Level2Out226[10] , \Level2Out226[9] , 
        \Level2Out226[8] , \Level2Out226[7] , \Level2Out226[6] , 
        \Level2Out226[5] , \Level2Out226[4] , \Level2Out226[3] , 
        \Level2Out226[2] , \Level2Out226[1] , \Level2Out226[0] }), .In1({
        \Level1Out226[31] , \Level1Out226[30] , \Level1Out226[29] , 
        \Level1Out226[28] , \Level1Out226[27] , \Level1Out226[26] , 
        \Level1Out226[25] , \Level1Out226[24] , \Level1Out226[23] , 
        \Level1Out226[22] , \Level1Out226[21] , \Level1Out226[20] , 
        \Level1Out226[19] , \Level1Out226[18] , \Level1Out226[17] , 
        \Level1Out226[16] , \Level1Out226[15] , \Level1Out226[14] , 
        \Level1Out226[13] , \Level1Out226[12] , \Level1Out226[11] , 
        \Level1Out226[10] , \Level1Out226[9] , \Level1Out226[8] , 
        \Level1Out226[7] , \Level1Out226[6] , \Level1Out226[5] , 
        \Level1Out226[4] , \Level1Out226[3] , \Level1Out226[2] , 
        \Level1Out226[1] , \Level1Out226[0] }), .In2({\Level1Out227[31] , 
        \Level1Out227[30] , \Level1Out227[29] , \Level1Out227[28] , 
        \Level1Out227[27] , \Level1Out227[26] , \Level1Out227[25] , 
        \Level1Out227[24] , \Level1Out227[23] , \Level1Out227[22] , 
        \Level1Out227[21] , \Level1Out227[20] , \Level1Out227[19] , 
        \Level1Out227[18] , \Level1Out227[17] , \Level1Out227[16] , 
        \Level1Out227[15] , \Level1Out227[14] , \Level1Out227[13] , 
        \Level1Out227[12] , \Level1Out227[11] , \Level1Out227[10] , 
        \Level1Out227[9] , \Level1Out227[8] , \Level1Out227[7] , 
        \Level1Out227[6] , \Level1Out227[5] , \Level1Out227[4] , 
        \Level1Out227[3] , \Level1Out227[2] , \Level1Out227[1] , 
        \Level1Out227[0] }), .Read1(\Level1Load226[0] ), .Read2(
        \Level1Load227[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_124_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load124[0] ), .Out({\Level4Out124[31] , \Level4Out124[30] , 
        \Level4Out124[29] , \Level4Out124[28] , \Level4Out124[27] , 
        \Level4Out124[26] , \Level4Out124[25] , \Level4Out124[24] , 
        \Level4Out124[23] , \Level4Out124[22] , \Level4Out124[21] , 
        \Level4Out124[20] , \Level4Out124[19] , \Level4Out124[18] , 
        \Level4Out124[17] , \Level4Out124[16] , \Level4Out124[15] , 
        \Level4Out124[14] , \Level4Out124[13] , \Level4Out124[12] , 
        \Level4Out124[11] , \Level4Out124[10] , \Level4Out124[9] , 
        \Level4Out124[8] , \Level4Out124[7] , \Level4Out124[6] , 
        \Level4Out124[5] , \Level4Out124[4] , \Level4Out124[3] , 
        \Level4Out124[2] , \Level4Out124[1] , \Level4Out124[0] }), .In1({
        \Level2Out124[31] , \Level2Out124[30] , \Level2Out124[29] , 
        \Level2Out124[28] , \Level2Out124[27] , \Level2Out124[26] , 
        \Level2Out124[25] , \Level2Out124[24] , \Level2Out124[23] , 
        \Level2Out124[22] , \Level2Out124[21] , \Level2Out124[20] , 
        \Level2Out124[19] , \Level2Out124[18] , \Level2Out124[17] , 
        \Level2Out124[16] , \Level2Out124[15] , \Level2Out124[14] , 
        \Level2Out124[13] , \Level2Out124[12] , \Level2Out124[11] , 
        \Level2Out124[10] , \Level2Out124[9] , \Level2Out124[8] , 
        \Level2Out124[7] , \Level2Out124[6] , \Level2Out124[5] , 
        \Level2Out124[4] , \Level2Out124[3] , \Level2Out124[2] , 
        \Level2Out124[1] , \Level2Out124[0] }), .In2({\Level2Out126[31] , 
        \Level2Out126[30] , \Level2Out126[29] , \Level2Out126[28] , 
        \Level2Out126[27] , \Level2Out126[26] , \Level2Out126[25] , 
        \Level2Out126[24] , \Level2Out126[23] , \Level2Out126[22] , 
        \Level2Out126[21] , \Level2Out126[20] , \Level2Out126[19] , 
        \Level2Out126[18] , \Level2Out126[17] , \Level2Out126[16] , 
        \Level2Out126[15] , \Level2Out126[14] , \Level2Out126[13] , 
        \Level2Out126[12] , \Level2Out126[11] , \Level2Out126[10] , 
        \Level2Out126[9] , \Level2Out126[8] , \Level2Out126[7] , 
        \Level2Out126[6] , \Level2Out126[5] , \Level2Out126[4] , 
        \Level2Out126[3] , \Level2Out126[2] , \Level2Out126[1] , 
        \Level2Out126[0] }), .Read1(\Level2Load124[0] ), .Read2(
        \Level2Load126[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load64[0] ), .Out({\Level32Out64[31] , \Level32Out64[30] , 
        \Level32Out64[29] , \Level32Out64[28] , \Level32Out64[27] , 
        \Level32Out64[26] , \Level32Out64[25] , \Level32Out64[24] , 
        \Level32Out64[23] , \Level32Out64[22] , \Level32Out64[21] , 
        \Level32Out64[20] , \Level32Out64[19] , \Level32Out64[18] , 
        \Level32Out64[17] , \Level32Out64[16] , \Level32Out64[15] , 
        \Level32Out64[14] , \Level32Out64[13] , \Level32Out64[12] , 
        \Level32Out64[11] , \Level32Out64[10] , \Level32Out64[9] , 
        \Level32Out64[8] , \Level32Out64[7] , \Level32Out64[6] , 
        \Level32Out64[5] , \Level32Out64[4] , \Level32Out64[3] , 
        \Level32Out64[2] , \Level32Out64[1] , \Level32Out64[0] }), .In1({
        \Level16Out64[31] , \Level16Out64[30] , \Level16Out64[29] , 
        \Level16Out64[28] , \Level16Out64[27] , \Level16Out64[26] , 
        \Level16Out64[25] , \Level16Out64[24] , \Level16Out64[23] , 
        \Level16Out64[22] , \Level16Out64[21] , \Level16Out64[20] , 
        \Level16Out64[19] , \Level16Out64[18] , \Level16Out64[17] , 
        \Level16Out64[16] , \Level16Out64[15] , \Level16Out64[14] , 
        \Level16Out64[13] , \Level16Out64[12] , \Level16Out64[11] , 
        \Level16Out64[10] , \Level16Out64[9] , \Level16Out64[8] , 
        \Level16Out64[7] , \Level16Out64[6] , \Level16Out64[5] , 
        \Level16Out64[4] , \Level16Out64[3] , \Level16Out64[2] , 
        \Level16Out64[1] , \Level16Out64[0] }), .In2({\Level16Out80[31] , 
        \Level16Out80[30] , \Level16Out80[29] , \Level16Out80[28] , 
        \Level16Out80[27] , \Level16Out80[26] , \Level16Out80[25] , 
        \Level16Out80[24] , \Level16Out80[23] , \Level16Out80[22] , 
        \Level16Out80[21] , \Level16Out80[20] , \Level16Out80[19] , 
        \Level16Out80[18] , \Level16Out80[17] , \Level16Out80[16] , 
        \Level16Out80[15] , \Level16Out80[14] , \Level16Out80[13] , 
        \Level16Out80[12] , \Level16Out80[11] , \Level16Out80[10] , 
        \Level16Out80[9] , \Level16Out80[8] , \Level16Out80[7] , 
        \Level16Out80[6] , \Level16Out80[5] , \Level16Out80[4] , 
        \Level16Out80[3] , \Level16Out80[2] , \Level16Out80[1] , 
        \Level16Out80[0] }), .Read1(\Level16Load64[0] ), .Read2(
        \Level16Load80[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_254 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink254[31] , \ScanLink254[30] , 
        \ScanLink254[29] , \ScanLink254[28] , \ScanLink254[27] , 
        \ScanLink254[26] , \ScanLink254[25] , \ScanLink254[24] , 
        \ScanLink254[23] , \ScanLink254[22] , \ScanLink254[21] , 
        \ScanLink254[20] , \ScanLink254[19] , \ScanLink254[18] , 
        \ScanLink254[17] , \ScanLink254[16] , \ScanLink254[15] , 
        \ScanLink254[14] , \ScanLink254[13] , \ScanLink254[12] , 
        \ScanLink254[11] , \ScanLink254[10] , \ScanLink254[9] , 
        \ScanLink254[8] , \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , 
        \ScanLink254[4] , \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , 
        \ScanLink254[0] }), .ScanOut({\ScanLink255[31] , \ScanLink255[30] , 
        \ScanLink255[29] , \ScanLink255[28] , \ScanLink255[27] , 
        \ScanLink255[26] , \ScanLink255[25] , \ScanLink255[24] , 
        \ScanLink255[23] , \ScanLink255[22] , \ScanLink255[21] , 
        \ScanLink255[20] , \ScanLink255[19] , \ScanLink255[18] , 
        \ScanLink255[17] , \ScanLink255[16] , \ScanLink255[15] , 
        \ScanLink255[14] , \ScanLink255[13] , \ScanLink255[12] , 
        \ScanLink255[11] , \ScanLink255[10] , \ScanLink255[9] , 
        \ScanLink255[8] , \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , 
        \ScanLink255[4] , \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , 
        \ScanLink255[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load254[0] ), .Out({\Level1Out254[31] , \Level1Out254[30] , 
        \Level1Out254[29] , \Level1Out254[28] , \Level1Out254[27] , 
        \Level1Out254[26] , \Level1Out254[25] , \Level1Out254[24] , 
        \Level1Out254[23] , \Level1Out254[22] , \Level1Out254[21] , 
        \Level1Out254[20] , \Level1Out254[19] , \Level1Out254[18] , 
        \Level1Out254[17] , \Level1Out254[16] , \Level1Out254[15] , 
        \Level1Out254[14] , \Level1Out254[13] , \Level1Out254[12] , 
        \Level1Out254[11] , \Level1Out254[10] , \Level1Out254[9] , 
        \Level1Out254[8] , \Level1Out254[7] , \Level1Out254[6] , 
        \Level1Out254[5] , \Level1Out254[4] , \Level1Out254[3] , 
        \Level1Out254[2] , \Level1Out254[1] , \Level1Out254[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanOut({\ScanLink14[31] , 
        \ScanLink14[30] , \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , 
        \ScanLink14[26] , \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , 
        \ScanLink14[22] , \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , 
        \ScanLink14[18] , \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , 
        \ScanLink14[14] , \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , 
        \ScanLink14[10] , \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , 
        \ScanLink14[6] , \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , 
        \ScanLink14[2] , \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load13[0] ), .Out({
        \Level1Out13[31] , \Level1Out13[30] , \Level1Out13[29] , 
        \Level1Out13[28] , \Level1Out13[27] , \Level1Out13[26] , 
        \Level1Out13[25] , \Level1Out13[24] , \Level1Out13[23] , 
        \Level1Out13[22] , \Level1Out13[21] , \Level1Out13[20] , 
        \Level1Out13[19] , \Level1Out13[18] , \Level1Out13[17] , 
        \Level1Out13[16] , \Level1Out13[15] , \Level1Out13[14] , 
        \Level1Out13[13] , \Level1Out13[12] , \Level1Out13[11] , 
        \Level1Out13[10] , \Level1Out13[9] , \Level1Out13[8] , 
        \Level1Out13[7] , \Level1Out13[6] , \Level1Out13[5] , \Level1Out13[4] , 
        \Level1Out13[3] , \Level1Out13[2] , \Level1Out13[1] , \Level1Out13[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanOut({\ScanLink15[31] , 
        \ScanLink15[30] , \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , 
        \ScanLink15[26] , \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , 
        \ScanLink15[22] , \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , 
        \ScanLink15[18] , \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , 
        \ScanLink15[14] , \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , 
        \ScanLink15[10] , \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , 
        \ScanLink15[6] , \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , 
        \ScanLink15[2] , \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load14[0] ), .Out({
        \Level1Out14[31] , \Level1Out14[30] , \Level1Out14[29] , 
        \Level1Out14[28] , \Level1Out14[27] , \Level1Out14[26] , 
        \Level1Out14[25] , \Level1Out14[24] , \Level1Out14[23] , 
        \Level1Out14[22] , \Level1Out14[21] , \Level1Out14[20] , 
        \Level1Out14[19] , \Level1Out14[18] , \Level1Out14[17] , 
        \Level1Out14[16] , \Level1Out14[15] , \Level1Out14[14] , 
        \Level1Out14[13] , \Level1Out14[12] , \Level1Out14[11] , 
        \Level1Out14[10] , \Level1Out14[9] , \Level1Out14[8] , 
        \Level1Out14[7] , \Level1Out14[6] , \Level1Out14[5] , \Level1Out14[4] , 
        \Level1Out14[3] , \Level1Out14[2] , \Level1Out14[1] , \Level1Out14[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_143 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink143[31] , \ScanLink143[30] , 
        \ScanLink143[29] , \ScanLink143[28] , \ScanLink143[27] , 
        \ScanLink143[26] , \ScanLink143[25] , \ScanLink143[24] , 
        \ScanLink143[23] , \ScanLink143[22] , \ScanLink143[21] , 
        \ScanLink143[20] , \ScanLink143[19] , \ScanLink143[18] , 
        \ScanLink143[17] , \ScanLink143[16] , \ScanLink143[15] , 
        \ScanLink143[14] , \ScanLink143[13] , \ScanLink143[12] , 
        \ScanLink143[11] , \ScanLink143[10] , \ScanLink143[9] , 
        \ScanLink143[8] , \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , 
        \ScanLink143[4] , \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , 
        \ScanLink143[0] }), .ScanOut({\ScanLink144[31] , \ScanLink144[30] , 
        \ScanLink144[29] , \ScanLink144[28] , \ScanLink144[27] , 
        \ScanLink144[26] , \ScanLink144[25] , \ScanLink144[24] , 
        \ScanLink144[23] , \ScanLink144[22] , \ScanLink144[21] , 
        \ScanLink144[20] , \ScanLink144[19] , \ScanLink144[18] , 
        \ScanLink144[17] , \ScanLink144[16] , \ScanLink144[15] , 
        \ScanLink144[14] , \ScanLink144[13] , \ScanLink144[12] , 
        \ScanLink144[11] , \ScanLink144[10] , \ScanLink144[9] , 
        \ScanLink144[8] , \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , 
        \ScanLink144[4] , \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , 
        \ScanLink144[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load143[0] ), .Out({\Level1Out143[31] , \Level1Out143[30] , 
        \Level1Out143[29] , \Level1Out143[28] , \Level1Out143[27] , 
        \Level1Out143[26] , \Level1Out143[25] , \Level1Out143[24] , 
        \Level1Out143[23] , \Level1Out143[22] , \Level1Out143[21] , 
        \Level1Out143[20] , \Level1Out143[19] , \Level1Out143[18] , 
        \Level1Out143[17] , \Level1Out143[16] , \Level1Out143[15] , 
        \Level1Out143[14] , \Level1Out143[13] , \Level1Out143[12] , 
        \Level1Out143[11] , \Level1Out143[10] , \Level1Out143[9] , 
        \Level1Out143[8] , \Level1Out143[7] , \Level1Out143[6] , 
        \Level1Out143[5] , \Level1Out143[4] , \Level1Out143[3] , 
        \Level1Out143[2] , \Level1Out143[1] , \Level1Out143[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_164 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink164[31] , \ScanLink164[30] , 
        \ScanLink164[29] , \ScanLink164[28] , \ScanLink164[27] , 
        \ScanLink164[26] , \ScanLink164[25] , \ScanLink164[24] , 
        \ScanLink164[23] , \ScanLink164[22] , \ScanLink164[21] , 
        \ScanLink164[20] , \ScanLink164[19] , \ScanLink164[18] , 
        \ScanLink164[17] , \ScanLink164[16] , \ScanLink164[15] , 
        \ScanLink164[14] , \ScanLink164[13] , \ScanLink164[12] , 
        \ScanLink164[11] , \ScanLink164[10] , \ScanLink164[9] , 
        \ScanLink164[8] , \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , 
        \ScanLink164[4] , \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , 
        \ScanLink164[0] }), .ScanOut({\ScanLink165[31] , \ScanLink165[30] , 
        \ScanLink165[29] , \ScanLink165[28] , \ScanLink165[27] , 
        \ScanLink165[26] , \ScanLink165[25] , \ScanLink165[24] , 
        \ScanLink165[23] , \ScanLink165[22] , \ScanLink165[21] , 
        \ScanLink165[20] , \ScanLink165[19] , \ScanLink165[18] , 
        \ScanLink165[17] , \ScanLink165[16] , \ScanLink165[15] , 
        \ScanLink165[14] , \ScanLink165[13] , \ScanLink165[12] , 
        \ScanLink165[11] , \ScanLink165[10] , \ScanLink165[9] , 
        \ScanLink165[8] , \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , 
        \ScanLink165[4] , \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , 
        \ScanLink165[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load164[0] ), .Out({\Level1Out164[31] , \Level1Out164[30] , 
        \Level1Out164[29] , \Level1Out164[28] , \Level1Out164[27] , 
        \Level1Out164[26] , \Level1Out164[25] , \Level1Out164[24] , 
        \Level1Out164[23] , \Level1Out164[22] , \Level1Out164[21] , 
        \Level1Out164[20] , \Level1Out164[19] , \Level1Out164[18] , 
        \Level1Out164[17] , \Level1Out164[16] , \Level1Out164[15] , 
        \Level1Out164[14] , \Level1Out164[13] , \Level1Out164[12] , 
        \Level1Out164[11] , \Level1Out164[10] , \Level1Out164[9] , 
        \Level1Out164[8] , \Level1Out164[7] , \Level1Out164[6] , 
        \Level1Out164[5] , \Level1Out164[4] , \Level1Out164[3] , 
        \Level1Out164[2] , \Level1Out164[1] , \Level1Out164[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_158 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink158[31] , \ScanLink158[30] , 
        \ScanLink158[29] , \ScanLink158[28] , \ScanLink158[27] , 
        \ScanLink158[26] , \ScanLink158[25] , \ScanLink158[24] , 
        \ScanLink158[23] , \ScanLink158[22] , \ScanLink158[21] , 
        \ScanLink158[20] , \ScanLink158[19] , \ScanLink158[18] , 
        \ScanLink158[17] , \ScanLink158[16] , \ScanLink158[15] , 
        \ScanLink158[14] , \ScanLink158[13] , \ScanLink158[12] , 
        \ScanLink158[11] , \ScanLink158[10] , \ScanLink158[9] , 
        \ScanLink158[8] , \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , 
        \ScanLink158[4] , \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , 
        \ScanLink158[0] }), .ScanOut({\ScanLink159[31] , \ScanLink159[30] , 
        \ScanLink159[29] , \ScanLink159[28] , \ScanLink159[27] , 
        \ScanLink159[26] , \ScanLink159[25] , \ScanLink159[24] , 
        \ScanLink159[23] , \ScanLink159[22] , \ScanLink159[21] , 
        \ScanLink159[20] , \ScanLink159[19] , \ScanLink159[18] , 
        \ScanLink159[17] , \ScanLink159[16] , \ScanLink159[15] , 
        \ScanLink159[14] , \ScanLink159[13] , \ScanLink159[12] , 
        \ScanLink159[11] , \ScanLink159[10] , \ScanLink159[9] , 
        \ScanLink159[8] , \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , 
        \ScanLink159[4] , \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , 
        \ScanLink159[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load158[0] ), .Out({\Level1Out158[31] , \Level1Out158[30] , 
        \Level1Out158[29] , \Level1Out158[28] , \Level1Out158[27] , 
        \Level1Out158[26] , \Level1Out158[25] , \Level1Out158[24] , 
        \Level1Out158[23] , \Level1Out158[22] , \Level1Out158[21] , 
        \Level1Out158[20] , \Level1Out158[19] , \Level1Out158[18] , 
        \Level1Out158[17] , \Level1Out158[16] , \Level1Out158[15] , 
        \Level1Out158[14] , \Level1Out158[13] , \Level1Out158[12] , 
        \Level1Out158[11] , \Level1Out158[10] , \Level1Out158[9] , 
        \Level1Out158[8] , \Level1Out158[7] , \Level1Out158[6] , 
        \Level1Out158[5] , \Level1Out158[4] , \Level1Out158[3] , 
        \Level1Out158[2] , \Level1Out158[1] , \Level1Out158[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load8[0] ), .Out({\Level4Out8[31] , \Level4Out8[30] , 
        \Level4Out8[29] , \Level4Out8[28] , \Level4Out8[27] , \Level4Out8[26] , 
        \Level4Out8[25] , \Level4Out8[24] , \Level4Out8[23] , \Level4Out8[22] , 
        \Level4Out8[21] , \Level4Out8[20] , \Level4Out8[19] , \Level4Out8[18] , 
        \Level4Out8[17] , \Level4Out8[16] , \Level4Out8[15] , \Level4Out8[14] , 
        \Level4Out8[13] , \Level4Out8[12] , \Level4Out8[11] , \Level4Out8[10] , 
        \Level4Out8[9] , \Level4Out8[8] , \Level4Out8[7] , \Level4Out8[6] , 
        \Level4Out8[5] , \Level4Out8[4] , \Level4Out8[3] , \Level4Out8[2] , 
        \Level4Out8[1] , \Level4Out8[0] }), .In1({\Level2Out8[31] , 
        \Level2Out8[30] , \Level2Out8[29] , \Level2Out8[28] , \Level2Out8[27] , 
        \Level2Out8[26] , \Level2Out8[25] , \Level2Out8[24] , \Level2Out8[23] , 
        \Level2Out8[22] , \Level2Out8[21] , \Level2Out8[20] , \Level2Out8[19] , 
        \Level2Out8[18] , \Level2Out8[17] , \Level2Out8[16] , \Level2Out8[15] , 
        \Level2Out8[14] , \Level2Out8[13] , \Level2Out8[12] , \Level2Out8[11] , 
        \Level2Out8[10] , \Level2Out8[9] , \Level2Out8[8] , \Level2Out8[7] , 
        \Level2Out8[6] , \Level2Out8[5] , \Level2Out8[4] , \Level2Out8[3] , 
        \Level2Out8[2] , \Level2Out8[1] , \Level2Out8[0] }), .In2({
        \Level2Out10[31] , \Level2Out10[30] , \Level2Out10[29] , 
        \Level2Out10[28] , \Level2Out10[27] , \Level2Out10[26] , 
        \Level2Out10[25] , \Level2Out10[24] , \Level2Out10[23] , 
        \Level2Out10[22] , \Level2Out10[21] , \Level2Out10[20] , 
        \Level2Out10[19] , \Level2Out10[18] , \Level2Out10[17] , 
        \Level2Out10[16] , \Level2Out10[15] , \Level2Out10[14] , 
        \Level2Out10[13] , \Level2Out10[12] , \Level2Out10[11] , 
        \Level2Out10[10] , \Level2Out10[9] , \Level2Out10[8] , 
        \Level2Out10[7] , \Level2Out10[6] , \Level2Out10[5] , \Level2Out10[4] , 
        \Level2Out10[3] , \Level2Out10[2] , \Level2Out10[1] , \Level2Out10[0] 
        }), .Read1(\Level2Load8[0] ), .Read2(\Level2Load10[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_33 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanOut({\ScanLink34[31] , 
        \ScanLink34[30] , \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , 
        \ScanLink34[26] , \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , 
        \ScanLink34[22] , \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , 
        \ScanLink34[18] , \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , 
        \ScanLink34[14] , \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , 
        \ScanLink34[10] , \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , 
        \ScanLink34[6] , \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , 
        \ScanLink34[2] , \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load33[0] ), .Out({
        \Level1Out33[31] , \Level1Out33[30] , \Level1Out33[29] , 
        \Level1Out33[28] , \Level1Out33[27] , \Level1Out33[26] , 
        \Level1Out33[25] , \Level1Out33[24] , \Level1Out33[23] , 
        \Level1Out33[22] , \Level1Out33[21] , \Level1Out33[20] , 
        \Level1Out33[19] , \Level1Out33[18] , \Level1Out33[17] , 
        \Level1Out33[16] , \Level1Out33[15] , \Level1Out33[14] , 
        \Level1Out33[13] , \Level1Out33[12] , \Level1Out33[11] , 
        \Level1Out33[10] , \Level1Out33[9] , \Level1Out33[8] , 
        \Level1Out33[7] , \Level1Out33[6] , \Level1Out33[5] , \Level1Out33[4] , 
        \Level1Out33[3] , \Level1Out33[2] , \Level1Out33[1] , \Level1Out33[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_180_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load180[0] ), .Out({\Level4Out180[31] , \Level4Out180[30] , 
        \Level4Out180[29] , \Level4Out180[28] , \Level4Out180[27] , 
        \Level4Out180[26] , \Level4Out180[25] , \Level4Out180[24] , 
        \Level4Out180[23] , \Level4Out180[22] , \Level4Out180[21] , 
        \Level4Out180[20] , \Level4Out180[19] , \Level4Out180[18] , 
        \Level4Out180[17] , \Level4Out180[16] , \Level4Out180[15] , 
        \Level4Out180[14] , \Level4Out180[13] , \Level4Out180[12] , 
        \Level4Out180[11] , \Level4Out180[10] , \Level4Out180[9] , 
        \Level4Out180[8] , \Level4Out180[7] , \Level4Out180[6] , 
        \Level4Out180[5] , \Level4Out180[4] , \Level4Out180[3] , 
        \Level4Out180[2] , \Level4Out180[1] , \Level4Out180[0] }), .In1({
        \Level2Out180[31] , \Level2Out180[30] , \Level2Out180[29] , 
        \Level2Out180[28] , \Level2Out180[27] , \Level2Out180[26] , 
        \Level2Out180[25] , \Level2Out180[24] , \Level2Out180[23] , 
        \Level2Out180[22] , \Level2Out180[21] , \Level2Out180[20] , 
        \Level2Out180[19] , \Level2Out180[18] , \Level2Out180[17] , 
        \Level2Out180[16] , \Level2Out180[15] , \Level2Out180[14] , 
        \Level2Out180[13] , \Level2Out180[12] , \Level2Out180[11] , 
        \Level2Out180[10] , \Level2Out180[9] , \Level2Out180[8] , 
        \Level2Out180[7] , \Level2Out180[6] , \Level2Out180[5] , 
        \Level2Out180[4] , \Level2Out180[3] , \Level2Out180[2] , 
        \Level2Out180[1] , \Level2Out180[0] }), .In2({\Level2Out182[31] , 
        \Level2Out182[30] , \Level2Out182[29] , \Level2Out182[28] , 
        \Level2Out182[27] , \Level2Out182[26] , \Level2Out182[25] , 
        \Level2Out182[24] , \Level2Out182[23] , \Level2Out182[22] , 
        \Level2Out182[21] , \Level2Out182[20] , \Level2Out182[19] , 
        \Level2Out182[18] , \Level2Out182[17] , \Level2Out182[16] , 
        \Level2Out182[15] , \Level2Out182[14] , \Level2Out182[13] , 
        \Level2Out182[12] , \Level2Out182[11] , \Level2Out182[10] , 
        \Level2Out182[9] , \Level2Out182[8] , \Level2Out182[7] , 
        \Level2Out182[6] , \Level2Out182[5] , \Level2Out182[4] , 
        \Level2Out182[3] , \Level2Out182[2] , \Level2Out182[1] , 
        \Level2Out182[0] }), .Read1(\Level2Load180[0] ), .Read2(
        \Level2Load182[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_34 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanOut({\ScanLink35[31] , 
        \ScanLink35[30] , \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , 
        \ScanLink35[26] , \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , 
        \ScanLink35[22] , \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , 
        \ScanLink35[18] , \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , 
        \ScanLink35[14] , \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , 
        \ScanLink35[10] , \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , 
        \ScanLink35[6] , \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , 
        \ScanLink35[2] , \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load34[0] ), .Out({
        \Level1Out34[31] , \Level1Out34[30] , \Level1Out34[29] , 
        \Level1Out34[28] , \Level1Out34[27] , \Level1Out34[26] , 
        \Level1Out34[25] , \Level1Out34[24] , \Level1Out34[23] , 
        \Level1Out34[22] , \Level1Out34[21] , \Level1Out34[20] , 
        \Level1Out34[19] , \Level1Out34[18] , \Level1Out34[17] , 
        \Level1Out34[16] , \Level1Out34[15] , \Level1Out34[14] , 
        \Level1Out34[13] , \Level1Out34[12] , \Level1Out34[11] , 
        \Level1Out34[10] , \Level1Out34[9] , \Level1Out34[8] , 
        \Level1Out34[7] , \Level1Out34[6] , \Level1Out34[5] , \Level1Out34[4] , 
        \Level1Out34[3] , \Level1Out34[2] , \Level1Out34[1] , \Level1Out34[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_111 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink111[31] , \ScanLink111[30] , 
        \ScanLink111[29] , \ScanLink111[28] , \ScanLink111[27] , 
        \ScanLink111[26] , \ScanLink111[25] , \ScanLink111[24] , 
        \ScanLink111[23] , \ScanLink111[22] , \ScanLink111[21] , 
        \ScanLink111[20] , \ScanLink111[19] , \ScanLink111[18] , 
        \ScanLink111[17] , \ScanLink111[16] , \ScanLink111[15] , 
        \ScanLink111[14] , \ScanLink111[13] , \ScanLink111[12] , 
        \ScanLink111[11] , \ScanLink111[10] , \ScanLink111[9] , 
        \ScanLink111[8] , \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , 
        \ScanLink111[4] , \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , 
        \ScanLink111[0] }), .ScanOut({\ScanLink112[31] , \ScanLink112[30] , 
        \ScanLink112[29] , \ScanLink112[28] , \ScanLink112[27] , 
        \ScanLink112[26] , \ScanLink112[25] , \ScanLink112[24] , 
        \ScanLink112[23] , \ScanLink112[22] , \ScanLink112[21] , 
        \ScanLink112[20] , \ScanLink112[19] , \ScanLink112[18] , 
        \ScanLink112[17] , \ScanLink112[16] , \ScanLink112[15] , 
        \ScanLink112[14] , \ScanLink112[13] , \ScanLink112[12] , 
        \ScanLink112[11] , \ScanLink112[10] , \ScanLink112[9] , 
        \ScanLink112[8] , \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , 
        \ScanLink112[4] , \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , 
        \ScanLink112[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load111[0] ), .Out({\Level1Out111[31] , \Level1Out111[30] , 
        \Level1Out111[29] , \Level1Out111[28] , \Level1Out111[27] , 
        \Level1Out111[26] , \Level1Out111[25] , \Level1Out111[24] , 
        \Level1Out111[23] , \Level1Out111[22] , \Level1Out111[21] , 
        \Level1Out111[20] , \Level1Out111[19] , \Level1Out111[18] , 
        \Level1Out111[17] , \Level1Out111[16] , \Level1Out111[15] , 
        \Level1Out111[14] , \Level1Out111[13] , \Level1Out111[12] , 
        \Level1Out111[11] , \Level1Out111[10] , \Level1Out111[9] , 
        \Level1Out111[8] , \Level1Out111[7] , \Level1Out111[6] , 
        \Level1Out111[5] , \Level1Out111[4] , \Level1Out111[3] , 
        \Level1Out111[2] , \Level1Out111[1] , \Level1Out111[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_136 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink136[31] , \ScanLink136[30] , 
        \ScanLink136[29] , \ScanLink136[28] , \ScanLink136[27] , 
        \ScanLink136[26] , \ScanLink136[25] , \ScanLink136[24] , 
        \ScanLink136[23] , \ScanLink136[22] , \ScanLink136[21] , 
        \ScanLink136[20] , \ScanLink136[19] , \ScanLink136[18] , 
        \ScanLink136[17] , \ScanLink136[16] , \ScanLink136[15] , 
        \ScanLink136[14] , \ScanLink136[13] , \ScanLink136[12] , 
        \ScanLink136[11] , \ScanLink136[10] , \ScanLink136[9] , 
        \ScanLink136[8] , \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , 
        \ScanLink136[4] , \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , 
        \ScanLink136[0] }), .ScanOut({\ScanLink137[31] , \ScanLink137[30] , 
        \ScanLink137[29] , \ScanLink137[28] , \ScanLink137[27] , 
        \ScanLink137[26] , \ScanLink137[25] , \ScanLink137[24] , 
        \ScanLink137[23] , \ScanLink137[22] , \ScanLink137[21] , 
        \ScanLink137[20] , \ScanLink137[19] , \ScanLink137[18] , 
        \ScanLink137[17] , \ScanLink137[16] , \ScanLink137[15] , 
        \ScanLink137[14] , \ScanLink137[13] , \ScanLink137[12] , 
        \ScanLink137[11] , \ScanLink137[10] , \ScanLink137[9] , 
        \ScanLink137[8] , \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , 
        \ScanLink137[4] , \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , 
        \ScanLink137[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load136[0] ), .Out({\Level1Out136[31] , \Level1Out136[30] , 
        \Level1Out136[29] , \Level1Out136[28] , \Level1Out136[27] , 
        \Level1Out136[26] , \Level1Out136[25] , \Level1Out136[24] , 
        \Level1Out136[23] , \Level1Out136[22] , \Level1Out136[21] , 
        \Level1Out136[20] , \Level1Out136[19] , \Level1Out136[18] , 
        \Level1Out136[17] , \Level1Out136[16] , \Level1Out136[15] , 
        \Level1Out136[14] , \Level1Out136[13] , \Level1Out136[12] , 
        \Level1Out136[11] , \Level1Out136[10] , \Level1Out136[9] , 
        \Level1Out136[8] , \Level1Out136[7] , \Level1Out136[6] , 
        \Level1Out136[5] , \Level1Out136[4] , \Level1Out136[3] , 
        \Level1Out136[2] , \Level1Out136[1] , \Level1Out136[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_206 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink206[31] , \ScanLink206[30] , 
        \ScanLink206[29] , \ScanLink206[28] , \ScanLink206[27] , 
        \ScanLink206[26] , \ScanLink206[25] , \ScanLink206[24] , 
        \ScanLink206[23] , \ScanLink206[22] , \ScanLink206[21] , 
        \ScanLink206[20] , \ScanLink206[19] , \ScanLink206[18] , 
        \ScanLink206[17] , \ScanLink206[16] , \ScanLink206[15] , 
        \ScanLink206[14] , \ScanLink206[13] , \ScanLink206[12] , 
        \ScanLink206[11] , \ScanLink206[10] , \ScanLink206[9] , 
        \ScanLink206[8] , \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , 
        \ScanLink206[4] , \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , 
        \ScanLink206[0] }), .ScanOut({\ScanLink207[31] , \ScanLink207[30] , 
        \ScanLink207[29] , \ScanLink207[28] , \ScanLink207[27] , 
        \ScanLink207[26] , \ScanLink207[25] , \ScanLink207[24] , 
        \ScanLink207[23] , \ScanLink207[22] , \ScanLink207[21] , 
        \ScanLink207[20] , \ScanLink207[19] , \ScanLink207[18] , 
        \ScanLink207[17] , \ScanLink207[16] , \ScanLink207[15] , 
        \ScanLink207[14] , \ScanLink207[13] , \ScanLink207[12] , 
        \ScanLink207[11] , \ScanLink207[10] , \ScanLink207[9] , 
        \ScanLink207[8] , \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , 
        \ScanLink207[4] , \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , 
        \ScanLink207[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load206[0] ), .Out({\Level1Out206[31] , \Level1Out206[30] , 
        \Level1Out206[29] , \Level1Out206[28] , \Level1Out206[27] , 
        \Level1Out206[26] , \Level1Out206[25] , \Level1Out206[24] , 
        \Level1Out206[23] , \Level1Out206[22] , \Level1Out206[21] , 
        \Level1Out206[20] , \Level1Out206[19] , \Level1Out206[18] , 
        \Level1Out206[17] , \Level1Out206[16] , \Level1Out206[15] , 
        \Level1Out206[14] , \Level1Out206[13] , \Level1Out206[12] , 
        \Level1Out206[11] , \Level1Out206[10] , \Level1Out206[9] , 
        \Level1Out206[8] , \Level1Out206[7] , \Level1Out206[6] , 
        \Level1Out206[5] , \Level1Out206[4] , \Level1Out206[3] , 
        \Level1Out206[2] , \Level1Out206[1] , \Level1Out206[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_221 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink221[31] , \ScanLink221[30] , 
        \ScanLink221[29] , \ScanLink221[28] , \ScanLink221[27] , 
        \ScanLink221[26] , \ScanLink221[25] , \ScanLink221[24] , 
        \ScanLink221[23] , \ScanLink221[22] , \ScanLink221[21] , 
        \ScanLink221[20] , \ScanLink221[19] , \ScanLink221[18] , 
        \ScanLink221[17] , \ScanLink221[16] , \ScanLink221[15] , 
        \ScanLink221[14] , \ScanLink221[13] , \ScanLink221[12] , 
        \ScanLink221[11] , \ScanLink221[10] , \ScanLink221[9] , 
        \ScanLink221[8] , \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , 
        \ScanLink221[4] , \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , 
        \ScanLink221[0] }), .ScanOut({\ScanLink222[31] , \ScanLink222[30] , 
        \ScanLink222[29] , \ScanLink222[28] , \ScanLink222[27] , 
        \ScanLink222[26] , \ScanLink222[25] , \ScanLink222[24] , 
        \ScanLink222[23] , \ScanLink222[22] , \ScanLink222[21] , 
        \ScanLink222[20] , \ScanLink222[19] , \ScanLink222[18] , 
        \ScanLink222[17] , \ScanLink222[16] , \ScanLink222[15] , 
        \ScanLink222[14] , \ScanLink222[13] , \ScanLink222[12] , 
        \ScanLink222[11] , \ScanLink222[10] , \ScanLink222[9] , 
        \ScanLink222[8] , \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , 
        \ScanLink222[4] , \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , 
        \ScanLink222[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load221[0] ), .Out({\Level1Out221[31] , \Level1Out221[30] , 
        \Level1Out221[29] , \Level1Out221[28] , \Level1Out221[27] , 
        \Level1Out221[26] , \Level1Out221[25] , \Level1Out221[24] , 
        \Level1Out221[23] , \Level1Out221[22] , \Level1Out221[21] , 
        \Level1Out221[20] , \Level1Out221[19] , \Level1Out221[18] , 
        \Level1Out221[17] , \Level1Out221[16] , \Level1Out221[15] , 
        \Level1Out221[14] , \Level1Out221[13] , \Level1Out221[12] , 
        \Level1Out221[11] , \Level1Out221[10] , \Level1Out221[9] , 
        \Level1Out221[8] , \Level1Out221[7] , \Level1Out221[6] , 
        \Level1Out221[5] , \Level1Out221[4] , \Level1Out221[3] , 
        \Level1Out221[2] , \Level1Out221[1] , \Level1Out221[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_120_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load120[0] ), .Out({\Level2Out120[31] , \Level2Out120[30] , 
        \Level2Out120[29] , \Level2Out120[28] , \Level2Out120[27] , 
        \Level2Out120[26] , \Level2Out120[25] , \Level2Out120[24] , 
        \Level2Out120[23] , \Level2Out120[22] , \Level2Out120[21] , 
        \Level2Out120[20] , \Level2Out120[19] , \Level2Out120[18] , 
        \Level2Out120[17] , \Level2Out120[16] , \Level2Out120[15] , 
        \Level2Out120[14] , \Level2Out120[13] , \Level2Out120[12] , 
        \Level2Out120[11] , \Level2Out120[10] , \Level2Out120[9] , 
        \Level2Out120[8] , \Level2Out120[7] , \Level2Out120[6] , 
        \Level2Out120[5] , \Level2Out120[4] , \Level2Out120[3] , 
        \Level2Out120[2] , \Level2Out120[1] , \Level2Out120[0] }), .In1({
        \Level1Out120[31] , \Level1Out120[30] , \Level1Out120[29] , 
        \Level1Out120[28] , \Level1Out120[27] , \Level1Out120[26] , 
        \Level1Out120[25] , \Level1Out120[24] , \Level1Out120[23] , 
        \Level1Out120[22] , \Level1Out120[21] , \Level1Out120[20] , 
        \Level1Out120[19] , \Level1Out120[18] , \Level1Out120[17] , 
        \Level1Out120[16] , \Level1Out120[15] , \Level1Out120[14] , 
        \Level1Out120[13] , \Level1Out120[12] , \Level1Out120[11] , 
        \Level1Out120[10] , \Level1Out120[9] , \Level1Out120[8] , 
        \Level1Out120[7] , \Level1Out120[6] , \Level1Out120[5] , 
        \Level1Out120[4] , \Level1Out120[3] , \Level1Out120[2] , 
        \Level1Out120[1] , \Level1Out120[0] }), .In2({\Level1Out121[31] , 
        \Level1Out121[30] , \Level1Out121[29] , \Level1Out121[28] , 
        \Level1Out121[27] , \Level1Out121[26] , \Level1Out121[25] , 
        \Level1Out121[24] , \Level1Out121[23] , \Level1Out121[22] , 
        \Level1Out121[21] , \Level1Out121[20] , \Level1Out121[19] , 
        \Level1Out121[18] , \Level1Out121[17] , \Level1Out121[16] , 
        \Level1Out121[15] , \Level1Out121[14] , \Level1Out121[13] , 
        \Level1Out121[12] , \Level1Out121[11] , \Level1Out121[10] , 
        \Level1Out121[9] , \Level1Out121[8] , \Level1Out121[7] , 
        \Level1Out121[6] , \Level1Out121[5] , \Level1Out121[4] , 
        \Level1Out121[3] , \Level1Out121[2] , \Level1Out121[1] , 
        \Level1Out121[0] }), .Read1(\Level1Load120[0] ), .Read2(
        \Level1Load121[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_66_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load66[0] ), .Out({\Level2Out66[31] , \Level2Out66[30] , 
        \Level2Out66[29] , \Level2Out66[28] , \Level2Out66[27] , 
        \Level2Out66[26] , \Level2Out66[25] , \Level2Out66[24] , 
        \Level2Out66[23] , \Level2Out66[22] , \Level2Out66[21] , 
        \Level2Out66[20] , \Level2Out66[19] , \Level2Out66[18] , 
        \Level2Out66[17] , \Level2Out66[16] , \Level2Out66[15] , 
        \Level2Out66[14] , \Level2Out66[13] , \Level2Out66[12] , 
        \Level2Out66[11] , \Level2Out66[10] , \Level2Out66[9] , 
        \Level2Out66[8] , \Level2Out66[7] , \Level2Out66[6] , \Level2Out66[5] , 
        \Level2Out66[4] , \Level2Out66[3] , \Level2Out66[2] , \Level2Out66[1] , 
        \Level2Out66[0] }), .In1({\Level1Out66[31] , \Level1Out66[30] , 
        \Level1Out66[29] , \Level1Out66[28] , \Level1Out66[27] , 
        \Level1Out66[26] , \Level1Out66[25] , \Level1Out66[24] , 
        \Level1Out66[23] , \Level1Out66[22] , \Level1Out66[21] , 
        \Level1Out66[20] , \Level1Out66[19] , \Level1Out66[18] , 
        \Level1Out66[17] , \Level1Out66[16] , \Level1Out66[15] , 
        \Level1Out66[14] , \Level1Out66[13] , \Level1Out66[12] , 
        \Level1Out66[11] , \Level1Out66[10] , \Level1Out66[9] , 
        \Level1Out66[8] , \Level1Out66[7] , \Level1Out66[6] , \Level1Out66[5] , 
        \Level1Out66[4] , \Level1Out66[3] , \Level1Out66[2] , \Level1Out66[1] , 
        \Level1Out66[0] }), .In2({\Level1Out67[31] , \Level1Out67[30] , 
        \Level1Out67[29] , \Level1Out67[28] , \Level1Out67[27] , 
        \Level1Out67[26] , \Level1Out67[25] , \Level1Out67[24] , 
        \Level1Out67[23] , \Level1Out67[22] , \Level1Out67[21] , 
        \Level1Out67[20] , \Level1Out67[19] , \Level1Out67[18] , 
        \Level1Out67[17] , \Level1Out67[16] , \Level1Out67[15] , 
        \Level1Out67[14] , \Level1Out67[13] , \Level1Out67[12] , 
        \Level1Out67[11] , \Level1Out67[10] , \Level1Out67[9] , 
        \Level1Out67[8] , \Level1Out67[7] , \Level1Out67[6] , \Level1Out67[5] , 
        \Level1Out67[4] , \Level1Out67[3] , \Level1Out67[2] , \Level1Out67[1] , 
        \Level1Out67[0] }), .Read1(\Level1Load66[0] ), .Read2(
        \Level1Load67[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_214_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load214[0] ), .Out({\Level2Out214[31] , \Level2Out214[30] , 
        \Level2Out214[29] , \Level2Out214[28] , \Level2Out214[27] , 
        \Level2Out214[26] , \Level2Out214[25] , \Level2Out214[24] , 
        \Level2Out214[23] , \Level2Out214[22] , \Level2Out214[21] , 
        \Level2Out214[20] , \Level2Out214[19] , \Level2Out214[18] , 
        \Level2Out214[17] , \Level2Out214[16] , \Level2Out214[15] , 
        \Level2Out214[14] , \Level2Out214[13] , \Level2Out214[12] , 
        \Level2Out214[11] , \Level2Out214[10] , \Level2Out214[9] , 
        \Level2Out214[8] , \Level2Out214[7] , \Level2Out214[6] , 
        \Level2Out214[5] , \Level2Out214[4] , \Level2Out214[3] , 
        \Level2Out214[2] , \Level2Out214[1] , \Level2Out214[0] }), .In1({
        \Level1Out214[31] , \Level1Out214[30] , \Level1Out214[29] , 
        \Level1Out214[28] , \Level1Out214[27] , \Level1Out214[26] , 
        \Level1Out214[25] , \Level1Out214[24] , \Level1Out214[23] , 
        \Level1Out214[22] , \Level1Out214[21] , \Level1Out214[20] , 
        \Level1Out214[19] , \Level1Out214[18] , \Level1Out214[17] , 
        \Level1Out214[16] , \Level1Out214[15] , \Level1Out214[14] , 
        \Level1Out214[13] , \Level1Out214[12] , \Level1Out214[11] , 
        \Level1Out214[10] , \Level1Out214[9] , \Level1Out214[8] , 
        \Level1Out214[7] , \Level1Out214[6] , \Level1Out214[5] , 
        \Level1Out214[4] , \Level1Out214[3] , \Level1Out214[2] , 
        \Level1Out214[1] , \Level1Out214[0] }), .In2({\Level1Out215[31] , 
        \Level1Out215[30] , \Level1Out215[29] , \Level1Out215[28] , 
        \Level1Out215[27] , \Level1Out215[26] , \Level1Out215[25] , 
        \Level1Out215[24] , \Level1Out215[23] , \Level1Out215[22] , 
        \Level1Out215[21] , \Level1Out215[20] , \Level1Out215[19] , 
        \Level1Out215[18] , \Level1Out215[17] , \Level1Out215[16] , 
        \Level1Out215[15] , \Level1Out215[14] , \Level1Out215[13] , 
        \Level1Out215[12] , \Level1Out215[11] , \Level1Out215[10] , 
        \Level1Out215[9] , \Level1Out215[8] , \Level1Out215[7] , 
        \Level1Out215[6] , \Level1Out215[5] , \Level1Out215[4] , 
        \Level1Out215[3] , \Level1Out215[2] , \Level1Out215[1] , 
        \Level1Out215[0] }), .Read1(\Level1Load214[0] ), .Read2(
        \Level1Load215[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_116_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load116[0] ), .Out({\Level4Out116[31] , \Level4Out116[30] , 
        \Level4Out116[29] , \Level4Out116[28] , \Level4Out116[27] , 
        \Level4Out116[26] , \Level4Out116[25] , \Level4Out116[24] , 
        \Level4Out116[23] , \Level4Out116[22] , \Level4Out116[21] , 
        \Level4Out116[20] , \Level4Out116[19] , \Level4Out116[18] , 
        \Level4Out116[17] , \Level4Out116[16] , \Level4Out116[15] , 
        \Level4Out116[14] , \Level4Out116[13] , \Level4Out116[12] , 
        \Level4Out116[11] , \Level4Out116[10] , \Level4Out116[9] , 
        \Level4Out116[8] , \Level4Out116[7] , \Level4Out116[6] , 
        \Level4Out116[5] , \Level4Out116[4] , \Level4Out116[3] , 
        \Level4Out116[2] , \Level4Out116[1] , \Level4Out116[0] }), .In1({
        \Level2Out116[31] , \Level2Out116[30] , \Level2Out116[29] , 
        \Level2Out116[28] , \Level2Out116[27] , \Level2Out116[26] , 
        \Level2Out116[25] , \Level2Out116[24] , \Level2Out116[23] , 
        \Level2Out116[22] , \Level2Out116[21] , \Level2Out116[20] , 
        \Level2Out116[19] , \Level2Out116[18] , \Level2Out116[17] , 
        \Level2Out116[16] , \Level2Out116[15] , \Level2Out116[14] , 
        \Level2Out116[13] , \Level2Out116[12] , \Level2Out116[11] , 
        \Level2Out116[10] , \Level2Out116[9] , \Level2Out116[8] , 
        \Level2Out116[7] , \Level2Out116[6] , \Level2Out116[5] , 
        \Level2Out116[4] , \Level2Out116[3] , \Level2Out116[2] , 
        \Level2Out116[1] , \Level2Out116[0] }), .In2({\Level2Out118[31] , 
        \Level2Out118[30] , \Level2Out118[29] , \Level2Out118[28] , 
        \Level2Out118[27] , \Level2Out118[26] , \Level2Out118[25] , 
        \Level2Out118[24] , \Level2Out118[23] , \Level2Out118[22] , 
        \Level2Out118[21] , \Level2Out118[20] , \Level2Out118[19] , 
        \Level2Out118[18] , \Level2Out118[17] , \Level2Out118[16] , 
        \Level2Out118[15] , \Level2Out118[14] , \Level2Out118[13] , 
        \Level2Out118[12] , \Level2Out118[11] , \Level2Out118[10] , 
        \Level2Out118[9] , \Level2Out118[8] , \Level2Out118[7] , 
        \Level2Out118[6] , \Level2Out118[5] , \Level2Out118[4] , 
        \Level2Out118[3] , \Level2Out118[2] , \Level2Out118[1] , 
        \Level2Out118[0] }), .Read1(\Level2Load116[0] ), .Read2(
        \Level2Load118[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_208_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load208[0] ), .Out({\Level4Out208[31] , \Level4Out208[30] , 
        \Level4Out208[29] , \Level4Out208[28] , \Level4Out208[27] , 
        \Level4Out208[26] , \Level4Out208[25] , \Level4Out208[24] , 
        \Level4Out208[23] , \Level4Out208[22] , \Level4Out208[21] , 
        \Level4Out208[20] , \Level4Out208[19] , \Level4Out208[18] , 
        \Level4Out208[17] , \Level4Out208[16] , \Level4Out208[15] , 
        \Level4Out208[14] , \Level4Out208[13] , \Level4Out208[12] , 
        \Level4Out208[11] , \Level4Out208[10] , \Level4Out208[9] , 
        \Level4Out208[8] , \Level4Out208[7] , \Level4Out208[6] , 
        \Level4Out208[5] , \Level4Out208[4] , \Level4Out208[3] , 
        \Level4Out208[2] , \Level4Out208[1] , \Level4Out208[0] }), .In1({
        \Level2Out208[31] , \Level2Out208[30] , \Level2Out208[29] , 
        \Level2Out208[28] , \Level2Out208[27] , \Level2Out208[26] , 
        \Level2Out208[25] , \Level2Out208[24] , \Level2Out208[23] , 
        \Level2Out208[22] , \Level2Out208[21] , \Level2Out208[20] , 
        \Level2Out208[19] , \Level2Out208[18] , \Level2Out208[17] , 
        \Level2Out208[16] , \Level2Out208[15] , \Level2Out208[14] , 
        \Level2Out208[13] , \Level2Out208[12] , \Level2Out208[11] , 
        \Level2Out208[10] , \Level2Out208[9] , \Level2Out208[8] , 
        \Level2Out208[7] , \Level2Out208[6] , \Level2Out208[5] , 
        \Level2Out208[4] , \Level2Out208[3] , \Level2Out208[2] , 
        \Level2Out208[1] , \Level2Out208[0] }), .In2({\Level2Out210[31] , 
        \Level2Out210[30] , \Level2Out210[29] , \Level2Out210[28] , 
        \Level2Out210[27] , \Level2Out210[26] , \Level2Out210[25] , 
        \Level2Out210[24] , \Level2Out210[23] , \Level2Out210[22] , 
        \Level2Out210[21] , \Level2Out210[20] , \Level2Out210[19] , 
        \Level2Out210[18] , \Level2Out210[17] , \Level2Out210[16] , 
        \Level2Out210[15] , \Level2Out210[14] , \Level2Out210[13] , 
        \Level2Out210[12] , \Level2Out210[11] , \Level2Out210[10] , 
        \Level2Out210[9] , \Level2Out210[8] , \Level2Out210[7] , 
        \Level2Out210[6] , \Level2Out210[5] , \Level2Out210[4] , 
        \Level2Out210[3] , \Level2Out210[2] , \Level2Out210[1] , 
        \Level2Out210[0] }), .Read1(\Level2Load208[0] ), .Read2(
        \Level2Load210[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load0[0] ), .Out({\Level32Out0[31] , \Level32Out0[30] , 
        \Level32Out0[29] , \Level32Out0[28] , \Level32Out0[27] , 
        \Level32Out0[26] , \Level32Out0[25] , \Level32Out0[24] , 
        \Level32Out0[23] , \Level32Out0[22] , \Level32Out0[21] , 
        \Level32Out0[20] , \Level32Out0[19] , \Level32Out0[18] , 
        \Level32Out0[17] , \Level32Out0[16] , \Level32Out0[15] , 
        \Level32Out0[14] , \Level32Out0[13] , \Level32Out0[12] , 
        \Level32Out0[11] , \Level32Out0[10] , \Level32Out0[9] , 
        \Level32Out0[8] , \Level32Out0[7] , \Level32Out0[6] , \Level32Out0[5] , 
        \Level32Out0[4] , \Level32Out0[3] , \Level32Out0[2] , \Level32Out0[1] , 
        \Level32Out0[0] }), .In1({\Level16Out0[31] , \Level16Out0[30] , 
        \Level16Out0[29] , \Level16Out0[28] , \Level16Out0[27] , 
        \Level16Out0[26] , \Level16Out0[25] , \Level16Out0[24] , 
        \Level16Out0[23] , \Level16Out0[22] , \Level16Out0[21] , 
        \Level16Out0[20] , \Level16Out0[19] , \Level16Out0[18] , 
        \Level16Out0[17] , \Level16Out0[16] , \Level16Out0[15] , 
        \Level16Out0[14] , \Level16Out0[13] , \Level16Out0[12] , 
        \Level16Out0[11] , \Level16Out0[10] , \Level16Out0[9] , 
        \Level16Out0[8] , \Level16Out0[7] , \Level16Out0[6] , \Level16Out0[5] , 
        \Level16Out0[4] , \Level16Out0[3] , \Level16Out0[2] , \Level16Out0[1] , 
        \Level16Out0[0] }), .In2({\Level16Out16[31] , \Level16Out16[30] , 
        \Level16Out16[29] , \Level16Out16[28] , \Level16Out16[27] , 
        \Level16Out16[26] , \Level16Out16[25] , \Level16Out16[24] , 
        \Level16Out16[23] , \Level16Out16[22] , \Level16Out16[21] , 
        \Level16Out16[20] , \Level16Out16[19] , \Level16Out16[18] , 
        \Level16Out16[17] , \Level16Out16[16] , \Level16Out16[15] , 
        \Level16Out16[14] , \Level16Out16[13] , \Level16Out16[12] , 
        \Level16Out16[11] , \Level16Out16[10] , \Level16Out16[9] , 
        \Level16Out16[8] , \Level16Out16[7] , \Level16Out16[6] , 
        \Level16Out16[5] , \Level16Out16[4] , \Level16Out16[3] , 
        \Level16Out16[2] , \Level16Out16[1] , \Level16Out16[0] }), .Read1(
        \Level16Load0[0] ), .Read2(\Level16Load16[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_41 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanOut({\ScanLink42[31] , 
        \ScanLink42[30] , \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , 
        \ScanLink42[26] , \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , 
        \ScanLink42[22] , \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , 
        \ScanLink42[18] , \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , 
        \ScanLink42[14] , \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , 
        \ScanLink42[10] , \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , 
        \ScanLink42[6] , \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , 
        \ScanLink42[2] , \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load41[0] ), .Out({
        \Level1Out41[31] , \Level1Out41[30] , \Level1Out41[29] , 
        \Level1Out41[28] , \Level1Out41[27] , \Level1Out41[26] , 
        \Level1Out41[25] , \Level1Out41[24] , \Level1Out41[23] , 
        \Level1Out41[22] , \Level1Out41[21] , \Level1Out41[20] , 
        \Level1Out41[19] , \Level1Out41[18] , \Level1Out41[17] , 
        \Level1Out41[16] , \Level1Out41[15] , \Level1Out41[14] , 
        \Level1Out41[13] , \Level1Out41[12] , \Level1Out41[11] , 
        \Level1Out41[10] , \Level1Out41[9] , \Level1Out41[8] , 
        \Level1Out41[7] , \Level1Out41[6] , \Level1Out41[5] , \Level1Out41[4] , 
        \Level1Out41[3] , \Level1Out41[2] , \Level1Out41[1] , \Level1Out41[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_98 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink98[31] , \ScanLink98[30] , 
        \ScanLink98[29] , \ScanLink98[28] , \ScanLink98[27] , \ScanLink98[26] , 
        \ScanLink98[25] , \ScanLink98[24] , \ScanLink98[23] , \ScanLink98[22] , 
        \ScanLink98[21] , \ScanLink98[20] , \ScanLink98[19] , \ScanLink98[18] , 
        \ScanLink98[17] , \ScanLink98[16] , \ScanLink98[15] , \ScanLink98[14] , 
        \ScanLink98[13] , \ScanLink98[12] , \ScanLink98[11] , \ScanLink98[10] , 
        \ScanLink98[9] , \ScanLink98[8] , \ScanLink98[7] , \ScanLink98[6] , 
        \ScanLink98[5] , \ScanLink98[4] , \ScanLink98[3] , \ScanLink98[2] , 
        \ScanLink98[1] , \ScanLink98[0] }), .ScanOut({\ScanLink99[31] , 
        \ScanLink99[30] , \ScanLink99[29] , \ScanLink99[28] , \ScanLink99[27] , 
        \ScanLink99[26] , \ScanLink99[25] , \ScanLink99[24] , \ScanLink99[23] , 
        \ScanLink99[22] , \ScanLink99[21] , \ScanLink99[20] , \ScanLink99[19] , 
        \ScanLink99[18] , \ScanLink99[17] , \ScanLink99[16] , \ScanLink99[15] , 
        \ScanLink99[14] , \ScanLink99[13] , \ScanLink99[12] , \ScanLink99[11] , 
        \ScanLink99[10] , \ScanLink99[9] , \ScanLink99[8] , \ScanLink99[7] , 
        \ScanLink99[6] , \ScanLink99[5] , \ScanLink99[4] , \ScanLink99[3] , 
        \ScanLink99[2] , \ScanLink99[1] , \ScanLink99[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load98[0] ), .Out({
        \Level1Out98[31] , \Level1Out98[30] , \Level1Out98[29] , 
        \Level1Out98[28] , \Level1Out98[27] , \Level1Out98[26] , 
        \Level1Out98[25] , \Level1Out98[24] , \Level1Out98[23] , 
        \Level1Out98[22] , \Level1Out98[21] , \Level1Out98[20] , 
        \Level1Out98[19] , \Level1Out98[18] , \Level1Out98[17] , 
        \Level1Out98[16] , \Level1Out98[15] , \Level1Out98[14] , 
        \Level1Out98[13] , \Level1Out98[12] , \Level1Out98[11] , 
        \Level1Out98[10] , \Level1Out98[9] , \Level1Out98[8] , 
        \Level1Out98[7] , \Level1Out98[6] , \Level1Out98[5] , \Level1Out98[4] , 
        \Level1Out98[3] , \Level1Out98[2] , \Level1Out98[1] , \Level1Out98[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_116 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink116[31] , \ScanLink116[30] , 
        \ScanLink116[29] , \ScanLink116[28] , \ScanLink116[27] , 
        \ScanLink116[26] , \ScanLink116[25] , \ScanLink116[24] , 
        \ScanLink116[23] , \ScanLink116[22] , \ScanLink116[21] , 
        \ScanLink116[20] , \ScanLink116[19] , \ScanLink116[18] , 
        \ScanLink116[17] , \ScanLink116[16] , \ScanLink116[15] , 
        \ScanLink116[14] , \ScanLink116[13] , \ScanLink116[12] , 
        \ScanLink116[11] , \ScanLink116[10] , \ScanLink116[9] , 
        \ScanLink116[8] , \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , 
        \ScanLink116[4] , \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , 
        \ScanLink116[0] }), .ScanOut({\ScanLink117[31] , \ScanLink117[30] , 
        \ScanLink117[29] , \ScanLink117[28] , \ScanLink117[27] , 
        \ScanLink117[26] , \ScanLink117[25] , \ScanLink117[24] , 
        \ScanLink117[23] , \ScanLink117[22] , \ScanLink117[21] , 
        \ScanLink117[20] , \ScanLink117[19] , \ScanLink117[18] , 
        \ScanLink117[17] , \ScanLink117[16] , \ScanLink117[15] , 
        \ScanLink117[14] , \ScanLink117[13] , \ScanLink117[12] , 
        \ScanLink117[11] , \ScanLink117[10] , \ScanLink117[9] , 
        \ScanLink117[8] , \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , 
        \ScanLink117[4] , \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , 
        \ScanLink117[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load116[0] ), .Out({\Level1Out116[31] , \Level1Out116[30] , 
        \Level1Out116[29] , \Level1Out116[28] , \Level1Out116[27] , 
        \Level1Out116[26] , \Level1Out116[25] , \Level1Out116[24] , 
        \Level1Out116[23] , \Level1Out116[22] , \Level1Out116[21] , 
        \Level1Out116[20] , \Level1Out116[19] , \Level1Out116[18] , 
        \Level1Out116[17] , \Level1Out116[16] , \Level1Out116[15] , 
        \Level1Out116[14] , \Level1Out116[13] , \Level1Out116[12] , 
        \Level1Out116[11] , \Level1Out116[10] , \Level1Out116[9] , 
        \Level1Out116[8] , \Level1Out116[7] , \Level1Out116[6] , 
        \Level1Out116[5] , \Level1Out116[4] , \Level1Out116[3] , 
        \Level1Out116[2] , \Level1Out116[1] , \Level1Out116[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_131 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink131[31] , \ScanLink131[30] , 
        \ScanLink131[29] , \ScanLink131[28] , \ScanLink131[27] , 
        \ScanLink131[26] , \ScanLink131[25] , \ScanLink131[24] , 
        \ScanLink131[23] , \ScanLink131[22] , \ScanLink131[21] , 
        \ScanLink131[20] , \ScanLink131[19] , \ScanLink131[18] , 
        \ScanLink131[17] , \ScanLink131[16] , \ScanLink131[15] , 
        \ScanLink131[14] , \ScanLink131[13] , \ScanLink131[12] , 
        \ScanLink131[11] , \ScanLink131[10] , \ScanLink131[9] , 
        \ScanLink131[8] , \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , 
        \ScanLink131[4] , \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , 
        \ScanLink131[0] }), .ScanOut({\ScanLink132[31] , \ScanLink132[30] , 
        \ScanLink132[29] , \ScanLink132[28] , \ScanLink132[27] , 
        \ScanLink132[26] , \ScanLink132[25] , \ScanLink132[24] , 
        \ScanLink132[23] , \ScanLink132[22] , \ScanLink132[21] , 
        \ScanLink132[20] , \ScanLink132[19] , \ScanLink132[18] , 
        \ScanLink132[17] , \ScanLink132[16] , \ScanLink132[15] , 
        \ScanLink132[14] , \ScanLink132[13] , \ScanLink132[12] , 
        \ScanLink132[11] , \ScanLink132[10] , \ScanLink132[9] , 
        \ScanLink132[8] , \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , 
        \ScanLink132[4] , \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , 
        \ScanLink132[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load131[0] ), .Out({\Level1Out131[31] , \Level1Out131[30] , 
        \Level1Out131[29] , \Level1Out131[28] , \Level1Out131[27] , 
        \Level1Out131[26] , \Level1Out131[25] , \Level1Out131[24] , 
        \Level1Out131[23] , \Level1Out131[22] , \Level1Out131[21] , 
        \Level1Out131[20] , \Level1Out131[19] , \Level1Out131[18] , 
        \Level1Out131[17] , \Level1Out131[16] , \Level1Out131[15] , 
        \Level1Out131[14] , \Level1Out131[13] , \Level1Out131[12] , 
        \Level1Out131[11] , \Level1Out131[10] , \Level1Out131[9] , 
        \Level1Out131[8] , \Level1Out131[7] , \Level1Out131[6] , 
        \Level1Out131[5] , \Level1Out131[4] , \Level1Out131[3] , 
        \Level1Out131[2] , \Level1Out131[1] , \Level1Out131[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_201 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink201[31] , \ScanLink201[30] , 
        \ScanLink201[29] , \ScanLink201[28] , \ScanLink201[27] , 
        \ScanLink201[26] , \ScanLink201[25] , \ScanLink201[24] , 
        \ScanLink201[23] , \ScanLink201[22] , \ScanLink201[21] , 
        \ScanLink201[20] , \ScanLink201[19] , \ScanLink201[18] , 
        \ScanLink201[17] , \ScanLink201[16] , \ScanLink201[15] , 
        \ScanLink201[14] , \ScanLink201[13] , \ScanLink201[12] , 
        \ScanLink201[11] , \ScanLink201[10] , \ScanLink201[9] , 
        \ScanLink201[8] , \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , 
        \ScanLink201[4] , \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , 
        \ScanLink201[0] }), .ScanOut({\ScanLink202[31] , \ScanLink202[30] , 
        \ScanLink202[29] , \ScanLink202[28] , \ScanLink202[27] , 
        \ScanLink202[26] , \ScanLink202[25] , \ScanLink202[24] , 
        \ScanLink202[23] , \ScanLink202[22] , \ScanLink202[21] , 
        \ScanLink202[20] , \ScanLink202[19] , \ScanLink202[18] , 
        \ScanLink202[17] , \ScanLink202[16] , \ScanLink202[15] , 
        \ScanLink202[14] , \ScanLink202[13] , \ScanLink202[12] , 
        \ScanLink202[11] , \ScanLink202[10] , \ScanLink202[9] , 
        \ScanLink202[8] , \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , 
        \ScanLink202[4] , \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , 
        \ScanLink202[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load201[0] ), .Out({\Level1Out201[31] , \Level1Out201[30] , 
        \Level1Out201[29] , \Level1Out201[28] , \Level1Out201[27] , 
        \Level1Out201[26] , \Level1Out201[25] , \Level1Out201[24] , 
        \Level1Out201[23] , \Level1Out201[22] , \Level1Out201[21] , 
        \Level1Out201[20] , \Level1Out201[19] , \Level1Out201[18] , 
        \Level1Out201[17] , \Level1Out201[16] , \Level1Out201[15] , 
        \Level1Out201[14] , \Level1Out201[13] , \Level1Out201[12] , 
        \Level1Out201[11] , \Level1Out201[10] , \Level1Out201[9] , 
        \Level1Out201[8] , \Level1Out201[7] , \Level1Out201[6] , 
        \Level1Out201[5] , \Level1Out201[4] , \Level1Out201[3] , 
        \Level1Out201[2] , \Level1Out201[1] , \Level1Out201[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_226 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink226[31] , \ScanLink226[30] , 
        \ScanLink226[29] , \ScanLink226[28] , \ScanLink226[27] , 
        \ScanLink226[26] , \ScanLink226[25] , \ScanLink226[24] , 
        \ScanLink226[23] , \ScanLink226[22] , \ScanLink226[21] , 
        \ScanLink226[20] , \ScanLink226[19] , \ScanLink226[18] , 
        \ScanLink226[17] , \ScanLink226[16] , \ScanLink226[15] , 
        \ScanLink226[14] , \ScanLink226[13] , \ScanLink226[12] , 
        \ScanLink226[11] , \ScanLink226[10] , \ScanLink226[9] , 
        \ScanLink226[8] , \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , 
        \ScanLink226[4] , \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , 
        \ScanLink226[0] }), .ScanOut({\ScanLink227[31] , \ScanLink227[30] , 
        \ScanLink227[29] , \ScanLink227[28] , \ScanLink227[27] , 
        \ScanLink227[26] , \ScanLink227[25] , \ScanLink227[24] , 
        \ScanLink227[23] , \ScanLink227[22] , \ScanLink227[21] , 
        \ScanLink227[20] , \ScanLink227[19] , \ScanLink227[18] , 
        \ScanLink227[17] , \ScanLink227[16] , \ScanLink227[15] , 
        \ScanLink227[14] , \ScanLink227[13] , \ScanLink227[12] , 
        \ScanLink227[11] , \ScanLink227[10] , \ScanLink227[9] , 
        \ScanLink227[8] , \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , 
        \ScanLink227[4] , \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , 
        \ScanLink227[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load226[0] ), .Out({\Level1Out226[31] , \Level1Out226[30] , 
        \Level1Out226[29] , \Level1Out226[28] , \Level1Out226[27] , 
        \Level1Out226[26] , \Level1Out226[25] , \Level1Out226[24] , 
        \Level1Out226[23] , \Level1Out226[22] , \Level1Out226[21] , 
        \Level1Out226[20] , \Level1Out226[19] , \Level1Out226[18] , 
        \Level1Out226[17] , \Level1Out226[16] , \Level1Out226[15] , 
        \Level1Out226[14] , \Level1Out226[13] , \Level1Out226[12] , 
        \Level1Out226[11] , \Level1Out226[10] , \Level1Out226[9] , 
        \Level1Out226[8] , \Level1Out226[7] , \Level1Out226[6] , 
        \Level1Out226[5] , \Level1Out226[4] , \Level1Out226[3] , 
        \Level1Out226[2] , \Level1Out226[1] , \Level1Out226[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load0[0] ), .Out({\Level2Out0[31] , \Level2Out0[30] , 
        \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , \Level2Out0[26] , 
        \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , \Level2Out0[22] , 
        \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , \Level2Out0[18] , 
        \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , \Level2Out0[14] , 
        \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , \Level2Out0[10] , 
        \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , \Level2Out0[6] , 
        \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , \Level2Out0[2] , 
        \Level2Out0[1] , \Level2Out0[0] }), .In1({\Level1Out0[31] , 
        \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , \Level1Out0[27] , 
        \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , \Level1Out0[23] , 
        \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , \Level1Out0[19] , 
        \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , \Level1Out0[15] , 
        \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , \Level1Out0[11] , 
        \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , \Level1Out0[7] , 
        \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , \Level1Out0[3] , 
        \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] }), .In2({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] }), 
        .Read1(\Level1Load0[0] ), .Read2(\Level1Load1[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_178 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink178[31] , \ScanLink178[30] , 
        \ScanLink178[29] , \ScanLink178[28] , \ScanLink178[27] , 
        \ScanLink178[26] , \ScanLink178[25] , \ScanLink178[24] , 
        \ScanLink178[23] , \ScanLink178[22] , \ScanLink178[21] , 
        \ScanLink178[20] , \ScanLink178[19] , \ScanLink178[18] , 
        \ScanLink178[17] , \ScanLink178[16] , \ScanLink178[15] , 
        \ScanLink178[14] , \ScanLink178[13] , \ScanLink178[12] , 
        \ScanLink178[11] , \ScanLink178[10] , \ScanLink178[9] , 
        \ScanLink178[8] , \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , 
        \ScanLink178[4] , \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , 
        \ScanLink178[0] }), .ScanOut({\ScanLink179[31] , \ScanLink179[30] , 
        \ScanLink179[29] , \ScanLink179[28] , \ScanLink179[27] , 
        \ScanLink179[26] , \ScanLink179[25] , \ScanLink179[24] , 
        \ScanLink179[23] , \ScanLink179[22] , \ScanLink179[21] , 
        \ScanLink179[20] , \ScanLink179[19] , \ScanLink179[18] , 
        \ScanLink179[17] , \ScanLink179[16] , \ScanLink179[15] , 
        \ScanLink179[14] , \ScanLink179[13] , \ScanLink179[12] , 
        \ScanLink179[11] , \ScanLink179[10] , \ScanLink179[9] , 
        \ScanLink179[8] , \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , 
        \ScanLink179[4] , \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , 
        \ScanLink179[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load178[0] ), .Out({\Level1Out178[31] , \Level1Out178[30] , 
        \Level1Out178[29] , \Level1Out178[28] , \Level1Out178[27] , 
        \Level1Out178[26] , \Level1Out178[25] , \Level1Out178[24] , 
        \Level1Out178[23] , \Level1Out178[22] , \Level1Out178[21] , 
        \Level1Out178[20] , \Level1Out178[19] , \Level1Out178[18] , 
        \Level1Out178[17] , \Level1Out178[16] , \Level1Out178[15] , 
        \Level1Out178[14] , \Level1Out178[13] , \Level1Out178[12] , 
        \Level1Out178[11] , \Level1Out178[10] , \Level1Out178[9] , 
        \Level1Out178[8] , \Level1Out178[7] , \Level1Out178[6] , 
        \Level1Out178[5] , \Level1Out178[4] , \Level1Out178[3] , 
        \Level1Out178[2] , \Level1Out178[1] , \Level1Out178[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_248 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink248[31] , \ScanLink248[30] , 
        \ScanLink248[29] , \ScanLink248[28] , \ScanLink248[27] , 
        \ScanLink248[26] , \ScanLink248[25] , \ScanLink248[24] , 
        \ScanLink248[23] , \ScanLink248[22] , \ScanLink248[21] , 
        \ScanLink248[20] , \ScanLink248[19] , \ScanLink248[18] , 
        \ScanLink248[17] , \ScanLink248[16] , \ScanLink248[15] , 
        \ScanLink248[14] , \ScanLink248[13] , \ScanLink248[12] , 
        \ScanLink248[11] , \ScanLink248[10] , \ScanLink248[9] , 
        \ScanLink248[8] , \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , 
        \ScanLink248[4] , \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , 
        \ScanLink248[0] }), .ScanOut({\ScanLink249[31] , \ScanLink249[30] , 
        \ScanLink249[29] , \ScanLink249[28] , \ScanLink249[27] , 
        \ScanLink249[26] , \ScanLink249[25] , \ScanLink249[24] , 
        \ScanLink249[23] , \ScanLink249[22] , \ScanLink249[21] , 
        \ScanLink249[20] , \ScanLink249[19] , \ScanLink249[18] , 
        \ScanLink249[17] , \ScanLink249[16] , \ScanLink249[15] , 
        \ScanLink249[14] , \ScanLink249[13] , \ScanLink249[12] , 
        \ScanLink249[11] , \ScanLink249[10] , \ScanLink249[9] , 
        \ScanLink249[8] , \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , 
        \ScanLink249[4] , \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , 
        \ScanLink249[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load248[0] ), .Out({\Level1Out248[31] , \Level1Out248[30] , 
        \Level1Out248[29] , \Level1Out248[28] , \Level1Out248[27] , 
        \Level1Out248[26] , \Level1Out248[25] , \Level1Out248[24] , 
        \Level1Out248[23] , \Level1Out248[22] , \Level1Out248[21] , 
        \Level1Out248[20] , \Level1Out248[19] , \Level1Out248[18] , 
        \Level1Out248[17] , \Level1Out248[16] , \Level1Out248[15] , 
        \Level1Out248[14] , \Level1Out248[13] , \Level1Out248[12] , 
        \Level1Out248[11] , \Level1Out248[10] , \Level1Out248[9] , 
        \Level1Out248[8] , \Level1Out248[7] , \Level1Out248[6] , 
        \Level1Out248[5] , \Level1Out248[4] , \Level1Out248[3] , 
        \Level1Out248[2] , \Level1Out248[1] , \Level1Out248[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_188_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load188[0] ), .Out({\Level2Out188[31] , \Level2Out188[30] , 
        \Level2Out188[29] , \Level2Out188[28] , \Level2Out188[27] , 
        \Level2Out188[26] , \Level2Out188[25] , \Level2Out188[24] , 
        \Level2Out188[23] , \Level2Out188[22] , \Level2Out188[21] , 
        \Level2Out188[20] , \Level2Out188[19] , \Level2Out188[18] , 
        \Level2Out188[17] , \Level2Out188[16] , \Level2Out188[15] , 
        \Level2Out188[14] , \Level2Out188[13] , \Level2Out188[12] , 
        \Level2Out188[11] , \Level2Out188[10] , \Level2Out188[9] , 
        \Level2Out188[8] , \Level2Out188[7] , \Level2Out188[6] , 
        \Level2Out188[5] , \Level2Out188[4] , \Level2Out188[3] , 
        \Level2Out188[2] , \Level2Out188[1] , \Level2Out188[0] }), .In1({
        \Level1Out188[31] , \Level1Out188[30] , \Level1Out188[29] , 
        \Level1Out188[28] , \Level1Out188[27] , \Level1Out188[26] , 
        \Level1Out188[25] , \Level1Out188[24] , \Level1Out188[23] , 
        \Level1Out188[22] , \Level1Out188[21] , \Level1Out188[20] , 
        \Level1Out188[19] , \Level1Out188[18] , \Level1Out188[17] , 
        \Level1Out188[16] , \Level1Out188[15] , \Level1Out188[14] , 
        \Level1Out188[13] , \Level1Out188[12] , \Level1Out188[11] , 
        \Level1Out188[10] , \Level1Out188[9] , \Level1Out188[8] , 
        \Level1Out188[7] , \Level1Out188[6] , \Level1Out188[5] , 
        \Level1Out188[4] , \Level1Out188[3] , \Level1Out188[2] , 
        \Level1Out188[1] , \Level1Out188[0] }), .In2({\Level1Out189[31] , 
        \Level1Out189[30] , \Level1Out189[29] , \Level1Out189[28] , 
        \Level1Out189[27] , \Level1Out189[26] , \Level1Out189[25] , 
        \Level1Out189[24] , \Level1Out189[23] , \Level1Out189[22] , 
        \Level1Out189[21] , \Level1Out189[20] , \Level1Out189[19] , 
        \Level1Out189[18] , \Level1Out189[17] , \Level1Out189[16] , 
        \Level1Out189[15] , \Level1Out189[14] , \Level1Out189[13] , 
        \Level1Out189[12] , \Level1Out189[11] , \Level1Out189[10] , 
        \Level1Out189[9] , \Level1Out189[8] , \Level1Out189[7] , 
        \Level1Out189[6] , \Level1Out189[5] , \Level1Out189[4] , 
        \Level1Out189[3] , \Level1Out189[2] , \Level1Out189[1] , 
        \Level1Out189[0] }), .Read1(\Level1Load188[0] ), .Read2(
        \Level1Load189[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_58_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load58[0] ), .Out({\Level2Out58[31] , \Level2Out58[30] , 
        \Level2Out58[29] , \Level2Out58[28] , \Level2Out58[27] , 
        \Level2Out58[26] , \Level2Out58[25] , \Level2Out58[24] , 
        \Level2Out58[23] , \Level2Out58[22] , \Level2Out58[21] , 
        \Level2Out58[20] , \Level2Out58[19] , \Level2Out58[18] , 
        \Level2Out58[17] , \Level2Out58[16] , \Level2Out58[15] , 
        \Level2Out58[14] , \Level2Out58[13] , \Level2Out58[12] , 
        \Level2Out58[11] , \Level2Out58[10] , \Level2Out58[9] , 
        \Level2Out58[8] , \Level2Out58[7] , \Level2Out58[6] , \Level2Out58[5] , 
        \Level2Out58[4] , \Level2Out58[3] , \Level2Out58[2] , \Level2Out58[1] , 
        \Level2Out58[0] }), .In1({\Level1Out58[31] , \Level1Out58[30] , 
        \Level1Out58[29] , \Level1Out58[28] , \Level1Out58[27] , 
        \Level1Out58[26] , \Level1Out58[25] , \Level1Out58[24] , 
        \Level1Out58[23] , \Level1Out58[22] , \Level1Out58[21] , 
        \Level1Out58[20] , \Level1Out58[19] , \Level1Out58[18] , 
        \Level1Out58[17] , \Level1Out58[16] , \Level1Out58[15] , 
        \Level1Out58[14] , \Level1Out58[13] , \Level1Out58[12] , 
        \Level1Out58[11] , \Level1Out58[10] , \Level1Out58[9] , 
        \Level1Out58[8] , \Level1Out58[7] , \Level1Out58[6] , \Level1Out58[5] , 
        \Level1Out58[4] , \Level1Out58[3] , \Level1Out58[2] , \Level1Out58[1] , 
        \Level1Out58[0] }), .In2({\Level1Out59[31] , \Level1Out59[30] , 
        \Level1Out59[29] , \Level1Out59[28] , \Level1Out59[27] , 
        \Level1Out59[26] , \Level1Out59[25] , \Level1Out59[24] , 
        \Level1Out59[23] , \Level1Out59[22] , \Level1Out59[21] , 
        \Level1Out59[20] , \Level1Out59[19] , \Level1Out59[18] , 
        \Level1Out59[17] , \Level1Out59[16] , \Level1Out59[15] , 
        \Level1Out59[14] , \Level1Out59[13] , \Level1Out59[12] , 
        \Level1Out59[11] , \Level1Out59[10] , \Level1Out59[9] , 
        \Level1Out59[8] , \Level1Out59[7] , \Level1Out59[6] , \Level1Out59[5] , 
        \Level1Out59[4] , \Level1Out59[3] , \Level1Out59[2] , \Level1Out59[1] , 
        \Level1Out59[0] }), .Read1(\Level1Load58[0] ), .Read2(
        \Level1Load59[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_72_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load72[0] ), .Out({\Level2Out72[31] , \Level2Out72[30] , 
        \Level2Out72[29] , \Level2Out72[28] , \Level2Out72[27] , 
        \Level2Out72[26] , \Level2Out72[25] , \Level2Out72[24] , 
        \Level2Out72[23] , \Level2Out72[22] , \Level2Out72[21] , 
        \Level2Out72[20] , \Level2Out72[19] , \Level2Out72[18] , 
        \Level2Out72[17] , \Level2Out72[16] , \Level2Out72[15] , 
        \Level2Out72[14] , \Level2Out72[13] , \Level2Out72[12] , 
        \Level2Out72[11] , \Level2Out72[10] , \Level2Out72[9] , 
        \Level2Out72[8] , \Level2Out72[7] , \Level2Out72[6] , \Level2Out72[5] , 
        \Level2Out72[4] , \Level2Out72[3] , \Level2Out72[2] , \Level2Out72[1] , 
        \Level2Out72[0] }), .In1({\Level1Out72[31] , \Level1Out72[30] , 
        \Level1Out72[29] , \Level1Out72[28] , \Level1Out72[27] , 
        \Level1Out72[26] , \Level1Out72[25] , \Level1Out72[24] , 
        \Level1Out72[23] , \Level1Out72[22] , \Level1Out72[21] , 
        \Level1Out72[20] , \Level1Out72[19] , \Level1Out72[18] , 
        \Level1Out72[17] , \Level1Out72[16] , \Level1Out72[15] , 
        \Level1Out72[14] , \Level1Out72[13] , \Level1Out72[12] , 
        \Level1Out72[11] , \Level1Out72[10] , \Level1Out72[9] , 
        \Level1Out72[8] , \Level1Out72[7] , \Level1Out72[6] , \Level1Out72[5] , 
        \Level1Out72[4] , \Level1Out72[3] , \Level1Out72[2] , \Level1Out72[1] , 
        \Level1Out72[0] }), .In2({\Level1Out73[31] , \Level1Out73[30] , 
        \Level1Out73[29] , \Level1Out73[28] , \Level1Out73[27] , 
        \Level1Out73[26] , \Level1Out73[25] , \Level1Out73[24] , 
        \Level1Out73[23] , \Level1Out73[22] , \Level1Out73[21] , 
        \Level1Out73[20] , \Level1Out73[19] , \Level1Out73[18] , 
        \Level1Out73[17] , \Level1Out73[16] , \Level1Out73[15] , 
        \Level1Out73[14] , \Level1Out73[13] , \Level1Out73[12] , 
        \Level1Out73[11] , \Level1Out73[10] , \Level1Out73[9] , 
        \Level1Out73[8] , \Level1Out73[7] , \Level1Out73[6] , \Level1Out73[5] , 
        \Level1Out73[4] , \Level1Out73[3] , \Level1Out73[2] , \Level1Out73[1] , 
        \Level1Out73[0] }), .Read1(\Level1Load72[0] ), .Read2(
        \Level1Load73[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_200_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load200[0] ), .Out({\Level2Out200[31] , \Level2Out200[30] , 
        \Level2Out200[29] , \Level2Out200[28] , \Level2Out200[27] , 
        \Level2Out200[26] , \Level2Out200[25] , \Level2Out200[24] , 
        \Level2Out200[23] , \Level2Out200[22] , \Level2Out200[21] , 
        \Level2Out200[20] , \Level2Out200[19] , \Level2Out200[18] , 
        \Level2Out200[17] , \Level2Out200[16] , \Level2Out200[15] , 
        \Level2Out200[14] , \Level2Out200[13] , \Level2Out200[12] , 
        \Level2Out200[11] , \Level2Out200[10] , \Level2Out200[9] , 
        \Level2Out200[8] , \Level2Out200[7] , \Level2Out200[6] , 
        \Level2Out200[5] , \Level2Out200[4] , \Level2Out200[3] , 
        \Level2Out200[2] , \Level2Out200[1] , \Level2Out200[0] }), .In1({
        \Level1Out200[31] , \Level1Out200[30] , \Level1Out200[29] , 
        \Level1Out200[28] , \Level1Out200[27] , \Level1Out200[26] , 
        \Level1Out200[25] , \Level1Out200[24] , \Level1Out200[23] , 
        \Level1Out200[22] , \Level1Out200[21] , \Level1Out200[20] , 
        \Level1Out200[19] , \Level1Out200[18] , \Level1Out200[17] , 
        \Level1Out200[16] , \Level1Out200[15] , \Level1Out200[14] , 
        \Level1Out200[13] , \Level1Out200[12] , \Level1Out200[11] , 
        \Level1Out200[10] , \Level1Out200[9] , \Level1Out200[8] , 
        \Level1Out200[7] , \Level1Out200[6] , \Level1Out200[5] , 
        \Level1Out200[4] , \Level1Out200[3] , \Level1Out200[2] , 
        \Level1Out200[1] , \Level1Out200[0] }), .In2({\Level1Out201[31] , 
        \Level1Out201[30] , \Level1Out201[29] , \Level1Out201[28] , 
        \Level1Out201[27] , \Level1Out201[26] , \Level1Out201[25] , 
        \Level1Out201[24] , \Level1Out201[23] , \Level1Out201[22] , 
        \Level1Out201[21] , \Level1Out201[20] , \Level1Out201[19] , 
        \Level1Out201[18] , \Level1Out201[17] , \Level1Out201[16] , 
        \Level1Out201[15] , \Level1Out201[14] , \Level1Out201[13] , 
        \Level1Out201[12] , \Level1Out201[11] , \Level1Out201[10] , 
        \Level1Out201[9] , \Level1Out201[8] , \Level1Out201[7] , 
        \Level1Out201[6] , \Level1Out201[5] , \Level1Out201[4] , 
        \Level1Out201[3] , \Level1Out201[2] , \Level1Out201[1] , 
        \Level1Out201[0] }), .Read1(\Level1Load200[0] ), .Read2(
        \Level1Load201[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_44_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load44[0] ), .Out({\Level4Out44[31] , \Level4Out44[30] , 
        \Level4Out44[29] , \Level4Out44[28] , \Level4Out44[27] , 
        \Level4Out44[26] , \Level4Out44[25] , \Level4Out44[24] , 
        \Level4Out44[23] , \Level4Out44[22] , \Level4Out44[21] , 
        \Level4Out44[20] , \Level4Out44[19] , \Level4Out44[18] , 
        \Level4Out44[17] , \Level4Out44[16] , \Level4Out44[15] , 
        \Level4Out44[14] , \Level4Out44[13] , \Level4Out44[12] , 
        \Level4Out44[11] , \Level4Out44[10] , \Level4Out44[9] , 
        \Level4Out44[8] , \Level4Out44[7] , \Level4Out44[6] , \Level4Out44[5] , 
        \Level4Out44[4] , \Level4Out44[3] , \Level4Out44[2] , \Level4Out44[1] , 
        \Level4Out44[0] }), .In1({\Level2Out44[31] , \Level2Out44[30] , 
        \Level2Out44[29] , \Level2Out44[28] , \Level2Out44[27] , 
        \Level2Out44[26] , \Level2Out44[25] , \Level2Out44[24] , 
        \Level2Out44[23] , \Level2Out44[22] , \Level2Out44[21] , 
        \Level2Out44[20] , \Level2Out44[19] , \Level2Out44[18] , 
        \Level2Out44[17] , \Level2Out44[16] , \Level2Out44[15] , 
        \Level2Out44[14] , \Level2Out44[13] , \Level2Out44[12] , 
        \Level2Out44[11] , \Level2Out44[10] , \Level2Out44[9] , 
        \Level2Out44[8] , \Level2Out44[7] , \Level2Out44[6] , \Level2Out44[5] , 
        \Level2Out44[4] , \Level2Out44[3] , \Level2Out44[2] , \Level2Out44[1] , 
        \Level2Out44[0] }), .In2({\Level2Out46[31] , \Level2Out46[30] , 
        \Level2Out46[29] , \Level2Out46[28] , \Level2Out46[27] , 
        \Level2Out46[26] , \Level2Out46[25] , \Level2Out46[24] , 
        \Level2Out46[23] , \Level2Out46[22] , \Level2Out46[21] , 
        \Level2Out46[20] , \Level2Out46[19] , \Level2Out46[18] , 
        \Level2Out46[17] , \Level2Out46[16] , \Level2Out46[15] , 
        \Level2Out46[14] , \Level2Out46[13] , \Level2Out46[12] , 
        \Level2Out46[11] , \Level2Out46[10] , \Level2Out46[9] , 
        \Level2Out46[8] , \Level2Out46[7] , \Level2Out46[6] , \Level2Out46[5] , 
        \Level2Out46[4] , \Level2Out46[3] , \Level2Out46[2] , \Level2Out46[1] , 
        \Level2Out46[0] }), .Read1(\Level2Load44[0] ), .Read2(
        \Level2Load46[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_134_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load134[0] ), .Out({\Level2Out134[31] , \Level2Out134[30] , 
        \Level2Out134[29] , \Level2Out134[28] , \Level2Out134[27] , 
        \Level2Out134[26] , \Level2Out134[25] , \Level2Out134[24] , 
        \Level2Out134[23] , \Level2Out134[22] , \Level2Out134[21] , 
        \Level2Out134[20] , \Level2Out134[19] , \Level2Out134[18] , 
        \Level2Out134[17] , \Level2Out134[16] , \Level2Out134[15] , 
        \Level2Out134[14] , \Level2Out134[13] , \Level2Out134[12] , 
        \Level2Out134[11] , \Level2Out134[10] , \Level2Out134[9] , 
        \Level2Out134[8] , \Level2Out134[7] , \Level2Out134[6] , 
        \Level2Out134[5] , \Level2Out134[4] , \Level2Out134[3] , 
        \Level2Out134[2] , \Level2Out134[1] , \Level2Out134[0] }), .In1({
        \Level1Out134[31] , \Level1Out134[30] , \Level1Out134[29] , 
        \Level1Out134[28] , \Level1Out134[27] , \Level1Out134[26] , 
        \Level1Out134[25] , \Level1Out134[24] , \Level1Out134[23] , 
        \Level1Out134[22] , \Level1Out134[21] , \Level1Out134[20] , 
        \Level1Out134[19] , \Level1Out134[18] , \Level1Out134[17] , 
        \Level1Out134[16] , \Level1Out134[15] , \Level1Out134[14] , 
        \Level1Out134[13] , \Level1Out134[12] , \Level1Out134[11] , 
        \Level1Out134[10] , \Level1Out134[9] , \Level1Out134[8] , 
        \Level1Out134[7] , \Level1Out134[6] , \Level1Out134[5] , 
        \Level1Out134[4] , \Level1Out134[3] , \Level1Out134[2] , 
        \Level1Out134[1] , \Level1Out134[0] }), .In2({\Level1Out135[31] , 
        \Level1Out135[30] , \Level1Out135[29] , \Level1Out135[28] , 
        \Level1Out135[27] , \Level1Out135[26] , \Level1Out135[25] , 
        \Level1Out135[24] , \Level1Out135[23] , \Level1Out135[22] , 
        \Level1Out135[21] , \Level1Out135[20] , \Level1Out135[19] , 
        \Level1Out135[18] , \Level1Out135[17] , \Level1Out135[16] , 
        \Level1Out135[15] , \Level1Out135[14] , \Level1Out135[13] , 
        \Level1Out135[12] , \Level1Out135[11] , \Level1Out135[10] , 
        \Level1Out135[9] , \Level1Out135[8] , \Level1Out135[7] , 
        \Level1Out135[6] , \Level1Out135[5] , \Level1Out135[4] , 
        \Level1Out135[3] , \Level1Out135[2] , \Level1Out135[1] , 
        \Level1Out135[0] }), .Read1(\Level1Load134[0] ), .Read2(
        \Level1Load135[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_190_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load190[0] ), .Out({\Level2Out190[31] , \Level2Out190[30] , 
        \Level2Out190[29] , \Level2Out190[28] , \Level2Out190[27] , 
        \Level2Out190[26] , \Level2Out190[25] , \Level2Out190[24] , 
        \Level2Out190[23] , \Level2Out190[22] , \Level2Out190[21] , 
        \Level2Out190[20] , \Level2Out190[19] , \Level2Out190[18] , 
        \Level2Out190[17] , \Level2Out190[16] , \Level2Out190[15] , 
        \Level2Out190[14] , \Level2Out190[13] , \Level2Out190[12] , 
        \Level2Out190[11] , \Level2Out190[10] , \Level2Out190[9] , 
        \Level2Out190[8] , \Level2Out190[7] , \Level2Out190[6] , 
        \Level2Out190[5] , \Level2Out190[4] , \Level2Out190[3] , 
        \Level2Out190[2] , \Level2Out190[1] , \Level2Out190[0] }), .In1({
        \Level1Out190[31] , \Level1Out190[30] , \Level1Out190[29] , 
        \Level1Out190[28] , \Level1Out190[27] , \Level1Out190[26] , 
        \Level1Out190[25] , \Level1Out190[24] , \Level1Out190[23] , 
        \Level1Out190[22] , \Level1Out190[21] , \Level1Out190[20] , 
        \Level1Out190[19] , \Level1Out190[18] , \Level1Out190[17] , 
        \Level1Out190[16] , \Level1Out190[15] , \Level1Out190[14] , 
        \Level1Out190[13] , \Level1Out190[12] , \Level1Out190[11] , 
        \Level1Out190[10] , \Level1Out190[9] , \Level1Out190[8] , 
        \Level1Out190[7] , \Level1Out190[6] , \Level1Out190[5] , 
        \Level1Out190[4] , \Level1Out190[3] , \Level1Out190[2] , 
        \Level1Out190[1] , \Level1Out190[0] }), .In2({\Level1Out191[31] , 
        \Level1Out191[30] , \Level1Out191[29] , \Level1Out191[28] , 
        \Level1Out191[27] , \Level1Out191[26] , \Level1Out191[25] , 
        \Level1Out191[24] , \Level1Out191[23] , \Level1Out191[22] , 
        \Level1Out191[21] , \Level1Out191[20] , \Level1Out191[19] , 
        \Level1Out191[18] , \Level1Out191[17] , \Level1Out191[16] , 
        \Level1Out191[15] , \Level1Out191[14] , \Level1Out191[13] , 
        \Level1Out191[12] , \Level1Out191[11] , \Level1Out191[10] , 
        \Level1Out191[9] , \Level1Out191[8] , \Level1Out191[7] , 
        \Level1Out191[6] , \Level1Out191[5] , \Level1Out191[4] , 
        \Level1Out191[3] , \Level1Out191[2] , \Level1Out191[1] , 
        \Level1Out191[0] }), .Read1(\Level1Load190[0] ), .Read2(
        \Level1Load191[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load128[0] ), .Out({\Level4Out128[31] , \Level4Out128[30] , 
        \Level4Out128[29] , \Level4Out128[28] , \Level4Out128[27] , 
        \Level4Out128[26] , \Level4Out128[25] , \Level4Out128[24] , 
        \Level4Out128[23] , \Level4Out128[22] , \Level4Out128[21] , 
        \Level4Out128[20] , \Level4Out128[19] , \Level4Out128[18] , 
        \Level4Out128[17] , \Level4Out128[16] , \Level4Out128[15] , 
        \Level4Out128[14] , \Level4Out128[13] , \Level4Out128[12] , 
        \Level4Out128[11] , \Level4Out128[10] , \Level4Out128[9] , 
        \Level4Out128[8] , \Level4Out128[7] , \Level4Out128[6] , 
        \Level4Out128[5] , \Level4Out128[4] , \Level4Out128[3] , 
        \Level4Out128[2] , \Level4Out128[1] , \Level4Out128[0] }), .In1({
        \Level2Out128[31] , \Level2Out128[30] , \Level2Out128[29] , 
        \Level2Out128[28] , \Level2Out128[27] , \Level2Out128[26] , 
        \Level2Out128[25] , \Level2Out128[24] , \Level2Out128[23] , 
        \Level2Out128[22] , \Level2Out128[21] , \Level2Out128[20] , 
        \Level2Out128[19] , \Level2Out128[18] , \Level2Out128[17] , 
        \Level2Out128[16] , \Level2Out128[15] , \Level2Out128[14] , 
        \Level2Out128[13] , \Level2Out128[12] , \Level2Out128[11] , 
        \Level2Out128[10] , \Level2Out128[9] , \Level2Out128[8] , 
        \Level2Out128[7] , \Level2Out128[6] , \Level2Out128[5] , 
        \Level2Out128[4] , \Level2Out128[3] , \Level2Out128[2] , 
        \Level2Out128[1] , \Level2Out128[0] }), .In2({\Level2Out130[31] , 
        \Level2Out130[30] , \Level2Out130[29] , \Level2Out130[28] , 
        \Level2Out130[27] , \Level2Out130[26] , \Level2Out130[25] , 
        \Level2Out130[24] , \Level2Out130[23] , \Level2Out130[22] , 
        \Level2Out130[21] , \Level2Out130[20] , \Level2Out130[19] , 
        \Level2Out130[18] , \Level2Out130[17] , \Level2Out130[16] , 
        \Level2Out130[15] , \Level2Out130[14] , \Level2Out130[13] , 
        \Level2Out130[12] , \Level2Out130[11] , \Level2Out130[10] , 
        \Level2Out130[9] , \Level2Out130[8] , \Level2Out130[7] , 
        \Level2Out130[6] , \Level2Out130[5] , \Level2Out130[4] , 
        \Level2Out130[3] , \Level2Out130[2] , \Level2Out130[1] , 
        \Level2Out130[0] }), .Read1(\Level2Load128[0] ), .Read2(
        \Level2Load130[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_236_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load236[0] ), .Out({\Level4Out236[31] , \Level4Out236[30] , 
        \Level4Out236[29] , \Level4Out236[28] , \Level4Out236[27] , 
        \Level4Out236[26] , \Level4Out236[25] , \Level4Out236[24] , 
        \Level4Out236[23] , \Level4Out236[22] , \Level4Out236[21] , 
        \Level4Out236[20] , \Level4Out236[19] , \Level4Out236[18] , 
        \Level4Out236[17] , \Level4Out236[16] , \Level4Out236[15] , 
        \Level4Out236[14] , \Level4Out236[13] , \Level4Out236[12] , 
        \Level4Out236[11] , \Level4Out236[10] , \Level4Out236[9] , 
        \Level4Out236[8] , \Level4Out236[7] , \Level4Out236[6] , 
        \Level4Out236[5] , \Level4Out236[4] , \Level4Out236[3] , 
        \Level4Out236[2] , \Level4Out236[1] , \Level4Out236[0] }), .In1({
        \Level2Out236[31] , \Level2Out236[30] , \Level2Out236[29] , 
        \Level2Out236[28] , \Level2Out236[27] , \Level2Out236[26] , 
        \Level2Out236[25] , \Level2Out236[24] , \Level2Out236[23] , 
        \Level2Out236[22] , \Level2Out236[21] , \Level2Out236[20] , 
        \Level2Out236[19] , \Level2Out236[18] , \Level2Out236[17] , 
        \Level2Out236[16] , \Level2Out236[15] , \Level2Out236[14] , 
        \Level2Out236[13] , \Level2Out236[12] , \Level2Out236[11] , 
        \Level2Out236[10] , \Level2Out236[9] , \Level2Out236[8] , 
        \Level2Out236[7] , \Level2Out236[6] , \Level2Out236[5] , 
        \Level2Out236[4] , \Level2Out236[3] , \Level2Out236[2] , 
        \Level2Out236[1] , \Level2Out236[0] }), .In2({\Level2Out238[31] , 
        \Level2Out238[30] , \Level2Out238[29] , \Level2Out238[28] , 
        \Level2Out238[27] , \Level2Out238[26] , \Level2Out238[25] , 
        \Level2Out238[24] , \Level2Out238[23] , \Level2Out238[22] , 
        \Level2Out238[21] , \Level2Out238[20] , \Level2Out238[19] , 
        \Level2Out238[18] , \Level2Out238[17] , \Level2Out238[16] , 
        \Level2Out238[15] , \Level2Out238[14] , \Level2Out238[13] , 
        \Level2Out238[12] , \Level2Out238[11] , \Level2Out238[10] , 
        \Level2Out238[9] , \Level2Out238[8] , \Level2Out238[7] , 
        \Level2Out238[6] , \Level2Out238[5] , \Level2Out238[4] , 
        \Level2Out238[3] , \Level2Out238[2] , \Level2Out238[1] , 
        \Level2Out238[0] }), .Read1(\Level2Load236[0] ), .Read2(
        \Level2Load238[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_48 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanOut({\ScanLink49[31] , 
        \ScanLink49[30] , \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , 
        \ScanLink49[26] , \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , 
        \ScanLink49[22] , \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , 
        \ScanLink49[18] , \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , 
        \ScanLink49[14] , \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , 
        \ScanLink49[10] , \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , 
        \ScanLink49[6] , \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , 
        \ScanLink49[2] , \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load48[0] ), .Out({
        \Level1Out48[31] , \Level1Out48[30] , \Level1Out48[29] , 
        \Level1Out48[28] , \Level1Out48[27] , \Level1Out48[26] , 
        \Level1Out48[25] , \Level1Out48[24] , \Level1Out48[23] , 
        \Level1Out48[22] , \Level1Out48[21] , \Level1Out48[20] , 
        \Level1Out48[19] , \Level1Out48[18] , \Level1Out48[17] , 
        \Level1Out48[16] , \Level1Out48[15] , \Level1Out48[14] , 
        \Level1Out48[13] , \Level1Out48[12] , \Level1Out48[11] , 
        \Level1Out48[10] , \Level1Out48[9] , \Level1Out48[8] , 
        \Level1Out48[7] , \Level1Out48[6] , \Level1Out48[5] , \Level1Out48[4] , 
        \Level1Out48[3] , \Level1Out48[2] , \Level1Out48[1] , \Level1Out48[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_53 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanOut({\ScanLink54[31] , 
        \ScanLink54[30] , \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , 
        \ScanLink54[26] , \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , 
        \ScanLink54[22] , \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , 
        \ScanLink54[18] , \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , 
        \ScanLink54[14] , \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , 
        \ScanLink54[10] , \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , 
        \ScanLink54[6] , \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , 
        \ScanLink54[2] , \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load53[0] ), .Out({
        \Level1Out53[31] , \Level1Out53[30] , \Level1Out53[29] , 
        \Level1Out53[28] , \Level1Out53[27] , \Level1Out53[26] , 
        \Level1Out53[25] , \Level1Out53[24] , \Level1Out53[23] , 
        \Level1Out53[22] , \Level1Out53[21] , \Level1Out53[20] , 
        \Level1Out53[19] , \Level1Out53[18] , \Level1Out53[17] , 
        \Level1Out53[16] , \Level1Out53[15] , \Level1Out53[14] , 
        \Level1Out53[13] , \Level1Out53[12] , \Level1Out53[11] , 
        \Level1Out53[10] , \Level1Out53[9] , \Level1Out53[8] , 
        \Level1Out53[7] , \Level1Out53[6] , \Level1Out53[5] , \Level1Out53[4] , 
        \Level1Out53[3] , \Level1Out53[2] , \Level1Out53[1] , \Level1Out53[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_66 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink66[31] , \ScanLink66[30] , 
        \ScanLink66[29] , \ScanLink66[28] , \ScanLink66[27] , \ScanLink66[26] , 
        \ScanLink66[25] , \ScanLink66[24] , \ScanLink66[23] , \ScanLink66[22] , 
        \ScanLink66[21] , \ScanLink66[20] , \ScanLink66[19] , \ScanLink66[18] , 
        \ScanLink66[17] , \ScanLink66[16] , \ScanLink66[15] , \ScanLink66[14] , 
        \ScanLink66[13] , \ScanLink66[12] , \ScanLink66[11] , \ScanLink66[10] , 
        \ScanLink66[9] , \ScanLink66[8] , \ScanLink66[7] , \ScanLink66[6] , 
        \ScanLink66[5] , \ScanLink66[4] , \ScanLink66[3] , \ScanLink66[2] , 
        \ScanLink66[1] , \ScanLink66[0] }), .ScanOut({\ScanLink67[31] , 
        \ScanLink67[30] , \ScanLink67[29] , \ScanLink67[28] , \ScanLink67[27] , 
        \ScanLink67[26] , \ScanLink67[25] , \ScanLink67[24] , \ScanLink67[23] , 
        \ScanLink67[22] , \ScanLink67[21] , \ScanLink67[20] , \ScanLink67[19] , 
        \ScanLink67[18] , \ScanLink67[17] , \ScanLink67[16] , \ScanLink67[15] , 
        \ScanLink67[14] , \ScanLink67[13] , \ScanLink67[12] , \ScanLink67[11] , 
        \ScanLink67[10] , \ScanLink67[9] , \ScanLink67[8] , \ScanLink67[7] , 
        \ScanLink67[6] , \ScanLink67[5] , \ScanLink67[4] , \ScanLink67[3] , 
        \ScanLink67[2] , \ScanLink67[1] , \ScanLink67[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load66[0] ), .Out({
        \Level1Out66[31] , \Level1Out66[30] , \Level1Out66[29] , 
        \Level1Out66[28] , \Level1Out66[27] , \Level1Out66[26] , 
        \Level1Out66[25] , \Level1Out66[24] , \Level1Out66[23] , 
        \Level1Out66[22] , \Level1Out66[21] , \Level1Out66[20] , 
        \Level1Out66[19] , \Level1Out66[18] , \Level1Out66[17] , 
        \Level1Out66[16] , \Level1Out66[15] , \Level1Out66[14] , 
        \Level1Out66[13] , \Level1Out66[12] , \Level1Out66[11] , 
        \Level1Out66[10] , \Level1Out66[9] , \Level1Out66[8] , 
        \Level1Out66[7] , \Level1Out66[6] , \Level1Out66[5] , \Level1Out66[4] , 
        \Level1Out66[3] , \Level1Out66[2] , \Level1Out66[1] , \Level1Out66[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_83 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink83[31] , \ScanLink83[30] , 
        \ScanLink83[29] , \ScanLink83[28] , \ScanLink83[27] , \ScanLink83[26] , 
        \ScanLink83[25] , \ScanLink83[24] , \ScanLink83[23] , \ScanLink83[22] , 
        \ScanLink83[21] , \ScanLink83[20] , \ScanLink83[19] , \ScanLink83[18] , 
        \ScanLink83[17] , \ScanLink83[16] , \ScanLink83[15] , \ScanLink83[14] , 
        \ScanLink83[13] , \ScanLink83[12] , \ScanLink83[11] , \ScanLink83[10] , 
        \ScanLink83[9] , \ScanLink83[8] , \ScanLink83[7] , \ScanLink83[6] , 
        \ScanLink83[5] , \ScanLink83[4] , \ScanLink83[3] , \ScanLink83[2] , 
        \ScanLink83[1] , \ScanLink83[0] }), .ScanOut({\ScanLink84[31] , 
        \ScanLink84[30] , \ScanLink84[29] , \ScanLink84[28] , \ScanLink84[27] , 
        \ScanLink84[26] , \ScanLink84[25] , \ScanLink84[24] , \ScanLink84[23] , 
        \ScanLink84[22] , \ScanLink84[21] , \ScanLink84[20] , \ScanLink84[19] , 
        \ScanLink84[18] , \ScanLink84[17] , \ScanLink84[16] , \ScanLink84[15] , 
        \ScanLink84[14] , \ScanLink84[13] , \ScanLink84[12] , \ScanLink84[11] , 
        \ScanLink84[10] , \ScanLink84[9] , \ScanLink84[8] , \ScanLink84[7] , 
        \ScanLink84[6] , \ScanLink84[5] , \ScanLink84[4] , \ScanLink84[3] , 
        \ScanLink84[2] , \ScanLink84[1] , \ScanLink84[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load83[0] ), .Out({
        \Level1Out83[31] , \Level1Out83[30] , \Level1Out83[29] , 
        \Level1Out83[28] , \Level1Out83[27] , \Level1Out83[26] , 
        \Level1Out83[25] , \Level1Out83[24] , \Level1Out83[23] , 
        \Level1Out83[22] , \Level1Out83[21] , \Level1Out83[20] , 
        \Level1Out83[19] , \Level1Out83[18] , \Level1Out83[17] , 
        \Level1Out83[16] , \Level1Out83[15] , \Level1Out83[14] , 
        \Level1Out83[13] , \Level1Out83[12] , \Level1Out83[11] , 
        \Level1Out83[10] , \Level1Out83[9] , \Level1Out83[8] , 
        \Level1Out83[7] , \Level1Out83[6] , \Level1Out83[5] , \Level1Out83[4] , 
        \Level1Out83[3] , \Level1Out83[2] , \Level1Out83[1] , \Level1Out83[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_144 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink144[31] , \ScanLink144[30] , 
        \ScanLink144[29] , \ScanLink144[28] , \ScanLink144[27] , 
        \ScanLink144[26] , \ScanLink144[25] , \ScanLink144[24] , 
        \ScanLink144[23] , \ScanLink144[22] , \ScanLink144[21] , 
        \ScanLink144[20] , \ScanLink144[19] , \ScanLink144[18] , 
        \ScanLink144[17] , \ScanLink144[16] , \ScanLink144[15] , 
        \ScanLink144[14] , \ScanLink144[13] , \ScanLink144[12] , 
        \ScanLink144[11] , \ScanLink144[10] , \ScanLink144[9] , 
        \ScanLink144[8] , \ScanLink144[7] , \ScanLink144[6] , \ScanLink144[5] , 
        \ScanLink144[4] , \ScanLink144[3] , \ScanLink144[2] , \ScanLink144[1] , 
        \ScanLink144[0] }), .ScanOut({\ScanLink145[31] , \ScanLink145[30] , 
        \ScanLink145[29] , \ScanLink145[28] , \ScanLink145[27] , 
        \ScanLink145[26] , \ScanLink145[25] , \ScanLink145[24] , 
        \ScanLink145[23] , \ScanLink145[22] , \ScanLink145[21] , 
        \ScanLink145[20] , \ScanLink145[19] , \ScanLink145[18] , 
        \ScanLink145[17] , \ScanLink145[16] , \ScanLink145[15] , 
        \ScanLink145[14] , \ScanLink145[13] , \ScanLink145[12] , 
        \ScanLink145[11] , \ScanLink145[10] , \ScanLink145[9] , 
        \ScanLink145[8] , \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , 
        \ScanLink145[4] , \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , 
        \ScanLink145[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load144[0] ), .Out({\Level1Out144[31] , \Level1Out144[30] , 
        \Level1Out144[29] , \Level1Out144[28] , \Level1Out144[27] , 
        \Level1Out144[26] , \Level1Out144[25] , \Level1Out144[24] , 
        \Level1Out144[23] , \Level1Out144[22] , \Level1Out144[21] , 
        \Level1Out144[20] , \Level1Out144[19] , \Level1Out144[18] , 
        \Level1Out144[17] , \Level1Out144[16] , \Level1Out144[15] , 
        \Level1Out144[14] , \Level1Out144[13] , \Level1Out144[12] , 
        \Level1Out144[11] , \Level1Out144[10] , \Level1Out144[9] , 
        \Level1Out144[8] , \Level1Out144[7] , \Level1Out144[6] , 
        \Level1Out144[5] , \Level1Out144[4] , \Level1Out144[3] , 
        \Level1Out144[2] , \Level1Out144[1] , \Level1Out144[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_76_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load76[0] ), .Out({\Level4Out76[31] , \Level4Out76[30] , 
        \Level4Out76[29] , \Level4Out76[28] , \Level4Out76[27] , 
        \Level4Out76[26] , \Level4Out76[25] , \Level4Out76[24] , 
        \Level4Out76[23] , \Level4Out76[22] , \Level4Out76[21] , 
        \Level4Out76[20] , \Level4Out76[19] , \Level4Out76[18] , 
        \Level4Out76[17] , \Level4Out76[16] , \Level4Out76[15] , 
        \Level4Out76[14] , \Level4Out76[13] , \Level4Out76[12] , 
        \Level4Out76[11] , \Level4Out76[10] , \Level4Out76[9] , 
        \Level4Out76[8] , \Level4Out76[7] , \Level4Out76[6] , \Level4Out76[5] , 
        \Level4Out76[4] , \Level4Out76[3] , \Level4Out76[2] , \Level4Out76[1] , 
        \Level4Out76[0] }), .In1({\Level2Out76[31] , \Level2Out76[30] , 
        \Level2Out76[29] , \Level2Out76[28] , \Level2Out76[27] , 
        \Level2Out76[26] , \Level2Out76[25] , \Level2Out76[24] , 
        \Level2Out76[23] , \Level2Out76[22] , \Level2Out76[21] , 
        \Level2Out76[20] , \Level2Out76[19] , \Level2Out76[18] , 
        \Level2Out76[17] , \Level2Out76[16] , \Level2Out76[15] , 
        \Level2Out76[14] , \Level2Out76[13] , \Level2Out76[12] , 
        \Level2Out76[11] , \Level2Out76[10] , \Level2Out76[9] , 
        \Level2Out76[8] , \Level2Out76[7] , \Level2Out76[6] , \Level2Out76[5] , 
        \Level2Out76[4] , \Level2Out76[3] , \Level2Out76[2] , \Level2Out76[1] , 
        \Level2Out76[0] }), .In2({\Level2Out78[31] , \Level2Out78[30] , 
        \Level2Out78[29] , \Level2Out78[28] , \Level2Out78[27] , 
        \Level2Out78[26] , \Level2Out78[25] , \Level2Out78[24] , 
        \Level2Out78[23] , \Level2Out78[22] , \Level2Out78[21] , 
        \Level2Out78[20] , \Level2Out78[19] , \Level2Out78[18] , 
        \Level2Out78[17] , \Level2Out78[16] , \Level2Out78[15] , 
        \Level2Out78[14] , \Level2Out78[13] , \Level2Out78[12] , 
        \Level2Out78[11] , \Level2Out78[10] , \Level2Out78[9] , 
        \Level2Out78[8] , \Level2Out78[7] , \Level2Out78[6] , \Level2Out78[5] , 
        \Level2Out78[4] , \Level2Out78[3] , \Level2Out78[2] , \Level2Out78[1] , 
        \Level2Out78[0] }), .Read1(\Level2Load76[0] ), .Read2(
        \Level2Load78[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_163 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink163[31] , \ScanLink163[30] , 
        \ScanLink163[29] , \ScanLink163[28] , \ScanLink163[27] , 
        \ScanLink163[26] , \ScanLink163[25] , \ScanLink163[24] , 
        \ScanLink163[23] , \ScanLink163[22] , \ScanLink163[21] , 
        \ScanLink163[20] , \ScanLink163[19] , \ScanLink163[18] , 
        \ScanLink163[17] , \ScanLink163[16] , \ScanLink163[15] , 
        \ScanLink163[14] , \ScanLink163[13] , \ScanLink163[12] , 
        \ScanLink163[11] , \ScanLink163[10] , \ScanLink163[9] , 
        \ScanLink163[8] , \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , 
        \ScanLink163[4] , \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , 
        \ScanLink163[0] }), .ScanOut({\ScanLink164[31] , \ScanLink164[30] , 
        \ScanLink164[29] , \ScanLink164[28] , \ScanLink164[27] , 
        \ScanLink164[26] , \ScanLink164[25] , \ScanLink164[24] , 
        \ScanLink164[23] , \ScanLink164[22] , \ScanLink164[21] , 
        \ScanLink164[20] , \ScanLink164[19] , \ScanLink164[18] , 
        \ScanLink164[17] , \ScanLink164[16] , \ScanLink164[15] , 
        \ScanLink164[14] , \ScanLink164[13] , \ScanLink164[12] , 
        \ScanLink164[11] , \ScanLink164[10] , \ScanLink164[9] , 
        \ScanLink164[8] , \ScanLink164[7] , \ScanLink164[6] , \ScanLink164[5] , 
        \ScanLink164[4] , \ScanLink164[3] , \ScanLink164[2] , \ScanLink164[1] , 
        \ScanLink164[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load163[0] ), .Out({\Level1Out163[31] , \Level1Out163[30] , 
        \Level1Out163[29] , \Level1Out163[28] , \Level1Out163[27] , 
        \Level1Out163[26] , \Level1Out163[25] , \Level1Out163[24] , 
        \Level1Out163[23] , \Level1Out163[22] , \Level1Out163[21] , 
        \Level1Out163[20] , \Level1Out163[19] , \Level1Out163[18] , 
        \Level1Out163[17] , \Level1Out163[16] , \Level1Out163[15] , 
        \Level1Out163[14] , \Level1Out163[13] , \Level1Out163[12] , 
        \Level1Out163[11] , \Level1Out163[10] , \Level1Out163[9] , 
        \Level1Out163[8] , \Level1Out163[7] , \Level1Out163[6] , 
        \Level1Out163[5] , \Level1Out163[4] , \Level1Out163[3] , 
        \Level1Out163[2] , \Level1Out163[1] , \Level1Out163[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_106_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load106[0] ), .Out({\Level2Out106[31] , \Level2Out106[30] , 
        \Level2Out106[29] , \Level2Out106[28] , \Level2Out106[27] , 
        \Level2Out106[26] , \Level2Out106[25] , \Level2Out106[24] , 
        \Level2Out106[23] , \Level2Out106[22] , \Level2Out106[21] , 
        \Level2Out106[20] , \Level2Out106[19] , \Level2Out106[18] , 
        \Level2Out106[17] , \Level2Out106[16] , \Level2Out106[15] , 
        \Level2Out106[14] , \Level2Out106[13] , \Level2Out106[12] , 
        \Level2Out106[11] , \Level2Out106[10] , \Level2Out106[9] , 
        \Level2Out106[8] , \Level2Out106[7] , \Level2Out106[6] , 
        \Level2Out106[5] , \Level2Out106[4] , \Level2Out106[3] , 
        \Level2Out106[2] , \Level2Out106[1] , \Level2Out106[0] }), .In1({
        \Level1Out106[31] , \Level1Out106[30] , \Level1Out106[29] , 
        \Level1Out106[28] , \Level1Out106[27] , \Level1Out106[26] , 
        \Level1Out106[25] , \Level1Out106[24] , \Level1Out106[23] , 
        \Level1Out106[22] , \Level1Out106[21] , \Level1Out106[20] , 
        \Level1Out106[19] , \Level1Out106[18] , \Level1Out106[17] , 
        \Level1Out106[16] , \Level1Out106[15] , \Level1Out106[14] , 
        \Level1Out106[13] , \Level1Out106[12] , \Level1Out106[11] , 
        \Level1Out106[10] , \Level1Out106[9] , \Level1Out106[8] , 
        \Level1Out106[7] , \Level1Out106[6] , \Level1Out106[5] , 
        \Level1Out106[4] , \Level1Out106[3] , \Level1Out106[2] , 
        \Level1Out106[1] , \Level1Out106[0] }), .In2({\Level1Out107[31] , 
        \Level1Out107[30] , \Level1Out107[29] , \Level1Out107[28] , 
        \Level1Out107[27] , \Level1Out107[26] , \Level1Out107[25] , 
        \Level1Out107[24] , \Level1Out107[23] , \Level1Out107[22] , 
        \Level1Out107[21] , \Level1Out107[20] , \Level1Out107[19] , 
        \Level1Out107[18] , \Level1Out107[17] , \Level1Out107[16] , 
        \Level1Out107[15] , \Level1Out107[14] , \Level1Out107[13] , 
        \Level1Out107[12] , \Level1Out107[11] , \Level1Out107[10] , 
        \Level1Out107[9] , \Level1Out107[8] , \Level1Out107[7] , 
        \Level1Out107[6] , \Level1Out107[5] , \Level1Out107[4] , 
        \Level1Out107[3] , \Level1Out107[2] , \Level1Out107[1] , 
        \Level1Out107[0] }), .Read1(\Level1Load106[0] ), .Read2(
        \Level1Load107[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_218_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load218[0] ), .Out({\Level2Out218[31] , \Level2Out218[30] , 
        \Level2Out218[29] , \Level2Out218[28] , \Level2Out218[27] , 
        \Level2Out218[26] , \Level2Out218[25] , \Level2Out218[24] , 
        \Level2Out218[23] , \Level2Out218[22] , \Level2Out218[21] , 
        \Level2Out218[20] , \Level2Out218[19] , \Level2Out218[18] , 
        \Level2Out218[17] , \Level2Out218[16] , \Level2Out218[15] , 
        \Level2Out218[14] , \Level2Out218[13] , \Level2Out218[12] , 
        \Level2Out218[11] , \Level2Out218[10] , \Level2Out218[9] , 
        \Level2Out218[8] , \Level2Out218[7] , \Level2Out218[6] , 
        \Level2Out218[5] , \Level2Out218[4] , \Level2Out218[3] , 
        \Level2Out218[2] , \Level2Out218[1] , \Level2Out218[0] }), .In1({
        \Level1Out218[31] , \Level1Out218[30] , \Level1Out218[29] , 
        \Level1Out218[28] , \Level1Out218[27] , \Level1Out218[26] , 
        \Level1Out218[25] , \Level1Out218[24] , \Level1Out218[23] , 
        \Level1Out218[22] , \Level1Out218[21] , \Level1Out218[20] , 
        \Level1Out218[19] , \Level1Out218[18] , \Level1Out218[17] , 
        \Level1Out218[16] , \Level1Out218[15] , \Level1Out218[14] , 
        \Level1Out218[13] , \Level1Out218[12] , \Level1Out218[11] , 
        \Level1Out218[10] , \Level1Out218[9] , \Level1Out218[8] , 
        \Level1Out218[7] , \Level1Out218[6] , \Level1Out218[5] , 
        \Level1Out218[4] , \Level1Out218[3] , \Level1Out218[2] , 
        \Level1Out218[1] , \Level1Out218[0] }), .In2({\Level1Out219[31] , 
        \Level1Out219[30] , \Level1Out219[29] , \Level1Out219[28] , 
        \Level1Out219[27] , \Level1Out219[26] , \Level1Out219[25] , 
        \Level1Out219[24] , \Level1Out219[23] , \Level1Out219[22] , 
        \Level1Out219[21] , \Level1Out219[20] , \Level1Out219[19] , 
        \Level1Out219[18] , \Level1Out219[17] , \Level1Out219[16] , 
        \Level1Out219[15] , \Level1Out219[14] , \Level1Out219[13] , 
        \Level1Out219[12] , \Level1Out219[11] , \Level1Out219[10] , 
        \Level1Out219[9] , \Level1Out219[8] , \Level1Out219[7] , 
        \Level1Out219[6] , \Level1Out219[5] , \Level1Out219[4] , 
        \Level1Out219[3] , \Level1Out219[2] , \Level1Out219[1] , 
        \Level1Out219[0] }), .Read1(\Level1Load218[0] ), .Read2(
        \Level1Load219[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_204_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load204[0] ), .Out({\Level4Out204[31] , \Level4Out204[30] , 
        \Level4Out204[29] , \Level4Out204[28] , \Level4Out204[27] , 
        \Level4Out204[26] , \Level4Out204[25] , \Level4Out204[24] , 
        \Level4Out204[23] , \Level4Out204[22] , \Level4Out204[21] , 
        \Level4Out204[20] , \Level4Out204[19] , \Level4Out204[18] , 
        \Level4Out204[17] , \Level4Out204[16] , \Level4Out204[15] , 
        \Level4Out204[14] , \Level4Out204[13] , \Level4Out204[12] , 
        \Level4Out204[11] , \Level4Out204[10] , \Level4Out204[9] , 
        \Level4Out204[8] , \Level4Out204[7] , \Level4Out204[6] , 
        \Level4Out204[5] , \Level4Out204[4] , \Level4Out204[3] , 
        \Level4Out204[2] , \Level4Out204[1] , \Level4Out204[0] }), .In1({
        \Level2Out204[31] , \Level2Out204[30] , \Level2Out204[29] , 
        \Level2Out204[28] , \Level2Out204[27] , \Level2Out204[26] , 
        \Level2Out204[25] , \Level2Out204[24] , \Level2Out204[23] , 
        \Level2Out204[22] , \Level2Out204[21] , \Level2Out204[20] , 
        \Level2Out204[19] , \Level2Out204[18] , \Level2Out204[17] , 
        \Level2Out204[16] , \Level2Out204[15] , \Level2Out204[14] , 
        \Level2Out204[13] , \Level2Out204[12] , \Level2Out204[11] , 
        \Level2Out204[10] , \Level2Out204[9] , \Level2Out204[8] , 
        \Level2Out204[7] , \Level2Out204[6] , \Level2Out204[5] , 
        \Level2Out204[4] , \Level2Out204[3] , \Level2Out204[2] , 
        \Level2Out204[1] , \Level2Out204[0] }), .In2({\Level2Out206[31] , 
        \Level2Out206[30] , \Level2Out206[29] , \Level2Out206[28] , 
        \Level2Out206[27] , \Level2Out206[26] , \Level2Out206[25] , 
        \Level2Out206[24] , \Level2Out206[23] , \Level2Out206[22] , 
        \Level2Out206[21] , \Level2Out206[20] , \Level2Out206[19] , 
        \Level2Out206[18] , \Level2Out206[17] , \Level2Out206[16] , 
        \Level2Out206[15] , \Level2Out206[14] , \Level2Out206[13] , 
        \Level2Out206[12] , \Level2Out206[11] , \Level2Out206[10] , 
        \Level2Out206[9] , \Level2Out206[8] , \Level2Out206[7] , 
        \Level2Out206[6] , \Level2Out206[5] , \Level2Out206[4] , 
        \Level2Out206[3] , \Level2Out206[2] , \Level2Out206[1] , 
        \Level2Out206[0] }), .Read1(\Level2Load204[0] ), .Read2(
        \Level2Load206[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_253 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink253[31] , \ScanLink253[30] , 
        \ScanLink253[29] , \ScanLink253[28] , \ScanLink253[27] , 
        \ScanLink253[26] , \ScanLink253[25] , \ScanLink253[24] , 
        \ScanLink253[23] , \ScanLink253[22] , \ScanLink253[21] , 
        \ScanLink253[20] , \ScanLink253[19] , \ScanLink253[18] , 
        \ScanLink253[17] , \ScanLink253[16] , \ScanLink253[15] , 
        \ScanLink253[14] , \ScanLink253[13] , \ScanLink253[12] , 
        \ScanLink253[11] , \ScanLink253[10] , \ScanLink253[9] , 
        \ScanLink253[8] , \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , 
        \ScanLink253[4] , \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , 
        \ScanLink253[0] }), .ScanOut({\ScanLink254[31] , \ScanLink254[30] , 
        \ScanLink254[29] , \ScanLink254[28] , \ScanLink254[27] , 
        \ScanLink254[26] , \ScanLink254[25] , \ScanLink254[24] , 
        \ScanLink254[23] , \ScanLink254[22] , \ScanLink254[21] , 
        \ScanLink254[20] , \ScanLink254[19] , \ScanLink254[18] , 
        \ScanLink254[17] , \ScanLink254[16] , \ScanLink254[15] , 
        \ScanLink254[14] , \ScanLink254[13] , \ScanLink254[12] , 
        \ScanLink254[11] , \ScanLink254[10] , \ScanLink254[9] , 
        \ScanLink254[8] , \ScanLink254[7] , \ScanLink254[6] , \ScanLink254[5] , 
        \ScanLink254[4] , \ScanLink254[3] , \ScanLink254[2] , \ScanLink254[1] , 
        \ScanLink254[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load253[0] ), .Out({\Level1Out253[31] , \Level1Out253[30] , 
        \Level1Out253[29] , \Level1Out253[28] , \Level1Out253[27] , 
        \Level1Out253[26] , \Level1Out253[25] , \Level1Out253[24] , 
        \Level1Out253[23] , \Level1Out253[22] , \Level1Out253[21] , 
        \Level1Out253[20] , \Level1Out253[19] , \Level1Out253[18] , 
        \Level1Out253[17] , \Level1Out253[16] , \Level1Out253[15] , 
        \Level1Out253[14] , \Level1Out253[13] , \Level1Out253[12] , 
        \Level1Out253[11] , \Level1Out253[10] , \Level1Out253[9] , 
        \Level1Out253[8] , \Level1Out253[7] , \Level1Out253[6] , 
        \Level1Out253[5] , \Level1Out253[4] , \Level1Out253[3] , 
        \Level1Out253[2] , \Level1Out253[1] , \Level1Out253[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load40[0] ), .Out({\Level2Out40[31] , \Level2Out40[30] , 
        \Level2Out40[29] , \Level2Out40[28] , \Level2Out40[27] , 
        \Level2Out40[26] , \Level2Out40[25] , \Level2Out40[24] , 
        \Level2Out40[23] , \Level2Out40[22] , \Level2Out40[21] , 
        \Level2Out40[20] , \Level2Out40[19] , \Level2Out40[18] , 
        \Level2Out40[17] , \Level2Out40[16] , \Level2Out40[15] , 
        \Level2Out40[14] , \Level2Out40[13] , \Level2Out40[12] , 
        \Level2Out40[11] , \Level2Out40[10] , \Level2Out40[9] , 
        \Level2Out40[8] , \Level2Out40[7] , \Level2Out40[6] , \Level2Out40[5] , 
        \Level2Out40[4] , \Level2Out40[3] , \Level2Out40[2] , \Level2Out40[1] , 
        \Level2Out40[0] }), .In1({\Level1Out40[31] , \Level1Out40[30] , 
        \Level1Out40[29] , \Level1Out40[28] , \Level1Out40[27] , 
        \Level1Out40[26] , \Level1Out40[25] , \Level1Out40[24] , 
        \Level1Out40[23] , \Level1Out40[22] , \Level1Out40[21] , 
        \Level1Out40[20] , \Level1Out40[19] , \Level1Out40[18] , 
        \Level1Out40[17] , \Level1Out40[16] , \Level1Out40[15] , 
        \Level1Out40[14] , \Level1Out40[13] , \Level1Out40[12] , 
        \Level1Out40[11] , \Level1Out40[10] , \Level1Out40[9] , 
        \Level1Out40[8] , \Level1Out40[7] , \Level1Out40[6] , \Level1Out40[5] , 
        \Level1Out40[4] , \Level1Out40[3] , \Level1Out40[2] , \Level1Out40[1] , 
        \Level1Out40[0] }), .In2({\Level1Out41[31] , \Level1Out41[30] , 
        \Level1Out41[29] , \Level1Out41[28] , \Level1Out41[27] , 
        \Level1Out41[26] , \Level1Out41[25] , \Level1Out41[24] , 
        \Level1Out41[23] , \Level1Out41[22] , \Level1Out41[21] , 
        \Level1Out41[20] , \Level1Out41[19] , \Level1Out41[18] , 
        \Level1Out41[17] , \Level1Out41[16] , \Level1Out41[15] , 
        \Level1Out41[14] , \Level1Out41[13] , \Level1Out41[12] , 
        \Level1Out41[11] , \Level1Out41[10] , \Level1Out41[9] , 
        \Level1Out41[8] , \Level1Out41[7] , \Level1Out41[6] , \Level1Out41[5] , 
        \Level1Out41[4] , \Level1Out41[3] , \Level1Out41[2] , \Level1Out41[1] , 
        \Level1Out41[0] }), .Read1(\Level1Load40[0] ), .Read2(
        \Level1Load41[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_232_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load232[0] ), .Out({\Level2Out232[31] , \Level2Out232[30] , 
        \Level2Out232[29] , \Level2Out232[28] , \Level2Out232[27] , 
        \Level2Out232[26] , \Level2Out232[25] , \Level2Out232[24] , 
        \Level2Out232[23] , \Level2Out232[22] , \Level2Out232[21] , 
        \Level2Out232[20] , \Level2Out232[19] , \Level2Out232[18] , 
        \Level2Out232[17] , \Level2Out232[16] , \Level2Out232[15] , 
        \Level2Out232[14] , \Level2Out232[13] , \Level2Out232[12] , 
        \Level2Out232[11] , \Level2Out232[10] , \Level2Out232[9] , 
        \Level2Out232[8] , \Level2Out232[7] , \Level2Out232[6] , 
        \Level2Out232[5] , \Level2Out232[4] , \Level2Out232[3] , 
        \Level2Out232[2] , \Level2Out232[1] , \Level2Out232[0] }), .In1({
        \Level1Out232[31] , \Level1Out232[30] , \Level1Out232[29] , 
        \Level1Out232[28] , \Level1Out232[27] , \Level1Out232[26] , 
        \Level1Out232[25] , \Level1Out232[24] , \Level1Out232[23] , 
        \Level1Out232[22] , \Level1Out232[21] , \Level1Out232[20] , 
        \Level1Out232[19] , \Level1Out232[18] , \Level1Out232[17] , 
        \Level1Out232[16] , \Level1Out232[15] , \Level1Out232[14] , 
        \Level1Out232[13] , \Level1Out232[12] , \Level1Out232[11] , 
        \Level1Out232[10] , \Level1Out232[9] , \Level1Out232[8] , 
        \Level1Out232[7] , \Level1Out232[6] , \Level1Out232[5] , 
        \Level1Out232[4] , \Level1Out232[3] , \Level1Out232[2] , 
        \Level1Out232[1] , \Level1Out232[0] }), .In2({\Level1Out233[31] , 
        \Level1Out233[30] , \Level1Out233[29] , \Level1Out233[28] , 
        \Level1Out233[27] , \Level1Out233[26] , \Level1Out233[25] , 
        \Level1Out233[24] , \Level1Out233[23] , \Level1Out233[22] , 
        \Level1Out233[21] , \Level1Out233[20] , \Level1Out233[19] , 
        \Level1Out233[18] , \Level1Out233[17] , \Level1Out233[16] , 
        \Level1Out233[15] , \Level1Out233[14] , \Level1Out233[13] , 
        \Level1Out233[12] , \Level1Out233[11] , \Level1Out233[10] , 
        \Level1Out233[9] , \Level1Out233[8] , \Level1Out233[7] , 
        \Level1Out233[6] , \Level1Out233[5] , \Level1Out233[4] , 
        \Level1Out233[3] , \Level1Out233[2] , \Level1Out233[1] , 
        \Level1Out233[0] }), .Read1(\Level1Load232[0] ), .Read2(
        \Level1Load233[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_91 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink91[31] , \ScanLink91[30] , 
        \ScanLink91[29] , \ScanLink91[28] , \ScanLink91[27] , \ScanLink91[26] , 
        \ScanLink91[25] , \ScanLink91[24] , \ScanLink91[23] , \ScanLink91[22] , 
        \ScanLink91[21] , \ScanLink91[20] , \ScanLink91[19] , \ScanLink91[18] , 
        \ScanLink91[17] , \ScanLink91[16] , \ScanLink91[15] , \ScanLink91[14] , 
        \ScanLink91[13] , \ScanLink91[12] , \ScanLink91[11] , \ScanLink91[10] , 
        \ScanLink91[9] , \ScanLink91[8] , \ScanLink91[7] , \ScanLink91[6] , 
        \ScanLink91[5] , \ScanLink91[4] , \ScanLink91[3] , \ScanLink91[2] , 
        \ScanLink91[1] , \ScanLink91[0] }), .ScanOut({\ScanLink92[31] , 
        \ScanLink92[30] , \ScanLink92[29] , \ScanLink92[28] , \ScanLink92[27] , 
        \ScanLink92[26] , \ScanLink92[25] , \ScanLink92[24] , \ScanLink92[23] , 
        \ScanLink92[22] , \ScanLink92[21] , \ScanLink92[20] , \ScanLink92[19] , 
        \ScanLink92[18] , \ScanLink92[17] , \ScanLink92[16] , \ScanLink92[15] , 
        \ScanLink92[14] , \ScanLink92[13] , \ScanLink92[12] , \ScanLink92[11] , 
        \ScanLink92[10] , \ScanLink92[9] , \ScanLink92[8] , \ScanLink92[7] , 
        \ScanLink92[6] , \ScanLink92[5] , \ScanLink92[4] , \ScanLink92[3] , 
        \ScanLink92[2] , \ScanLink92[1] , \ScanLink92[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load91[0] ), .Out({
        \Level1Out91[31] , \Level1Out91[30] , \Level1Out91[29] , 
        \Level1Out91[28] , \Level1Out91[27] , \Level1Out91[26] , 
        \Level1Out91[25] , \Level1Out91[24] , \Level1Out91[23] , 
        \Level1Out91[22] , \Level1Out91[21] , \Level1Out91[20] , 
        \Level1Out91[19] , \Level1Out91[18] , \Level1Out91[17] , 
        \Level1Out91[16] , \Level1Out91[15] , \Level1Out91[14] , 
        \Level1Out91[13] , \Level1Out91[12] , \Level1Out91[11] , 
        \Level1Out91[10] , \Level1Out91[9] , \Level1Out91[8] , 
        \Level1Out91[7] , \Level1Out91[6] , \Level1Out91[5] , \Level1Out91[4] , 
        \Level1Out91[3] , \Level1Out91[2] , \Level1Out91[1] , \Level1Out91[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_186 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink186[31] , \ScanLink186[30] , 
        \ScanLink186[29] , \ScanLink186[28] , \ScanLink186[27] , 
        \ScanLink186[26] , \ScanLink186[25] , \ScanLink186[24] , 
        \ScanLink186[23] , \ScanLink186[22] , \ScanLink186[21] , 
        \ScanLink186[20] , \ScanLink186[19] , \ScanLink186[18] , 
        \ScanLink186[17] , \ScanLink186[16] , \ScanLink186[15] , 
        \ScanLink186[14] , \ScanLink186[13] , \ScanLink186[12] , 
        \ScanLink186[11] , \ScanLink186[10] , \ScanLink186[9] , 
        \ScanLink186[8] , \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , 
        \ScanLink186[4] , \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , 
        \ScanLink186[0] }), .ScanOut({\ScanLink187[31] , \ScanLink187[30] , 
        \ScanLink187[29] , \ScanLink187[28] , \ScanLink187[27] , 
        \ScanLink187[26] , \ScanLink187[25] , \ScanLink187[24] , 
        \ScanLink187[23] , \ScanLink187[22] , \ScanLink187[21] , 
        \ScanLink187[20] , \ScanLink187[19] , \ScanLink187[18] , 
        \ScanLink187[17] , \ScanLink187[16] , \ScanLink187[15] , 
        \ScanLink187[14] , \ScanLink187[13] , \ScanLink187[12] , 
        \ScanLink187[11] , \ScanLink187[10] , \ScanLink187[9] , 
        \ScanLink187[8] , \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , 
        \ScanLink187[4] , \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , 
        \ScanLink187[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load186[0] ), .Out({\Level1Out186[31] , \Level1Out186[30] , 
        \Level1Out186[29] , \Level1Out186[28] , \Level1Out186[27] , 
        \Level1Out186[26] , \Level1Out186[25] , \Level1Out186[24] , 
        \Level1Out186[23] , \Level1Out186[22] , \Level1Out186[21] , 
        \Level1Out186[20] , \Level1Out186[19] , \Level1Out186[18] , 
        \Level1Out186[17] , \Level1Out186[16] , \Level1Out186[15] , 
        \Level1Out186[14] , \Level1Out186[13] , \Level1Out186[12] , 
        \Level1Out186[11] , \Level1Out186[10] , \Level1Out186[9] , 
        \Level1Out186[8] , \Level1Out186[7] , \Level1Out186[6] , 
        \Level1Out186[5] , \Level1Out186[4] , \Level1Out186[3] , 
        \Level1Out186[2] , \Level1Out186[1] , \Level1Out186[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_128 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level128Load128[0] ), .Out({\Level128Out128[31] , 
        \Level128Out128[30] , \Level128Out128[29] , \Level128Out128[28] , 
        \Level128Out128[27] , \Level128Out128[26] , \Level128Out128[25] , 
        \Level128Out128[24] , \Level128Out128[23] , \Level128Out128[22] , 
        \Level128Out128[21] , \Level128Out128[20] , \Level128Out128[19] , 
        \Level128Out128[18] , \Level128Out128[17] , \Level128Out128[16] , 
        \Level128Out128[15] , \Level128Out128[14] , \Level128Out128[13] , 
        \Level128Out128[12] , \Level128Out128[11] , \Level128Out128[10] , 
        \Level128Out128[9] , \Level128Out128[8] , \Level128Out128[7] , 
        \Level128Out128[6] , \Level128Out128[5] , \Level128Out128[4] , 
        \Level128Out128[3] , \Level128Out128[2] , \Level128Out128[1] , 
        \Level128Out128[0] }), .In1({\Level64Out128[31] , \Level64Out128[30] , 
        \Level64Out128[29] , \Level64Out128[28] , \Level64Out128[27] , 
        \Level64Out128[26] , \Level64Out128[25] , \Level64Out128[24] , 
        \Level64Out128[23] , \Level64Out128[22] , \Level64Out128[21] , 
        \Level64Out128[20] , \Level64Out128[19] , \Level64Out128[18] , 
        \Level64Out128[17] , \Level64Out128[16] , \Level64Out128[15] , 
        \Level64Out128[14] , \Level64Out128[13] , \Level64Out128[12] , 
        \Level64Out128[11] , \Level64Out128[10] , \Level64Out128[9] , 
        \Level64Out128[8] , \Level64Out128[7] , \Level64Out128[6] , 
        \Level64Out128[5] , \Level64Out128[4] , \Level64Out128[3] , 
        \Level64Out128[2] , \Level64Out128[1] , \Level64Out128[0] }), .In2({
        \Level64Out192[31] , \Level64Out192[30] , \Level64Out192[29] , 
        \Level64Out192[28] , \Level64Out192[27] , \Level64Out192[26] , 
        \Level64Out192[25] , \Level64Out192[24] , \Level64Out192[23] , 
        \Level64Out192[22] , \Level64Out192[21] , \Level64Out192[20] , 
        \Level64Out192[19] , \Level64Out192[18] , \Level64Out192[17] , 
        \Level64Out192[16] , \Level64Out192[15] , \Level64Out192[14] , 
        \Level64Out192[13] , \Level64Out192[12] , \Level64Out192[11] , 
        \Level64Out192[10] , \Level64Out192[9] , \Level64Out192[8] , 
        \Level64Out192[7] , \Level64Out192[6] , \Level64Out192[5] , 
        \Level64Out192[4] , \Level64Out192[3] , \Level64Out192[2] , 
        \Level64Out192[1] , \Level64Out192[0] }), .Read1(\Level64Load128[0] ), 
        .Read2(\Level64Load192[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_194 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink194[31] , \ScanLink194[30] , 
        \ScanLink194[29] , \ScanLink194[28] , \ScanLink194[27] , 
        \ScanLink194[26] , \ScanLink194[25] , \ScanLink194[24] , 
        \ScanLink194[23] , \ScanLink194[22] , \ScanLink194[21] , 
        \ScanLink194[20] , \ScanLink194[19] , \ScanLink194[18] , 
        \ScanLink194[17] , \ScanLink194[16] , \ScanLink194[15] , 
        \ScanLink194[14] , \ScanLink194[13] , \ScanLink194[12] , 
        \ScanLink194[11] , \ScanLink194[10] , \ScanLink194[9] , 
        \ScanLink194[8] , \ScanLink194[7] , \ScanLink194[6] , \ScanLink194[5] , 
        \ScanLink194[4] , \ScanLink194[3] , \ScanLink194[2] , \ScanLink194[1] , 
        \ScanLink194[0] }), .ScanOut({\ScanLink195[31] , \ScanLink195[30] , 
        \ScanLink195[29] , \ScanLink195[28] , \ScanLink195[27] , 
        \ScanLink195[26] , \ScanLink195[25] , \ScanLink195[24] , 
        \ScanLink195[23] , \ScanLink195[22] , \ScanLink195[21] , 
        \ScanLink195[20] , \ScanLink195[19] , \ScanLink195[18] , 
        \ScanLink195[17] , \ScanLink195[16] , \ScanLink195[15] , 
        \ScanLink195[14] , \ScanLink195[13] , \ScanLink195[12] , 
        \ScanLink195[11] , \ScanLink195[10] , \ScanLink195[9] , 
        \ScanLink195[8] , \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , 
        \ScanLink195[4] , \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , 
        \ScanLink195[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load194[0] ), .Out({\Level1Out194[31] , \Level1Out194[30] , 
        \Level1Out194[29] , \Level1Out194[28] , \Level1Out194[27] , 
        \Level1Out194[26] , \Level1Out194[25] , \Level1Out194[24] , 
        \Level1Out194[23] , \Level1Out194[22] , \Level1Out194[21] , 
        \Level1Out194[20] , \Level1Out194[19] , \Level1Out194[18] , 
        \Level1Out194[17] , \Level1Out194[16] , \Level1Out194[15] , 
        \Level1Out194[14] , \Level1Out194[13] , \Level1Out194[12] , 
        \Level1Out194[11] , \Level1Out194[10] , \Level1Out194[9] , 
        \Level1Out194[8] , \Level1Out194[7] , \Level1Out194[6] , 
        \Level1Out194[5] , \Level1Out194[4] , \Level1Out194[3] , 
        \Level1Out194[2] , \Level1Out194[1] , \Level1Out194[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_10_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load10[0] ), .Out({\Level2Out10[31] , \Level2Out10[30] , 
        \Level2Out10[29] , \Level2Out10[28] , \Level2Out10[27] , 
        \Level2Out10[26] , \Level2Out10[25] , \Level2Out10[24] , 
        \Level2Out10[23] , \Level2Out10[22] , \Level2Out10[21] , 
        \Level2Out10[20] , \Level2Out10[19] , \Level2Out10[18] , 
        \Level2Out10[17] , \Level2Out10[16] , \Level2Out10[15] , 
        \Level2Out10[14] , \Level2Out10[13] , \Level2Out10[12] , 
        \Level2Out10[11] , \Level2Out10[10] , \Level2Out10[9] , 
        \Level2Out10[8] , \Level2Out10[7] , \Level2Out10[6] , \Level2Out10[5] , 
        \Level2Out10[4] , \Level2Out10[3] , \Level2Out10[2] , \Level2Out10[1] , 
        \Level2Out10[0] }), .In1({\Level1Out10[31] , \Level1Out10[30] , 
        \Level1Out10[29] , \Level1Out10[28] , \Level1Out10[27] , 
        \Level1Out10[26] , \Level1Out10[25] , \Level1Out10[24] , 
        \Level1Out10[23] , \Level1Out10[22] , \Level1Out10[21] , 
        \Level1Out10[20] , \Level1Out10[19] , \Level1Out10[18] , 
        \Level1Out10[17] , \Level1Out10[16] , \Level1Out10[15] , 
        \Level1Out10[14] , \Level1Out10[13] , \Level1Out10[12] , 
        \Level1Out10[11] , \Level1Out10[10] , \Level1Out10[9] , 
        \Level1Out10[8] , \Level1Out10[7] , \Level1Out10[6] , \Level1Out10[5] , 
        \Level1Out10[4] , \Level1Out10[3] , \Level1Out10[2] , \Level1Out10[1] , 
        \Level1Out10[0] }), .In2({\Level1Out11[31] , \Level1Out11[30] , 
        \Level1Out11[29] , \Level1Out11[28] , \Level1Out11[27] , 
        \Level1Out11[26] , \Level1Out11[25] , \Level1Out11[24] , 
        \Level1Out11[23] , \Level1Out11[22] , \Level1Out11[21] , 
        \Level1Out11[20] , \Level1Out11[19] , \Level1Out11[18] , 
        \Level1Out11[17] , \Level1Out11[16] , \Level1Out11[15] , 
        \Level1Out11[14] , \Level1Out11[13] , \Level1Out11[12] , 
        \Level1Out11[11] , \Level1Out11[10] , \Level1Out11[9] , 
        \Level1Out11[8] , \Level1Out11[7] , \Level1Out11[6] , \Level1Out11[5] , 
        \Level1Out11[4] , \Level1Out11[3] , \Level1Out11[2] , \Level1Out11[1] , 
        \Level1Out11[0] }), .Read1(\Level1Load10[0] ), .Read2(
        \Level1Load11[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load4[0] ), .Out({\Level4Out4[31] , \Level4Out4[30] , 
        \Level4Out4[29] , \Level4Out4[28] , \Level4Out4[27] , \Level4Out4[26] , 
        \Level4Out4[25] , \Level4Out4[24] , \Level4Out4[23] , \Level4Out4[22] , 
        \Level4Out4[21] , \Level4Out4[20] , \Level4Out4[19] , \Level4Out4[18] , 
        \Level4Out4[17] , \Level4Out4[16] , \Level4Out4[15] , \Level4Out4[14] , 
        \Level4Out4[13] , \Level4Out4[12] , \Level4Out4[11] , \Level4Out4[10] , 
        \Level4Out4[9] , \Level4Out4[8] , \Level4Out4[7] , \Level4Out4[6] , 
        \Level4Out4[5] , \Level4Out4[4] , \Level4Out4[3] , \Level4Out4[2] , 
        \Level4Out4[1] , \Level4Out4[0] }), .In1({\Level2Out4[31] , 
        \Level2Out4[30] , \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , 
        \Level2Out4[26] , \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , 
        \Level2Out4[22] , \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , 
        \Level2Out4[18] , \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , 
        \Level2Out4[14] , \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , 
        \Level2Out4[10] , \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , 
        \Level2Out4[6] , \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , 
        \Level2Out4[2] , \Level2Out4[1] , \Level2Out4[0] }), .In2({
        \Level2Out6[31] , \Level2Out6[30] , \Level2Out6[29] , \Level2Out6[28] , 
        \Level2Out6[27] , \Level2Out6[26] , \Level2Out6[25] , \Level2Out6[24] , 
        \Level2Out6[23] , \Level2Out6[22] , \Level2Out6[21] , \Level2Out6[20] , 
        \Level2Out6[19] , \Level2Out6[18] , \Level2Out6[17] , \Level2Out6[16] , 
        \Level2Out6[15] , \Level2Out6[14] , \Level2Out6[13] , \Level2Out6[12] , 
        \Level2Out6[11] , \Level2Out6[10] , \Level2Out6[9] , \Level2Out6[8] , 
        \Level2Out6[7] , \Level2Out6[6] , \Level2Out6[5] , \Level2Out6[4] , 
        \Level2Out6[3] , \Level2Out6[2] , \Level2Out6[1] , \Level2Out6[0] }), 
        .Read1(\Level2Load4[0] ), .Read2(\Level2Load6[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_160_32 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load160[0] ), .Out({\Level32Out160[31] , \Level32Out160[30] , 
        \Level32Out160[29] , \Level32Out160[28] , \Level32Out160[27] , 
        \Level32Out160[26] , \Level32Out160[25] , \Level32Out160[24] , 
        \Level32Out160[23] , \Level32Out160[22] , \Level32Out160[21] , 
        \Level32Out160[20] , \Level32Out160[19] , \Level32Out160[18] , 
        \Level32Out160[17] , \Level32Out160[16] , \Level32Out160[15] , 
        \Level32Out160[14] , \Level32Out160[13] , \Level32Out160[12] , 
        \Level32Out160[11] , \Level32Out160[10] , \Level32Out160[9] , 
        \Level32Out160[8] , \Level32Out160[7] , \Level32Out160[6] , 
        \Level32Out160[5] , \Level32Out160[4] , \Level32Out160[3] , 
        \Level32Out160[2] , \Level32Out160[1] , \Level32Out160[0] }), .In1({
        \Level16Out160[31] , \Level16Out160[30] , \Level16Out160[29] , 
        \Level16Out160[28] , \Level16Out160[27] , \Level16Out160[26] , 
        \Level16Out160[25] , \Level16Out160[24] , \Level16Out160[23] , 
        \Level16Out160[22] , \Level16Out160[21] , \Level16Out160[20] , 
        \Level16Out160[19] , \Level16Out160[18] , \Level16Out160[17] , 
        \Level16Out160[16] , \Level16Out160[15] , \Level16Out160[14] , 
        \Level16Out160[13] , \Level16Out160[12] , \Level16Out160[11] , 
        \Level16Out160[10] , \Level16Out160[9] , \Level16Out160[8] , 
        \Level16Out160[7] , \Level16Out160[6] , \Level16Out160[5] , 
        \Level16Out160[4] , \Level16Out160[3] , \Level16Out160[2] , 
        \Level16Out160[1] , \Level16Out160[0] }), .In2({\Level16Out176[31] , 
        \Level16Out176[30] , \Level16Out176[29] , \Level16Out176[28] , 
        \Level16Out176[27] , \Level16Out176[26] , \Level16Out176[25] , 
        \Level16Out176[24] , \Level16Out176[23] , \Level16Out176[22] , 
        \Level16Out176[21] , \Level16Out176[20] , \Level16Out176[19] , 
        \Level16Out176[18] , \Level16Out176[17] , \Level16Out176[16] , 
        \Level16Out176[15] , \Level16Out176[14] , \Level16Out176[13] , 
        \Level16Out176[12] , \Level16Out176[11] , \Level16Out176[10] , 
        \Level16Out176[9] , \Level16Out176[8] , \Level16Out176[7] , 
        \Level16Out176[6] , \Level16Out176[5] , \Level16Out176[4] , 
        \Level16Out176[3] , \Level16Out176[2] , \Level16Out176[1] , 
        \Level16Out176[0] }), .Read1(\Level16Load160[0] ), .Read2(
        \Level16Load176[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_156_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load156[0] ), .Out({\Level2Out156[31] , \Level2Out156[30] , 
        \Level2Out156[29] , \Level2Out156[28] , \Level2Out156[27] , 
        \Level2Out156[26] , \Level2Out156[25] , \Level2Out156[24] , 
        \Level2Out156[23] , \Level2Out156[22] , \Level2Out156[21] , 
        \Level2Out156[20] , \Level2Out156[19] , \Level2Out156[18] , 
        \Level2Out156[17] , \Level2Out156[16] , \Level2Out156[15] , 
        \Level2Out156[14] , \Level2Out156[13] , \Level2Out156[12] , 
        \Level2Out156[11] , \Level2Out156[10] , \Level2Out156[9] , 
        \Level2Out156[8] , \Level2Out156[7] , \Level2Out156[6] , 
        \Level2Out156[5] , \Level2Out156[4] , \Level2Out156[3] , 
        \Level2Out156[2] , \Level2Out156[1] , \Level2Out156[0] }), .In1({
        \Level1Out156[31] , \Level1Out156[30] , \Level1Out156[29] , 
        \Level1Out156[28] , \Level1Out156[27] , \Level1Out156[26] , 
        \Level1Out156[25] , \Level1Out156[24] , \Level1Out156[23] , 
        \Level1Out156[22] , \Level1Out156[21] , \Level1Out156[20] , 
        \Level1Out156[19] , \Level1Out156[18] , \Level1Out156[17] , 
        \Level1Out156[16] , \Level1Out156[15] , \Level1Out156[14] , 
        \Level1Out156[13] , \Level1Out156[12] , \Level1Out156[11] , 
        \Level1Out156[10] , \Level1Out156[9] , \Level1Out156[8] , 
        \Level1Out156[7] , \Level1Out156[6] , \Level1Out156[5] , 
        \Level1Out156[4] , \Level1Out156[3] , \Level1Out156[2] , 
        \Level1Out156[1] , \Level1Out156[0] }), .In2({\Level1Out157[31] , 
        \Level1Out157[30] , \Level1Out157[29] , \Level1Out157[28] , 
        \Level1Out157[27] , \Level1Out157[26] , \Level1Out157[25] , 
        \Level1Out157[24] , \Level1Out157[23] , \Level1Out157[22] , 
        \Level1Out157[21] , \Level1Out157[20] , \Level1Out157[19] , 
        \Level1Out157[18] , \Level1Out157[17] , \Level1Out157[16] , 
        \Level1Out157[15] , \Level1Out157[14] , \Level1Out157[13] , 
        \Level1Out157[12] , \Level1Out157[11] , \Level1Out157[10] , 
        \Level1Out157[9] , \Level1Out157[8] , \Level1Out157[7] , 
        \Level1Out157[6] , \Level1Out157[5] , \Level1Out157[4] , 
        \Level1Out157[3] , \Level1Out157[2] , \Level1Out157[1] , 
        \Level1Out157[0] }), .Read1(\Level1Load156[0] ), .Read2(
        \Level1Load157[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_248_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load248[0] ), .Out({\Level2Out248[31] , \Level2Out248[30] , 
        \Level2Out248[29] , \Level2Out248[28] , \Level2Out248[27] , 
        \Level2Out248[26] , \Level2Out248[25] , \Level2Out248[24] , 
        \Level2Out248[23] , \Level2Out248[22] , \Level2Out248[21] , 
        \Level2Out248[20] , \Level2Out248[19] , \Level2Out248[18] , 
        \Level2Out248[17] , \Level2Out248[16] , \Level2Out248[15] , 
        \Level2Out248[14] , \Level2Out248[13] , \Level2Out248[12] , 
        \Level2Out248[11] , \Level2Out248[10] , \Level2Out248[9] , 
        \Level2Out248[8] , \Level2Out248[7] , \Level2Out248[6] , 
        \Level2Out248[5] , \Level2Out248[4] , \Level2Out248[3] , 
        \Level2Out248[2] , \Level2Out248[1] , \Level2Out248[0] }), .In1({
        \Level1Out248[31] , \Level1Out248[30] , \Level1Out248[29] , 
        \Level1Out248[28] , \Level1Out248[27] , \Level1Out248[26] , 
        \Level1Out248[25] , \Level1Out248[24] , \Level1Out248[23] , 
        \Level1Out248[22] , \Level1Out248[21] , \Level1Out248[20] , 
        \Level1Out248[19] , \Level1Out248[18] , \Level1Out248[17] , 
        \Level1Out248[16] , \Level1Out248[15] , \Level1Out248[14] , 
        \Level1Out248[13] , \Level1Out248[12] , \Level1Out248[11] , 
        \Level1Out248[10] , \Level1Out248[9] , \Level1Out248[8] , 
        \Level1Out248[7] , \Level1Out248[6] , \Level1Out248[5] , 
        \Level1Out248[4] , \Level1Out248[3] , \Level1Out248[2] , 
        \Level1Out248[1] , \Level1Out248[0] }), .In2({\Level1Out249[31] , 
        \Level1Out249[30] , \Level1Out249[29] , \Level1Out249[28] , 
        \Level1Out249[27] , \Level1Out249[26] , \Level1Out249[25] , 
        \Level1Out249[24] , \Level1Out249[23] , \Level1Out249[22] , 
        \Level1Out249[21] , \Level1Out249[20] , \Level1Out249[19] , 
        \Level1Out249[18] , \Level1Out249[17] , \Level1Out249[16] , 
        \Level1Out249[15] , \Level1Out249[14] , \Level1Out249[13] , 
        \Level1Out249[12] , \Level1Out249[11] , \Level1Out249[10] , 
        \Level1Out249[9] , \Level1Out249[8] , \Level1Out249[7] , 
        \Level1Out249[6] , \Level1Out249[5] , \Level1Out249[4] , 
        \Level1Out249[3] , \Level1Out249[2] , \Level1Out249[1] , 
        \Level1Out249[0] }), .Read1(\Level1Load248[0] ), .Read2(
        \Level1Load249[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_160_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load160[0] ), .Out({\Level4Out160[31] , \Level4Out160[30] , 
        \Level4Out160[29] , \Level4Out160[28] , \Level4Out160[27] , 
        \Level4Out160[26] , \Level4Out160[25] , \Level4Out160[24] , 
        \Level4Out160[23] , \Level4Out160[22] , \Level4Out160[21] , 
        \Level4Out160[20] , \Level4Out160[19] , \Level4Out160[18] , 
        \Level4Out160[17] , \Level4Out160[16] , \Level4Out160[15] , 
        \Level4Out160[14] , \Level4Out160[13] , \Level4Out160[12] , 
        \Level4Out160[11] , \Level4Out160[10] , \Level4Out160[9] , 
        \Level4Out160[8] , \Level4Out160[7] , \Level4Out160[6] , 
        \Level4Out160[5] , \Level4Out160[4] , \Level4Out160[3] , 
        \Level4Out160[2] , \Level4Out160[1] , \Level4Out160[0] }), .In1({
        \Level2Out160[31] , \Level2Out160[30] , \Level2Out160[29] , 
        \Level2Out160[28] , \Level2Out160[27] , \Level2Out160[26] , 
        \Level2Out160[25] , \Level2Out160[24] , \Level2Out160[23] , 
        \Level2Out160[22] , \Level2Out160[21] , \Level2Out160[20] , 
        \Level2Out160[19] , \Level2Out160[18] , \Level2Out160[17] , 
        \Level2Out160[16] , \Level2Out160[15] , \Level2Out160[14] , 
        \Level2Out160[13] , \Level2Out160[12] , \Level2Out160[11] , 
        \Level2Out160[10] , \Level2Out160[9] , \Level2Out160[8] , 
        \Level2Out160[7] , \Level2Out160[6] , \Level2Out160[5] , 
        \Level2Out160[4] , \Level2Out160[3] , \Level2Out160[2] , 
        \Level2Out160[1] , \Level2Out160[0] }), .In2({\Level2Out162[31] , 
        \Level2Out162[30] , \Level2Out162[29] , \Level2Out162[28] , 
        \Level2Out162[27] , \Level2Out162[26] , \Level2Out162[25] , 
        \Level2Out162[24] , \Level2Out162[23] , \Level2Out162[22] , 
        \Level2Out162[21] , \Level2Out162[20] , \Level2Out162[19] , 
        \Level2Out162[18] , \Level2Out162[17] , \Level2Out162[16] , 
        \Level2Out162[15] , \Level2Out162[14] , \Level2Out162[13] , 
        \Level2Out162[12] , \Level2Out162[11] , \Level2Out162[10] , 
        \Level2Out162[9] , \Level2Out162[8] , \Level2Out162[7] , 
        \Level2Out162[6] , \Level2Out162[5] , \Level2Out162[4] , 
        \Level2Out162[3] , \Level2Out162[2] , \Level2Out162[1] , 
        \Level2Out162[0] }), .Read1(\Level2Load160[0] ), .Read2(
        \Level2Load162[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_138 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink138[31] , \ScanLink138[30] , 
        \ScanLink138[29] , \ScanLink138[28] , \ScanLink138[27] , 
        \ScanLink138[26] , \ScanLink138[25] , \ScanLink138[24] , 
        \ScanLink138[23] , \ScanLink138[22] , \ScanLink138[21] , 
        \ScanLink138[20] , \ScanLink138[19] , \ScanLink138[18] , 
        \ScanLink138[17] , \ScanLink138[16] , \ScanLink138[15] , 
        \ScanLink138[14] , \ScanLink138[13] , \ScanLink138[12] , 
        \ScanLink138[11] , \ScanLink138[10] , \ScanLink138[9] , 
        \ScanLink138[8] , \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , 
        \ScanLink138[4] , \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , 
        \ScanLink138[0] }), .ScanOut({\ScanLink139[31] , \ScanLink139[30] , 
        \ScanLink139[29] , \ScanLink139[28] , \ScanLink139[27] , 
        \ScanLink139[26] , \ScanLink139[25] , \ScanLink139[24] , 
        \ScanLink139[23] , \ScanLink139[22] , \ScanLink139[21] , 
        \ScanLink139[20] , \ScanLink139[19] , \ScanLink139[18] , 
        \ScanLink139[17] , \ScanLink139[16] , \ScanLink139[15] , 
        \ScanLink139[14] , \ScanLink139[13] , \ScanLink139[12] , 
        \ScanLink139[11] , \ScanLink139[10] , \ScanLink139[9] , 
        \ScanLink139[8] , \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , 
        \ScanLink139[4] , \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , 
        \ScanLink139[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load138[0] ), .Out({\Level1Out138[31] , \Level1Out138[30] , 
        \Level1Out138[29] , \Level1Out138[28] , \Level1Out138[27] , 
        \Level1Out138[26] , \Level1Out138[25] , \Level1Out138[24] , 
        \Level1Out138[23] , \Level1Out138[22] , \Level1Out138[21] , 
        \Level1Out138[20] , \Level1Out138[19] , \Level1Out138[18] , 
        \Level1Out138[17] , \Level1Out138[16] , \Level1Out138[15] , 
        \Level1Out138[14] , \Level1Out138[13] , \Level1Out138[12] , 
        \Level1Out138[11] , \Level1Out138[10] , \Level1Out138[9] , 
        \Level1Out138[8] , \Level1Out138[7] , \Level1Out138[6] , 
        \Level1Out138[5] , \Level1Out138[4] , \Level1Out138[3] , 
        \Level1Out138[2] , \Level1Out138[1] , \Level1Out138[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_208 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink208[31] , \ScanLink208[30] , 
        \ScanLink208[29] , \ScanLink208[28] , \ScanLink208[27] , 
        \ScanLink208[26] , \ScanLink208[25] , \ScanLink208[24] , 
        \ScanLink208[23] , \ScanLink208[22] , \ScanLink208[21] , 
        \ScanLink208[20] , \ScanLink208[19] , \ScanLink208[18] , 
        \ScanLink208[17] , \ScanLink208[16] , \ScanLink208[15] , 
        \ScanLink208[14] , \ScanLink208[13] , \ScanLink208[12] , 
        \ScanLink208[11] , \ScanLink208[10] , \ScanLink208[9] , 
        \ScanLink208[8] , \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , 
        \ScanLink208[4] , \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , 
        \ScanLink208[0] }), .ScanOut({\ScanLink209[31] , \ScanLink209[30] , 
        \ScanLink209[29] , \ScanLink209[28] , \ScanLink209[27] , 
        \ScanLink209[26] , \ScanLink209[25] , \ScanLink209[24] , 
        \ScanLink209[23] , \ScanLink209[22] , \ScanLink209[21] , 
        \ScanLink209[20] , \ScanLink209[19] , \ScanLink209[18] , 
        \ScanLink209[17] , \ScanLink209[16] , \ScanLink209[15] , 
        \ScanLink209[14] , \ScanLink209[13] , \ScanLink209[12] , 
        \ScanLink209[11] , \ScanLink209[10] , \ScanLink209[9] , 
        \ScanLink209[8] , \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , 
        \ScanLink209[4] , \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , 
        \ScanLink209[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load208[0] ), .Out({\Level1Out208[31] , \Level1Out208[30] , 
        \Level1Out208[29] , \Level1Out208[28] , \Level1Out208[27] , 
        \Level1Out208[26] , \Level1Out208[25] , \Level1Out208[24] , 
        \Level1Out208[23] , \Level1Out208[22] , \Level1Out208[21] , 
        \Level1Out208[20] , \Level1Out208[19] , \Level1Out208[18] , 
        \Level1Out208[17] , \Level1Out208[16] , \Level1Out208[15] , 
        \Level1Out208[14] , \Level1Out208[13] , \Level1Out208[12] , 
        \Level1Out208[11] , \Level1Out208[10] , \Level1Out208[9] , 
        \Level1Out208[8] , \Level1Out208[7] , \Level1Out208[6] , 
        \Level1Out208[5] , \Level1Out208[4] , \Level1Out208[3] , 
        \Level1Out208[2] , \Level1Out208[1] , \Level1Out208[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_86_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load86[0] ), .Out({\Level2Out86[31] , \Level2Out86[30] , 
        \Level2Out86[29] , \Level2Out86[28] , \Level2Out86[27] , 
        \Level2Out86[26] , \Level2Out86[25] , \Level2Out86[24] , 
        \Level2Out86[23] , \Level2Out86[22] , \Level2Out86[21] , 
        \Level2Out86[20] , \Level2Out86[19] , \Level2Out86[18] , 
        \Level2Out86[17] , \Level2Out86[16] , \Level2Out86[15] , 
        \Level2Out86[14] , \Level2Out86[13] , \Level2Out86[12] , 
        \Level2Out86[11] , \Level2Out86[10] , \Level2Out86[9] , 
        \Level2Out86[8] , \Level2Out86[7] , \Level2Out86[6] , \Level2Out86[5] , 
        \Level2Out86[4] , \Level2Out86[3] , \Level2Out86[2] , \Level2Out86[1] , 
        \Level2Out86[0] }), .In1({\Level1Out86[31] , \Level1Out86[30] , 
        \Level1Out86[29] , \Level1Out86[28] , \Level1Out86[27] , 
        \Level1Out86[26] , \Level1Out86[25] , \Level1Out86[24] , 
        \Level1Out86[23] , \Level1Out86[22] , \Level1Out86[21] , 
        \Level1Out86[20] , \Level1Out86[19] , \Level1Out86[18] , 
        \Level1Out86[17] , \Level1Out86[16] , \Level1Out86[15] , 
        \Level1Out86[14] , \Level1Out86[13] , \Level1Out86[12] , 
        \Level1Out86[11] , \Level1Out86[10] , \Level1Out86[9] , 
        \Level1Out86[8] , \Level1Out86[7] , \Level1Out86[6] , \Level1Out86[5] , 
        \Level1Out86[4] , \Level1Out86[3] , \Level1Out86[2] , \Level1Out86[1] , 
        \Level1Out86[0] }), .In2({\Level1Out87[31] , \Level1Out87[30] , 
        \Level1Out87[29] , \Level1Out87[28] , \Level1Out87[27] , 
        \Level1Out87[26] , \Level1Out87[25] , \Level1Out87[24] , 
        \Level1Out87[23] , \Level1Out87[22] , \Level1Out87[21] , 
        \Level1Out87[20] , \Level1Out87[19] , \Level1Out87[18] , 
        \Level1Out87[17] , \Level1Out87[16] , \Level1Out87[15] , 
        \Level1Out87[14] , \Level1Out87[13] , \Level1Out87[12] , 
        \Level1Out87[11] , \Level1Out87[10] , \Level1Out87[9] , 
        \Level1Out87[8] , \Level1Out87[7] , \Level1Out87[6] , \Level1Out87[5] , 
        \Level1Out87[4] , \Level1Out87[3] , \Level1Out87[2] , \Level1Out87[1] , 
        \Level1Out87[0] }), .Read1(\Level1Load86[0] ), .Read2(
        \Level1Load87[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load24[0] ), .Out({\Level8Out24[31] , \Level8Out24[30] , 
        \Level8Out24[29] , \Level8Out24[28] , \Level8Out24[27] , 
        \Level8Out24[26] , \Level8Out24[25] , \Level8Out24[24] , 
        \Level8Out24[23] , \Level8Out24[22] , \Level8Out24[21] , 
        \Level8Out24[20] , \Level8Out24[19] , \Level8Out24[18] , 
        \Level8Out24[17] , \Level8Out24[16] , \Level8Out24[15] , 
        \Level8Out24[14] , \Level8Out24[13] , \Level8Out24[12] , 
        \Level8Out24[11] , \Level8Out24[10] , \Level8Out24[9] , 
        \Level8Out24[8] , \Level8Out24[7] , \Level8Out24[6] , \Level8Out24[5] , 
        \Level8Out24[4] , \Level8Out24[3] , \Level8Out24[2] , \Level8Out24[1] , 
        \Level8Out24[0] }), .In1({\Level4Out24[31] , \Level4Out24[30] , 
        \Level4Out24[29] , \Level4Out24[28] , \Level4Out24[27] , 
        \Level4Out24[26] , \Level4Out24[25] , \Level4Out24[24] , 
        \Level4Out24[23] , \Level4Out24[22] , \Level4Out24[21] , 
        \Level4Out24[20] , \Level4Out24[19] , \Level4Out24[18] , 
        \Level4Out24[17] , \Level4Out24[16] , \Level4Out24[15] , 
        \Level4Out24[14] , \Level4Out24[13] , \Level4Out24[12] , 
        \Level4Out24[11] , \Level4Out24[10] , \Level4Out24[9] , 
        \Level4Out24[8] , \Level4Out24[7] , \Level4Out24[6] , \Level4Out24[5] , 
        \Level4Out24[4] , \Level4Out24[3] , \Level4Out24[2] , \Level4Out24[1] , 
        \Level4Out24[0] }), .In2({\Level4Out28[31] , \Level4Out28[30] , 
        \Level4Out28[29] , \Level4Out28[28] , \Level4Out28[27] , 
        \Level4Out28[26] , \Level4Out28[25] , \Level4Out28[24] , 
        \Level4Out28[23] , \Level4Out28[22] , \Level4Out28[21] , 
        \Level4Out28[20] , \Level4Out28[19] , \Level4Out28[18] , 
        \Level4Out28[17] , \Level4Out28[16] , \Level4Out28[15] , 
        \Level4Out28[14] , \Level4Out28[13] , \Level4Out28[12] , 
        \Level4Out28[11] , \Level4Out28[10] , \Level4Out28[9] , 
        \Level4Out28[8] , \Level4Out28[7] , \Level4Out28[6] , \Level4Out28[5] , 
        \Level4Out28[4] , \Level4Out28[3] , \Level4Out28[2] , \Level4Out28[1] , 
        \Level4Out28[0] }), .Read1(\Level4Load24[0] ), .Read2(
        \Level4Load28[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_156 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink156[31] , \ScanLink156[30] , 
        \ScanLink156[29] , \ScanLink156[28] , \ScanLink156[27] , 
        \ScanLink156[26] , \ScanLink156[25] , \ScanLink156[24] , 
        \ScanLink156[23] , \ScanLink156[22] , \ScanLink156[21] , 
        \ScanLink156[20] , \ScanLink156[19] , \ScanLink156[18] , 
        \ScanLink156[17] , \ScanLink156[16] , \ScanLink156[15] , 
        \ScanLink156[14] , \ScanLink156[13] , \ScanLink156[12] , 
        \ScanLink156[11] , \ScanLink156[10] , \ScanLink156[9] , 
        \ScanLink156[8] , \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , 
        \ScanLink156[4] , \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , 
        \ScanLink156[0] }), .ScanOut({\ScanLink157[31] , \ScanLink157[30] , 
        \ScanLink157[29] , \ScanLink157[28] , \ScanLink157[27] , 
        \ScanLink157[26] , \ScanLink157[25] , \ScanLink157[24] , 
        \ScanLink157[23] , \ScanLink157[22] , \ScanLink157[21] , 
        \ScanLink157[20] , \ScanLink157[19] , \ScanLink157[18] , 
        \ScanLink157[17] , \ScanLink157[16] , \ScanLink157[15] , 
        \ScanLink157[14] , \ScanLink157[13] , \ScanLink157[12] , 
        \ScanLink157[11] , \ScanLink157[10] , \ScanLink157[9] , 
        \ScanLink157[8] , \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , 
        \ScanLink157[4] , \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , 
        \ScanLink157[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load156[0] ), .Out({\Level1Out156[31] , \Level1Out156[30] , 
        \Level1Out156[29] , \Level1Out156[28] , \Level1Out156[27] , 
        \Level1Out156[26] , \Level1Out156[25] , \Level1Out156[24] , 
        \Level1Out156[23] , \Level1Out156[22] , \Level1Out156[21] , 
        \Level1Out156[20] , \Level1Out156[19] , \Level1Out156[18] , 
        \Level1Out156[17] , \Level1Out156[16] , \Level1Out156[15] , 
        \Level1Out156[14] , \Level1Out156[13] , \Level1Out156[12] , 
        \Level1Out156[11] , \Level1Out156[10] , \Level1Out156[9] , 
        \Level1Out156[8] , \Level1Out156[7] , \Level1Out156[6] , 
        \Level1Out156[5] , \Level1Out156[4] , \Level1Out156[3] , 
        \Level1Out156[2] , \Level1Out156[1] , \Level1Out156[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_171 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink171[31] , \ScanLink171[30] , 
        \ScanLink171[29] , \ScanLink171[28] , \ScanLink171[27] , 
        \ScanLink171[26] , \ScanLink171[25] , \ScanLink171[24] , 
        \ScanLink171[23] , \ScanLink171[22] , \ScanLink171[21] , 
        \ScanLink171[20] , \ScanLink171[19] , \ScanLink171[18] , 
        \ScanLink171[17] , \ScanLink171[16] , \ScanLink171[15] , 
        \ScanLink171[14] , \ScanLink171[13] , \ScanLink171[12] , 
        \ScanLink171[11] , \ScanLink171[10] , \ScanLink171[9] , 
        \ScanLink171[8] , \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , 
        \ScanLink171[4] , \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , 
        \ScanLink171[0] }), .ScanOut({\ScanLink172[31] , \ScanLink172[30] , 
        \ScanLink172[29] , \ScanLink172[28] , \ScanLink172[27] , 
        \ScanLink172[26] , \ScanLink172[25] , \ScanLink172[24] , 
        \ScanLink172[23] , \ScanLink172[22] , \ScanLink172[21] , 
        \ScanLink172[20] , \ScanLink172[19] , \ScanLink172[18] , 
        \ScanLink172[17] , \ScanLink172[16] , \ScanLink172[15] , 
        \ScanLink172[14] , \ScanLink172[13] , \ScanLink172[12] , 
        \ScanLink172[11] , \ScanLink172[10] , \ScanLink172[9] , 
        \ScanLink172[8] , \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , 
        \ScanLink172[4] , \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , 
        \ScanLink172[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load171[0] ), .Out({\Level1Out171[31] , \Level1Out171[30] , 
        \Level1Out171[29] , \Level1Out171[28] , \Level1Out171[27] , 
        \Level1Out171[26] , \Level1Out171[25] , \Level1Out171[24] , 
        \Level1Out171[23] , \Level1Out171[22] , \Level1Out171[21] , 
        \Level1Out171[20] , \Level1Out171[19] , \Level1Out171[18] , 
        \Level1Out171[17] , \Level1Out171[16] , \Level1Out171[15] , 
        \Level1Out171[14] , \Level1Out171[13] , \Level1Out171[12] , 
        \Level1Out171[11] , \Level1Out171[10] , \Level1Out171[9] , 
        \Level1Out171[8] , \Level1Out171[7] , \Level1Out171[6] , 
        \Level1Out171[5] , \Level1Out171[4] , \Level1Out171[3] , 
        \Level1Out171[2] , \Level1Out171[1] , \Level1Out171[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_241 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink241[31] , \ScanLink241[30] , 
        \ScanLink241[29] , \ScanLink241[28] , \ScanLink241[27] , 
        \ScanLink241[26] , \ScanLink241[25] , \ScanLink241[24] , 
        \ScanLink241[23] , \ScanLink241[22] , \ScanLink241[21] , 
        \ScanLink241[20] , \ScanLink241[19] , \ScanLink241[18] , 
        \ScanLink241[17] , \ScanLink241[16] , \ScanLink241[15] , 
        \ScanLink241[14] , \ScanLink241[13] , \ScanLink241[12] , 
        \ScanLink241[11] , \ScanLink241[10] , \ScanLink241[9] , 
        \ScanLink241[8] , \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , 
        \ScanLink241[4] , \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , 
        \ScanLink241[0] }), .ScanOut({\ScanLink242[31] , \ScanLink242[30] , 
        \ScanLink242[29] , \ScanLink242[28] , \ScanLink242[27] , 
        \ScanLink242[26] , \ScanLink242[25] , \ScanLink242[24] , 
        \ScanLink242[23] , \ScanLink242[22] , \ScanLink242[21] , 
        \ScanLink242[20] , \ScanLink242[19] , \ScanLink242[18] , 
        \ScanLink242[17] , \ScanLink242[16] , \ScanLink242[15] , 
        \ScanLink242[14] , \ScanLink242[13] , \ScanLink242[12] , 
        \ScanLink242[11] , \ScanLink242[10] , \ScanLink242[9] , 
        \ScanLink242[8] , \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , 
        \ScanLink242[4] , \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , 
        \ScanLink242[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load241[0] ), .Out({\Level1Out241[31] , \Level1Out241[30] , 
        \Level1Out241[29] , \Level1Out241[28] , \Level1Out241[27] , 
        \Level1Out241[26] , \Level1Out241[25] , \Level1Out241[24] , 
        \Level1Out241[23] , \Level1Out241[22] , \Level1Out241[21] , 
        \Level1Out241[20] , \Level1Out241[19] , \Level1Out241[18] , 
        \Level1Out241[17] , \Level1Out241[16] , \Level1Out241[15] , 
        \Level1Out241[14] , \Level1Out241[13] , \Level1Out241[12] , 
        \Level1Out241[11] , \Level1Out241[10] , \Level1Out241[9] , 
        \Level1Out241[8] , \Level1Out241[7] , \Level1Out241[6] , 
        \Level1Out241[5] , \Level1Out241[4] , \Level1Out241[3] , 
        \Level1Out241[2] , \Level1Out241[1] , \Level1Out241[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_74 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink74[31] , \ScanLink74[30] , 
        \ScanLink74[29] , \ScanLink74[28] , \ScanLink74[27] , \ScanLink74[26] , 
        \ScanLink74[25] , \ScanLink74[24] , \ScanLink74[23] , \ScanLink74[22] , 
        \ScanLink74[21] , \ScanLink74[20] , \ScanLink74[19] , \ScanLink74[18] , 
        \ScanLink74[17] , \ScanLink74[16] , \ScanLink74[15] , \ScanLink74[14] , 
        \ScanLink74[13] , \ScanLink74[12] , \ScanLink74[11] , \ScanLink74[10] , 
        \ScanLink74[9] , \ScanLink74[8] , \ScanLink74[7] , \ScanLink74[6] , 
        \ScanLink74[5] , \ScanLink74[4] , \ScanLink74[3] , \ScanLink74[2] , 
        \ScanLink74[1] , \ScanLink74[0] }), .ScanOut({\ScanLink75[31] , 
        \ScanLink75[30] , \ScanLink75[29] , \ScanLink75[28] , \ScanLink75[27] , 
        \ScanLink75[26] , \ScanLink75[25] , \ScanLink75[24] , \ScanLink75[23] , 
        \ScanLink75[22] , \ScanLink75[21] , \ScanLink75[20] , \ScanLink75[19] , 
        \ScanLink75[18] , \ScanLink75[17] , \ScanLink75[16] , \ScanLink75[15] , 
        \ScanLink75[14] , \ScanLink75[13] , \ScanLink75[12] , \ScanLink75[11] , 
        \ScanLink75[10] , \ScanLink75[9] , \ScanLink75[8] , \ScanLink75[7] , 
        \ScanLink75[6] , \ScanLink75[5] , \ScanLink75[4] , \ScanLink75[3] , 
        \ScanLink75[2] , \ScanLink75[1] , \ScanLink75[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load74[0] ), .Out({
        \Level1Out74[31] , \Level1Out74[30] , \Level1Out74[29] , 
        \Level1Out74[28] , \Level1Out74[27] , \Level1Out74[26] , 
        \Level1Out74[25] , \Level1Out74[24] , \Level1Out74[23] , 
        \Level1Out74[22] , \Level1Out74[21] , \Level1Out74[20] , 
        \Level1Out74[19] , \Level1Out74[18] , \Level1Out74[17] , 
        \Level1Out74[16] , \Level1Out74[15] , \Level1Out74[14] , 
        \Level1Out74[13] , \Level1Out74[12] , \Level1Out74[11] , 
        \Level1Out74[10] , \Level1Out74[9] , \Level1Out74[8] , 
        \Level1Out74[7] , \Level1Out74[6] , \Level1Out74[5] , \Level1Out74[4] , 
        \Level1Out74[3] , \Level1Out74[2] , \Level1Out74[1] , \Level1Out74[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanOut({\ScanLink8[31] , 
        \ScanLink8[30] , \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , 
        \ScanLink8[26] , \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , 
        \ScanLink8[22] , \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , 
        \ScanLink8[18] , \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , 
        \ScanLink8[14] , \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , 
        \ScanLink8[10] , \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , 
        \ScanLink8[6] , \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , 
        \ScanLink8[2] , \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load7[0] ), .Out({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanOut({\ScanLink13[31] , 
        \ScanLink13[30] , \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , 
        \ScanLink13[26] , \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , 
        \ScanLink13[22] , \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , 
        \ScanLink13[18] , \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , 
        \ScanLink13[14] , \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , 
        \ScanLink13[10] , \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , 
        \ScanLink13[6] , \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , 
        \ScanLink13[2] , \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load12[0] ), .Out({
        \Level1Out12[31] , \Level1Out12[30] , \Level1Out12[29] , 
        \Level1Out12[28] , \Level1Out12[27] , \Level1Out12[26] , 
        \Level1Out12[25] , \Level1Out12[24] , \Level1Out12[23] , 
        \Level1Out12[22] , \Level1Out12[21] , \Level1Out12[20] , 
        \Level1Out12[19] , \Level1Out12[18] , \Level1Out12[17] , 
        \Level1Out12[16] , \Level1Out12[15] , \Level1Out12[14] , 
        \Level1Out12[13] , \Level1Out12[12] , \Level1Out12[11] , 
        \Level1Out12[10] , \Level1Out12[9] , \Level1Out12[8] , 
        \Level1Out12[7] , \Level1Out12[6] , \Level1Out12[5] , \Level1Out12[4] , 
        \Level1Out12[3] , \Level1Out12[2] , \Level1Out12[1] , \Level1Out12[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_26 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanOut({\ScanLink27[31] , 
        \ScanLink27[30] , \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , 
        \ScanLink27[26] , \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , 
        \ScanLink27[22] , \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , 
        \ScanLink27[18] , \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , 
        \ScanLink27[14] , \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , 
        \ScanLink27[10] , \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , 
        \ScanLink27[6] , \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , 
        \ScanLink27[2] , \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load26[0] ), .Out({
        \Level1Out26[31] , \Level1Out26[30] , \Level1Out26[29] , 
        \Level1Out26[28] , \Level1Out26[27] , \Level1Out26[26] , 
        \Level1Out26[25] , \Level1Out26[24] , \Level1Out26[23] , 
        \Level1Out26[22] , \Level1Out26[21] , \Level1Out26[20] , 
        \Level1Out26[19] , \Level1Out26[18] , \Level1Out26[17] , 
        \Level1Out26[16] , \Level1Out26[15] , \Level1Out26[14] , 
        \Level1Out26[13] , \Level1Out26[12] , \Level1Out26[11] , 
        \Level1Out26[10] , \Level1Out26[9] , \Level1Out26[8] , 
        \Level1Out26[7] , \Level1Out26[6] , \Level1Out26[5] , \Level1Out26[4] , 
        \Level1Out26[3] , \Level1Out26[2] , \Level1Out26[1] , \Level1Out26[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_104 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink104[31] , \ScanLink104[30] , 
        \ScanLink104[29] , \ScanLink104[28] , \ScanLink104[27] , 
        \ScanLink104[26] , \ScanLink104[25] , \ScanLink104[24] , 
        \ScanLink104[23] , \ScanLink104[22] , \ScanLink104[21] , 
        \ScanLink104[20] , \ScanLink104[19] , \ScanLink104[18] , 
        \ScanLink104[17] , \ScanLink104[16] , \ScanLink104[15] , 
        \ScanLink104[14] , \ScanLink104[13] , \ScanLink104[12] , 
        \ScanLink104[11] , \ScanLink104[10] , \ScanLink104[9] , 
        \ScanLink104[8] , \ScanLink104[7] , \ScanLink104[6] , \ScanLink104[5] , 
        \ScanLink104[4] , \ScanLink104[3] , \ScanLink104[2] , \ScanLink104[1] , 
        \ScanLink104[0] }), .ScanOut({\ScanLink105[31] , \ScanLink105[30] , 
        \ScanLink105[29] , \ScanLink105[28] , \ScanLink105[27] , 
        \ScanLink105[26] , \ScanLink105[25] , \ScanLink105[24] , 
        \ScanLink105[23] , \ScanLink105[22] , \ScanLink105[21] , 
        \ScanLink105[20] , \ScanLink105[19] , \ScanLink105[18] , 
        \ScanLink105[17] , \ScanLink105[16] , \ScanLink105[15] , 
        \ScanLink105[14] , \ScanLink105[13] , \ScanLink105[12] , 
        \ScanLink105[11] , \ScanLink105[10] , \ScanLink105[9] , 
        \ScanLink105[8] , \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , 
        \ScanLink105[4] , \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , 
        \ScanLink105[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load104[0] ), .Out({\Level1Out104[31] , \Level1Out104[30] , 
        \Level1Out104[29] , \Level1Out104[28] , \Level1Out104[27] , 
        \Level1Out104[26] , \Level1Out104[25] , \Level1Out104[24] , 
        \Level1Out104[23] , \Level1Out104[22] , \Level1Out104[21] , 
        \Level1Out104[20] , \Level1Out104[19] , \Level1Out104[18] , 
        \Level1Out104[17] , \Level1Out104[16] , \Level1Out104[15] , 
        \Level1Out104[14] , \Level1Out104[13] , \Level1Out104[12] , 
        \Level1Out104[11] , \Level1Out104[10] , \Level1Out104[9] , 
        \Level1Out104[8] , \Level1Out104[7] , \Level1Out104[6] , 
        \Level1Out104[5] , \Level1Out104[4] , \Level1Out104[3] , 
        \Level1Out104[2] , \Level1Out104[1] , \Level1Out104[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_123 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink123[31] , \ScanLink123[30] , 
        \ScanLink123[29] , \ScanLink123[28] , \ScanLink123[27] , 
        \ScanLink123[26] , \ScanLink123[25] , \ScanLink123[24] , 
        \ScanLink123[23] , \ScanLink123[22] , \ScanLink123[21] , 
        \ScanLink123[20] , \ScanLink123[19] , \ScanLink123[18] , 
        \ScanLink123[17] , \ScanLink123[16] , \ScanLink123[15] , 
        \ScanLink123[14] , \ScanLink123[13] , \ScanLink123[12] , 
        \ScanLink123[11] , \ScanLink123[10] , \ScanLink123[9] , 
        \ScanLink123[8] , \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , 
        \ScanLink123[4] , \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , 
        \ScanLink123[0] }), .ScanOut({\ScanLink124[31] , \ScanLink124[30] , 
        \ScanLink124[29] , \ScanLink124[28] , \ScanLink124[27] , 
        \ScanLink124[26] , \ScanLink124[25] , \ScanLink124[24] , 
        \ScanLink124[23] , \ScanLink124[22] , \ScanLink124[21] , 
        \ScanLink124[20] , \ScanLink124[19] , \ScanLink124[18] , 
        \ScanLink124[17] , \ScanLink124[16] , \ScanLink124[15] , 
        \ScanLink124[14] , \ScanLink124[13] , \ScanLink124[12] , 
        \ScanLink124[11] , \ScanLink124[10] , \ScanLink124[9] , 
        \ScanLink124[8] , \ScanLink124[7] , \ScanLink124[6] , \ScanLink124[5] , 
        \ScanLink124[4] , \ScanLink124[3] , \ScanLink124[2] , \ScanLink124[1] , 
        \ScanLink124[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load123[0] ), .Out({\Level1Out123[31] , \Level1Out123[30] , 
        \Level1Out123[29] , \Level1Out123[28] , \Level1Out123[27] , 
        \Level1Out123[26] , \Level1Out123[25] , \Level1Out123[24] , 
        \Level1Out123[23] , \Level1Out123[22] , \Level1Out123[21] , 
        \Level1Out123[20] , \Level1Out123[19] , \Level1Out123[18] , 
        \Level1Out123[17] , \Level1Out123[16] , \Level1Out123[15] , 
        \Level1Out123[14] , \Level1Out123[13] , \Level1Out123[12] , 
        \Level1Out123[11] , \Level1Out123[10] , \Level1Out123[9] , 
        \Level1Out123[8] , \Level1Out123[7] , \Level1Out123[6] , 
        \Level1Out123[5] , \Level1Out123[4] , \Level1Out123[3] , 
        \Level1Out123[2] , \Level1Out123[1] , \Level1Out123[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_164_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load164[0] ), .Out({\Level2Out164[31] , \Level2Out164[30] , 
        \Level2Out164[29] , \Level2Out164[28] , \Level2Out164[27] , 
        \Level2Out164[26] , \Level2Out164[25] , \Level2Out164[24] , 
        \Level2Out164[23] , \Level2Out164[22] , \Level2Out164[21] , 
        \Level2Out164[20] , \Level2Out164[19] , \Level2Out164[18] , 
        \Level2Out164[17] , \Level2Out164[16] , \Level2Out164[15] , 
        \Level2Out164[14] , \Level2Out164[13] , \Level2Out164[12] , 
        \Level2Out164[11] , \Level2Out164[10] , \Level2Out164[9] , 
        \Level2Out164[8] , \Level2Out164[7] , \Level2Out164[6] , 
        \Level2Out164[5] , \Level2Out164[4] , \Level2Out164[3] , 
        \Level2Out164[2] , \Level2Out164[1] , \Level2Out164[0] }), .In1({
        \Level1Out164[31] , \Level1Out164[30] , \Level1Out164[29] , 
        \Level1Out164[28] , \Level1Out164[27] , \Level1Out164[26] , 
        \Level1Out164[25] , \Level1Out164[24] , \Level1Out164[23] , 
        \Level1Out164[22] , \Level1Out164[21] , \Level1Out164[20] , 
        \Level1Out164[19] , \Level1Out164[18] , \Level1Out164[17] , 
        \Level1Out164[16] , \Level1Out164[15] , \Level1Out164[14] , 
        \Level1Out164[13] , \Level1Out164[12] , \Level1Out164[11] , 
        \Level1Out164[10] , \Level1Out164[9] , \Level1Out164[8] , 
        \Level1Out164[7] , \Level1Out164[6] , \Level1Out164[5] , 
        \Level1Out164[4] , \Level1Out164[3] , \Level1Out164[2] , 
        \Level1Out164[1] , \Level1Out164[0] }), .In2({\Level1Out165[31] , 
        \Level1Out165[30] , \Level1Out165[29] , \Level1Out165[28] , 
        \Level1Out165[27] , \Level1Out165[26] , \Level1Out165[25] , 
        \Level1Out165[24] , \Level1Out165[23] , \Level1Out165[22] , 
        \Level1Out165[21] , \Level1Out165[20] , \Level1Out165[19] , 
        \Level1Out165[18] , \Level1Out165[17] , \Level1Out165[16] , 
        \Level1Out165[15] , \Level1Out165[14] , \Level1Out165[13] , 
        \Level1Out165[12] , \Level1Out165[11] , \Level1Out165[10] , 
        \Level1Out165[9] , \Level1Out165[8] , \Level1Out165[7] , 
        \Level1Out165[6] , \Level1Out165[5] , \Level1Out165[4] , 
        \Level1Out165[3] , \Level1Out165[2] , \Level1Out165[1] , 
        \Level1Out165[0] }), .Read1(\Level1Load164[0] ), .Read2(
        \Level1Load165[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load32[0] ), .Out({\Level32Out32[31] , \Level32Out32[30] , 
        \Level32Out32[29] , \Level32Out32[28] , \Level32Out32[27] , 
        \Level32Out32[26] , \Level32Out32[25] , \Level32Out32[24] , 
        \Level32Out32[23] , \Level32Out32[22] , \Level32Out32[21] , 
        \Level32Out32[20] , \Level32Out32[19] , \Level32Out32[18] , 
        \Level32Out32[17] , \Level32Out32[16] , \Level32Out32[15] , 
        \Level32Out32[14] , \Level32Out32[13] , \Level32Out32[12] , 
        \Level32Out32[11] , \Level32Out32[10] , \Level32Out32[9] , 
        \Level32Out32[8] , \Level32Out32[7] , \Level32Out32[6] , 
        \Level32Out32[5] , \Level32Out32[4] , \Level32Out32[3] , 
        \Level32Out32[2] , \Level32Out32[1] , \Level32Out32[0] }), .In1({
        \Level16Out32[31] , \Level16Out32[30] , \Level16Out32[29] , 
        \Level16Out32[28] , \Level16Out32[27] , \Level16Out32[26] , 
        \Level16Out32[25] , \Level16Out32[24] , \Level16Out32[23] , 
        \Level16Out32[22] , \Level16Out32[21] , \Level16Out32[20] , 
        \Level16Out32[19] , \Level16Out32[18] , \Level16Out32[17] , 
        \Level16Out32[16] , \Level16Out32[15] , \Level16Out32[14] , 
        \Level16Out32[13] , \Level16Out32[12] , \Level16Out32[11] , 
        \Level16Out32[10] , \Level16Out32[9] , \Level16Out32[8] , 
        \Level16Out32[7] , \Level16Out32[6] , \Level16Out32[5] , 
        \Level16Out32[4] , \Level16Out32[3] , \Level16Out32[2] , 
        \Level16Out32[1] , \Level16Out32[0] }), .In2({\Level16Out48[31] , 
        \Level16Out48[30] , \Level16Out48[29] , \Level16Out48[28] , 
        \Level16Out48[27] , \Level16Out48[26] , \Level16Out48[25] , 
        \Level16Out48[24] , \Level16Out48[23] , \Level16Out48[22] , 
        \Level16Out48[21] , \Level16Out48[20] , \Level16Out48[19] , 
        \Level16Out48[18] , \Level16Out48[17] , \Level16Out48[16] , 
        \Level16Out48[15] , \Level16Out48[14] , \Level16Out48[13] , 
        \Level16Out48[12] , \Level16Out48[11] , \Level16Out48[10] , 
        \Level16Out48[9] , \Level16Out48[8] , \Level16Out48[7] , 
        \Level16Out48[6] , \Level16Out48[5] , \Level16Out48[4] , 
        \Level16Out48[3] , \Level16Out48[2] , \Level16Out48[1] , 
        \Level16Out48[0] }), .Read1(\Level16Load32[0] ), .Read2(
        \Level16Load48[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_213 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink213[31] , \ScanLink213[30] , 
        \ScanLink213[29] , \ScanLink213[28] , \ScanLink213[27] , 
        \ScanLink213[26] , \ScanLink213[25] , \ScanLink213[24] , 
        \ScanLink213[23] , \ScanLink213[22] , \ScanLink213[21] , 
        \ScanLink213[20] , \ScanLink213[19] , \ScanLink213[18] , 
        \ScanLink213[17] , \ScanLink213[16] , \ScanLink213[15] , 
        \ScanLink213[14] , \ScanLink213[13] , \ScanLink213[12] , 
        \ScanLink213[11] , \ScanLink213[10] , \ScanLink213[9] , 
        \ScanLink213[8] , \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , 
        \ScanLink213[4] , \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , 
        \ScanLink213[0] }), .ScanOut({\ScanLink214[31] , \ScanLink214[30] , 
        \ScanLink214[29] , \ScanLink214[28] , \ScanLink214[27] , 
        \ScanLink214[26] , \ScanLink214[25] , \ScanLink214[24] , 
        \ScanLink214[23] , \ScanLink214[22] , \ScanLink214[21] , 
        \ScanLink214[20] , \ScanLink214[19] , \ScanLink214[18] , 
        \ScanLink214[17] , \ScanLink214[16] , \ScanLink214[15] , 
        \ScanLink214[14] , \ScanLink214[13] , \ScanLink214[12] , 
        \ScanLink214[11] , \ScanLink214[10] , \ScanLink214[9] , 
        \ScanLink214[8] , \ScanLink214[7] , \ScanLink214[6] , \ScanLink214[5] , 
        \ScanLink214[4] , \ScanLink214[3] , \ScanLink214[2] , \ScanLink214[1] , 
        \ScanLink214[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load213[0] ), .Out({\Level1Out213[31] , \Level1Out213[30] , 
        \Level1Out213[29] , \Level1Out213[28] , \Level1Out213[27] , 
        \Level1Out213[26] , \Level1Out213[25] , \Level1Out213[24] , 
        \Level1Out213[23] , \Level1Out213[22] , \Level1Out213[21] , 
        \Level1Out213[20] , \Level1Out213[19] , \Level1Out213[18] , 
        \Level1Out213[17] , \Level1Out213[16] , \Level1Out213[15] , 
        \Level1Out213[14] , \Level1Out213[13] , \Level1Out213[12] , 
        \Level1Out213[11] , \Level1Out213[10] , \Level1Out213[9] , 
        \Level1Out213[8] , \Level1Out213[7] , \Level1Out213[6] , 
        \Level1Out213[5] , \Level1Out213[4] , \Level1Out213[3] , 
        \Level1Out213[2] , \Level1Out213[1] , \Level1Out213[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_234 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink234[31] , \ScanLink234[30] , 
        \ScanLink234[29] , \ScanLink234[28] , \ScanLink234[27] , 
        \ScanLink234[26] , \ScanLink234[25] , \ScanLink234[24] , 
        \ScanLink234[23] , \ScanLink234[22] , \ScanLink234[21] , 
        \ScanLink234[20] , \ScanLink234[19] , \ScanLink234[18] , 
        \ScanLink234[17] , \ScanLink234[16] , \ScanLink234[15] , 
        \ScanLink234[14] , \ScanLink234[13] , \ScanLink234[12] , 
        \ScanLink234[11] , \ScanLink234[10] , \ScanLink234[9] , 
        \ScanLink234[8] , \ScanLink234[7] , \ScanLink234[6] , \ScanLink234[5] , 
        \ScanLink234[4] , \ScanLink234[3] , \ScanLink234[2] , \ScanLink234[1] , 
        \ScanLink234[0] }), .ScanOut({\ScanLink235[31] , \ScanLink235[30] , 
        \ScanLink235[29] , \ScanLink235[28] , \ScanLink235[27] , 
        \ScanLink235[26] , \ScanLink235[25] , \ScanLink235[24] , 
        \ScanLink235[23] , \ScanLink235[22] , \ScanLink235[21] , 
        \ScanLink235[20] , \ScanLink235[19] , \ScanLink235[18] , 
        \ScanLink235[17] , \ScanLink235[16] , \ScanLink235[15] , 
        \ScanLink235[14] , \ScanLink235[13] , \ScanLink235[12] , 
        \ScanLink235[11] , \ScanLink235[10] , \ScanLink235[9] , 
        \ScanLink235[8] , \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , 
        \ScanLink235[4] , \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , 
        \ScanLink235[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load234[0] ), .Out({\Level1Out234[31] , \Level1Out234[30] , 
        \Level1Out234[29] , \Level1Out234[28] , \Level1Out234[27] , 
        \Level1Out234[26] , \Level1Out234[25] , \Level1Out234[24] , 
        \Level1Out234[23] , \Level1Out234[22] , \Level1Out234[21] , 
        \Level1Out234[20] , \Level1Out234[19] , \Level1Out234[18] , 
        \Level1Out234[17] , \Level1Out234[16] , \Level1Out234[15] , 
        \Level1Out234[14] , \Level1Out234[13] , \Level1Out234[12] , 
        \Level1Out234[11] , \Level1Out234[10] , \Level1Out234[9] , 
        \Level1Out234[8] , \Level1Out234[7] , \Level1Out234[6] , 
        \Level1Out234[5] , \Level1Out234[4] , \Level1Out234[3] , 
        \Level1Out234[2] , \Level1Out234[1] , \Level1Out234[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_22_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load22[0] ), .Out({\Level2Out22[31] , \Level2Out22[30] , 
        \Level2Out22[29] , \Level2Out22[28] , \Level2Out22[27] , 
        \Level2Out22[26] , \Level2Out22[25] , \Level2Out22[24] , 
        \Level2Out22[23] , \Level2Out22[22] , \Level2Out22[21] , 
        \Level2Out22[20] , \Level2Out22[19] , \Level2Out22[18] , 
        \Level2Out22[17] , \Level2Out22[16] , \Level2Out22[15] , 
        \Level2Out22[14] , \Level2Out22[13] , \Level2Out22[12] , 
        \Level2Out22[11] , \Level2Out22[10] , \Level2Out22[9] , 
        \Level2Out22[8] , \Level2Out22[7] , \Level2Out22[6] , \Level2Out22[5] , 
        \Level2Out22[4] , \Level2Out22[3] , \Level2Out22[2] , \Level2Out22[1] , 
        \Level2Out22[0] }), .In1({\Level1Out22[31] , \Level1Out22[30] , 
        \Level1Out22[29] , \Level1Out22[28] , \Level1Out22[27] , 
        \Level1Out22[26] , \Level1Out22[25] , \Level1Out22[24] , 
        \Level1Out22[23] , \Level1Out22[22] , \Level1Out22[21] , 
        \Level1Out22[20] , \Level1Out22[19] , \Level1Out22[18] , 
        \Level1Out22[17] , \Level1Out22[16] , \Level1Out22[15] , 
        \Level1Out22[14] , \Level1Out22[13] , \Level1Out22[12] , 
        \Level1Out22[11] , \Level1Out22[10] , \Level1Out22[9] , 
        \Level1Out22[8] , \Level1Out22[7] , \Level1Out22[6] , \Level1Out22[5] , 
        \Level1Out22[4] , \Level1Out22[3] , \Level1Out22[2] , \Level1Out22[1] , 
        \Level1Out22[0] }), .In2({\Level1Out23[31] , \Level1Out23[30] , 
        \Level1Out23[29] , \Level1Out23[28] , \Level1Out23[27] , 
        \Level1Out23[26] , \Level1Out23[25] , \Level1Out23[24] , 
        \Level1Out23[23] , \Level1Out23[22] , \Level1Out23[21] , 
        \Level1Out23[20] , \Level1Out23[19] , \Level1Out23[18] , 
        \Level1Out23[17] , \Level1Out23[16] , \Level1Out23[15] , 
        \Level1Out23[14] , \Level1Out23[13] , \Level1Out23[12] , 
        \Level1Out23[11] , \Level1Out23[10] , \Level1Out23[9] , 
        \Level1Out23[8] , \Level1Out23[7] , \Level1Out23[6] , \Level1Out23[5] , 
        \Level1Out23[4] , \Level1Out23[3] , \Level1Out23[2] , \Level1Out23[1] , 
        \Level1Out23[0] }), .Read1(\Level1Load22[0] ), .Read2(
        \Level1Load23[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_250_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load250[0] ), .Out({\Level2Out250[31] , \Level2Out250[30] , 
        \Level2Out250[29] , \Level2Out250[28] , \Level2Out250[27] , 
        \Level2Out250[26] , \Level2Out250[25] , \Level2Out250[24] , 
        \Level2Out250[23] , \Level2Out250[22] , \Level2Out250[21] , 
        \Level2Out250[20] , \Level2Out250[19] , \Level2Out250[18] , 
        \Level2Out250[17] , \Level2Out250[16] , \Level2Out250[15] , 
        \Level2Out250[14] , \Level2Out250[13] , \Level2Out250[12] , 
        \Level2Out250[11] , \Level2Out250[10] , \Level2Out250[9] , 
        \Level2Out250[8] , \Level2Out250[7] , \Level2Out250[6] , 
        \Level2Out250[5] , \Level2Out250[4] , \Level2Out250[3] , 
        \Level2Out250[2] , \Level2Out250[1] , \Level2Out250[0] }), .In1({
        \Level1Out250[31] , \Level1Out250[30] , \Level1Out250[29] , 
        \Level1Out250[28] , \Level1Out250[27] , \Level1Out250[26] , 
        \Level1Out250[25] , \Level1Out250[24] , \Level1Out250[23] , 
        \Level1Out250[22] , \Level1Out250[21] , \Level1Out250[20] , 
        \Level1Out250[19] , \Level1Out250[18] , \Level1Out250[17] , 
        \Level1Out250[16] , \Level1Out250[15] , \Level1Out250[14] , 
        \Level1Out250[13] , \Level1Out250[12] , \Level1Out250[11] , 
        \Level1Out250[10] , \Level1Out250[9] , \Level1Out250[8] , 
        \Level1Out250[7] , \Level1Out250[6] , \Level1Out250[5] , 
        \Level1Out250[4] , \Level1Out250[3] , \Level1Out250[2] , 
        \Level1Out250[1] , \Level1Out250[0] }), .In2({\Level1Out251[31] , 
        \Level1Out251[30] , \Level1Out251[29] , \Level1Out251[28] , 
        \Level1Out251[27] , \Level1Out251[26] , \Level1Out251[25] , 
        \Level1Out251[24] , \Level1Out251[23] , \Level1Out251[22] , 
        \Level1Out251[21] , \Level1Out251[20] , \Level1Out251[19] , 
        \Level1Out251[18] , \Level1Out251[17] , \Level1Out251[16] , 
        \Level1Out251[15] , \Level1Out251[14] , \Level1Out251[13] , 
        \Level1Out251[12] , \Level1Out251[11] , \Level1Out251[10] , 
        \Level1Out251[9] , \Level1Out251[8] , \Level1Out251[7] , 
        \Level1Out251[6] , \Level1Out251[5] , \Level1Out251[4] , 
        \Level1Out251[3] , \Level1Out251[2] , \Level1Out251[1] , 
        \Level1Out251[0] }), .Read1(\Level1Load250[0] ), .Read2(
        \Level1Load251[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_80_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load80[0] ), .Out({\Level8Out80[31] , \Level8Out80[30] , 
        \Level8Out80[29] , \Level8Out80[28] , \Level8Out80[27] , 
        \Level8Out80[26] , \Level8Out80[25] , \Level8Out80[24] , 
        \Level8Out80[23] , \Level8Out80[22] , \Level8Out80[21] , 
        \Level8Out80[20] , \Level8Out80[19] , \Level8Out80[18] , 
        \Level8Out80[17] , \Level8Out80[16] , \Level8Out80[15] , 
        \Level8Out80[14] , \Level8Out80[13] , \Level8Out80[12] , 
        \Level8Out80[11] , \Level8Out80[10] , \Level8Out80[9] , 
        \Level8Out80[8] , \Level8Out80[7] , \Level8Out80[6] , \Level8Out80[5] , 
        \Level8Out80[4] , \Level8Out80[3] , \Level8Out80[2] , \Level8Out80[1] , 
        \Level8Out80[0] }), .In1({\Level4Out80[31] , \Level4Out80[30] , 
        \Level4Out80[29] , \Level4Out80[28] , \Level4Out80[27] , 
        \Level4Out80[26] , \Level4Out80[25] , \Level4Out80[24] , 
        \Level4Out80[23] , \Level4Out80[22] , \Level4Out80[21] , 
        \Level4Out80[20] , \Level4Out80[19] , \Level4Out80[18] , 
        \Level4Out80[17] , \Level4Out80[16] , \Level4Out80[15] , 
        \Level4Out80[14] , \Level4Out80[13] , \Level4Out80[12] , 
        \Level4Out80[11] , \Level4Out80[10] , \Level4Out80[9] , 
        \Level4Out80[8] , \Level4Out80[7] , \Level4Out80[6] , \Level4Out80[5] , 
        \Level4Out80[4] , \Level4Out80[3] , \Level4Out80[2] , \Level4Out80[1] , 
        \Level4Out80[0] }), .In2({\Level4Out84[31] , \Level4Out84[30] , 
        \Level4Out84[29] , \Level4Out84[28] , \Level4Out84[27] , 
        \Level4Out84[26] , \Level4Out84[25] , \Level4Out84[24] , 
        \Level4Out84[23] , \Level4Out84[22] , \Level4Out84[21] , 
        \Level4Out84[20] , \Level4Out84[19] , \Level4Out84[18] , 
        \Level4Out84[17] , \Level4Out84[16] , \Level4Out84[15] , 
        \Level4Out84[14] , \Level4Out84[13] , \Level4Out84[12] , 
        \Level4Out84[11] , \Level4Out84[10] , \Level4Out84[9] , 
        \Level4Out84[8] , \Level4Out84[7] , \Level4Out84[6] , \Level4Out84[5] , 
        \Level4Out84[4] , \Level4Out84[3] , \Level4Out84[2] , \Level4Out84[1] , 
        \Level4Out84[0] }), .Read1(\Level4Load80[0] ), .Read2(
        \Level4Load84[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_152_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load152[0] ), .Out({\Level4Out152[31] , \Level4Out152[30] , 
        \Level4Out152[29] , \Level4Out152[28] , \Level4Out152[27] , 
        \Level4Out152[26] , \Level4Out152[25] , \Level4Out152[24] , 
        \Level4Out152[23] , \Level4Out152[22] , \Level4Out152[21] , 
        \Level4Out152[20] , \Level4Out152[19] , \Level4Out152[18] , 
        \Level4Out152[17] , \Level4Out152[16] , \Level4Out152[15] , 
        \Level4Out152[14] , \Level4Out152[13] , \Level4Out152[12] , 
        \Level4Out152[11] , \Level4Out152[10] , \Level4Out152[9] , 
        \Level4Out152[8] , \Level4Out152[7] , \Level4Out152[6] , 
        \Level4Out152[5] , \Level4Out152[4] , \Level4Out152[3] , 
        \Level4Out152[2] , \Level4Out152[1] , \Level4Out152[0] }), .In1({
        \Level2Out152[31] , \Level2Out152[30] , \Level2Out152[29] , 
        \Level2Out152[28] , \Level2Out152[27] , \Level2Out152[26] , 
        \Level2Out152[25] , \Level2Out152[24] , \Level2Out152[23] , 
        \Level2Out152[22] , \Level2Out152[21] , \Level2Out152[20] , 
        \Level2Out152[19] , \Level2Out152[18] , \Level2Out152[17] , 
        \Level2Out152[16] , \Level2Out152[15] , \Level2Out152[14] , 
        \Level2Out152[13] , \Level2Out152[12] , \Level2Out152[11] , 
        \Level2Out152[10] , \Level2Out152[9] , \Level2Out152[8] , 
        \Level2Out152[7] , \Level2Out152[6] , \Level2Out152[5] , 
        \Level2Out152[4] , \Level2Out152[3] , \Level2Out152[2] , 
        \Level2Out152[1] , \Level2Out152[0] }), .In2({\Level2Out154[31] , 
        \Level2Out154[30] , \Level2Out154[29] , \Level2Out154[28] , 
        \Level2Out154[27] , \Level2Out154[26] , \Level2Out154[25] , 
        \Level2Out154[24] , \Level2Out154[23] , \Level2Out154[22] , 
        \Level2Out154[21] , \Level2Out154[20] , \Level2Out154[19] , 
        \Level2Out154[18] , \Level2Out154[17] , \Level2Out154[16] , 
        \Level2Out154[15] , \Level2Out154[14] , \Level2Out154[13] , 
        \Level2Out154[12] , \Level2Out154[11] , \Level2Out154[10] , 
        \Level2Out154[9] , \Level2Out154[8] , \Level2Out154[7] , 
        \Level2Out154[6] , \Level2Out154[5] , \Level2Out154[4] , 
        \Level2Out154[3] , \Level2Out154[2] , \Level2Out154[1] , 
        \Level2Out154[0] }), .Read1(\Level2Load152[0] ), .Read2(
        \Level2Load154[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_35 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanOut({\ScanLink36[31] , 
        \ScanLink36[30] , \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , 
        \ScanLink36[26] , \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , 
        \ScanLink36[22] , \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , 
        \ScanLink36[18] , \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , 
        \ScanLink36[14] , \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , 
        \ScanLink36[10] , \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , 
        \ScanLink36[6] , \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , 
        \ScanLink36[2] , \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load35[0] ), .Out({
        \Level1Out35[31] , \Level1Out35[30] , \Level1Out35[29] , 
        \Level1Out35[28] , \Level1Out35[27] , \Level1Out35[26] , 
        \Level1Out35[25] , \Level1Out35[24] , \Level1Out35[23] , 
        \Level1Out35[22] , \Level1Out35[21] , \Level1Out35[20] , 
        \Level1Out35[19] , \Level1Out35[18] , \Level1Out35[17] , 
        \Level1Out35[16] , \Level1Out35[15] , \Level1Out35[14] , 
        \Level1Out35[13] , \Level1Out35[12] , \Level1Out35[11] , 
        \Level1Out35[10] , \Level1Out35[9] , \Level1Out35[8] , 
        \Level1Out35[7] , \Level1Out35[6] , \Level1Out35[5] , \Level1Out35[4] , 
        \Level1Out35[3] , \Level1Out35[2] , \Level1Out35[1] , \Level1Out35[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_40 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanOut({\ScanLink41[31] , 
        \ScanLink41[30] , \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , 
        \ScanLink41[26] , \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , 
        \ScanLink41[22] , \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , 
        \ScanLink41[18] , \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , 
        \ScanLink41[14] , \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , 
        \ScanLink41[10] , \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , 
        \ScanLink41[6] , \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , 
        \ScanLink41[2] , \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load40[0] ), .Out({
        \Level1Out40[31] , \Level1Out40[30] , \Level1Out40[29] , 
        \Level1Out40[28] , \Level1Out40[27] , \Level1Out40[26] , 
        \Level1Out40[25] , \Level1Out40[24] , \Level1Out40[23] , 
        \Level1Out40[22] , \Level1Out40[21] , \Level1Out40[20] , 
        \Level1Out40[19] , \Level1Out40[18] , \Level1Out40[17] , 
        \Level1Out40[16] , \Level1Out40[15] , \Level1Out40[14] , 
        \Level1Out40[13] , \Level1Out40[12] , \Level1Out40[11] , 
        \Level1Out40[10] , \Level1Out40[9] , \Level1Out40[8] , 
        \Level1Out40[7] , \Level1Out40[6] , \Level1Out40[5] , \Level1Out40[4] , 
        \Level1Out40[3] , \Level1Out40[2] , \Level1Out40[1] , \Level1Out40[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_82 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink82[31] , \ScanLink82[30] , 
        \ScanLink82[29] , \ScanLink82[28] , \ScanLink82[27] , \ScanLink82[26] , 
        \ScanLink82[25] , \ScanLink82[24] , \ScanLink82[23] , \ScanLink82[22] , 
        \ScanLink82[21] , \ScanLink82[20] , \ScanLink82[19] , \ScanLink82[18] , 
        \ScanLink82[17] , \ScanLink82[16] , \ScanLink82[15] , \ScanLink82[14] , 
        \ScanLink82[13] , \ScanLink82[12] , \ScanLink82[11] , \ScanLink82[10] , 
        \ScanLink82[9] , \ScanLink82[8] , \ScanLink82[7] , \ScanLink82[6] , 
        \ScanLink82[5] , \ScanLink82[4] , \ScanLink82[3] , \ScanLink82[2] , 
        \ScanLink82[1] , \ScanLink82[0] }), .ScanOut({\ScanLink83[31] , 
        \ScanLink83[30] , \ScanLink83[29] , \ScanLink83[28] , \ScanLink83[27] , 
        \ScanLink83[26] , \ScanLink83[25] , \ScanLink83[24] , \ScanLink83[23] , 
        \ScanLink83[22] , \ScanLink83[21] , \ScanLink83[20] , \ScanLink83[19] , 
        \ScanLink83[18] , \ScanLink83[17] , \ScanLink83[16] , \ScanLink83[15] , 
        \ScanLink83[14] , \ScanLink83[13] , \ScanLink83[12] , \ScanLink83[11] , 
        \ScanLink83[10] , \ScanLink83[9] , \ScanLink83[8] , \ScanLink83[7] , 
        \ScanLink83[6] , \ScanLink83[5] , \ScanLink83[4] , \ScanLink83[3] , 
        \ScanLink83[2] , \ScanLink83[1] , \ScanLink83[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load82[0] ), .Out({
        \Level1Out82[31] , \Level1Out82[30] , \Level1Out82[29] , 
        \Level1Out82[28] , \Level1Out82[27] , \Level1Out82[26] , 
        \Level1Out82[25] , \Level1Out82[24] , \Level1Out82[23] , 
        \Level1Out82[22] , \Level1Out82[21] , \Level1Out82[20] , 
        \Level1Out82[19] , \Level1Out82[18] , \Level1Out82[17] , 
        \Level1Out82[16] , \Level1Out82[15] , \Level1Out82[14] , 
        \Level1Out82[13] , \Level1Out82[12] , \Level1Out82[11] , 
        \Level1Out82[10] , \Level1Out82[9] , \Level1Out82[8] , 
        \Level1Out82[7] , \Level1Out82[6] , \Level1Out82[5] , \Level1Out82[4] , 
        \Level1Out82[3] , \Level1Out82[2] , \Level1Out82[1] , \Level1Out82[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_184_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load184[0] ), .Out({\Level4Out184[31] , \Level4Out184[30] , 
        \Level4Out184[29] , \Level4Out184[28] , \Level4Out184[27] , 
        \Level4Out184[26] , \Level4Out184[25] , \Level4Out184[24] , 
        \Level4Out184[23] , \Level4Out184[22] , \Level4Out184[21] , 
        \Level4Out184[20] , \Level4Out184[19] , \Level4Out184[18] , 
        \Level4Out184[17] , \Level4Out184[16] , \Level4Out184[15] , 
        \Level4Out184[14] , \Level4Out184[13] , \Level4Out184[12] , 
        \Level4Out184[11] , \Level4Out184[10] , \Level4Out184[9] , 
        \Level4Out184[8] , \Level4Out184[7] , \Level4Out184[6] , 
        \Level4Out184[5] , \Level4Out184[4] , \Level4Out184[3] , 
        \Level4Out184[2] , \Level4Out184[1] , \Level4Out184[0] }), .In1({
        \Level2Out184[31] , \Level2Out184[30] , \Level2Out184[29] , 
        \Level2Out184[28] , \Level2Out184[27] , \Level2Out184[26] , 
        \Level2Out184[25] , \Level2Out184[24] , \Level2Out184[23] , 
        \Level2Out184[22] , \Level2Out184[21] , \Level2Out184[20] , 
        \Level2Out184[19] , \Level2Out184[18] , \Level2Out184[17] , 
        \Level2Out184[16] , \Level2Out184[15] , \Level2Out184[14] , 
        \Level2Out184[13] , \Level2Out184[12] , \Level2Out184[11] , 
        \Level2Out184[10] , \Level2Out184[9] , \Level2Out184[8] , 
        \Level2Out184[7] , \Level2Out184[6] , \Level2Out184[5] , 
        \Level2Out184[4] , \Level2Out184[3] , \Level2Out184[2] , 
        \Level2Out184[1] , \Level2Out184[0] }), .In2({\Level2Out186[31] , 
        \Level2Out186[30] , \Level2Out186[29] , \Level2Out186[28] , 
        \Level2Out186[27] , \Level2Out186[26] , \Level2Out186[25] , 
        \Level2Out186[24] , \Level2Out186[23] , \Level2Out186[22] , 
        \Level2Out186[21] , \Level2Out186[20] , \Level2Out186[19] , 
        \Level2Out186[18] , \Level2Out186[17] , \Level2Out186[16] , 
        \Level2Out186[15] , \Level2Out186[14] , \Level2Out186[13] , 
        \Level2Out186[12] , \Level2Out186[11] , \Level2Out186[10] , 
        \Level2Out186[9] , \Level2Out186[8] , \Level2Out186[7] , 
        \Level2Out186[6] , \Level2Out186[5] , \Level2Out186[4] , 
        \Level2Out186[3] , \Level2Out186[2] , \Level2Out186[1] , 
        \Level2Out186[0] }), .Read1(\Level2Load184[0] ), .Read2(
        \Level2Load186[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load16[0] ), .Out({\Level8Out16[31] , \Level8Out16[30] , 
        \Level8Out16[29] , \Level8Out16[28] , \Level8Out16[27] , 
        \Level8Out16[26] , \Level8Out16[25] , \Level8Out16[24] , 
        \Level8Out16[23] , \Level8Out16[22] , \Level8Out16[21] , 
        \Level8Out16[20] , \Level8Out16[19] , \Level8Out16[18] , 
        \Level8Out16[17] , \Level8Out16[16] , \Level8Out16[15] , 
        \Level8Out16[14] , \Level8Out16[13] , \Level8Out16[12] , 
        \Level8Out16[11] , \Level8Out16[10] , \Level8Out16[9] , 
        \Level8Out16[8] , \Level8Out16[7] , \Level8Out16[6] , \Level8Out16[5] , 
        \Level8Out16[4] , \Level8Out16[3] , \Level8Out16[2] , \Level8Out16[1] , 
        \Level8Out16[0] }), .In1({\Level4Out16[31] , \Level4Out16[30] , 
        \Level4Out16[29] , \Level4Out16[28] , \Level4Out16[27] , 
        \Level4Out16[26] , \Level4Out16[25] , \Level4Out16[24] , 
        \Level4Out16[23] , \Level4Out16[22] , \Level4Out16[21] , 
        \Level4Out16[20] , \Level4Out16[19] , \Level4Out16[18] , 
        \Level4Out16[17] , \Level4Out16[16] , \Level4Out16[15] , 
        \Level4Out16[14] , \Level4Out16[13] , \Level4Out16[12] , 
        \Level4Out16[11] , \Level4Out16[10] , \Level4Out16[9] , 
        \Level4Out16[8] , \Level4Out16[7] , \Level4Out16[6] , \Level4Out16[5] , 
        \Level4Out16[4] , \Level4Out16[3] , \Level4Out16[2] , \Level4Out16[1] , 
        \Level4Out16[0] }), .In2({\Level4Out20[31] , \Level4Out20[30] , 
        \Level4Out20[29] , \Level4Out20[28] , \Level4Out20[27] , 
        \Level4Out20[26] , \Level4Out20[25] , \Level4Out20[24] , 
        \Level4Out20[23] , \Level4Out20[22] , \Level4Out20[21] , 
        \Level4Out20[20] , \Level4Out20[19] , \Level4Out20[18] , 
        \Level4Out20[17] , \Level4Out20[16] , \Level4Out20[15] , 
        \Level4Out20[14] , \Level4Out20[13] , \Level4Out20[12] , 
        \Level4Out20[11] , \Level4Out20[10] , \Level4Out20[9] , 
        \Level4Out20[8] , \Level4Out20[7] , \Level4Out20[6] , \Level4Out20[5] , 
        \Level4Out20[4] , \Level4Out20[3] , \Level4Out20[2] , \Level4Out20[1] , 
        \Level4Out20[0] }), .Read1(\Level4Load16[0] ), .Read2(
        \Level4Load20[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_187 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink187[31] , \ScanLink187[30] , 
        \ScanLink187[29] , \ScanLink187[28] , \ScanLink187[27] , 
        \ScanLink187[26] , \ScanLink187[25] , \ScanLink187[24] , 
        \ScanLink187[23] , \ScanLink187[22] , \ScanLink187[21] , 
        \ScanLink187[20] , \ScanLink187[19] , \ScanLink187[18] , 
        \ScanLink187[17] , \ScanLink187[16] , \ScanLink187[15] , 
        \ScanLink187[14] , \ScanLink187[13] , \ScanLink187[12] , 
        \ScanLink187[11] , \ScanLink187[10] , \ScanLink187[9] , 
        \ScanLink187[8] , \ScanLink187[7] , \ScanLink187[6] , \ScanLink187[5] , 
        \ScanLink187[4] , \ScanLink187[3] , \ScanLink187[2] , \ScanLink187[1] , 
        \ScanLink187[0] }), .ScanOut({\ScanLink188[31] , \ScanLink188[30] , 
        \ScanLink188[29] , \ScanLink188[28] , \ScanLink188[27] , 
        \ScanLink188[26] , \ScanLink188[25] , \ScanLink188[24] , 
        \ScanLink188[23] , \ScanLink188[22] , \ScanLink188[21] , 
        \ScanLink188[20] , \ScanLink188[19] , \ScanLink188[18] , 
        \ScanLink188[17] , \ScanLink188[16] , \ScanLink188[15] , 
        \ScanLink188[14] , \ScanLink188[13] , \ScanLink188[12] , 
        \ScanLink188[11] , \ScanLink188[10] , \ScanLink188[9] , 
        \ScanLink188[8] , \ScanLink188[7] , \ScanLink188[6] , \ScanLink188[5] , 
        \ScanLink188[4] , \ScanLink188[3] , \ScanLink188[2] , \ScanLink188[1] , 
        \ScanLink188[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load187[0] ), .Out({\Level1Out187[31] , \Level1Out187[30] , 
        \Level1Out187[29] , \Level1Out187[28] , \Level1Out187[27] , 
        \Level1Out187[26] , \Level1Out187[25] , \Level1Out187[24] , 
        \Level1Out187[23] , \Level1Out187[22] , \Level1Out187[21] , 
        \Level1Out187[20] , \Level1Out187[19] , \Level1Out187[18] , 
        \Level1Out187[17] , \Level1Out187[16] , \Level1Out187[15] , 
        \Level1Out187[14] , \Level1Out187[13] , \Level1Out187[12] , 
        \Level1Out187[11] , \Level1Out187[10] , \Level1Out187[9] , 
        \Level1Out187[8] , \Level1Out187[7] , \Level1Out187[6] , 
        \Level1Out187[5] , \Level1Out187[4] , \Level1Out187[3] , 
        \Level1Out187[2] , \Level1Out187[1] , \Level1Out187[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_198_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load198[0] ), .Out({\Level2Out198[31] , \Level2Out198[30] , 
        \Level2Out198[29] , \Level2Out198[28] , \Level2Out198[27] , 
        \Level2Out198[26] , \Level2Out198[25] , \Level2Out198[24] , 
        \Level2Out198[23] , \Level2Out198[22] , \Level2Out198[21] , 
        \Level2Out198[20] , \Level2Out198[19] , \Level2Out198[18] , 
        \Level2Out198[17] , \Level2Out198[16] , \Level2Out198[15] , 
        \Level2Out198[14] , \Level2Out198[13] , \Level2Out198[12] , 
        \Level2Out198[11] , \Level2Out198[10] , \Level2Out198[9] , 
        \Level2Out198[8] , \Level2Out198[7] , \Level2Out198[6] , 
        \Level2Out198[5] , \Level2Out198[4] , \Level2Out198[3] , 
        \Level2Out198[2] , \Level2Out198[1] , \Level2Out198[0] }), .In1({
        \Level1Out198[31] , \Level1Out198[30] , \Level1Out198[29] , 
        \Level1Out198[28] , \Level1Out198[27] , \Level1Out198[26] , 
        \Level1Out198[25] , \Level1Out198[24] , \Level1Out198[23] , 
        \Level1Out198[22] , \Level1Out198[21] , \Level1Out198[20] , 
        \Level1Out198[19] , \Level1Out198[18] , \Level1Out198[17] , 
        \Level1Out198[16] , \Level1Out198[15] , \Level1Out198[14] , 
        \Level1Out198[13] , \Level1Out198[12] , \Level1Out198[11] , 
        \Level1Out198[10] , \Level1Out198[9] , \Level1Out198[8] , 
        \Level1Out198[7] , \Level1Out198[6] , \Level1Out198[5] , 
        \Level1Out198[4] , \Level1Out198[3] , \Level1Out198[2] , 
        \Level1Out198[1] , \Level1Out198[0] }), .In2({\Level1Out199[31] , 
        \Level1Out199[30] , \Level1Out199[29] , \Level1Out199[28] , 
        \Level1Out199[27] , \Level1Out199[26] , \Level1Out199[25] , 
        \Level1Out199[24] , \Level1Out199[23] , \Level1Out199[22] , 
        \Level1Out199[21] , \Level1Out199[20] , \Level1Out199[19] , 
        \Level1Out199[18] , \Level1Out199[17] , \Level1Out199[16] , 
        \Level1Out199[15] , \Level1Out199[14] , \Level1Out199[13] , 
        \Level1Out199[12] , \Level1Out199[11] , \Level1Out199[10] , 
        \Level1Out199[9] , \Level1Out199[8] , \Level1Out199[7] , 
        \Level1Out199[6] , \Level1Out199[5] , \Level1Out199[4] , 
        \Level1Out199[3] , \Level1Out199[2] , \Level1Out199[1] , 
        \Level1Out199[0] }), .Read1(\Level1Load198[0] ), .Read2(
        \Level1Load199[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load56[0] ), .Out({\Level8Out56[31] , \Level8Out56[30] , 
        \Level8Out56[29] , \Level8Out56[28] , \Level8Out56[27] , 
        \Level8Out56[26] , \Level8Out56[25] , \Level8Out56[24] , 
        \Level8Out56[23] , \Level8Out56[22] , \Level8Out56[21] , 
        \Level8Out56[20] , \Level8Out56[19] , \Level8Out56[18] , 
        \Level8Out56[17] , \Level8Out56[16] , \Level8Out56[15] , 
        \Level8Out56[14] , \Level8Out56[13] , \Level8Out56[12] , 
        \Level8Out56[11] , \Level8Out56[10] , \Level8Out56[9] , 
        \Level8Out56[8] , \Level8Out56[7] , \Level8Out56[6] , \Level8Out56[5] , 
        \Level8Out56[4] , \Level8Out56[3] , \Level8Out56[2] , \Level8Out56[1] , 
        \Level8Out56[0] }), .In1({\Level4Out56[31] , \Level4Out56[30] , 
        \Level4Out56[29] , \Level4Out56[28] , \Level4Out56[27] , 
        \Level4Out56[26] , \Level4Out56[25] , \Level4Out56[24] , 
        \Level4Out56[23] , \Level4Out56[22] , \Level4Out56[21] , 
        \Level4Out56[20] , \Level4Out56[19] , \Level4Out56[18] , 
        \Level4Out56[17] , \Level4Out56[16] , \Level4Out56[15] , 
        \Level4Out56[14] , \Level4Out56[13] , \Level4Out56[12] , 
        \Level4Out56[11] , \Level4Out56[10] , \Level4Out56[9] , 
        \Level4Out56[8] , \Level4Out56[7] , \Level4Out56[6] , \Level4Out56[5] , 
        \Level4Out56[4] , \Level4Out56[3] , \Level4Out56[2] , \Level4Out56[1] , 
        \Level4Out56[0] }), .In2({\Level4Out60[31] , \Level4Out60[30] , 
        \Level4Out60[29] , \Level4Out60[28] , \Level4Out60[27] , 
        \Level4Out60[26] , \Level4Out60[25] , \Level4Out60[24] , 
        \Level4Out60[23] , \Level4Out60[22] , \Level4Out60[21] , 
        \Level4Out60[20] , \Level4Out60[19] , \Level4Out60[18] , 
        \Level4Out60[17] , \Level4Out60[16] , \Level4Out60[15] , 
        \Level4Out60[14] , \Level4Out60[13] , \Level4Out60[12] , 
        \Level4Out60[11] , \Level4Out60[10] , \Level4Out60[9] , 
        \Level4Out60[8] , \Level4Out60[7] , \Level4Out60[6] , \Level4Out60[5] , 
        \Level4Out60[4] , \Level4Out60[3] , \Level4Out60[2] , \Level4Out60[1] , 
        \Level4Out60[0] }), .Read1(\Level4Load56[0] ), .Read2(
        \Level4Load60[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_224_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load224[0] ), .Out({\Level8Out224[31] , \Level8Out224[30] , 
        \Level8Out224[29] , \Level8Out224[28] , \Level8Out224[27] , 
        \Level8Out224[26] , \Level8Out224[25] , \Level8Out224[24] , 
        \Level8Out224[23] , \Level8Out224[22] , \Level8Out224[21] , 
        \Level8Out224[20] , \Level8Out224[19] , \Level8Out224[18] , 
        \Level8Out224[17] , \Level8Out224[16] , \Level8Out224[15] , 
        \Level8Out224[14] , \Level8Out224[13] , \Level8Out224[12] , 
        \Level8Out224[11] , \Level8Out224[10] , \Level8Out224[9] , 
        \Level8Out224[8] , \Level8Out224[7] , \Level8Out224[6] , 
        \Level8Out224[5] , \Level8Out224[4] , \Level8Out224[3] , 
        \Level8Out224[2] , \Level8Out224[1] , \Level8Out224[0] }), .In1({
        \Level4Out224[31] , \Level4Out224[30] , \Level4Out224[29] , 
        \Level4Out224[28] , \Level4Out224[27] , \Level4Out224[26] , 
        \Level4Out224[25] , \Level4Out224[24] , \Level4Out224[23] , 
        \Level4Out224[22] , \Level4Out224[21] , \Level4Out224[20] , 
        \Level4Out224[19] , \Level4Out224[18] , \Level4Out224[17] , 
        \Level4Out224[16] , \Level4Out224[15] , \Level4Out224[14] , 
        \Level4Out224[13] , \Level4Out224[12] , \Level4Out224[11] , 
        \Level4Out224[10] , \Level4Out224[9] , \Level4Out224[8] , 
        \Level4Out224[7] , \Level4Out224[6] , \Level4Out224[5] , 
        \Level4Out224[4] , \Level4Out224[3] , \Level4Out224[2] , 
        \Level4Out224[1] , \Level4Out224[0] }), .In2({\Level4Out228[31] , 
        \Level4Out228[30] , \Level4Out228[29] , \Level4Out228[28] , 
        \Level4Out228[27] , \Level4Out228[26] , \Level4Out228[25] , 
        \Level4Out228[24] , \Level4Out228[23] , \Level4Out228[22] , 
        \Level4Out228[21] , \Level4Out228[20] , \Level4Out228[19] , 
        \Level4Out228[18] , \Level4Out228[17] , \Level4Out228[16] , 
        \Level4Out228[15] , \Level4Out228[14] , \Level4Out228[13] , 
        \Level4Out228[12] , \Level4Out228[11] , \Level4Out228[10] , 
        \Level4Out228[9] , \Level4Out228[8] , \Level4Out228[7] , 
        \Level4Out228[6] , \Level4Out228[5] , \Level4Out228[4] , 
        \Level4Out228[3] , \Level4Out228[2] , \Level4Out228[1] , 
        \Level4Out228[0] }), .Read1(\Level4Load224[0] ), .Read2(
        \Level4Load228[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load48[0] ), .Out({\Level2Out48[31] , \Level2Out48[30] , 
        \Level2Out48[29] , \Level2Out48[28] , \Level2Out48[27] , 
        \Level2Out48[26] , \Level2Out48[25] , \Level2Out48[24] , 
        \Level2Out48[23] , \Level2Out48[22] , \Level2Out48[21] , 
        \Level2Out48[20] , \Level2Out48[19] , \Level2Out48[18] , 
        \Level2Out48[17] , \Level2Out48[16] , \Level2Out48[15] , 
        \Level2Out48[14] , \Level2Out48[13] , \Level2Out48[12] , 
        \Level2Out48[11] , \Level2Out48[10] , \Level2Out48[9] , 
        \Level2Out48[8] , \Level2Out48[7] , \Level2Out48[6] , \Level2Out48[5] , 
        \Level2Out48[4] , \Level2Out48[3] , \Level2Out48[2] , \Level2Out48[1] , 
        \Level2Out48[0] }), .In1({\Level1Out48[31] , \Level1Out48[30] , 
        \Level1Out48[29] , \Level1Out48[28] , \Level1Out48[27] , 
        \Level1Out48[26] , \Level1Out48[25] , \Level1Out48[24] , 
        \Level1Out48[23] , \Level1Out48[22] , \Level1Out48[21] , 
        \Level1Out48[20] , \Level1Out48[19] , \Level1Out48[18] , 
        \Level1Out48[17] , \Level1Out48[16] , \Level1Out48[15] , 
        \Level1Out48[14] , \Level1Out48[13] , \Level1Out48[12] , 
        \Level1Out48[11] , \Level1Out48[10] , \Level1Out48[9] , 
        \Level1Out48[8] , \Level1Out48[7] , \Level1Out48[6] , \Level1Out48[5] , 
        \Level1Out48[4] , \Level1Out48[3] , \Level1Out48[2] , \Level1Out48[1] , 
        \Level1Out48[0] }), .In2({\Level1Out49[31] , \Level1Out49[30] , 
        \Level1Out49[29] , \Level1Out49[28] , \Level1Out49[27] , 
        \Level1Out49[26] , \Level1Out49[25] , \Level1Out49[24] , 
        \Level1Out49[23] , \Level1Out49[22] , \Level1Out49[21] , 
        \Level1Out49[20] , \Level1Out49[19] , \Level1Out49[18] , 
        \Level1Out49[17] , \Level1Out49[16] , \Level1Out49[15] , 
        \Level1Out49[14] , \Level1Out49[13] , \Level1Out49[12] , 
        \Level1Out49[11] , \Level1Out49[10] , \Level1Out49[9] , 
        \Level1Out49[8] , \Level1Out49[7] , \Level1Out49[6] , \Level1Out49[5] , 
        \Level1Out49[4] , \Level1Out49[3] , \Level1Out49[2] , \Level1Out49[1] , 
        \Level1Out49[0] }), .Read1(\Level1Load48[0] ), .Read2(
        \Level1Load49[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_62_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load62[0] ), .Out({\Level2Out62[31] , \Level2Out62[30] , 
        \Level2Out62[29] , \Level2Out62[28] , \Level2Out62[27] , 
        \Level2Out62[26] , \Level2Out62[25] , \Level2Out62[24] , 
        \Level2Out62[23] , \Level2Out62[22] , \Level2Out62[21] , 
        \Level2Out62[20] , \Level2Out62[19] , \Level2Out62[18] , 
        \Level2Out62[17] , \Level2Out62[16] , \Level2Out62[15] , 
        \Level2Out62[14] , \Level2Out62[13] , \Level2Out62[12] , 
        \Level2Out62[11] , \Level2Out62[10] , \Level2Out62[9] , 
        \Level2Out62[8] , \Level2Out62[7] , \Level2Out62[6] , \Level2Out62[5] , 
        \Level2Out62[4] , \Level2Out62[3] , \Level2Out62[2] , \Level2Out62[1] , 
        \Level2Out62[0] }), .In1({\Level1Out62[31] , \Level1Out62[30] , 
        \Level1Out62[29] , \Level1Out62[28] , \Level1Out62[27] , 
        \Level1Out62[26] , \Level1Out62[25] , \Level1Out62[24] , 
        \Level1Out62[23] , \Level1Out62[22] , \Level1Out62[21] , 
        \Level1Out62[20] , \Level1Out62[19] , \Level1Out62[18] , 
        \Level1Out62[17] , \Level1Out62[16] , \Level1Out62[15] , 
        \Level1Out62[14] , \Level1Out62[13] , \Level1Out62[12] , 
        \Level1Out62[11] , \Level1Out62[10] , \Level1Out62[9] , 
        \Level1Out62[8] , \Level1Out62[7] , \Level1Out62[6] , \Level1Out62[5] , 
        \Level1Out62[4] , \Level1Out62[3] , \Level1Out62[2] , \Level1Out62[1] , 
        \Level1Out62[0] }), .In2({\Level1Out63[31] , \Level1Out63[30] , 
        \Level1Out63[29] , \Level1Out63[28] , \Level1Out63[27] , 
        \Level1Out63[26] , \Level1Out63[25] , \Level1Out63[24] , 
        \Level1Out63[23] , \Level1Out63[22] , \Level1Out63[21] , 
        \Level1Out63[20] , \Level1Out63[19] , \Level1Out63[18] , 
        \Level1Out63[17] , \Level1Out63[16] , \Level1Out63[15] , 
        \Level1Out63[14] , \Level1Out63[13] , \Level1Out63[12] , 
        \Level1Out63[11] , \Level1Out63[10] , \Level1Out63[9] , 
        \Level1Out63[8] , \Level1Out63[7] , \Level1Out63[6] , \Level1Out63[5] , 
        \Level1Out63[4] , \Level1Out63[3] , \Level1Out63[2] , \Level1Out63[1] , 
        \Level1Out63[0] }), .Read1(\Level1Load62[0] ), .Read2(
        \Level1Load63[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_124_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load124[0] ), .Out({\Level2Out124[31] , \Level2Out124[30] , 
        \Level2Out124[29] , \Level2Out124[28] , \Level2Out124[27] , 
        \Level2Out124[26] , \Level2Out124[25] , \Level2Out124[24] , 
        \Level2Out124[23] , \Level2Out124[22] , \Level2Out124[21] , 
        \Level2Out124[20] , \Level2Out124[19] , \Level2Out124[18] , 
        \Level2Out124[17] , \Level2Out124[16] , \Level2Out124[15] , 
        \Level2Out124[14] , \Level2Out124[13] , \Level2Out124[12] , 
        \Level2Out124[11] , \Level2Out124[10] , \Level2Out124[9] , 
        \Level2Out124[8] , \Level2Out124[7] , \Level2Out124[6] , 
        \Level2Out124[5] , \Level2Out124[4] , \Level2Out124[3] , 
        \Level2Out124[2] , \Level2Out124[1] , \Level2Out124[0] }), .In1({
        \Level1Out124[31] , \Level1Out124[30] , \Level1Out124[29] , 
        \Level1Out124[28] , \Level1Out124[27] , \Level1Out124[26] , 
        \Level1Out124[25] , \Level1Out124[24] , \Level1Out124[23] , 
        \Level1Out124[22] , \Level1Out124[21] , \Level1Out124[20] , 
        \Level1Out124[19] , \Level1Out124[18] , \Level1Out124[17] , 
        \Level1Out124[16] , \Level1Out124[15] , \Level1Out124[14] , 
        \Level1Out124[13] , \Level1Out124[12] , \Level1Out124[11] , 
        \Level1Out124[10] , \Level1Out124[9] , \Level1Out124[8] , 
        \Level1Out124[7] , \Level1Out124[6] , \Level1Out124[5] , 
        \Level1Out124[4] , \Level1Out124[3] , \Level1Out124[2] , 
        \Level1Out124[1] , \Level1Out124[0] }), .In2({\Level1Out125[31] , 
        \Level1Out125[30] , \Level1Out125[29] , \Level1Out125[28] , 
        \Level1Out125[27] , \Level1Out125[26] , \Level1Out125[25] , 
        \Level1Out125[24] , \Level1Out125[23] , \Level1Out125[22] , 
        \Level1Out125[21] , \Level1Out125[20] , \Level1Out125[19] , 
        \Level1Out125[18] , \Level1Out125[17] , \Level1Out125[16] , 
        \Level1Out125[15] , \Level1Out125[14] , \Level1Out125[13] , 
        \Level1Out125[12] , \Level1Out125[11] , \Level1Out125[10] , 
        \Level1Out125[9] , \Level1Out125[8] , \Level1Out125[7] , 
        \Level1Out125[6] , \Level1Out125[5] , \Level1Out125[4] , 
        \Level1Out125[3] , \Level1Out125[2] , \Level1Out125[1] , 
        \Level1Out125[0] }), .Read1(\Level1Load124[0] ), .Read2(
        \Level1Load125[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_210_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load210[0] ), .Out({\Level2Out210[31] , \Level2Out210[30] , 
        \Level2Out210[29] , \Level2Out210[28] , \Level2Out210[27] , 
        \Level2Out210[26] , \Level2Out210[25] , \Level2Out210[24] , 
        \Level2Out210[23] , \Level2Out210[22] , \Level2Out210[21] , 
        \Level2Out210[20] , \Level2Out210[19] , \Level2Out210[18] , 
        \Level2Out210[17] , \Level2Out210[16] , \Level2Out210[15] , 
        \Level2Out210[14] , \Level2Out210[13] , \Level2Out210[12] , 
        \Level2Out210[11] , \Level2Out210[10] , \Level2Out210[9] , 
        \Level2Out210[8] , \Level2Out210[7] , \Level2Out210[6] , 
        \Level2Out210[5] , \Level2Out210[4] , \Level2Out210[3] , 
        \Level2Out210[2] , \Level2Out210[1] , \Level2Out210[0] }), .In1({
        \Level1Out210[31] , \Level1Out210[30] , \Level1Out210[29] , 
        \Level1Out210[28] , \Level1Out210[27] , \Level1Out210[26] , 
        \Level1Out210[25] , \Level1Out210[24] , \Level1Out210[23] , 
        \Level1Out210[22] , \Level1Out210[21] , \Level1Out210[20] , 
        \Level1Out210[19] , \Level1Out210[18] , \Level1Out210[17] , 
        \Level1Out210[16] , \Level1Out210[15] , \Level1Out210[14] , 
        \Level1Out210[13] , \Level1Out210[12] , \Level1Out210[11] , 
        \Level1Out210[10] , \Level1Out210[9] , \Level1Out210[8] , 
        \Level1Out210[7] , \Level1Out210[6] , \Level1Out210[5] , 
        \Level1Out210[4] , \Level1Out210[3] , \Level1Out210[2] , 
        \Level1Out210[1] , \Level1Out210[0] }), .In2({\Level1Out211[31] , 
        \Level1Out211[30] , \Level1Out211[29] , \Level1Out211[28] , 
        \Level1Out211[27] , \Level1Out211[26] , \Level1Out211[25] , 
        \Level1Out211[24] , \Level1Out211[23] , \Level1Out211[22] , 
        \Level1Out211[21] , \Level1Out211[20] , \Level1Out211[19] , 
        \Level1Out211[18] , \Level1Out211[17] , \Level1Out211[16] , 
        \Level1Out211[15] , \Level1Out211[14] , \Level1Out211[13] , 
        \Level1Out211[12] , \Level1Out211[11] , \Level1Out211[10] , 
        \Level1Out211[9] , \Level1Out211[8] , \Level1Out211[7] , 
        \Level1Out211[6] , \Level1Out211[5] , \Level1Out211[4] , 
        \Level1Out211[3] , \Level1Out211[2] , \Level1Out211[1] , 
        \Level1Out211[0] }), .Read1(\Level1Load210[0] ), .Read2(
        \Level1Load211[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_112_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load112[0] ), .Out({\Level4Out112[31] , \Level4Out112[30] , 
        \Level4Out112[29] , \Level4Out112[28] , \Level4Out112[27] , 
        \Level4Out112[26] , \Level4Out112[25] , \Level4Out112[24] , 
        \Level4Out112[23] , \Level4Out112[22] , \Level4Out112[21] , 
        \Level4Out112[20] , \Level4Out112[19] , \Level4Out112[18] , 
        \Level4Out112[17] , \Level4Out112[16] , \Level4Out112[15] , 
        \Level4Out112[14] , \Level4Out112[13] , \Level4Out112[12] , 
        \Level4Out112[11] , \Level4Out112[10] , \Level4Out112[9] , 
        \Level4Out112[8] , \Level4Out112[7] , \Level4Out112[6] , 
        \Level4Out112[5] , \Level4Out112[4] , \Level4Out112[3] , 
        \Level4Out112[2] , \Level4Out112[1] , \Level4Out112[0] }), .In1({
        \Level2Out112[31] , \Level2Out112[30] , \Level2Out112[29] , 
        \Level2Out112[28] , \Level2Out112[27] , \Level2Out112[26] , 
        \Level2Out112[25] , \Level2Out112[24] , \Level2Out112[23] , 
        \Level2Out112[22] , \Level2Out112[21] , \Level2Out112[20] , 
        \Level2Out112[19] , \Level2Out112[18] , \Level2Out112[17] , 
        \Level2Out112[16] , \Level2Out112[15] , \Level2Out112[14] , 
        \Level2Out112[13] , \Level2Out112[12] , \Level2Out112[11] , 
        \Level2Out112[10] , \Level2Out112[9] , \Level2Out112[8] , 
        \Level2Out112[7] , \Level2Out112[6] , \Level2Out112[5] , 
        \Level2Out112[4] , \Level2Out112[3] , \Level2Out112[2] , 
        \Level2Out112[1] , \Level2Out112[0] }), .In2({\Level2Out114[31] , 
        \Level2Out114[30] , \Level2Out114[29] , \Level2Out114[28] , 
        \Level2Out114[27] , \Level2Out114[26] , \Level2Out114[25] , 
        \Level2Out114[24] , \Level2Out114[23] , \Level2Out114[22] , 
        \Level2Out114[21] , \Level2Out114[20] , \Level2Out114[19] , 
        \Level2Out114[18] , \Level2Out114[17] , \Level2Out114[16] , 
        \Level2Out114[15] , \Level2Out114[14] , \Level2Out114[13] , 
        \Level2Out114[12] , \Level2Out114[11] , \Level2Out114[10] , 
        \Level2Out114[9] , \Level2Out114[8] , \Level2Out114[7] , 
        \Level2Out114[6] , \Level2Out114[5] , \Level2Out114[4] , 
        \Level2Out114[3] , \Level2Out114[2] , \Level2Out114[1] , 
        \Level2Out114[0] }), .Read1(\Level2Load112[0] ), .Read2(
        \Level2Load114[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load48[0] ), .Out({\Level16Out48[31] , \Level16Out48[30] , 
        \Level16Out48[29] , \Level16Out48[28] , \Level16Out48[27] , 
        \Level16Out48[26] , \Level16Out48[25] , \Level16Out48[24] , 
        \Level16Out48[23] , \Level16Out48[22] , \Level16Out48[21] , 
        \Level16Out48[20] , \Level16Out48[19] , \Level16Out48[18] , 
        \Level16Out48[17] , \Level16Out48[16] , \Level16Out48[15] , 
        \Level16Out48[14] , \Level16Out48[13] , \Level16Out48[12] , 
        \Level16Out48[11] , \Level16Out48[10] , \Level16Out48[9] , 
        \Level16Out48[8] , \Level16Out48[7] , \Level16Out48[6] , 
        \Level16Out48[5] , \Level16Out48[4] , \Level16Out48[3] , 
        \Level16Out48[2] , \Level16Out48[1] , \Level16Out48[0] }), .In1({
        \Level8Out48[31] , \Level8Out48[30] , \Level8Out48[29] , 
        \Level8Out48[28] , \Level8Out48[27] , \Level8Out48[26] , 
        \Level8Out48[25] , \Level8Out48[24] , \Level8Out48[23] , 
        \Level8Out48[22] , \Level8Out48[21] , \Level8Out48[20] , 
        \Level8Out48[19] , \Level8Out48[18] , \Level8Out48[17] , 
        \Level8Out48[16] , \Level8Out48[15] , \Level8Out48[14] , 
        \Level8Out48[13] , \Level8Out48[12] , \Level8Out48[11] , 
        \Level8Out48[10] , \Level8Out48[9] , \Level8Out48[8] , 
        \Level8Out48[7] , \Level8Out48[6] , \Level8Out48[5] , \Level8Out48[4] , 
        \Level8Out48[3] , \Level8Out48[2] , \Level8Out48[1] , \Level8Out48[0] 
        }), .In2({\Level8Out56[31] , \Level8Out56[30] , \Level8Out56[29] , 
        \Level8Out56[28] , \Level8Out56[27] , \Level8Out56[26] , 
        \Level8Out56[25] , \Level8Out56[24] , \Level8Out56[23] , 
        \Level8Out56[22] , \Level8Out56[21] , \Level8Out56[20] , 
        \Level8Out56[19] , \Level8Out56[18] , \Level8Out56[17] , 
        \Level8Out56[16] , \Level8Out56[15] , \Level8Out56[14] , 
        \Level8Out56[13] , \Level8Out56[12] , \Level8Out56[11] , 
        \Level8Out56[10] , \Level8Out56[9] , \Level8Out56[8] , 
        \Level8Out56[7] , \Level8Out56[6] , \Level8Out56[5] , \Level8Out56[4] , 
        \Level8Out56[3] , \Level8Out56[2] , \Level8Out56[1] , \Level8Out56[0] 
        }), .Read1(\Level8Load48[0] ), .Read2(\Level8Load56[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_67 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink67[31] , \ScanLink67[30] , 
        \ScanLink67[29] , \ScanLink67[28] , \ScanLink67[27] , \ScanLink67[26] , 
        \ScanLink67[25] , \ScanLink67[24] , \ScanLink67[23] , \ScanLink67[22] , 
        \ScanLink67[21] , \ScanLink67[20] , \ScanLink67[19] , \ScanLink67[18] , 
        \ScanLink67[17] , \ScanLink67[16] , \ScanLink67[15] , \ScanLink67[14] , 
        \ScanLink67[13] , \ScanLink67[12] , \ScanLink67[11] , \ScanLink67[10] , 
        \ScanLink67[9] , \ScanLink67[8] , \ScanLink67[7] , \ScanLink67[6] , 
        \ScanLink67[5] , \ScanLink67[4] , \ScanLink67[3] , \ScanLink67[2] , 
        \ScanLink67[1] , \ScanLink67[0] }), .ScanOut({\ScanLink68[31] , 
        \ScanLink68[30] , \ScanLink68[29] , \ScanLink68[28] , \ScanLink68[27] , 
        \ScanLink68[26] , \ScanLink68[25] , \ScanLink68[24] , \ScanLink68[23] , 
        \ScanLink68[22] , \ScanLink68[21] , \ScanLink68[20] , \ScanLink68[19] , 
        \ScanLink68[18] , \ScanLink68[17] , \ScanLink68[16] , \ScanLink68[15] , 
        \ScanLink68[14] , \ScanLink68[13] , \ScanLink68[12] , \ScanLink68[11] , 
        \ScanLink68[10] , \ScanLink68[9] , \ScanLink68[8] , \ScanLink68[7] , 
        \ScanLink68[6] , \ScanLink68[5] , \ScanLink68[4] , \ScanLink68[3] , 
        \ScanLink68[2] , \ScanLink68[1] , \ScanLink68[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load67[0] ), .Out({
        \Level1Out67[31] , \Level1Out67[30] , \Level1Out67[29] , 
        \Level1Out67[28] , \Level1Out67[27] , \Level1Out67[26] , 
        \Level1Out67[25] , \Level1Out67[24] , \Level1Out67[23] , 
        \Level1Out67[22] , \Level1Out67[21] , \Level1Out67[20] , 
        \Level1Out67[19] , \Level1Out67[18] , \Level1Out67[17] , 
        \Level1Out67[16] , \Level1Out67[15] , \Level1Out67[14] , 
        \Level1Out67[13] , \Level1Out67[12] , \Level1Out67[11] , 
        \Level1Out67[10] , \Level1Out67[9] , \Level1Out67[8] , 
        \Level1Out67[7] , \Level1Out67[6] , \Level1Out67[5] , \Level1Out67[4] , 
        \Level1Out67[3] , \Level1Out67[2] , \Level1Out67[1] , \Level1Out67[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_145 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink145[31] , \ScanLink145[30] , 
        \ScanLink145[29] , \ScanLink145[28] , \ScanLink145[27] , 
        \ScanLink145[26] , \ScanLink145[25] , \ScanLink145[24] , 
        \ScanLink145[23] , \ScanLink145[22] , \ScanLink145[21] , 
        \ScanLink145[20] , \ScanLink145[19] , \ScanLink145[18] , 
        \ScanLink145[17] , \ScanLink145[16] , \ScanLink145[15] , 
        \ScanLink145[14] , \ScanLink145[13] , \ScanLink145[12] , 
        \ScanLink145[11] , \ScanLink145[10] , \ScanLink145[9] , 
        \ScanLink145[8] , \ScanLink145[7] , \ScanLink145[6] , \ScanLink145[5] , 
        \ScanLink145[4] , \ScanLink145[3] , \ScanLink145[2] , \ScanLink145[1] , 
        \ScanLink145[0] }), .ScanOut({\ScanLink146[31] , \ScanLink146[30] , 
        \ScanLink146[29] , \ScanLink146[28] , \ScanLink146[27] , 
        \ScanLink146[26] , \ScanLink146[25] , \ScanLink146[24] , 
        \ScanLink146[23] , \ScanLink146[22] , \ScanLink146[21] , 
        \ScanLink146[20] , \ScanLink146[19] , \ScanLink146[18] , 
        \ScanLink146[17] , \ScanLink146[16] , \ScanLink146[15] , 
        \ScanLink146[14] , \ScanLink146[13] , \ScanLink146[12] , 
        \ScanLink146[11] , \ScanLink146[10] , \ScanLink146[9] , 
        \ScanLink146[8] , \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , 
        \ScanLink146[4] , \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , 
        \ScanLink146[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load145[0] ), .Out({\Level1Out145[31] , \Level1Out145[30] , 
        \Level1Out145[29] , \Level1Out145[28] , \Level1Out145[27] , 
        \Level1Out145[26] , \Level1Out145[25] , \Level1Out145[24] , 
        \Level1Out145[23] , \Level1Out145[22] , \Level1Out145[21] , 
        \Level1Out145[20] , \Level1Out145[19] , \Level1Out145[18] , 
        \Level1Out145[17] , \Level1Out145[16] , \Level1Out145[15] , 
        \Level1Out145[14] , \Level1Out145[13] , \Level1Out145[12] , 
        \Level1Out145[11] , \Level1Out145[10] , \Level1Out145[9] , 
        \Level1Out145[8] , \Level1Out145[7] , \Level1Out145[6] , 
        \Level1Out145[5] , \Level1Out145[4] , \Level1Out145[3] , 
        \Level1Out145[2] , \Level1Out145[1] , \Level1Out145[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_162 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink162[31] , \ScanLink162[30] , 
        \ScanLink162[29] , \ScanLink162[28] , \ScanLink162[27] , 
        \ScanLink162[26] , \ScanLink162[25] , \ScanLink162[24] , 
        \ScanLink162[23] , \ScanLink162[22] , \ScanLink162[21] , 
        \ScanLink162[20] , \ScanLink162[19] , \ScanLink162[18] , 
        \ScanLink162[17] , \ScanLink162[16] , \ScanLink162[15] , 
        \ScanLink162[14] , \ScanLink162[13] , \ScanLink162[12] , 
        \ScanLink162[11] , \ScanLink162[10] , \ScanLink162[9] , 
        \ScanLink162[8] , \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , 
        \ScanLink162[4] , \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , 
        \ScanLink162[0] }), .ScanOut({\ScanLink163[31] , \ScanLink163[30] , 
        \ScanLink163[29] , \ScanLink163[28] , \ScanLink163[27] , 
        \ScanLink163[26] , \ScanLink163[25] , \ScanLink163[24] , 
        \ScanLink163[23] , \ScanLink163[22] , \ScanLink163[21] , 
        \ScanLink163[20] , \ScanLink163[19] , \ScanLink163[18] , 
        \ScanLink163[17] , \ScanLink163[16] , \ScanLink163[15] , 
        \ScanLink163[14] , \ScanLink163[13] , \ScanLink163[12] , 
        \ScanLink163[11] , \ScanLink163[10] , \ScanLink163[9] , 
        \ScanLink163[8] , \ScanLink163[7] , \ScanLink163[6] , \ScanLink163[5] , 
        \ScanLink163[4] , \ScanLink163[3] , \ScanLink163[2] , \ScanLink163[1] , 
        \ScanLink163[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load162[0] ), .Out({\Level1Out162[31] , \Level1Out162[30] , 
        \Level1Out162[29] , \Level1Out162[28] , \Level1Out162[27] , 
        \Level1Out162[26] , \Level1Out162[25] , \Level1Out162[24] , 
        \Level1Out162[23] , \Level1Out162[22] , \Level1Out162[21] , 
        \Level1Out162[20] , \Level1Out162[19] , \Level1Out162[18] , 
        \Level1Out162[17] , \Level1Out162[16] , \Level1Out162[15] , 
        \Level1Out162[14] , \Level1Out162[13] , \Level1Out162[12] , 
        \Level1Out162[11] , \Level1Out162[10] , \Level1Out162[9] , 
        \Level1Out162[8] , \Level1Out162[7] , \Level1Out162[6] , 
        \Level1Out162[5] , \Level1Out162[4] , \Level1Out162[3] , 
        \Level1Out162[2] , \Level1Out162[1] , \Level1Out162[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_179 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink179[31] , \ScanLink179[30] , 
        \ScanLink179[29] , \ScanLink179[28] , \ScanLink179[27] , 
        \ScanLink179[26] , \ScanLink179[25] , \ScanLink179[24] , 
        \ScanLink179[23] , \ScanLink179[22] , \ScanLink179[21] , 
        \ScanLink179[20] , \ScanLink179[19] , \ScanLink179[18] , 
        \ScanLink179[17] , \ScanLink179[16] , \ScanLink179[15] , 
        \ScanLink179[14] , \ScanLink179[13] , \ScanLink179[12] , 
        \ScanLink179[11] , \ScanLink179[10] , \ScanLink179[9] , 
        \ScanLink179[8] , \ScanLink179[7] , \ScanLink179[6] , \ScanLink179[5] , 
        \ScanLink179[4] , \ScanLink179[3] , \ScanLink179[2] , \ScanLink179[1] , 
        \ScanLink179[0] }), .ScanOut({\ScanLink180[31] , \ScanLink180[30] , 
        \ScanLink180[29] , \ScanLink180[28] , \ScanLink180[27] , 
        \ScanLink180[26] , \ScanLink180[25] , \ScanLink180[24] , 
        \ScanLink180[23] , \ScanLink180[22] , \ScanLink180[21] , 
        \ScanLink180[20] , \ScanLink180[19] , \ScanLink180[18] , 
        \ScanLink180[17] , \ScanLink180[16] , \ScanLink180[15] , 
        \ScanLink180[14] , \ScanLink180[13] , \ScanLink180[12] , 
        \ScanLink180[11] , \ScanLink180[10] , \ScanLink180[9] , 
        \ScanLink180[8] , \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , 
        \ScanLink180[4] , \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , 
        \ScanLink180[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load179[0] ), .Out({\Level1Out179[31] , \Level1Out179[30] , 
        \Level1Out179[29] , \Level1Out179[28] , \Level1Out179[27] , 
        \Level1Out179[26] , \Level1Out179[25] , \Level1Out179[24] , 
        \Level1Out179[23] , \Level1Out179[22] , \Level1Out179[21] , 
        \Level1Out179[20] , \Level1Out179[19] , \Level1Out179[18] , 
        \Level1Out179[17] , \Level1Out179[16] , \Level1Out179[15] , 
        \Level1Out179[14] , \Level1Out179[13] , \Level1Out179[12] , 
        \Level1Out179[11] , \Level1Out179[10] , \Level1Out179[9] , 
        \Level1Out179[8] , \Level1Out179[7] , \Level1Out179[6] , 
        \Level1Out179[5] , \Level1Out179[4] , \Level1Out179[3] , 
        \Level1Out179[2] , \Level1Out179[1] , \Level1Out179[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_249 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink249[31] , \ScanLink249[30] , 
        \ScanLink249[29] , \ScanLink249[28] , \ScanLink249[27] , 
        \ScanLink249[26] , \ScanLink249[25] , \ScanLink249[24] , 
        \ScanLink249[23] , \ScanLink249[22] , \ScanLink249[21] , 
        \ScanLink249[20] , \ScanLink249[19] , \ScanLink249[18] , 
        \ScanLink249[17] , \ScanLink249[16] , \ScanLink249[15] , 
        \ScanLink249[14] , \ScanLink249[13] , \ScanLink249[12] , 
        \ScanLink249[11] , \ScanLink249[10] , \ScanLink249[9] , 
        \ScanLink249[8] , \ScanLink249[7] , \ScanLink249[6] , \ScanLink249[5] , 
        \ScanLink249[4] , \ScanLink249[3] , \ScanLink249[2] , \ScanLink249[1] , 
        \ScanLink249[0] }), .ScanOut({\ScanLink250[31] , \ScanLink250[30] , 
        \ScanLink250[29] , \ScanLink250[28] , \ScanLink250[27] , 
        \ScanLink250[26] , \ScanLink250[25] , \ScanLink250[24] , 
        \ScanLink250[23] , \ScanLink250[22] , \ScanLink250[21] , 
        \ScanLink250[20] , \ScanLink250[19] , \ScanLink250[18] , 
        \ScanLink250[17] , \ScanLink250[16] , \ScanLink250[15] , 
        \ScanLink250[14] , \ScanLink250[13] , \ScanLink250[12] , 
        \ScanLink250[11] , \ScanLink250[10] , \ScanLink250[9] , 
        \ScanLink250[8] , \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , 
        \ScanLink250[4] , \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , 
        \ScanLink250[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load249[0] ), .Out({\Level1Out249[31] , \Level1Out249[30] , 
        \Level1Out249[29] , \Level1Out249[28] , \Level1Out249[27] , 
        \Level1Out249[26] , \Level1Out249[25] , \Level1Out249[24] , 
        \Level1Out249[23] , \Level1Out249[22] , \Level1Out249[21] , 
        \Level1Out249[20] , \Level1Out249[19] , \Level1Out249[18] , 
        \Level1Out249[17] , \Level1Out249[16] , \Level1Out249[15] , 
        \Level1Out249[14] , \Level1Out249[13] , \Level1Out249[12] , 
        \Level1Out249[11] , \Level1Out249[10] , \Level1Out249[9] , 
        \Level1Out249[8] , \Level1Out249[7] , \Level1Out249[6] , 
        \Level1Out249[5] , \Level1Out249[4] , \Level1Out249[3] , 
        \Level1Out249[2] , \Level1Out249[1] , \Level1Out249[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_252 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink252[31] , \ScanLink252[30] , 
        \ScanLink252[29] , \ScanLink252[28] , \ScanLink252[27] , 
        \ScanLink252[26] , \ScanLink252[25] , \ScanLink252[24] , 
        \ScanLink252[23] , \ScanLink252[22] , \ScanLink252[21] , 
        \ScanLink252[20] , \ScanLink252[19] , \ScanLink252[18] , 
        \ScanLink252[17] , \ScanLink252[16] , \ScanLink252[15] , 
        \ScanLink252[14] , \ScanLink252[13] , \ScanLink252[12] , 
        \ScanLink252[11] , \ScanLink252[10] , \ScanLink252[9] , 
        \ScanLink252[8] , \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , 
        \ScanLink252[4] , \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , 
        \ScanLink252[0] }), .ScanOut({\ScanLink253[31] , \ScanLink253[30] , 
        \ScanLink253[29] , \ScanLink253[28] , \ScanLink253[27] , 
        \ScanLink253[26] , \ScanLink253[25] , \ScanLink253[24] , 
        \ScanLink253[23] , \ScanLink253[22] , \ScanLink253[21] , 
        \ScanLink253[20] , \ScanLink253[19] , \ScanLink253[18] , 
        \ScanLink253[17] , \ScanLink253[16] , \ScanLink253[15] , 
        \ScanLink253[14] , \ScanLink253[13] , \ScanLink253[12] , 
        \ScanLink253[11] , \ScanLink253[10] , \ScanLink253[9] , 
        \ScanLink253[8] , \ScanLink253[7] , \ScanLink253[6] , \ScanLink253[5] , 
        \ScanLink253[4] , \ScanLink253[3] , \ScanLink253[2] , \ScanLink253[1] , 
        \ScanLink253[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load252[0] ), .Out({\Level1Out252[31] , \Level1Out252[30] , 
        \Level1Out252[29] , \Level1Out252[28] , \Level1Out252[27] , 
        \Level1Out252[26] , \Level1Out252[25] , \Level1Out252[24] , 
        \Level1Out252[23] , \Level1Out252[22] , \Level1Out252[21] , 
        \Level1Out252[20] , \Level1Out252[19] , \Level1Out252[18] , 
        \Level1Out252[17] , \Level1Out252[16] , \Level1Out252[15] , 
        \Level1Out252[14] , \Level1Out252[13] , \Level1Out252[12] , 
        \Level1Out252[11] , \Level1Out252[10] , \Level1Out252[9] , 
        \Level1Out252[8] , \Level1Out252[7] , \Level1Out252[6] , 
        \Level1Out252[5] , \Level1Out252[4] , \Level1Out252[3] , 
        \Level1Out252[2] , \Level1Out252[1] , \Level1Out252[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load8[0] ), .Out({\Level2Out8[31] , \Level2Out8[30] , 
        \Level2Out8[29] , \Level2Out8[28] , \Level2Out8[27] , \Level2Out8[26] , 
        \Level2Out8[25] , \Level2Out8[24] , \Level2Out8[23] , \Level2Out8[22] , 
        \Level2Out8[21] , \Level2Out8[20] , \Level2Out8[19] , \Level2Out8[18] , 
        \Level2Out8[17] , \Level2Out8[16] , \Level2Out8[15] , \Level2Out8[14] , 
        \Level2Out8[13] , \Level2Out8[12] , \Level2Out8[11] , \Level2Out8[10] , 
        \Level2Out8[9] , \Level2Out8[8] , \Level2Out8[7] , \Level2Out8[6] , 
        \Level2Out8[5] , \Level2Out8[4] , \Level2Out8[3] , \Level2Out8[2] , 
        \Level2Out8[1] , \Level2Out8[0] }), .In1({\Level1Out8[31] , 
        \Level1Out8[30] , \Level1Out8[29] , \Level1Out8[28] , \Level1Out8[27] , 
        \Level1Out8[26] , \Level1Out8[25] , \Level1Out8[24] , \Level1Out8[23] , 
        \Level1Out8[22] , \Level1Out8[21] , \Level1Out8[20] , \Level1Out8[19] , 
        \Level1Out8[18] , \Level1Out8[17] , \Level1Out8[16] , \Level1Out8[15] , 
        \Level1Out8[14] , \Level1Out8[13] , \Level1Out8[12] , \Level1Out8[11] , 
        \Level1Out8[10] , \Level1Out8[9] , \Level1Out8[8] , \Level1Out8[7] , 
        \Level1Out8[6] , \Level1Out8[5] , \Level1Out8[4] , \Level1Out8[3] , 
        \Level1Out8[2] , \Level1Out8[1] , \Level1Out8[0] }), .In2({
        \Level1Out9[31] , \Level1Out9[30] , \Level1Out9[29] , \Level1Out9[28] , 
        \Level1Out9[27] , \Level1Out9[26] , \Level1Out9[25] , \Level1Out9[24] , 
        \Level1Out9[23] , \Level1Out9[22] , \Level1Out9[21] , \Level1Out9[20] , 
        \Level1Out9[19] , \Level1Out9[18] , \Level1Out9[17] , \Level1Out9[16] , 
        \Level1Out9[15] , \Level1Out9[14] , \Level1Out9[13] , \Level1Out9[12] , 
        \Level1Out9[11] , \Level1Out9[10] , \Level1Out9[9] , \Level1Out9[8] , 
        \Level1Out9[7] , \Level1Out9[6] , \Level1Out9[5] , \Level1Out9[4] , 
        \Level1Out9[3] , \Level1Out9[2] , \Level1Out9[1] , \Level1Out9[0] }), 
        .Read1(\Level1Load8[0] ), .Read2(\Level1Load9[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_180_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load180[0] ), .Out({\Level2Out180[31] , \Level2Out180[30] , 
        \Level2Out180[29] , \Level2Out180[28] , \Level2Out180[27] , 
        \Level2Out180[26] , \Level2Out180[25] , \Level2Out180[24] , 
        \Level2Out180[23] , \Level2Out180[22] , \Level2Out180[21] , 
        \Level2Out180[20] , \Level2Out180[19] , \Level2Out180[18] , 
        \Level2Out180[17] , \Level2Out180[16] , \Level2Out180[15] , 
        \Level2Out180[14] , \Level2Out180[13] , \Level2Out180[12] , 
        \Level2Out180[11] , \Level2Out180[10] , \Level2Out180[9] , 
        \Level2Out180[8] , \Level2Out180[7] , \Level2Out180[6] , 
        \Level2Out180[5] , \Level2Out180[4] , \Level2Out180[3] , 
        \Level2Out180[2] , \Level2Out180[1] , \Level2Out180[0] }), .In1({
        \Level1Out180[31] , \Level1Out180[30] , \Level1Out180[29] , 
        \Level1Out180[28] , \Level1Out180[27] , \Level1Out180[26] , 
        \Level1Out180[25] , \Level1Out180[24] , \Level1Out180[23] , 
        \Level1Out180[22] , \Level1Out180[21] , \Level1Out180[20] , 
        \Level1Out180[19] , \Level1Out180[18] , \Level1Out180[17] , 
        \Level1Out180[16] , \Level1Out180[15] , \Level1Out180[14] , 
        \Level1Out180[13] , \Level1Out180[12] , \Level1Out180[11] , 
        \Level1Out180[10] , \Level1Out180[9] , \Level1Out180[8] , 
        \Level1Out180[7] , \Level1Out180[6] , \Level1Out180[5] , 
        \Level1Out180[4] , \Level1Out180[3] , \Level1Out180[2] , 
        \Level1Out180[1] , \Level1Out180[0] }), .In2({\Level1Out181[31] , 
        \Level1Out181[30] , \Level1Out181[29] , \Level1Out181[28] , 
        \Level1Out181[27] , \Level1Out181[26] , \Level1Out181[25] , 
        \Level1Out181[24] , \Level1Out181[23] , \Level1Out181[22] , 
        \Level1Out181[21] , \Level1Out181[20] , \Level1Out181[19] , 
        \Level1Out181[18] , \Level1Out181[17] , \Level1Out181[16] , 
        \Level1Out181[15] , \Level1Out181[14] , \Level1Out181[13] , 
        \Level1Out181[12] , \Level1Out181[11] , \Level1Out181[10] , 
        \Level1Out181[9] , \Level1Out181[8] , \Level1Out181[7] , 
        \Level1Out181[6] , \Level1Out181[5] , \Level1Out181[4] , 
        \Level1Out181[3] , \Level1Out181[2] , \Level1Out181[1] , 
        \Level1Out181[0] }), .Read1(\Level1Load180[0] ), .Read2(
        \Level1Load181[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load64[0] ), .Out({\Level8Out64[31] , \Level8Out64[30] , 
        \Level8Out64[29] , \Level8Out64[28] , \Level8Out64[27] , 
        \Level8Out64[26] , \Level8Out64[25] , \Level8Out64[24] , 
        \Level8Out64[23] , \Level8Out64[22] , \Level8Out64[21] , 
        \Level8Out64[20] , \Level8Out64[19] , \Level8Out64[18] , 
        \Level8Out64[17] , \Level8Out64[16] , \Level8Out64[15] , 
        \Level8Out64[14] , \Level8Out64[13] , \Level8Out64[12] , 
        \Level8Out64[11] , \Level8Out64[10] , \Level8Out64[9] , 
        \Level8Out64[8] , \Level8Out64[7] , \Level8Out64[6] , \Level8Out64[5] , 
        \Level8Out64[4] , \Level8Out64[3] , \Level8Out64[2] , \Level8Out64[1] , 
        \Level8Out64[0] }), .In1({\Level4Out64[31] , \Level4Out64[30] , 
        \Level4Out64[29] , \Level4Out64[28] , \Level4Out64[27] , 
        \Level4Out64[26] , \Level4Out64[25] , \Level4Out64[24] , 
        \Level4Out64[23] , \Level4Out64[22] , \Level4Out64[21] , 
        \Level4Out64[20] , \Level4Out64[19] , \Level4Out64[18] , 
        \Level4Out64[17] , \Level4Out64[16] , \Level4Out64[15] , 
        \Level4Out64[14] , \Level4Out64[13] , \Level4Out64[12] , 
        \Level4Out64[11] , \Level4Out64[10] , \Level4Out64[9] , 
        \Level4Out64[8] , \Level4Out64[7] , \Level4Out64[6] , \Level4Out64[5] , 
        \Level4Out64[4] , \Level4Out64[3] , \Level4Out64[2] , \Level4Out64[1] , 
        \Level4Out64[0] }), .In2({\Level4Out68[31] , \Level4Out68[30] , 
        \Level4Out68[29] , \Level4Out68[28] , \Level4Out68[27] , 
        \Level4Out68[26] , \Level4Out68[25] , \Level4Out68[24] , 
        \Level4Out68[23] , \Level4Out68[22] , \Level4Out68[21] , 
        \Level4Out68[20] , \Level4Out68[19] , \Level4Out68[18] , 
        \Level4Out68[17] , \Level4Out68[16] , \Level4Out68[15] , 
        \Level4Out68[14] , \Level4Out68[13] , \Level4Out68[12] , 
        \Level4Out68[11] , \Level4Out68[10] , \Level4Out68[9] , 
        \Level4Out68[8] , \Level4Out68[7] , \Level4Out68[6] , \Level4Out68[5] , 
        \Level4Out68[4] , \Level4Out68[3] , \Level4Out68[2] , \Level4Out68[1] , 
        \Level4Out68[0] }), .Read1(\Level4Load64[0] ), .Read2(
        \Level4Load68[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_216_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load216[0] ), .Out({\Level8Out216[31] , \Level8Out216[30] , 
        \Level8Out216[29] , \Level8Out216[28] , \Level8Out216[27] , 
        \Level8Out216[26] , \Level8Out216[25] , \Level8Out216[24] , 
        \Level8Out216[23] , \Level8Out216[22] , \Level8Out216[21] , 
        \Level8Out216[20] , \Level8Out216[19] , \Level8Out216[18] , 
        \Level8Out216[17] , \Level8Out216[16] , \Level8Out216[15] , 
        \Level8Out216[14] , \Level8Out216[13] , \Level8Out216[12] , 
        \Level8Out216[11] , \Level8Out216[10] , \Level8Out216[9] , 
        \Level8Out216[8] , \Level8Out216[7] , \Level8Out216[6] , 
        \Level8Out216[5] , \Level8Out216[4] , \Level8Out216[3] , 
        \Level8Out216[2] , \Level8Out216[1] , \Level8Out216[0] }), .In1({
        \Level4Out216[31] , \Level4Out216[30] , \Level4Out216[29] , 
        \Level4Out216[28] , \Level4Out216[27] , \Level4Out216[26] , 
        \Level4Out216[25] , \Level4Out216[24] , \Level4Out216[23] , 
        \Level4Out216[22] , \Level4Out216[21] , \Level4Out216[20] , 
        \Level4Out216[19] , \Level4Out216[18] , \Level4Out216[17] , 
        \Level4Out216[16] , \Level4Out216[15] , \Level4Out216[14] , 
        \Level4Out216[13] , \Level4Out216[12] , \Level4Out216[11] , 
        \Level4Out216[10] , \Level4Out216[9] , \Level4Out216[8] , 
        \Level4Out216[7] , \Level4Out216[6] , \Level4Out216[5] , 
        \Level4Out216[4] , \Level4Out216[3] , \Level4Out216[2] , 
        \Level4Out216[1] , \Level4Out216[0] }), .In2({\Level4Out220[31] , 
        \Level4Out220[30] , \Level4Out220[29] , \Level4Out220[28] , 
        \Level4Out220[27] , \Level4Out220[26] , \Level4Out220[25] , 
        \Level4Out220[24] , \Level4Out220[23] , \Level4Out220[22] , 
        \Level4Out220[21] , \Level4Out220[20] , \Level4Out220[19] , 
        \Level4Out220[18] , \Level4Out220[17] , \Level4Out220[16] , 
        \Level4Out220[15] , \Level4Out220[14] , \Level4Out220[13] , 
        \Level4Out220[12] , \Level4Out220[11] , \Level4Out220[10] , 
        \Level4Out220[9] , \Level4Out220[8] , \Level4Out220[7] , 
        \Level4Out220[6] , \Level4Out220[5] , \Level4Out220[4] , 
        \Level4Out220[3] , \Level4Out220[2] , \Level4Out220[1] , 
        \Level4Out220[0] }), .Read1(\Level4Load216[0] ), .Read2(
        \Level4Load220[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_27 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanOut({\ScanLink28[31] , 
        \ScanLink28[30] , \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , 
        \ScanLink28[26] , \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , 
        \ScanLink28[22] , \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , 
        \ScanLink28[18] , \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , 
        \ScanLink28[14] , \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , 
        \ScanLink28[10] , \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , 
        \ScanLink28[6] , \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , 
        \ScanLink28[2] , \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load27[0] ), .Out({
        \Level1Out27[31] , \Level1Out27[30] , \Level1Out27[29] , 
        \Level1Out27[28] , \Level1Out27[27] , \Level1Out27[26] , 
        \Level1Out27[25] , \Level1Out27[24] , \Level1Out27[23] , 
        \Level1Out27[22] , \Level1Out27[21] , \Level1Out27[20] , 
        \Level1Out27[19] , \Level1Out27[18] , \Level1Out27[17] , 
        \Level1Out27[16] , \Level1Out27[15] , \Level1Out27[14] , 
        \Level1Out27[13] , \Level1Out27[12] , \Level1Out27[11] , 
        \Level1Out27[10] , \Level1Out27[9] , \Level1Out27[8] , 
        \Level1Out27[7] , \Level1Out27[6] , \Level1Out27[5] , \Level1Out27[4] , 
        \Level1Out27[3] , \Level1Out27[2] , \Level1Out27[1] , \Level1Out27[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_99 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink99[31] , \ScanLink99[30] , 
        \ScanLink99[29] , \ScanLink99[28] , \ScanLink99[27] , \ScanLink99[26] , 
        \ScanLink99[25] , \ScanLink99[24] , \ScanLink99[23] , \ScanLink99[22] , 
        \ScanLink99[21] , \ScanLink99[20] , \ScanLink99[19] , \ScanLink99[18] , 
        \ScanLink99[17] , \ScanLink99[16] , \ScanLink99[15] , \ScanLink99[14] , 
        \ScanLink99[13] , \ScanLink99[12] , \ScanLink99[11] , \ScanLink99[10] , 
        \ScanLink99[9] , \ScanLink99[8] , \ScanLink99[7] , \ScanLink99[6] , 
        \ScanLink99[5] , \ScanLink99[4] , \ScanLink99[3] , \ScanLink99[2] , 
        \ScanLink99[1] , \ScanLink99[0] }), .ScanOut({\ScanLink100[31] , 
        \ScanLink100[30] , \ScanLink100[29] , \ScanLink100[28] , 
        \ScanLink100[27] , \ScanLink100[26] , \ScanLink100[25] , 
        \ScanLink100[24] , \ScanLink100[23] , \ScanLink100[22] , 
        \ScanLink100[21] , \ScanLink100[20] , \ScanLink100[19] , 
        \ScanLink100[18] , \ScanLink100[17] , \ScanLink100[16] , 
        \ScanLink100[15] , \ScanLink100[14] , \ScanLink100[13] , 
        \ScanLink100[12] , \ScanLink100[11] , \ScanLink100[10] , 
        \ScanLink100[9] , \ScanLink100[8] , \ScanLink100[7] , \ScanLink100[6] , 
        \ScanLink100[5] , \ScanLink100[4] , \ScanLink100[3] , \ScanLink100[2] , 
        \ScanLink100[1] , \ScanLink100[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Id(1'b1), .Load(\Level1Load99[0] ), .Out({\Level1Out99[31] , 
        \Level1Out99[30] , \Level1Out99[29] , \Level1Out99[28] , 
        \Level1Out99[27] , \Level1Out99[26] , \Level1Out99[25] , 
        \Level1Out99[24] , \Level1Out99[23] , \Level1Out99[22] , 
        \Level1Out99[21] , \Level1Out99[20] , \Level1Out99[19] , 
        \Level1Out99[18] , \Level1Out99[17] , \Level1Out99[16] , 
        \Level1Out99[15] , \Level1Out99[14] , \Level1Out99[13] , 
        \Level1Out99[12] , \Level1Out99[11] , \Level1Out99[10] , 
        \Level1Out99[9] , \Level1Out99[8] , \Level1Out99[7] , \Level1Out99[6] , 
        \Level1Out99[5] , \Level1Out99[4] , \Level1Out99[3] , \Level1Out99[2] , 
        \Level1Out99[1] , \Level1Out99[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_130 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink130[31] , \ScanLink130[30] , 
        \ScanLink130[29] , \ScanLink130[28] , \ScanLink130[27] , 
        \ScanLink130[26] , \ScanLink130[25] , \ScanLink130[24] , 
        \ScanLink130[23] , \ScanLink130[22] , \ScanLink130[21] , 
        \ScanLink130[20] , \ScanLink130[19] , \ScanLink130[18] , 
        \ScanLink130[17] , \ScanLink130[16] , \ScanLink130[15] , 
        \ScanLink130[14] , \ScanLink130[13] , \ScanLink130[12] , 
        \ScanLink130[11] , \ScanLink130[10] , \ScanLink130[9] , 
        \ScanLink130[8] , \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , 
        \ScanLink130[4] , \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , 
        \ScanLink130[0] }), .ScanOut({\ScanLink131[31] , \ScanLink131[30] , 
        \ScanLink131[29] , \ScanLink131[28] , \ScanLink131[27] , 
        \ScanLink131[26] , \ScanLink131[25] , \ScanLink131[24] , 
        \ScanLink131[23] , \ScanLink131[22] , \ScanLink131[21] , 
        \ScanLink131[20] , \ScanLink131[19] , \ScanLink131[18] , 
        \ScanLink131[17] , \ScanLink131[16] , \ScanLink131[15] , 
        \ScanLink131[14] , \ScanLink131[13] , \ScanLink131[12] , 
        \ScanLink131[11] , \ScanLink131[10] , \ScanLink131[9] , 
        \ScanLink131[8] , \ScanLink131[7] , \ScanLink131[6] , \ScanLink131[5] , 
        \ScanLink131[4] , \ScanLink131[3] , \ScanLink131[2] , \ScanLink131[1] , 
        \ScanLink131[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load130[0] ), .Out({\Level1Out130[31] , \Level1Out130[30] , 
        \Level1Out130[29] , \Level1Out130[28] , \Level1Out130[27] , 
        \Level1Out130[26] , \Level1Out130[25] , \Level1Out130[24] , 
        \Level1Out130[23] , \Level1Out130[22] , \Level1Out130[21] , 
        \Level1Out130[20] , \Level1Out130[19] , \Level1Out130[18] , 
        \Level1Out130[17] , \Level1Out130[16] , \Level1Out130[15] , 
        \Level1Out130[14] , \Level1Out130[13] , \Level1Out130[12] , 
        \Level1Out130[11] , \Level1Out130[10] , \Level1Out130[9] , 
        \Level1Out130[8] , \Level1Out130[7] , \Level1Out130[6] , 
        \Level1Out130[5] , \Level1Out130[4] , \Level1Out130[3] , 
        \Level1Out130[2] , \Level1Out130[1] , \Level1Out130[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_200 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink200[31] , \ScanLink200[30] , 
        \ScanLink200[29] , \ScanLink200[28] , \ScanLink200[27] , 
        \ScanLink200[26] , \ScanLink200[25] , \ScanLink200[24] , 
        \ScanLink200[23] , \ScanLink200[22] , \ScanLink200[21] , 
        \ScanLink200[20] , \ScanLink200[19] , \ScanLink200[18] , 
        \ScanLink200[17] , \ScanLink200[16] , \ScanLink200[15] , 
        \ScanLink200[14] , \ScanLink200[13] , \ScanLink200[12] , 
        \ScanLink200[11] , \ScanLink200[10] , \ScanLink200[9] , 
        \ScanLink200[8] , \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , 
        \ScanLink200[4] , \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , 
        \ScanLink200[0] }), .ScanOut({\ScanLink201[31] , \ScanLink201[30] , 
        \ScanLink201[29] , \ScanLink201[28] , \ScanLink201[27] , 
        \ScanLink201[26] , \ScanLink201[25] , \ScanLink201[24] , 
        \ScanLink201[23] , \ScanLink201[22] , \ScanLink201[21] , 
        \ScanLink201[20] , \ScanLink201[19] , \ScanLink201[18] , 
        \ScanLink201[17] , \ScanLink201[16] , \ScanLink201[15] , 
        \ScanLink201[14] , \ScanLink201[13] , \ScanLink201[12] , 
        \ScanLink201[11] , \ScanLink201[10] , \ScanLink201[9] , 
        \ScanLink201[8] , \ScanLink201[7] , \ScanLink201[6] , \ScanLink201[5] , 
        \ScanLink201[4] , \ScanLink201[3] , \ScanLink201[2] , \ScanLink201[1] , 
        \ScanLink201[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load200[0] ), .Out({\Level1Out200[31] , \Level1Out200[30] , 
        \Level1Out200[29] , \Level1Out200[28] , \Level1Out200[27] , 
        \Level1Out200[26] , \Level1Out200[25] , \Level1Out200[24] , 
        \Level1Out200[23] , \Level1Out200[22] , \Level1Out200[21] , 
        \Level1Out200[20] , \Level1Out200[19] , \Level1Out200[18] , 
        \Level1Out200[17] , \Level1Out200[16] , \Level1Out200[15] , 
        \Level1Out200[14] , \Level1Out200[13] , \Level1Out200[12] , 
        \Level1Out200[11] , \Level1Out200[10] , \Level1Out200[9] , 
        \Level1Out200[8] , \Level1Out200[7] , \Level1Out200[6] , 
        \Level1Out200[5] , \Level1Out200[4] , \Level1Out200[3] , 
        \Level1Out200[2] , \Level1Out200[1] , \Level1Out200[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_116_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load116[0] ), .Out({\Level2Out116[31] , \Level2Out116[30] , 
        \Level2Out116[29] , \Level2Out116[28] , \Level2Out116[27] , 
        \Level2Out116[26] , \Level2Out116[25] , \Level2Out116[24] , 
        \Level2Out116[23] , \Level2Out116[22] , \Level2Out116[21] , 
        \Level2Out116[20] , \Level2Out116[19] , \Level2Out116[18] , 
        \Level2Out116[17] , \Level2Out116[16] , \Level2Out116[15] , 
        \Level2Out116[14] , \Level2Out116[13] , \Level2Out116[12] , 
        \Level2Out116[11] , \Level2Out116[10] , \Level2Out116[9] , 
        \Level2Out116[8] , \Level2Out116[7] , \Level2Out116[6] , 
        \Level2Out116[5] , \Level2Out116[4] , \Level2Out116[3] , 
        \Level2Out116[2] , \Level2Out116[1] , \Level2Out116[0] }), .In1({
        \Level1Out116[31] , \Level1Out116[30] , \Level1Out116[29] , 
        \Level1Out116[28] , \Level1Out116[27] , \Level1Out116[26] , 
        \Level1Out116[25] , \Level1Out116[24] , \Level1Out116[23] , 
        \Level1Out116[22] , \Level1Out116[21] , \Level1Out116[20] , 
        \Level1Out116[19] , \Level1Out116[18] , \Level1Out116[17] , 
        \Level1Out116[16] , \Level1Out116[15] , \Level1Out116[14] , 
        \Level1Out116[13] , \Level1Out116[12] , \Level1Out116[11] , 
        \Level1Out116[10] , \Level1Out116[9] , \Level1Out116[8] , 
        \Level1Out116[7] , \Level1Out116[6] , \Level1Out116[5] , 
        \Level1Out116[4] , \Level1Out116[3] , \Level1Out116[2] , 
        \Level1Out116[1] , \Level1Out116[0] }), .In2({\Level1Out117[31] , 
        \Level1Out117[30] , \Level1Out117[29] , \Level1Out117[28] , 
        \Level1Out117[27] , \Level1Out117[26] , \Level1Out117[25] , 
        \Level1Out117[24] , \Level1Out117[23] , \Level1Out117[22] , 
        \Level1Out117[21] , \Level1Out117[20] , \Level1Out117[19] , 
        \Level1Out117[18] , \Level1Out117[17] , \Level1Out117[16] , 
        \Level1Out117[15] , \Level1Out117[14] , \Level1Out117[13] , 
        \Level1Out117[12] , \Level1Out117[11] , \Level1Out117[10] , 
        \Level1Out117[9] , \Level1Out117[8] , \Level1Out117[7] , 
        \Level1Out117[6] , \Level1Out117[5] , \Level1Out117[4] , 
        \Level1Out117[3] , \Level1Out117[2] , \Level1Out117[1] , 
        \Level1Out117[0] }), .Read1(\Level1Load116[0] ), .Read2(
        \Level1Load117[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_208_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load208[0] ), .Out({\Level2Out208[31] , \Level2Out208[30] , 
        \Level2Out208[29] , \Level2Out208[28] , \Level2Out208[27] , 
        \Level2Out208[26] , \Level2Out208[25] , \Level2Out208[24] , 
        \Level2Out208[23] , \Level2Out208[22] , \Level2Out208[21] , 
        \Level2Out208[20] , \Level2Out208[19] , \Level2Out208[18] , 
        \Level2Out208[17] , \Level2Out208[16] , \Level2Out208[15] , 
        \Level2Out208[14] , \Level2Out208[13] , \Level2Out208[12] , 
        \Level2Out208[11] , \Level2Out208[10] , \Level2Out208[9] , 
        \Level2Out208[8] , \Level2Out208[7] , \Level2Out208[6] , 
        \Level2Out208[5] , \Level2Out208[4] , \Level2Out208[3] , 
        \Level2Out208[2] , \Level2Out208[1] , \Level2Out208[0] }), .In1({
        \Level1Out208[31] , \Level1Out208[30] , \Level1Out208[29] , 
        \Level1Out208[28] , \Level1Out208[27] , \Level1Out208[26] , 
        \Level1Out208[25] , \Level1Out208[24] , \Level1Out208[23] , 
        \Level1Out208[22] , \Level1Out208[21] , \Level1Out208[20] , 
        \Level1Out208[19] , \Level1Out208[18] , \Level1Out208[17] , 
        \Level1Out208[16] , \Level1Out208[15] , \Level1Out208[14] , 
        \Level1Out208[13] , \Level1Out208[12] , \Level1Out208[11] , 
        \Level1Out208[10] , \Level1Out208[9] , \Level1Out208[8] , 
        \Level1Out208[7] , \Level1Out208[6] , \Level1Out208[5] , 
        \Level1Out208[4] , \Level1Out208[3] , \Level1Out208[2] , 
        \Level1Out208[1] , \Level1Out208[0] }), .In2({\Level1Out209[31] , 
        \Level1Out209[30] , \Level1Out209[29] , \Level1Out209[28] , 
        \Level1Out209[27] , \Level1Out209[26] , \Level1Out209[25] , 
        \Level1Out209[24] , \Level1Out209[23] , \Level1Out209[22] , 
        \Level1Out209[21] , \Level1Out209[20] , \Level1Out209[19] , 
        \Level1Out209[18] , \Level1Out209[17] , \Level1Out209[16] , 
        \Level1Out209[15] , \Level1Out209[14] , \Level1Out209[13] , 
        \Level1Out209[12] , \Level1Out209[11] , \Level1Out209[10] , 
        \Level1Out209[9] , \Level1Out209[8] , \Level1Out209[7] , 
        \Level1Out209[6] , \Level1Out209[5] , \Level1Out209[4] , 
        \Level1Out209[3] , \Level1Out209[2] , \Level1Out209[1] , 
        \Level1Out209[0] }), .Read1(\Level1Load208[0] ), .Read2(
        \Level1Load209[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_227 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink227[31] , \ScanLink227[30] , 
        \ScanLink227[29] , \ScanLink227[28] , \ScanLink227[27] , 
        \ScanLink227[26] , \ScanLink227[25] , \ScanLink227[24] , 
        \ScanLink227[23] , \ScanLink227[22] , \ScanLink227[21] , 
        \ScanLink227[20] , \ScanLink227[19] , \ScanLink227[18] , 
        \ScanLink227[17] , \ScanLink227[16] , \ScanLink227[15] , 
        \ScanLink227[14] , \ScanLink227[13] , \ScanLink227[12] , 
        \ScanLink227[11] , \ScanLink227[10] , \ScanLink227[9] , 
        \ScanLink227[8] , \ScanLink227[7] , \ScanLink227[6] , \ScanLink227[5] , 
        \ScanLink227[4] , \ScanLink227[3] , \ScanLink227[2] , \ScanLink227[1] , 
        \ScanLink227[0] }), .ScanOut({\ScanLink228[31] , \ScanLink228[30] , 
        \ScanLink228[29] , \ScanLink228[28] , \ScanLink228[27] , 
        \ScanLink228[26] , \ScanLink228[25] , \ScanLink228[24] , 
        \ScanLink228[23] , \ScanLink228[22] , \ScanLink228[21] , 
        \ScanLink228[20] , \ScanLink228[19] , \ScanLink228[18] , 
        \ScanLink228[17] , \ScanLink228[16] , \ScanLink228[15] , 
        \ScanLink228[14] , \ScanLink228[13] , \ScanLink228[12] , 
        \ScanLink228[11] , \ScanLink228[10] , \ScanLink228[9] , 
        \ScanLink228[8] , \ScanLink228[7] , \ScanLink228[6] , \ScanLink228[5] , 
        \ScanLink228[4] , \ScanLink228[3] , \ScanLink228[2] , \ScanLink228[1] , 
        \ScanLink228[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load227[0] ), .Out({\Level1Out227[31] , \Level1Out227[30] , 
        \Level1Out227[29] , \Level1Out227[28] , \Level1Out227[27] , 
        \Level1Out227[26] , \Level1Out227[25] , \Level1Out227[24] , 
        \Level1Out227[23] , \Level1Out227[22] , \Level1Out227[21] , 
        \Level1Out227[20] , \Level1Out227[19] , \Level1Out227[18] , 
        \Level1Out227[17] , \Level1Out227[16] , \Level1Out227[15] , 
        \Level1Out227[14] , \Level1Out227[13] , \Level1Out227[12] , 
        \Level1Out227[11] , \Level1Out227[10] , \Level1Out227[9] , 
        \Level1Out227[8] , \Level1Out227[7] , \Level1Out227[6] , 
        \Level1Out227[5] , \Level1Out227[4] , \Level1Out227[3] , 
        \Level1Out227[2] , \Level1Out227[1] , \Level1Out227[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_50_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load50[0] ), .Out({\Level2Out50[31] , \Level2Out50[30] , 
        \Level2Out50[29] , \Level2Out50[28] , \Level2Out50[27] , 
        \Level2Out50[26] , \Level2Out50[25] , \Level2Out50[24] , 
        \Level2Out50[23] , \Level2Out50[22] , \Level2Out50[21] , 
        \Level2Out50[20] , \Level2Out50[19] , \Level2Out50[18] , 
        \Level2Out50[17] , \Level2Out50[16] , \Level2Out50[15] , 
        \Level2Out50[14] , \Level2Out50[13] , \Level2Out50[12] , 
        \Level2Out50[11] , \Level2Out50[10] , \Level2Out50[9] , 
        \Level2Out50[8] , \Level2Out50[7] , \Level2Out50[6] , \Level2Out50[5] , 
        \Level2Out50[4] , \Level2Out50[3] , \Level2Out50[2] , \Level2Out50[1] , 
        \Level2Out50[0] }), .In1({\Level1Out50[31] , \Level1Out50[30] , 
        \Level1Out50[29] , \Level1Out50[28] , \Level1Out50[27] , 
        \Level1Out50[26] , \Level1Out50[25] , \Level1Out50[24] , 
        \Level1Out50[23] , \Level1Out50[22] , \Level1Out50[21] , 
        \Level1Out50[20] , \Level1Out50[19] , \Level1Out50[18] , 
        \Level1Out50[17] , \Level1Out50[16] , \Level1Out50[15] , 
        \Level1Out50[14] , \Level1Out50[13] , \Level1Out50[12] , 
        \Level1Out50[11] , \Level1Out50[10] , \Level1Out50[9] , 
        \Level1Out50[8] , \Level1Out50[7] , \Level1Out50[6] , \Level1Out50[5] , 
        \Level1Out50[4] , \Level1Out50[3] , \Level1Out50[2] , \Level1Out50[1] , 
        \Level1Out50[0] }), .In2({\Level1Out51[31] , \Level1Out51[30] , 
        \Level1Out51[29] , \Level1Out51[28] , \Level1Out51[27] , 
        \Level1Out51[26] , \Level1Out51[25] , \Level1Out51[24] , 
        \Level1Out51[23] , \Level1Out51[22] , \Level1Out51[21] , 
        \Level1Out51[20] , \Level1Out51[19] , \Level1Out51[18] , 
        \Level1Out51[17] , \Level1Out51[16] , \Level1Out51[15] , 
        \Level1Out51[14] , \Level1Out51[13] , \Level1Out51[12] , 
        \Level1Out51[11] , \Level1Out51[10] , \Level1Out51[9] , 
        \Level1Out51[8] , \Level1Out51[7] , \Level1Out51[6] , \Level1Out51[5] , 
        \Level1Out51[4] , \Level1Out51[3] , \Level1Out51[2] , \Level1Out51[1] , 
        \Level1Out51[0] }), .Read1(\Level1Load50[0] ), .Read2(
        \Level1Load51[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_222_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load222[0] ), .Out({\Level2Out222[31] , \Level2Out222[30] , 
        \Level2Out222[29] , \Level2Out222[28] , \Level2Out222[27] , 
        \Level2Out222[26] , \Level2Out222[25] , \Level2Out222[24] , 
        \Level2Out222[23] , \Level2Out222[22] , \Level2Out222[21] , 
        \Level2Out222[20] , \Level2Out222[19] , \Level2Out222[18] , 
        \Level2Out222[17] , \Level2Out222[16] , \Level2Out222[15] , 
        \Level2Out222[14] , \Level2Out222[13] , \Level2Out222[12] , 
        \Level2Out222[11] , \Level2Out222[10] , \Level2Out222[9] , 
        \Level2Out222[8] , \Level2Out222[7] , \Level2Out222[6] , 
        \Level2Out222[5] , \Level2Out222[4] , \Level2Out222[3] , 
        \Level2Out222[2] , \Level2Out222[1] , \Level2Out222[0] }), .In1({
        \Level1Out222[31] , \Level1Out222[30] , \Level1Out222[29] , 
        \Level1Out222[28] , \Level1Out222[27] , \Level1Out222[26] , 
        \Level1Out222[25] , \Level1Out222[24] , \Level1Out222[23] , 
        \Level1Out222[22] , \Level1Out222[21] , \Level1Out222[20] , 
        \Level1Out222[19] , \Level1Out222[18] , \Level1Out222[17] , 
        \Level1Out222[16] , \Level1Out222[15] , \Level1Out222[14] , 
        \Level1Out222[13] , \Level1Out222[12] , \Level1Out222[11] , 
        \Level1Out222[10] , \Level1Out222[9] , \Level1Out222[8] , 
        \Level1Out222[7] , \Level1Out222[6] , \Level1Out222[5] , 
        \Level1Out222[4] , \Level1Out222[3] , \Level1Out222[2] , 
        \Level1Out222[1] , \Level1Out222[0] }), .In2({\Level1Out223[31] , 
        \Level1Out223[30] , \Level1Out223[29] , \Level1Out223[28] , 
        \Level1Out223[27] , \Level1Out223[26] , \Level1Out223[25] , 
        \Level1Out223[24] , \Level1Out223[23] , \Level1Out223[22] , 
        \Level1Out223[21] , \Level1Out223[20] , \Level1Out223[19] , 
        \Level1Out223[18] , \Level1Out223[17] , \Level1Out223[16] , 
        \Level1Out223[15] , \Level1Out223[14] , \Level1Out223[13] , 
        \Level1Out223[12] , \Level1Out223[11] , \Level1Out223[10] , 
        \Level1Out223[9] , \Level1Out223[8] , \Level1Out223[7] , 
        \Level1Out223[6] , \Level1Out223[5] , \Level1Out223[4] , 
        \Level1Out223[3] , \Level1Out223[2] , \Level1Out223[1] , 
        \Level1Out223[0] }), .Read1(\Level1Load222[0] ), .Read2(
        \Level1Load223[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_105 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink105[31] , \ScanLink105[30] , 
        \ScanLink105[29] , \ScanLink105[28] , \ScanLink105[27] , 
        \ScanLink105[26] , \ScanLink105[25] , \ScanLink105[24] , 
        \ScanLink105[23] , \ScanLink105[22] , \ScanLink105[21] , 
        \ScanLink105[20] , \ScanLink105[19] , \ScanLink105[18] , 
        \ScanLink105[17] , \ScanLink105[16] , \ScanLink105[15] , 
        \ScanLink105[14] , \ScanLink105[13] , \ScanLink105[12] , 
        \ScanLink105[11] , \ScanLink105[10] , \ScanLink105[9] , 
        \ScanLink105[8] , \ScanLink105[7] , \ScanLink105[6] , \ScanLink105[5] , 
        \ScanLink105[4] , \ScanLink105[3] , \ScanLink105[2] , \ScanLink105[1] , 
        \ScanLink105[0] }), .ScanOut({\ScanLink106[31] , \ScanLink106[30] , 
        \ScanLink106[29] , \ScanLink106[28] , \ScanLink106[27] , 
        \ScanLink106[26] , \ScanLink106[25] , \ScanLink106[24] , 
        \ScanLink106[23] , \ScanLink106[22] , \ScanLink106[21] , 
        \ScanLink106[20] , \ScanLink106[19] , \ScanLink106[18] , 
        \ScanLink106[17] , \ScanLink106[16] , \ScanLink106[15] , 
        \ScanLink106[14] , \ScanLink106[13] , \ScanLink106[12] , 
        \ScanLink106[11] , \ScanLink106[10] , \ScanLink106[9] , 
        \ScanLink106[8] , \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , 
        \ScanLink106[4] , \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , 
        \ScanLink106[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load105[0] ), .Out({\Level1Out105[31] , \Level1Out105[30] , 
        \Level1Out105[29] , \Level1Out105[28] , \Level1Out105[27] , 
        \Level1Out105[26] , \Level1Out105[25] , \Level1Out105[24] , 
        \Level1Out105[23] , \Level1Out105[22] , \Level1Out105[21] , 
        \Level1Out105[20] , \Level1Out105[19] , \Level1Out105[18] , 
        \Level1Out105[17] , \Level1Out105[16] , \Level1Out105[15] , 
        \Level1Out105[14] , \Level1Out105[13] , \Level1Out105[12] , 
        \Level1Out105[11] , \Level1Out105[10] , \Level1Out105[9] , 
        \Level1Out105[8] , \Level1Out105[7] , \Level1Out105[6] , 
        \Level1Out105[5] , \Level1Out105[4] , \Level1Out105[3] , 
        \Level1Out105[2] , \Level1Out105[1] , \Level1Out105[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_117 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink117[31] , \ScanLink117[30] , 
        \ScanLink117[29] , \ScanLink117[28] , \ScanLink117[27] , 
        \ScanLink117[26] , \ScanLink117[25] , \ScanLink117[24] , 
        \ScanLink117[23] , \ScanLink117[22] , \ScanLink117[21] , 
        \ScanLink117[20] , \ScanLink117[19] , \ScanLink117[18] , 
        \ScanLink117[17] , \ScanLink117[16] , \ScanLink117[15] , 
        \ScanLink117[14] , \ScanLink117[13] , \ScanLink117[12] , 
        \ScanLink117[11] , \ScanLink117[10] , \ScanLink117[9] , 
        \ScanLink117[8] , \ScanLink117[7] , \ScanLink117[6] , \ScanLink117[5] , 
        \ScanLink117[4] , \ScanLink117[3] , \ScanLink117[2] , \ScanLink117[1] , 
        \ScanLink117[0] }), .ScanOut({\ScanLink118[31] , \ScanLink118[30] , 
        \ScanLink118[29] , \ScanLink118[28] , \ScanLink118[27] , 
        \ScanLink118[26] , \ScanLink118[25] , \ScanLink118[24] , 
        \ScanLink118[23] , \ScanLink118[22] , \ScanLink118[21] , 
        \ScanLink118[20] , \ScanLink118[19] , \ScanLink118[18] , 
        \ScanLink118[17] , \ScanLink118[16] , \ScanLink118[15] , 
        \ScanLink118[14] , \ScanLink118[13] , \ScanLink118[12] , 
        \ScanLink118[11] , \ScanLink118[10] , \ScanLink118[9] , 
        \ScanLink118[8] , \ScanLink118[7] , \ScanLink118[6] , \ScanLink118[5] , 
        \ScanLink118[4] , \ScanLink118[3] , \ScanLink118[2] , \ScanLink118[1] , 
        \ScanLink118[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load117[0] ), .Out({\Level1Out117[31] , \Level1Out117[30] , 
        \Level1Out117[29] , \Level1Out117[28] , \Level1Out117[27] , 
        \Level1Out117[26] , \Level1Out117[25] , \Level1Out117[24] , 
        \Level1Out117[23] , \Level1Out117[22] , \Level1Out117[21] , 
        \Level1Out117[20] , \Level1Out117[19] , \Level1Out117[18] , 
        \Level1Out117[17] , \Level1Out117[16] , \Level1Out117[15] , 
        \Level1Out117[14] , \Level1Out117[13] , \Level1Out117[12] , 
        \Level1Out117[11] , \Level1Out117[10] , \Level1Out117[9] , 
        \Level1Out117[8] , \Level1Out117[7] , \Level1Out117[6] , 
        \Level1Out117[5] , \Level1Out117[4] , \Level1Out117[3] , 
        \Level1Out117[2] , \Level1Out117[1] , \Level1Out117[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_122 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink122[31] , \ScanLink122[30] , 
        \ScanLink122[29] , \ScanLink122[28] , \ScanLink122[27] , 
        \ScanLink122[26] , \ScanLink122[25] , \ScanLink122[24] , 
        \ScanLink122[23] , \ScanLink122[22] , \ScanLink122[21] , 
        \ScanLink122[20] , \ScanLink122[19] , \ScanLink122[18] , 
        \ScanLink122[17] , \ScanLink122[16] , \ScanLink122[15] , 
        \ScanLink122[14] , \ScanLink122[13] , \ScanLink122[12] , 
        \ScanLink122[11] , \ScanLink122[10] , \ScanLink122[9] , 
        \ScanLink122[8] , \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , 
        \ScanLink122[4] , \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , 
        \ScanLink122[0] }), .ScanOut({\ScanLink123[31] , \ScanLink123[30] , 
        \ScanLink123[29] , \ScanLink123[28] , \ScanLink123[27] , 
        \ScanLink123[26] , \ScanLink123[25] , \ScanLink123[24] , 
        \ScanLink123[23] , \ScanLink123[22] , \ScanLink123[21] , 
        \ScanLink123[20] , \ScanLink123[19] , \ScanLink123[18] , 
        \ScanLink123[17] , \ScanLink123[16] , \ScanLink123[15] , 
        \ScanLink123[14] , \ScanLink123[13] , \ScanLink123[12] , 
        \ScanLink123[11] , \ScanLink123[10] , \ScanLink123[9] , 
        \ScanLink123[8] , \ScanLink123[7] , \ScanLink123[6] , \ScanLink123[5] , 
        \ScanLink123[4] , \ScanLink123[3] , \ScanLink123[2] , \ScanLink123[1] , 
        \ScanLink123[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load122[0] ), .Out({\Level1Out122[31] , \Level1Out122[30] , 
        \Level1Out122[29] , \Level1Out122[28] , \Level1Out122[27] , 
        \Level1Out122[26] , \Level1Out122[25] , \Level1Out122[24] , 
        \Level1Out122[23] , \Level1Out122[22] , \Level1Out122[21] , 
        \Level1Out122[20] , \Level1Out122[19] , \Level1Out122[18] , 
        \Level1Out122[17] , \Level1Out122[16] , \Level1Out122[15] , 
        \Level1Out122[14] , \Level1Out122[13] , \Level1Out122[12] , 
        \Level1Out122[11] , \Level1Out122[10] , \Level1Out122[9] , 
        \Level1Out122[8] , \Level1Out122[7] , \Level1Out122[6] , 
        \Level1Out122[5] , \Level1Out122[4] , \Level1Out122[3] , 
        \Level1Out122[2] , \Level1Out122[1] , \Level1Out122[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_120_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load120[0] ), .Out({\Level4Out120[31] , \Level4Out120[30] , 
        \Level4Out120[29] , \Level4Out120[28] , \Level4Out120[27] , 
        \Level4Out120[26] , \Level4Out120[25] , \Level4Out120[24] , 
        \Level4Out120[23] , \Level4Out120[22] , \Level4Out120[21] , 
        \Level4Out120[20] , \Level4Out120[19] , \Level4Out120[18] , 
        \Level4Out120[17] , \Level4Out120[16] , \Level4Out120[15] , 
        \Level4Out120[14] , \Level4Out120[13] , \Level4Out120[12] , 
        \Level4Out120[11] , \Level4Out120[10] , \Level4Out120[9] , 
        \Level4Out120[8] , \Level4Out120[7] , \Level4Out120[6] , 
        \Level4Out120[5] , \Level4Out120[4] , \Level4Out120[3] , 
        \Level4Out120[2] , \Level4Out120[1] , \Level4Out120[0] }), .In1({
        \Level2Out120[31] , \Level2Out120[30] , \Level2Out120[29] , 
        \Level2Out120[28] , \Level2Out120[27] , \Level2Out120[26] , 
        \Level2Out120[25] , \Level2Out120[24] , \Level2Out120[23] , 
        \Level2Out120[22] , \Level2Out120[21] , \Level2Out120[20] , 
        \Level2Out120[19] , \Level2Out120[18] , \Level2Out120[17] , 
        \Level2Out120[16] , \Level2Out120[15] , \Level2Out120[14] , 
        \Level2Out120[13] , \Level2Out120[12] , \Level2Out120[11] , 
        \Level2Out120[10] , \Level2Out120[9] , \Level2Out120[8] , 
        \Level2Out120[7] , \Level2Out120[6] , \Level2Out120[5] , 
        \Level2Out120[4] , \Level2Out120[3] , \Level2Out120[2] , 
        \Level2Out120[1] , \Level2Out120[0] }), .In2({\Level2Out122[31] , 
        \Level2Out122[30] , \Level2Out122[29] , \Level2Out122[28] , 
        \Level2Out122[27] , \Level2Out122[26] , \Level2Out122[25] , 
        \Level2Out122[24] , \Level2Out122[23] , \Level2Out122[22] , 
        \Level2Out122[21] , \Level2Out122[20] , \Level2Out122[19] , 
        \Level2Out122[18] , \Level2Out122[17] , \Level2Out122[16] , 
        \Level2Out122[15] , \Level2Out122[14] , \Level2Out122[13] , 
        \Level2Out122[12] , \Level2Out122[11] , \Level2Out122[10] , 
        \Level2Out122[9] , \Level2Out122[8] , \Level2Out122[7] , 
        \Level2Out122[6] , \Level2Out122[5] , \Level2Out122[4] , 
        \Level2Out122[3] , \Level2Out122[2] , \Level2Out122[1] , 
        \Level2Out122[0] }), .Read1(\Level2Load120[0] ), .Read2(
        \Level2Load122[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_212 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink212[31] , \ScanLink212[30] , 
        \ScanLink212[29] , \ScanLink212[28] , \ScanLink212[27] , 
        \ScanLink212[26] , \ScanLink212[25] , \ScanLink212[24] , 
        \ScanLink212[23] , \ScanLink212[22] , \ScanLink212[21] , 
        \ScanLink212[20] , \ScanLink212[19] , \ScanLink212[18] , 
        \ScanLink212[17] , \ScanLink212[16] , \ScanLink212[15] , 
        \ScanLink212[14] , \ScanLink212[13] , \ScanLink212[12] , 
        \ScanLink212[11] , \ScanLink212[10] , \ScanLink212[9] , 
        \ScanLink212[8] , \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , 
        \ScanLink212[4] , \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , 
        \ScanLink212[0] }), .ScanOut({\ScanLink213[31] , \ScanLink213[30] , 
        \ScanLink213[29] , \ScanLink213[28] , \ScanLink213[27] , 
        \ScanLink213[26] , \ScanLink213[25] , \ScanLink213[24] , 
        \ScanLink213[23] , \ScanLink213[22] , \ScanLink213[21] , 
        \ScanLink213[20] , \ScanLink213[19] , \ScanLink213[18] , 
        \ScanLink213[17] , \ScanLink213[16] , \ScanLink213[15] , 
        \ScanLink213[14] , \ScanLink213[13] , \ScanLink213[12] , 
        \ScanLink213[11] , \ScanLink213[10] , \ScanLink213[9] , 
        \ScanLink213[8] , \ScanLink213[7] , \ScanLink213[6] , \ScanLink213[5] , 
        \ScanLink213[4] , \ScanLink213[3] , \ScanLink213[2] , \ScanLink213[1] , 
        \ScanLink213[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load212[0] ), .Out({\Level1Out212[31] , \Level1Out212[30] , 
        \Level1Out212[29] , \Level1Out212[28] , \Level1Out212[27] , 
        \Level1Out212[26] , \Level1Out212[25] , \Level1Out212[24] , 
        \Level1Out212[23] , \Level1Out212[22] , \Level1Out212[21] , 
        \Level1Out212[20] , \Level1Out212[19] , \Level1Out212[18] , 
        \Level1Out212[17] , \Level1Out212[16] , \Level1Out212[15] , 
        \Level1Out212[14] , \Level1Out212[13] , \Level1Out212[12] , 
        \Level1Out212[11] , \Level1Out212[10] , \Level1Out212[9] , 
        \Level1Out212[8] , \Level1Out212[7] , \Level1Out212[6] , 
        \Level1Out212[5] , \Level1Out212[4] , \Level1Out212[3] , 
        \Level1Out212[2] , \Level1Out212[1] , \Level1Out212[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_235 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink235[31] , \ScanLink235[30] , 
        \ScanLink235[29] , \ScanLink235[28] , \ScanLink235[27] , 
        \ScanLink235[26] , \ScanLink235[25] , \ScanLink235[24] , 
        \ScanLink235[23] , \ScanLink235[22] , \ScanLink235[21] , 
        \ScanLink235[20] , \ScanLink235[19] , \ScanLink235[18] , 
        \ScanLink235[17] , \ScanLink235[16] , \ScanLink235[15] , 
        \ScanLink235[14] , \ScanLink235[13] , \ScanLink235[12] , 
        \ScanLink235[11] , \ScanLink235[10] , \ScanLink235[9] , 
        \ScanLink235[8] , \ScanLink235[7] , \ScanLink235[6] , \ScanLink235[5] , 
        \ScanLink235[4] , \ScanLink235[3] , \ScanLink235[2] , \ScanLink235[1] , 
        \ScanLink235[0] }), .ScanOut({\ScanLink236[31] , \ScanLink236[30] , 
        \ScanLink236[29] , \ScanLink236[28] , \ScanLink236[27] , 
        \ScanLink236[26] , \ScanLink236[25] , \ScanLink236[24] , 
        \ScanLink236[23] , \ScanLink236[22] , \ScanLink236[21] , 
        \ScanLink236[20] , \ScanLink236[19] , \ScanLink236[18] , 
        \ScanLink236[17] , \ScanLink236[16] , \ScanLink236[15] , 
        \ScanLink236[14] , \ScanLink236[13] , \ScanLink236[12] , 
        \ScanLink236[11] , \ScanLink236[10] , \ScanLink236[9] , 
        \ScanLink236[8] , \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , 
        \ScanLink236[4] , \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , 
        \ScanLink236[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load235[0] ), .Out({\Level1Out235[31] , \Level1Out235[30] , 
        \Level1Out235[29] , \Level1Out235[28] , \Level1Out235[27] , 
        \Level1Out235[26] , \Level1Out235[25] , \Level1Out235[24] , 
        \Level1Out235[23] , \Level1Out235[22] , \Level1Out235[21] , 
        \Level1Out235[20] , \Level1Out235[19] , \Level1Out235[18] , 
        \Level1Out235[17] , \Level1Out235[16] , \Level1Out235[15] , 
        \Level1Out235[14] , \Level1Out235[13] , \Level1Out235[12] , 
        \Level1Out235[11] , \Level1Out235[10] , \Level1Out235[9] , 
        \Level1Out235[8] , \Level1Out235[7] , \Level1Out235[6] , 
        \Level1Out235[5] , \Level1Out235[4] , \Level1Out235[3] , 
        \Level1Out235[2] , \Level1Out235[1] , \Level1Out235[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_49 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanOut({\ScanLink50[31] , 
        \ScanLink50[30] , \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , 
        \ScanLink50[26] , \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , 
        \ScanLink50[22] , \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , 
        \ScanLink50[18] , \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , 
        \ScanLink50[14] , \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , 
        \ScanLink50[10] , \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , 
        \ScanLink50[6] , \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , 
        \ScanLink50[2] , \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load49[0] ), .Out({
        \Level1Out49[31] , \Level1Out49[30] , \Level1Out49[29] , 
        \Level1Out49[28] , \Level1Out49[27] , \Level1Out49[26] , 
        \Level1Out49[25] , \Level1Out49[24] , \Level1Out49[23] , 
        \Level1Out49[22] , \Level1Out49[21] , \Level1Out49[20] , 
        \Level1Out49[19] , \Level1Out49[18] , \Level1Out49[17] , 
        \Level1Out49[16] , \Level1Out49[15] , \Level1Out49[14] , 
        \Level1Out49[13] , \Level1Out49[12] , \Level1Out49[11] , 
        \Level1Out49[10] , \Level1Out49[9] , \Level1Out49[8] , 
        \Level1Out49[7] , \Level1Out49[6] , \Level1Out49[5] , \Level1Out49[4] , 
        \Level1Out49[3] , \Level1Out49[2] , \Level1Out49[1] , \Level1Out49[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_36_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load36[0] ), .Out({\Level4Out36[31] , \Level4Out36[30] , 
        \Level4Out36[29] , \Level4Out36[28] , \Level4Out36[27] , 
        \Level4Out36[26] , \Level4Out36[25] , \Level4Out36[24] , 
        \Level4Out36[23] , \Level4Out36[22] , \Level4Out36[21] , 
        \Level4Out36[20] , \Level4Out36[19] , \Level4Out36[18] , 
        \Level4Out36[17] , \Level4Out36[16] , \Level4Out36[15] , 
        \Level4Out36[14] , \Level4Out36[13] , \Level4Out36[12] , 
        \Level4Out36[11] , \Level4Out36[10] , \Level4Out36[9] , 
        \Level4Out36[8] , \Level4Out36[7] , \Level4Out36[6] , \Level4Out36[5] , 
        \Level4Out36[4] , \Level4Out36[3] , \Level4Out36[2] , \Level4Out36[1] , 
        \Level4Out36[0] }), .In1({\Level2Out36[31] , \Level2Out36[30] , 
        \Level2Out36[29] , \Level2Out36[28] , \Level2Out36[27] , 
        \Level2Out36[26] , \Level2Out36[25] , \Level2Out36[24] , 
        \Level2Out36[23] , \Level2Out36[22] , \Level2Out36[21] , 
        \Level2Out36[20] , \Level2Out36[19] , \Level2Out36[18] , 
        \Level2Out36[17] , \Level2Out36[16] , \Level2Out36[15] , 
        \Level2Out36[14] , \Level2Out36[13] , \Level2Out36[12] , 
        \Level2Out36[11] , \Level2Out36[10] , \Level2Out36[9] , 
        \Level2Out36[8] , \Level2Out36[7] , \Level2Out36[6] , \Level2Out36[5] , 
        \Level2Out36[4] , \Level2Out36[3] , \Level2Out36[2] , \Level2Out36[1] , 
        \Level2Out36[0] }), .In2({\Level2Out38[31] , \Level2Out38[30] , 
        \Level2Out38[29] , \Level2Out38[28] , \Level2Out38[27] , 
        \Level2Out38[26] , \Level2Out38[25] , \Level2Out38[24] , 
        \Level2Out38[23] , \Level2Out38[22] , \Level2Out38[21] , 
        \Level2Out38[20] , \Level2Out38[19] , \Level2Out38[18] , 
        \Level2Out38[17] , \Level2Out38[16] , \Level2Out38[15] , 
        \Level2Out38[14] , \Level2Out38[13] , \Level2Out38[12] , 
        \Level2Out38[11] , \Level2Out38[10] , \Level2Out38[9] , 
        \Level2Out38[8] , \Level2Out38[7] , \Level2Out38[6] , \Level2Out38[5] , 
        \Level2Out38[4] , \Level2Out38[3] , \Level2Out38[2] , \Level2Out38[1] , 
        \Level2Out38[0] }), .Read1(\Level2Load36[0] ), .Read2(
        \Level2Load38[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_32 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load192[0] ), .Out({\Level32Out192[31] , \Level32Out192[30] , 
        \Level32Out192[29] , \Level32Out192[28] , \Level32Out192[27] , 
        \Level32Out192[26] , \Level32Out192[25] , \Level32Out192[24] , 
        \Level32Out192[23] , \Level32Out192[22] , \Level32Out192[21] , 
        \Level32Out192[20] , \Level32Out192[19] , \Level32Out192[18] , 
        \Level32Out192[17] , \Level32Out192[16] , \Level32Out192[15] , 
        \Level32Out192[14] , \Level32Out192[13] , \Level32Out192[12] , 
        \Level32Out192[11] , \Level32Out192[10] , \Level32Out192[9] , 
        \Level32Out192[8] , \Level32Out192[7] , \Level32Out192[6] , 
        \Level32Out192[5] , \Level32Out192[4] , \Level32Out192[3] , 
        \Level32Out192[2] , \Level32Out192[1] , \Level32Out192[0] }), .In1({
        \Level16Out192[31] , \Level16Out192[30] , \Level16Out192[29] , 
        \Level16Out192[28] , \Level16Out192[27] , \Level16Out192[26] , 
        \Level16Out192[25] , \Level16Out192[24] , \Level16Out192[23] , 
        \Level16Out192[22] , \Level16Out192[21] , \Level16Out192[20] , 
        \Level16Out192[19] , \Level16Out192[18] , \Level16Out192[17] , 
        \Level16Out192[16] , \Level16Out192[15] , \Level16Out192[14] , 
        \Level16Out192[13] , \Level16Out192[12] , \Level16Out192[11] , 
        \Level16Out192[10] , \Level16Out192[9] , \Level16Out192[8] , 
        \Level16Out192[7] , \Level16Out192[6] , \Level16Out192[5] , 
        \Level16Out192[4] , \Level16Out192[3] , \Level16Out192[2] , 
        \Level16Out192[1] , \Level16Out192[0] }), .In2({\Level16Out208[31] , 
        \Level16Out208[30] , \Level16Out208[29] , \Level16Out208[28] , 
        \Level16Out208[27] , \Level16Out208[26] , \Level16Out208[25] , 
        \Level16Out208[24] , \Level16Out208[23] , \Level16Out208[22] , 
        \Level16Out208[21] , \Level16Out208[20] , \Level16Out208[19] , 
        \Level16Out208[18] , \Level16Out208[17] , \Level16Out208[16] , 
        \Level16Out208[15] , \Level16Out208[14] , \Level16Out208[13] , 
        \Level16Out208[12] , \Level16Out208[11] , \Level16Out208[10] , 
        \Level16Out208[9] , \Level16Out208[8] , \Level16Out208[7] , 
        \Level16Out208[6] , \Level16Out208[5] , \Level16Out208[4] , 
        \Level16Out208[3] , \Level16Out208[2] , \Level16Out208[1] , 
        \Level16Out208[0] }), .Read1(\Level16Load192[0] ), .Read2(
        \Level16Load208[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_88_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load88[0] ), .Out({\Level8Out88[31] , \Level8Out88[30] , 
        \Level8Out88[29] , \Level8Out88[28] , \Level8Out88[27] , 
        \Level8Out88[26] , \Level8Out88[25] , \Level8Out88[24] , 
        \Level8Out88[23] , \Level8Out88[22] , \Level8Out88[21] , 
        \Level8Out88[20] , \Level8Out88[19] , \Level8Out88[18] , 
        \Level8Out88[17] , \Level8Out88[16] , \Level8Out88[15] , 
        \Level8Out88[14] , \Level8Out88[13] , \Level8Out88[12] , 
        \Level8Out88[11] , \Level8Out88[10] , \Level8Out88[9] , 
        \Level8Out88[8] , \Level8Out88[7] , \Level8Out88[6] , \Level8Out88[5] , 
        \Level8Out88[4] , \Level8Out88[3] , \Level8Out88[2] , \Level8Out88[1] , 
        \Level8Out88[0] }), .In1({\Level4Out88[31] , \Level4Out88[30] , 
        \Level4Out88[29] , \Level4Out88[28] , \Level4Out88[27] , 
        \Level4Out88[26] , \Level4Out88[25] , \Level4Out88[24] , 
        \Level4Out88[23] , \Level4Out88[22] , \Level4Out88[21] , 
        \Level4Out88[20] , \Level4Out88[19] , \Level4Out88[18] , 
        \Level4Out88[17] , \Level4Out88[16] , \Level4Out88[15] , 
        \Level4Out88[14] , \Level4Out88[13] , \Level4Out88[12] , 
        \Level4Out88[11] , \Level4Out88[10] , \Level4Out88[9] , 
        \Level4Out88[8] , \Level4Out88[7] , \Level4Out88[6] , \Level4Out88[5] , 
        \Level4Out88[4] , \Level4Out88[3] , \Level4Out88[2] , \Level4Out88[1] , 
        \Level4Out88[0] }), .In2({\Level4Out92[31] , \Level4Out92[30] , 
        \Level4Out92[29] , \Level4Out92[28] , \Level4Out92[27] , 
        \Level4Out92[26] , \Level4Out92[25] , \Level4Out92[24] , 
        \Level4Out92[23] , \Level4Out92[22] , \Level4Out92[21] , 
        \Level4Out92[20] , \Level4Out92[19] , \Level4Out92[18] , 
        \Level4Out92[17] , \Level4Out92[16] , \Level4Out92[15] , 
        \Level4Out92[14] , \Level4Out92[13] , \Level4Out92[12] , 
        \Level4Out92[11] , \Level4Out92[10] , \Level4Out92[9] , 
        \Level4Out92[8] , \Level4Out92[7] , \Level4Out92[6] , \Level4Out92[5] , 
        \Level4Out92[4] , \Level4Out92[3] , \Level4Out92[2] , \Level4Out92[1] , 
        \Level4Out92[0] }), .Read1(\Level4Load88[0] ), .Read2(
        \Level4Load92[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_96_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load96[0] ), .Out({\Level2Out96[31] , \Level2Out96[30] , 
        \Level2Out96[29] , \Level2Out96[28] , \Level2Out96[27] , 
        \Level2Out96[26] , \Level2Out96[25] , \Level2Out96[24] , 
        \Level2Out96[23] , \Level2Out96[22] , \Level2Out96[21] , 
        \Level2Out96[20] , \Level2Out96[19] , \Level2Out96[18] , 
        \Level2Out96[17] , \Level2Out96[16] , \Level2Out96[15] , 
        \Level2Out96[14] , \Level2Out96[13] , \Level2Out96[12] , 
        \Level2Out96[11] , \Level2Out96[10] , \Level2Out96[9] , 
        \Level2Out96[8] , \Level2Out96[7] , \Level2Out96[6] , \Level2Out96[5] , 
        \Level2Out96[4] , \Level2Out96[3] , \Level2Out96[2] , \Level2Out96[1] , 
        \Level2Out96[0] }), .In1({\Level1Out96[31] , \Level1Out96[30] , 
        \Level1Out96[29] , \Level1Out96[28] , \Level1Out96[27] , 
        \Level1Out96[26] , \Level1Out96[25] , \Level1Out96[24] , 
        \Level1Out96[23] , \Level1Out96[22] , \Level1Out96[21] , 
        \Level1Out96[20] , \Level1Out96[19] , \Level1Out96[18] , 
        \Level1Out96[17] , \Level1Out96[16] , \Level1Out96[15] , 
        \Level1Out96[14] , \Level1Out96[13] , \Level1Out96[12] , 
        \Level1Out96[11] , \Level1Out96[10] , \Level1Out96[9] , 
        \Level1Out96[8] , \Level1Out96[7] , \Level1Out96[6] , \Level1Out96[5] , 
        \Level1Out96[4] , \Level1Out96[3] , \Level1Out96[2] , \Level1Out96[1] , 
        \Level1Out96[0] }), .In2({\Level1Out97[31] , \Level1Out97[30] , 
        \Level1Out97[29] , \Level1Out97[28] , \Level1Out97[27] , 
        \Level1Out97[26] , \Level1Out97[25] , \Level1Out97[24] , 
        \Level1Out97[23] , \Level1Out97[22] , \Level1Out97[21] , 
        \Level1Out97[20] , \Level1Out97[19] , \Level1Out97[18] , 
        \Level1Out97[17] , \Level1Out97[16] , \Level1Out97[15] , 
        \Level1Out97[14] , \Level1Out97[13] , \Level1Out97[12] , 
        \Level1Out97[11] , \Level1Out97[10] , \Level1Out97[9] , 
        \Level1Out97[8] , \Level1Out97[7] , \Level1Out97[6] , \Level1Out97[5] , 
        \Level1Out97[4] , \Level1Out97[3] , \Level1Out97[2] , \Level1Out97[1] , 
        \Level1Out97[0] }), .Read1(\Level1Load96[0] ), .Read2(
        \Level1Load97[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_146_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load146[0] ), .Out({\Level2Out146[31] , \Level2Out146[30] , 
        \Level2Out146[29] , \Level2Out146[28] , \Level2Out146[27] , 
        \Level2Out146[26] , \Level2Out146[25] , \Level2Out146[24] , 
        \Level2Out146[23] , \Level2Out146[22] , \Level2Out146[21] , 
        \Level2Out146[20] , \Level2Out146[19] , \Level2Out146[18] , 
        \Level2Out146[17] , \Level2Out146[16] , \Level2Out146[15] , 
        \Level2Out146[14] , \Level2Out146[13] , \Level2Out146[12] , 
        \Level2Out146[11] , \Level2Out146[10] , \Level2Out146[9] , 
        \Level2Out146[8] , \Level2Out146[7] , \Level2Out146[6] , 
        \Level2Out146[5] , \Level2Out146[4] , \Level2Out146[3] , 
        \Level2Out146[2] , \Level2Out146[1] , \Level2Out146[0] }), .In1({
        \Level1Out146[31] , \Level1Out146[30] , \Level1Out146[29] , 
        \Level1Out146[28] , \Level1Out146[27] , \Level1Out146[26] , 
        \Level1Out146[25] , \Level1Out146[24] , \Level1Out146[23] , 
        \Level1Out146[22] , \Level1Out146[21] , \Level1Out146[20] , 
        \Level1Out146[19] , \Level1Out146[18] , \Level1Out146[17] , 
        \Level1Out146[16] , \Level1Out146[15] , \Level1Out146[14] , 
        \Level1Out146[13] , \Level1Out146[12] , \Level1Out146[11] , 
        \Level1Out146[10] , \Level1Out146[9] , \Level1Out146[8] , 
        \Level1Out146[7] , \Level1Out146[6] , \Level1Out146[5] , 
        \Level1Out146[4] , \Level1Out146[3] , \Level1Out146[2] , 
        \Level1Out146[1] , \Level1Out146[0] }), .In2({\Level1Out147[31] , 
        \Level1Out147[30] , \Level1Out147[29] , \Level1Out147[28] , 
        \Level1Out147[27] , \Level1Out147[26] , \Level1Out147[25] , 
        \Level1Out147[24] , \Level1Out147[23] , \Level1Out147[22] , 
        \Level1Out147[21] , \Level1Out147[20] , \Level1Out147[19] , 
        \Level1Out147[18] , \Level1Out147[17] , \Level1Out147[16] , 
        \Level1Out147[15] , \Level1Out147[14] , \Level1Out147[13] , 
        \Level1Out147[12] , \Level1Out147[11] , \Level1Out147[10] , 
        \Level1Out147[9] , \Level1Out147[8] , \Level1Out147[7] , 
        \Level1Out147[6] , \Level1Out147[5] , \Level1Out147[4] , 
        \Level1Out147[3] , \Level1Out147[2] , \Level1Out147[1] , 
        \Level1Out147[0] }), .Read1(\Level1Load146[0] ), .Read2(
        \Level1Load147[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_244_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load244[0] ), .Out({\Level4Out244[31] , \Level4Out244[30] , 
        \Level4Out244[29] , \Level4Out244[28] , \Level4Out244[27] , 
        \Level4Out244[26] , \Level4Out244[25] , \Level4Out244[24] , 
        \Level4Out244[23] , \Level4Out244[22] , \Level4Out244[21] , 
        \Level4Out244[20] , \Level4Out244[19] , \Level4Out244[18] , 
        \Level4Out244[17] , \Level4Out244[16] , \Level4Out244[15] , 
        \Level4Out244[14] , \Level4Out244[13] , \Level4Out244[12] , 
        \Level4Out244[11] , \Level4Out244[10] , \Level4Out244[9] , 
        \Level4Out244[8] , \Level4Out244[7] , \Level4Out244[6] , 
        \Level4Out244[5] , \Level4Out244[4] , \Level4Out244[3] , 
        \Level4Out244[2] , \Level4Out244[1] , \Level4Out244[0] }), .In1({
        \Level2Out244[31] , \Level2Out244[30] , \Level2Out244[29] , 
        \Level2Out244[28] , \Level2Out244[27] , \Level2Out244[26] , 
        \Level2Out244[25] , \Level2Out244[24] , \Level2Out244[23] , 
        \Level2Out244[22] , \Level2Out244[21] , \Level2Out244[20] , 
        \Level2Out244[19] , \Level2Out244[18] , \Level2Out244[17] , 
        \Level2Out244[16] , \Level2Out244[15] , \Level2Out244[14] , 
        \Level2Out244[13] , \Level2Out244[12] , \Level2Out244[11] , 
        \Level2Out244[10] , \Level2Out244[9] , \Level2Out244[8] , 
        \Level2Out244[7] , \Level2Out244[6] , \Level2Out244[5] , 
        \Level2Out244[4] , \Level2Out244[3] , \Level2Out244[2] , 
        \Level2Out244[1] , \Level2Out244[0] }), .In2({\Level2Out246[31] , 
        \Level2Out246[30] , \Level2Out246[29] , \Level2Out246[28] , 
        \Level2Out246[27] , \Level2Out246[26] , \Level2Out246[25] , 
        \Level2Out246[24] , \Level2Out246[23] , \Level2Out246[22] , 
        \Level2Out246[21] , \Level2Out246[20] , \Level2Out246[19] , 
        \Level2Out246[18] , \Level2Out246[17] , \Level2Out246[16] , 
        \Level2Out246[15] , \Level2Out246[14] , \Level2Out246[13] , 
        \Level2Out246[12] , \Level2Out246[11] , \Level2Out246[10] , 
        \Level2Out246[9] , \Level2Out246[8] , \Level2Out246[7] , 
        \Level2Out246[6] , \Level2Out246[5] , \Level2Out246[4] , 
        \Level2Out246[3] , \Level2Out246[2] , \Level2Out246[1] , 
        \Level2Out246[0] }), .Read1(\Level2Load244[0] ), .Read2(
        \Level2Load246[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_52 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanOut({\ScanLink53[31] , 
        \ScanLink53[30] , \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , 
        \ScanLink53[26] , \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , 
        \ScanLink53[22] , \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , 
        \ScanLink53[18] , \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , 
        \ScanLink53[14] , \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , 
        \ScanLink53[10] , \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , 
        \ScanLink53[6] , \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , 
        \ScanLink53[2] , \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load52[0] ), .Out({
        \Level1Out52[31] , \Level1Out52[30] , \Level1Out52[29] , 
        \Level1Out52[28] , \Level1Out52[27] , \Level1Out52[26] , 
        \Level1Out52[25] , \Level1Out52[24] , \Level1Out52[23] , 
        \Level1Out52[22] , \Level1Out52[21] , \Level1Out52[20] , 
        \Level1Out52[19] , \Level1Out52[18] , \Level1Out52[17] , 
        \Level1Out52[16] , \Level1Out52[15] , \Level1Out52[14] , 
        \Level1Out52[13] , \Level1Out52[12] , \Level1Out52[11] , 
        \Level1Out52[10] , \Level1Out52[9] , \Level1Out52[8] , 
        \Level1Out52[7] , \Level1Out52[6] , \Level1Out52[5] , \Level1Out52[4] , 
        \Level1Out52[3] , \Level1Out52[2] , \Level1Out52[1] , \Level1Out52[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_157 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink157[31] , \ScanLink157[30] , 
        \ScanLink157[29] , \ScanLink157[28] , \ScanLink157[27] , 
        \ScanLink157[26] , \ScanLink157[25] , \ScanLink157[24] , 
        \ScanLink157[23] , \ScanLink157[22] , \ScanLink157[21] , 
        \ScanLink157[20] , \ScanLink157[19] , \ScanLink157[18] , 
        \ScanLink157[17] , \ScanLink157[16] , \ScanLink157[15] , 
        \ScanLink157[14] , \ScanLink157[13] , \ScanLink157[12] , 
        \ScanLink157[11] , \ScanLink157[10] , \ScanLink157[9] , 
        \ScanLink157[8] , \ScanLink157[7] , \ScanLink157[6] , \ScanLink157[5] , 
        \ScanLink157[4] , \ScanLink157[3] , \ScanLink157[2] , \ScanLink157[1] , 
        \ScanLink157[0] }), .ScanOut({\ScanLink158[31] , \ScanLink158[30] , 
        \ScanLink158[29] , \ScanLink158[28] , \ScanLink158[27] , 
        \ScanLink158[26] , \ScanLink158[25] , \ScanLink158[24] , 
        \ScanLink158[23] , \ScanLink158[22] , \ScanLink158[21] , 
        \ScanLink158[20] , \ScanLink158[19] , \ScanLink158[18] , 
        \ScanLink158[17] , \ScanLink158[16] , \ScanLink158[15] , 
        \ScanLink158[14] , \ScanLink158[13] , \ScanLink158[12] , 
        \ScanLink158[11] , \ScanLink158[10] , \ScanLink158[9] , 
        \ScanLink158[8] , \ScanLink158[7] , \ScanLink158[6] , \ScanLink158[5] , 
        \ScanLink158[4] , \ScanLink158[3] , \ScanLink158[2] , \ScanLink158[1] , 
        \ScanLink158[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load157[0] ), .Out({\Level1Out157[31] , \Level1Out157[30] , 
        \Level1Out157[29] , \Level1Out157[28] , \Level1Out157[27] , 
        \Level1Out157[26] , \Level1Out157[25] , \Level1Out157[24] , 
        \Level1Out157[23] , \Level1Out157[22] , \Level1Out157[21] , 
        \Level1Out157[20] , \Level1Out157[19] , \Level1Out157[18] , 
        \Level1Out157[17] , \Level1Out157[16] , \Level1Out157[15] , 
        \Level1Out157[14] , \Level1Out157[13] , \Level1Out157[12] , 
        \Level1Out157[11] , \Level1Out157[10] , \Level1Out157[9] , 
        \Level1Out157[8] , \Level1Out157[7] , \Level1Out157[6] , 
        \Level1Out157[5] , \Level1Out157[4] , \Level1Out157[3] , 
        \Level1Out157[2] , \Level1Out157[1] , \Level1Out157[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_18_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load18[0] ), .Out({\Level2Out18[31] , \Level2Out18[30] , 
        \Level2Out18[29] , \Level2Out18[28] , \Level2Out18[27] , 
        \Level2Out18[26] , \Level2Out18[25] , \Level2Out18[24] , 
        \Level2Out18[23] , \Level2Out18[22] , \Level2Out18[21] , 
        \Level2Out18[20] , \Level2Out18[19] , \Level2Out18[18] , 
        \Level2Out18[17] , \Level2Out18[16] , \Level2Out18[15] , 
        \Level2Out18[14] , \Level2Out18[13] , \Level2Out18[12] , 
        \Level2Out18[11] , \Level2Out18[10] , \Level2Out18[9] , 
        \Level2Out18[8] , \Level2Out18[7] , \Level2Out18[6] , \Level2Out18[5] , 
        \Level2Out18[4] , \Level2Out18[3] , \Level2Out18[2] , \Level2Out18[1] , 
        \Level2Out18[0] }), .In1({\Level1Out18[31] , \Level1Out18[30] , 
        \Level1Out18[29] , \Level1Out18[28] , \Level1Out18[27] , 
        \Level1Out18[26] , \Level1Out18[25] , \Level1Out18[24] , 
        \Level1Out18[23] , \Level1Out18[22] , \Level1Out18[21] , 
        \Level1Out18[20] , \Level1Out18[19] , \Level1Out18[18] , 
        \Level1Out18[17] , \Level1Out18[16] , \Level1Out18[15] , 
        \Level1Out18[14] , \Level1Out18[13] , \Level1Out18[12] , 
        \Level1Out18[11] , \Level1Out18[10] , \Level1Out18[9] , 
        \Level1Out18[8] , \Level1Out18[7] , \Level1Out18[6] , \Level1Out18[5] , 
        \Level1Out18[4] , \Level1Out18[3] , \Level1Out18[2] , \Level1Out18[1] , 
        \Level1Out18[0] }), .In2({\Level1Out19[31] , \Level1Out19[30] , 
        \Level1Out19[29] , \Level1Out19[28] , \Level1Out19[27] , 
        \Level1Out19[26] , \Level1Out19[25] , \Level1Out19[24] , 
        \Level1Out19[23] , \Level1Out19[22] , \Level1Out19[21] , 
        \Level1Out19[20] , \Level1Out19[19] , \Level1Out19[18] , 
        \Level1Out19[17] , \Level1Out19[16] , \Level1Out19[15] , 
        \Level1Out19[14] , \Level1Out19[13] , \Level1Out19[12] , 
        \Level1Out19[11] , \Level1Out19[10] , \Level1Out19[9] , 
        \Level1Out19[8] , \Level1Out19[7] , \Level1Out19[6] , \Level1Out19[5] , 
        \Level1Out19[4] , \Level1Out19[3] , \Level1Out19[2] , \Level1Out19[1] , 
        \Level1Out19[0] }), .Read1(\Level1Load18[0] ), .Read2(
        \Level1Load19[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_174_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load174[0] ), .Out({\Level2Out174[31] , \Level2Out174[30] , 
        \Level2Out174[29] , \Level2Out174[28] , \Level2Out174[27] , 
        \Level2Out174[26] , \Level2Out174[25] , \Level2Out174[24] , 
        \Level2Out174[23] , \Level2Out174[22] , \Level2Out174[21] , 
        \Level2Out174[20] , \Level2Out174[19] , \Level2Out174[18] , 
        \Level2Out174[17] , \Level2Out174[16] , \Level2Out174[15] , 
        \Level2Out174[14] , \Level2Out174[13] , \Level2Out174[12] , 
        \Level2Out174[11] , \Level2Out174[10] , \Level2Out174[9] , 
        \Level2Out174[8] , \Level2Out174[7] , \Level2Out174[6] , 
        \Level2Out174[5] , \Level2Out174[4] , \Level2Out174[3] , 
        \Level2Out174[2] , \Level2Out174[1] , \Level2Out174[0] }), .In1({
        \Level1Out174[31] , \Level1Out174[30] , \Level1Out174[29] , 
        \Level1Out174[28] , \Level1Out174[27] , \Level1Out174[26] , 
        \Level1Out174[25] , \Level1Out174[24] , \Level1Out174[23] , 
        \Level1Out174[22] , \Level1Out174[21] , \Level1Out174[20] , 
        \Level1Out174[19] , \Level1Out174[18] , \Level1Out174[17] , 
        \Level1Out174[16] , \Level1Out174[15] , \Level1Out174[14] , 
        \Level1Out174[13] , \Level1Out174[12] , \Level1Out174[11] , 
        \Level1Out174[10] , \Level1Out174[9] , \Level1Out174[8] , 
        \Level1Out174[7] , \Level1Out174[6] , \Level1Out174[5] , 
        \Level1Out174[4] , \Level1Out174[3] , \Level1Out174[2] , 
        \Level1Out174[1] , \Level1Out174[0] }), .In2({\Level1Out175[31] , 
        \Level1Out175[30] , \Level1Out175[29] , \Level1Out175[28] , 
        \Level1Out175[27] , \Level1Out175[26] , \Level1Out175[25] , 
        \Level1Out175[24] , \Level1Out175[23] , \Level1Out175[22] , 
        \Level1Out175[21] , \Level1Out175[20] , \Level1Out175[19] , 
        \Level1Out175[18] , \Level1Out175[17] , \Level1Out175[16] , 
        \Level1Out175[15] , \Level1Out175[14] , \Level1Out175[13] , 
        \Level1Out175[12] , \Level1Out175[11] , \Level1Out175[10] , 
        \Level1Out175[9] , \Level1Out175[8] , \Level1Out175[7] , 
        \Level1Out175[6] , \Level1Out175[5] , \Level1Out175[4] , 
        \Level1Out175[3] , \Level1Out175[2] , \Level1Out175[1] , 
        \Level1Out175[0] }), .Read1(\Level1Load174[0] ), .Read2(
        \Level1Load175[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_168_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load168[0] ), .Out({\Level4Out168[31] , \Level4Out168[30] , 
        \Level4Out168[29] , \Level4Out168[28] , \Level4Out168[27] , 
        \Level4Out168[26] , \Level4Out168[25] , \Level4Out168[24] , 
        \Level4Out168[23] , \Level4Out168[22] , \Level4Out168[21] , 
        \Level4Out168[20] , \Level4Out168[19] , \Level4Out168[18] , 
        \Level4Out168[17] , \Level4Out168[16] , \Level4Out168[15] , 
        \Level4Out168[14] , \Level4Out168[13] , \Level4Out168[12] , 
        \Level4Out168[11] , \Level4Out168[10] , \Level4Out168[9] , 
        \Level4Out168[8] , \Level4Out168[7] , \Level4Out168[6] , 
        \Level4Out168[5] , \Level4Out168[4] , \Level4Out168[3] , 
        \Level4Out168[2] , \Level4Out168[1] , \Level4Out168[0] }), .In1({
        \Level2Out168[31] , \Level2Out168[30] , \Level2Out168[29] , 
        \Level2Out168[28] , \Level2Out168[27] , \Level2Out168[26] , 
        \Level2Out168[25] , \Level2Out168[24] , \Level2Out168[23] , 
        \Level2Out168[22] , \Level2Out168[21] , \Level2Out168[20] , 
        \Level2Out168[19] , \Level2Out168[18] , \Level2Out168[17] , 
        \Level2Out168[16] , \Level2Out168[15] , \Level2Out168[14] , 
        \Level2Out168[13] , \Level2Out168[12] , \Level2Out168[11] , 
        \Level2Out168[10] , \Level2Out168[9] , \Level2Out168[8] , 
        \Level2Out168[7] , \Level2Out168[6] , \Level2Out168[5] , 
        \Level2Out168[4] , \Level2Out168[3] , \Level2Out168[2] , 
        \Level2Out168[1] , \Level2Out168[0] }), .In2({\Level2Out170[31] , 
        \Level2Out170[30] , \Level2Out170[29] , \Level2Out170[28] , 
        \Level2Out170[27] , \Level2Out170[26] , \Level2Out170[25] , 
        \Level2Out170[24] , \Level2Out170[23] , \Level2Out170[22] , 
        \Level2Out170[21] , \Level2Out170[20] , \Level2Out170[19] , 
        \Level2Out170[18] , \Level2Out170[17] , \Level2Out170[16] , 
        \Level2Out170[15] , \Level2Out170[14] , \Level2Out170[13] , 
        \Level2Out170[12] , \Level2Out170[11] , \Level2Out170[10] , 
        \Level2Out170[9] , \Level2Out170[8] , \Level2Out170[7] , 
        \Level2Out170[6] , \Level2Out170[5] , \Level2Out170[4] , 
        \Level2Out170[3] , \Level2Out170[2] , \Level2Out170[1] , 
        \Level2Out170[0] }), .Read1(\Level2Load168[0] ), .Read2(
        \Level2Load170[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_170 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink170[31] , \ScanLink170[30] , 
        \ScanLink170[29] , \ScanLink170[28] , \ScanLink170[27] , 
        \ScanLink170[26] , \ScanLink170[25] , \ScanLink170[24] , 
        \ScanLink170[23] , \ScanLink170[22] , \ScanLink170[21] , 
        \ScanLink170[20] , \ScanLink170[19] , \ScanLink170[18] , 
        \ScanLink170[17] , \ScanLink170[16] , \ScanLink170[15] , 
        \ScanLink170[14] , \ScanLink170[13] , \ScanLink170[12] , 
        \ScanLink170[11] , \ScanLink170[10] , \ScanLink170[9] , 
        \ScanLink170[8] , \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , 
        \ScanLink170[4] , \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , 
        \ScanLink170[0] }), .ScanOut({\ScanLink171[31] , \ScanLink171[30] , 
        \ScanLink171[29] , \ScanLink171[28] , \ScanLink171[27] , 
        \ScanLink171[26] , \ScanLink171[25] , \ScanLink171[24] , 
        \ScanLink171[23] , \ScanLink171[22] , \ScanLink171[21] , 
        \ScanLink171[20] , \ScanLink171[19] , \ScanLink171[18] , 
        \ScanLink171[17] , \ScanLink171[16] , \ScanLink171[15] , 
        \ScanLink171[14] , \ScanLink171[13] , \ScanLink171[12] , 
        \ScanLink171[11] , \ScanLink171[10] , \ScanLink171[9] , 
        \ScanLink171[8] , \ScanLink171[7] , \ScanLink171[6] , \ScanLink171[5] , 
        \ScanLink171[4] , \ScanLink171[3] , \ScanLink171[2] , \ScanLink171[1] , 
        \ScanLink171[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load170[0] ), .Out({\Level1Out170[31] , \Level1Out170[30] , 
        \Level1Out170[29] , \Level1Out170[28] , \Level1Out170[27] , 
        \Level1Out170[26] , \Level1Out170[25] , \Level1Out170[24] , 
        \Level1Out170[23] , \Level1Out170[22] , \Level1Out170[21] , 
        \Level1Out170[20] , \Level1Out170[19] , \Level1Out170[18] , 
        \Level1Out170[17] , \Level1Out170[16] , \Level1Out170[15] , 
        \Level1Out170[14] , \Level1Out170[13] , \Level1Out170[12] , 
        \Level1Out170[11] , \Level1Out170[10] , \Level1Out170[9] , 
        \Level1Out170[8] , \Level1Out170[7] , \Level1Out170[6] , 
        \Level1Out170[5] , \Level1Out170[4] , \Level1Out170[3] , 
        \Level1Out170[2] , \Level1Out170[1] , \Level1Out170[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_240_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load240[0] ), .Out({\Level2Out240[31] , \Level2Out240[30] , 
        \Level2Out240[29] , \Level2Out240[28] , \Level2Out240[27] , 
        \Level2Out240[26] , \Level2Out240[25] , \Level2Out240[24] , 
        \Level2Out240[23] , \Level2Out240[22] , \Level2Out240[21] , 
        \Level2Out240[20] , \Level2Out240[19] , \Level2Out240[18] , 
        \Level2Out240[17] , \Level2Out240[16] , \Level2Out240[15] , 
        \Level2Out240[14] , \Level2Out240[13] , \Level2Out240[12] , 
        \Level2Out240[11] , \Level2Out240[10] , \Level2Out240[9] , 
        \Level2Out240[8] , \Level2Out240[7] , \Level2Out240[6] , 
        \Level2Out240[5] , \Level2Out240[4] , \Level2Out240[3] , 
        \Level2Out240[2] , \Level2Out240[1] , \Level2Out240[0] }), .In1({
        \Level1Out240[31] , \Level1Out240[30] , \Level1Out240[29] , 
        \Level1Out240[28] , \Level1Out240[27] , \Level1Out240[26] , 
        \Level1Out240[25] , \Level1Out240[24] , \Level1Out240[23] , 
        \Level1Out240[22] , \Level1Out240[21] , \Level1Out240[20] , 
        \Level1Out240[19] , \Level1Out240[18] , \Level1Out240[17] , 
        \Level1Out240[16] , \Level1Out240[15] , \Level1Out240[14] , 
        \Level1Out240[13] , \Level1Out240[12] , \Level1Out240[11] , 
        \Level1Out240[10] , \Level1Out240[9] , \Level1Out240[8] , 
        \Level1Out240[7] , \Level1Out240[6] , \Level1Out240[5] , 
        \Level1Out240[4] , \Level1Out240[3] , \Level1Out240[2] , 
        \Level1Out240[1] , \Level1Out240[0] }), .In2({\Level1Out241[31] , 
        \Level1Out241[30] , \Level1Out241[29] , \Level1Out241[28] , 
        \Level1Out241[27] , \Level1Out241[26] , \Level1Out241[25] , 
        \Level1Out241[24] , \Level1Out241[23] , \Level1Out241[22] , 
        \Level1Out241[21] , \Level1Out241[20] , \Level1Out241[19] , 
        \Level1Out241[18] , \Level1Out241[17] , \Level1Out241[16] , 
        \Level1Out241[15] , \Level1Out241[14] , \Level1Out241[13] , 
        \Level1Out241[12] , \Level1Out241[11] , \Level1Out241[10] , 
        \Level1Out241[9] , \Level1Out241[8] , \Level1Out241[7] , 
        \Level1Out241[6] , \Level1Out241[5] , \Level1Out241[4] , 
        \Level1Out241[3] , \Level1Out241[2] , \Level1Out241[1] , 
        \Level1Out241[0] }), .Read1(\Level1Load240[0] ), .Read2(
        \Level1Load241[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_240 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink240[31] , \ScanLink240[30] , 
        \ScanLink240[29] , \ScanLink240[28] , \ScanLink240[27] , 
        \ScanLink240[26] , \ScanLink240[25] , \ScanLink240[24] , 
        \ScanLink240[23] , \ScanLink240[22] , \ScanLink240[21] , 
        \ScanLink240[20] , \ScanLink240[19] , \ScanLink240[18] , 
        \ScanLink240[17] , \ScanLink240[16] , \ScanLink240[15] , 
        \ScanLink240[14] , \ScanLink240[13] , \ScanLink240[12] , 
        \ScanLink240[11] , \ScanLink240[10] , \ScanLink240[9] , 
        \ScanLink240[8] , \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , 
        \ScanLink240[4] , \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , 
        \ScanLink240[0] }), .ScanOut({\ScanLink241[31] , \ScanLink241[30] , 
        \ScanLink241[29] , \ScanLink241[28] , \ScanLink241[27] , 
        \ScanLink241[26] , \ScanLink241[25] , \ScanLink241[24] , 
        \ScanLink241[23] , \ScanLink241[22] , \ScanLink241[21] , 
        \ScanLink241[20] , \ScanLink241[19] , \ScanLink241[18] , 
        \ScanLink241[17] , \ScanLink241[16] , \ScanLink241[15] , 
        \ScanLink241[14] , \ScanLink241[13] , \ScanLink241[12] , 
        \ScanLink241[11] , \ScanLink241[10] , \ScanLink241[9] , 
        \ScanLink241[8] , \ScanLink241[7] , \ScanLink241[6] , \ScanLink241[5] , 
        \ScanLink241[4] , \ScanLink241[3] , \ScanLink241[2] , \ScanLink241[1] , 
        \ScanLink241[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load240[0] ), .Out({\Level1Out240[31] , \Level1Out240[30] , 
        \Level1Out240[29] , \Level1Out240[28] , \Level1Out240[27] , 
        \Level1Out240[26] , \Level1Out240[25] , \Level1Out240[24] , 
        \Level1Out240[23] , \Level1Out240[22] , \Level1Out240[21] , 
        \Level1Out240[20] , \Level1Out240[19] , \Level1Out240[18] , 
        \Level1Out240[17] , \Level1Out240[16] , \Level1Out240[15] , 
        \Level1Out240[14] , \Level1Out240[13] , \Level1Out240[12] , 
        \Level1Out240[11] , \Level1Out240[10] , \Level1Out240[9] , 
        \Level1Out240[8] , \Level1Out240[7] , \Level1Out240[6] , 
        \Level1Out240[5] , \Level1Out240[4] , \Level1Out240[3] , 
        \Level1Out240[2] , \Level1Out240[1] , \Level1Out240[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load32[0] ), .Out({\Level2Out32[31] , \Level2Out32[30] , 
        \Level2Out32[29] , \Level2Out32[28] , \Level2Out32[27] , 
        \Level2Out32[26] , \Level2Out32[25] , \Level2Out32[24] , 
        \Level2Out32[23] , \Level2Out32[22] , \Level2Out32[21] , 
        \Level2Out32[20] , \Level2Out32[19] , \Level2Out32[18] , 
        \Level2Out32[17] , \Level2Out32[16] , \Level2Out32[15] , 
        \Level2Out32[14] , \Level2Out32[13] , \Level2Out32[12] , 
        \Level2Out32[11] , \Level2Out32[10] , \Level2Out32[9] , 
        \Level2Out32[8] , \Level2Out32[7] , \Level2Out32[6] , \Level2Out32[5] , 
        \Level2Out32[4] , \Level2Out32[3] , \Level2Out32[2] , \Level2Out32[1] , 
        \Level2Out32[0] }), .In1({\Level1Out32[31] , \Level1Out32[30] , 
        \Level1Out32[29] , \Level1Out32[28] , \Level1Out32[27] , 
        \Level1Out32[26] , \Level1Out32[25] , \Level1Out32[24] , 
        \Level1Out32[23] , \Level1Out32[22] , \Level1Out32[21] , 
        \Level1Out32[20] , \Level1Out32[19] , \Level1Out32[18] , 
        \Level1Out32[17] , \Level1Out32[16] , \Level1Out32[15] , 
        \Level1Out32[14] , \Level1Out32[13] , \Level1Out32[12] , 
        \Level1Out32[11] , \Level1Out32[10] , \Level1Out32[9] , 
        \Level1Out32[8] , \Level1Out32[7] , \Level1Out32[6] , \Level1Out32[5] , 
        \Level1Out32[4] , \Level1Out32[3] , \Level1Out32[2] , \Level1Out32[1] , 
        \Level1Out32[0] }), .In2({\Level1Out33[31] , \Level1Out33[30] , 
        \Level1Out33[29] , \Level1Out33[28] , \Level1Out33[27] , 
        \Level1Out33[26] , \Level1Out33[25] , \Level1Out33[24] , 
        \Level1Out33[23] , \Level1Out33[22] , \Level1Out33[21] , 
        \Level1Out33[20] , \Level1Out33[19] , \Level1Out33[18] , 
        \Level1Out33[17] , \Level1Out33[16] , \Level1Out33[15] , 
        \Level1Out33[14] , \Level1Out33[13] , \Level1Out33[12] , 
        \Level1Out33[11] , \Level1Out33[10] , \Level1Out33[9] , 
        \Level1Out33[8] , \Level1Out33[7] , \Level1Out33[6] , \Level1Out33[5] , 
        \Level1Out33[4] , \Level1Out33[3] , \Level1Out33[2] , \Level1Out33[1] , 
        \Level1Out33[0] }), .Read1(\Level1Load32[0] ), .Read2(
        \Level1Load33[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_55 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanOut({\ScanLink56[31] , 
        \ScanLink56[30] , \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , 
        \ScanLink56[26] , \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , 
        \ScanLink56[22] , \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , 
        \ScanLink56[18] , \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , 
        \ScanLink56[14] , \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , 
        \ScanLink56[10] , \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , 
        \ScanLink56[6] , \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , 
        \ScanLink56[2] , \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load55[0] ), .Out({
        \Level1Out55[31] , \Level1Out55[30] , \Level1Out55[29] , 
        \Level1Out55[28] , \Level1Out55[27] , \Level1Out55[26] , 
        \Level1Out55[25] , \Level1Out55[24] , \Level1Out55[23] , 
        \Level1Out55[22] , \Level1Out55[21] , \Level1Out55[20] , 
        \Level1Out55[19] , \Level1Out55[18] , \Level1Out55[17] , 
        \Level1Out55[16] , \Level1Out55[15] , \Level1Out55[14] , 
        \Level1Out55[13] , \Level1Out55[12] , \Level1Out55[11] , 
        \Level1Out55[10] , \Level1Out55[9] , \Level1Out55[8] , 
        \Level1Out55[7] , \Level1Out55[6] , \Level1Out55[5] , \Level1Out55[4] , 
        \Level1Out55[3] , \Level1Out55[2] , \Level1Out55[1] , \Level1Out55[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_72 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink72[31] , \ScanLink72[30] , 
        \ScanLink72[29] , \ScanLink72[28] , \ScanLink72[27] , \ScanLink72[26] , 
        \ScanLink72[25] , \ScanLink72[24] , \ScanLink72[23] , \ScanLink72[22] , 
        \ScanLink72[21] , \ScanLink72[20] , \ScanLink72[19] , \ScanLink72[18] , 
        \ScanLink72[17] , \ScanLink72[16] , \ScanLink72[15] , \ScanLink72[14] , 
        \ScanLink72[13] , \ScanLink72[12] , \ScanLink72[11] , \ScanLink72[10] , 
        \ScanLink72[9] , \ScanLink72[8] , \ScanLink72[7] , \ScanLink72[6] , 
        \ScanLink72[5] , \ScanLink72[4] , \ScanLink72[3] , \ScanLink72[2] , 
        \ScanLink72[1] , \ScanLink72[0] }), .ScanOut({\ScanLink73[31] , 
        \ScanLink73[30] , \ScanLink73[29] , \ScanLink73[28] , \ScanLink73[27] , 
        \ScanLink73[26] , \ScanLink73[25] , \ScanLink73[24] , \ScanLink73[23] , 
        \ScanLink73[22] , \ScanLink73[21] , \ScanLink73[20] , \ScanLink73[19] , 
        \ScanLink73[18] , \ScanLink73[17] , \ScanLink73[16] , \ScanLink73[15] , 
        \ScanLink73[14] , \ScanLink73[13] , \ScanLink73[12] , \ScanLink73[11] , 
        \ScanLink73[10] , \ScanLink73[9] , \ScanLink73[8] , \ScanLink73[7] , 
        \ScanLink73[6] , \ScanLink73[5] , \ScanLink73[4] , \ScanLink73[3] , 
        \ScanLink73[2] , \ScanLink73[1] , \ScanLink73[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load72[0] ), .Out({
        \Level1Out72[31] , \Level1Out72[30] , \Level1Out72[29] , 
        \Level1Out72[28] , \Level1Out72[27] , \Level1Out72[26] , 
        \Level1Out72[25] , \Level1Out72[24] , \Level1Out72[23] , 
        \Level1Out72[22] , \Level1Out72[21] , \Level1Out72[20] , 
        \Level1Out72[19] , \Level1Out72[18] , \Level1Out72[17] , 
        \Level1Out72[16] , \Level1Out72[15] , \Level1Out72[14] , 
        \Level1Out72[13] , \Level1Out72[12] , \Level1Out72[11] , 
        \Level1Out72[10] , \Level1Out72[9] , \Level1Out72[8] , 
        \Level1Out72[7] , \Level1Out72[6] , \Level1Out72[5] , \Level1Out72[4] , 
        \Level1Out72[3] , \Level1Out72[2] , \Level1Out72[1] , \Level1Out72[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_75 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink75[31] , \ScanLink75[30] , 
        \ScanLink75[29] , \ScanLink75[28] , \ScanLink75[27] , \ScanLink75[26] , 
        \ScanLink75[25] , \ScanLink75[24] , \ScanLink75[23] , \ScanLink75[22] , 
        \ScanLink75[21] , \ScanLink75[20] , \ScanLink75[19] , \ScanLink75[18] , 
        \ScanLink75[17] , \ScanLink75[16] , \ScanLink75[15] , \ScanLink75[14] , 
        \ScanLink75[13] , \ScanLink75[12] , \ScanLink75[11] , \ScanLink75[10] , 
        \ScanLink75[9] , \ScanLink75[8] , \ScanLink75[7] , \ScanLink75[6] , 
        \ScanLink75[5] , \ScanLink75[4] , \ScanLink75[3] , \ScanLink75[2] , 
        \ScanLink75[1] , \ScanLink75[0] }), .ScanOut({\ScanLink76[31] , 
        \ScanLink76[30] , \ScanLink76[29] , \ScanLink76[28] , \ScanLink76[27] , 
        \ScanLink76[26] , \ScanLink76[25] , \ScanLink76[24] , \ScanLink76[23] , 
        \ScanLink76[22] , \ScanLink76[21] , \ScanLink76[20] , \ScanLink76[19] , 
        \ScanLink76[18] , \ScanLink76[17] , \ScanLink76[16] , \ScanLink76[15] , 
        \ScanLink76[14] , \ScanLink76[13] , \ScanLink76[12] , \ScanLink76[11] , 
        \ScanLink76[10] , \ScanLink76[9] , \ScanLink76[8] , \ScanLink76[7] , 
        \ScanLink76[6] , \ScanLink76[5] , \ScanLink76[4] , \ScanLink76[3] , 
        \ScanLink76[2] , \ScanLink76[1] , \ScanLink76[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load75[0] ), .Out({
        \Level1Out75[31] , \Level1Out75[30] , \Level1Out75[29] , 
        \Level1Out75[28] , \Level1Out75[27] , \Level1Out75[26] , 
        \Level1Out75[25] , \Level1Out75[24] , \Level1Out75[23] , 
        \Level1Out75[22] , \Level1Out75[21] , \Level1Out75[20] , 
        \Level1Out75[19] , \Level1Out75[18] , \Level1Out75[17] , 
        \Level1Out75[16] , \Level1Out75[15] , \Level1Out75[14] , 
        \Level1Out75[13] , \Level1Out75[12] , \Level1Out75[11] , 
        \Level1Out75[10] , \Level1Out75[9] , \Level1Out75[8] , 
        \Level1Out75[7] , \Level1Out75[6] , \Level1Out75[5] , \Level1Out75[4] , 
        \Level1Out75[3] , \Level1Out75[2] , \Level1Out75[1] , \Level1Out75[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_92_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load92[0] ), .Out({\Level4Out92[31] , \Level4Out92[30] , 
        \Level4Out92[29] , \Level4Out92[28] , \Level4Out92[27] , 
        \Level4Out92[26] , \Level4Out92[25] , \Level4Out92[24] , 
        \Level4Out92[23] , \Level4Out92[22] , \Level4Out92[21] , 
        \Level4Out92[20] , \Level4Out92[19] , \Level4Out92[18] , 
        \Level4Out92[17] , \Level4Out92[16] , \Level4Out92[15] , 
        \Level4Out92[14] , \Level4Out92[13] , \Level4Out92[12] , 
        \Level4Out92[11] , \Level4Out92[10] , \Level4Out92[9] , 
        \Level4Out92[8] , \Level4Out92[7] , \Level4Out92[6] , \Level4Out92[5] , 
        \Level4Out92[4] , \Level4Out92[3] , \Level4Out92[2] , \Level4Out92[1] , 
        \Level4Out92[0] }), .In1({\Level2Out92[31] , \Level2Out92[30] , 
        \Level2Out92[29] , \Level2Out92[28] , \Level2Out92[27] , 
        \Level2Out92[26] , \Level2Out92[25] , \Level2Out92[24] , 
        \Level2Out92[23] , \Level2Out92[22] , \Level2Out92[21] , 
        \Level2Out92[20] , \Level2Out92[19] , \Level2Out92[18] , 
        \Level2Out92[17] , \Level2Out92[16] , \Level2Out92[15] , 
        \Level2Out92[14] , \Level2Out92[13] , \Level2Out92[12] , 
        \Level2Out92[11] , \Level2Out92[10] , \Level2Out92[9] , 
        \Level2Out92[8] , \Level2Out92[7] , \Level2Out92[6] , \Level2Out92[5] , 
        \Level2Out92[4] , \Level2Out92[3] , \Level2Out92[2] , \Level2Out92[1] , 
        \Level2Out92[0] }), .In2({\Level2Out94[31] , \Level2Out94[30] , 
        \Level2Out94[29] , \Level2Out94[28] , \Level2Out94[27] , 
        \Level2Out94[26] , \Level2Out94[25] , \Level2Out94[24] , 
        \Level2Out94[23] , \Level2Out94[22] , \Level2Out94[21] , 
        \Level2Out94[20] , \Level2Out94[19] , \Level2Out94[18] , 
        \Level2Out94[17] , \Level2Out94[16] , \Level2Out94[15] , 
        \Level2Out94[14] , \Level2Out94[13] , \Level2Out94[12] , 
        \Level2Out94[11] , \Level2Out94[10] , \Level2Out94[9] , 
        \Level2Out94[8] , \Level2Out94[7] , \Level2Out94[6] , \Level2Out94[5] , 
        \Level2Out94[4] , \Level2Out94[3] , \Level2Out94[2] , \Level2Out94[1] , 
        \Level2Out94[0] }), .Read1(\Level2Load92[0] ), .Read2(
        \Level2Load94[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_90 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink90[31] , \ScanLink90[30] , 
        \ScanLink90[29] , \ScanLink90[28] , \ScanLink90[27] , \ScanLink90[26] , 
        \ScanLink90[25] , \ScanLink90[24] , \ScanLink90[23] , \ScanLink90[22] , 
        \ScanLink90[21] , \ScanLink90[20] , \ScanLink90[19] , \ScanLink90[18] , 
        \ScanLink90[17] , \ScanLink90[16] , \ScanLink90[15] , \ScanLink90[14] , 
        \ScanLink90[13] , \ScanLink90[12] , \ScanLink90[11] , \ScanLink90[10] , 
        \ScanLink90[9] , \ScanLink90[8] , \ScanLink90[7] , \ScanLink90[6] , 
        \ScanLink90[5] , \ScanLink90[4] , \ScanLink90[3] , \ScanLink90[2] , 
        \ScanLink90[1] , \ScanLink90[0] }), .ScanOut({\ScanLink91[31] , 
        \ScanLink91[30] , \ScanLink91[29] , \ScanLink91[28] , \ScanLink91[27] , 
        \ScanLink91[26] , \ScanLink91[25] , \ScanLink91[24] , \ScanLink91[23] , 
        \ScanLink91[22] , \ScanLink91[21] , \ScanLink91[20] , \ScanLink91[19] , 
        \ScanLink91[18] , \ScanLink91[17] , \ScanLink91[16] , \ScanLink91[15] , 
        \ScanLink91[14] , \ScanLink91[13] , \ScanLink91[12] , \ScanLink91[11] , 
        \ScanLink91[10] , \ScanLink91[9] , \ScanLink91[8] , \ScanLink91[7] , 
        \ScanLink91[6] , \ScanLink91[5] , \ScanLink91[4] , \ScanLink91[3] , 
        \ScanLink91[2] , \ScanLink91[1] , \ScanLink91[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load90[0] ), .Out({
        \Level1Out90[31] , \Level1Out90[30] , \Level1Out90[29] , 
        \Level1Out90[28] , \Level1Out90[27] , \Level1Out90[26] , 
        \Level1Out90[25] , \Level1Out90[24] , \Level1Out90[23] , 
        \Level1Out90[22] , \Level1Out90[21] , \Level1Out90[20] , 
        \Level1Out90[19] , \Level1Out90[18] , \Level1Out90[17] , 
        \Level1Out90[16] , \Level1Out90[15] , \Level1Out90[14] , 
        \Level1Out90[13] , \Level1Out90[12] , \Level1Out90[11] , 
        \Level1Out90[10] , \Level1Out90[9] , \Level1Out90[8] , 
        \Level1Out90[7] , \Level1Out90[6] , \Level1Out90[5] , \Level1Out90[4] , 
        \Level1Out90[3] , \Level1Out90[2] , \Level1Out90[1] , \Level1Out90[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_195 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink195[31] , \ScanLink195[30] , 
        \ScanLink195[29] , \ScanLink195[28] , \ScanLink195[27] , 
        \ScanLink195[26] , \ScanLink195[25] , \ScanLink195[24] , 
        \ScanLink195[23] , \ScanLink195[22] , \ScanLink195[21] , 
        \ScanLink195[20] , \ScanLink195[19] , \ScanLink195[18] , 
        \ScanLink195[17] , \ScanLink195[16] , \ScanLink195[15] , 
        \ScanLink195[14] , \ScanLink195[13] , \ScanLink195[12] , 
        \ScanLink195[11] , \ScanLink195[10] , \ScanLink195[9] , 
        \ScanLink195[8] , \ScanLink195[7] , \ScanLink195[6] , \ScanLink195[5] , 
        \ScanLink195[4] , \ScanLink195[3] , \ScanLink195[2] , \ScanLink195[1] , 
        \ScanLink195[0] }), .ScanOut({\ScanLink196[31] , \ScanLink196[30] , 
        \ScanLink196[29] , \ScanLink196[28] , \ScanLink196[27] , 
        \ScanLink196[26] , \ScanLink196[25] , \ScanLink196[24] , 
        \ScanLink196[23] , \ScanLink196[22] , \ScanLink196[21] , 
        \ScanLink196[20] , \ScanLink196[19] , \ScanLink196[18] , 
        \ScanLink196[17] , \ScanLink196[16] , \ScanLink196[15] , 
        \ScanLink196[14] , \ScanLink196[13] , \ScanLink196[12] , 
        \ScanLink196[11] , \ScanLink196[10] , \ScanLink196[9] , 
        \ScanLink196[8] , \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , 
        \ScanLink196[4] , \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , 
        \ScanLink196[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load195[0] ), .Out({\Level1Out195[31] , \Level1Out195[30] , 
        \Level1Out195[29] , \Level1Out195[28] , \Level1Out195[27] , 
        \Level1Out195[26] , \Level1Out195[25] , \Level1Out195[24] , 
        \Level1Out195[23] , \Level1Out195[22] , \Level1Out195[21] , 
        \Level1Out195[20] , \Level1Out195[19] , \Level1Out195[18] , 
        \Level1Out195[17] , \Level1Out195[16] , \Level1Out195[15] , 
        \Level1Out195[14] , \Level1Out195[13] , \Level1Out195[12] , 
        \Level1Out195[11] , \Level1Out195[10] , \Level1Out195[9] , 
        \Level1Out195[8] , \Level1Out195[7] , \Level1Out195[6] , 
        \Level1Out195[5] , \Level1Out195[4] , \Level1Out195[3] , 
        \Level1Out195[2] , \Level1Out195[1] , \Level1Out195[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_64 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level64Load128[0] ), .Out({\Level64Out128[31] , \Level64Out128[30] , 
        \Level64Out128[29] , \Level64Out128[28] , \Level64Out128[27] , 
        \Level64Out128[26] , \Level64Out128[25] , \Level64Out128[24] , 
        \Level64Out128[23] , \Level64Out128[22] , \Level64Out128[21] , 
        \Level64Out128[20] , \Level64Out128[19] , \Level64Out128[18] , 
        \Level64Out128[17] , \Level64Out128[16] , \Level64Out128[15] , 
        \Level64Out128[14] , \Level64Out128[13] , \Level64Out128[12] , 
        \Level64Out128[11] , \Level64Out128[10] , \Level64Out128[9] , 
        \Level64Out128[8] , \Level64Out128[7] , \Level64Out128[6] , 
        \Level64Out128[5] , \Level64Out128[4] , \Level64Out128[3] , 
        \Level64Out128[2] , \Level64Out128[1] , \Level64Out128[0] }), .In1({
        \Level32Out128[31] , \Level32Out128[30] , \Level32Out128[29] , 
        \Level32Out128[28] , \Level32Out128[27] , \Level32Out128[26] , 
        \Level32Out128[25] , \Level32Out128[24] , \Level32Out128[23] , 
        \Level32Out128[22] , \Level32Out128[21] , \Level32Out128[20] , 
        \Level32Out128[19] , \Level32Out128[18] , \Level32Out128[17] , 
        \Level32Out128[16] , \Level32Out128[15] , \Level32Out128[14] , 
        \Level32Out128[13] , \Level32Out128[12] , \Level32Out128[11] , 
        \Level32Out128[10] , \Level32Out128[9] , \Level32Out128[8] , 
        \Level32Out128[7] , \Level32Out128[6] , \Level32Out128[5] , 
        \Level32Out128[4] , \Level32Out128[3] , \Level32Out128[2] , 
        \Level32Out128[1] , \Level32Out128[0] }), .In2({\Level32Out160[31] , 
        \Level32Out160[30] , \Level32Out160[29] , \Level32Out160[28] , 
        \Level32Out160[27] , \Level32Out160[26] , \Level32Out160[25] , 
        \Level32Out160[24] , \Level32Out160[23] , \Level32Out160[22] , 
        \Level32Out160[21] , \Level32Out160[20] , \Level32Out160[19] , 
        \Level32Out160[18] , \Level32Out160[17] , \Level32Out160[16] , 
        \Level32Out160[15] , \Level32Out160[14] , \Level32Out160[13] , 
        \Level32Out160[12] , \Level32Out160[11] , \Level32Out160[10] , 
        \Level32Out160[9] , \Level32Out160[8] , \Level32Out160[7] , 
        \Level32Out160[6] , \Level32Out160[5] , \Level32Out160[4] , 
        \Level32Out160[3] , \Level32Out160[2] , \Level32Out160[1] , 
        \Level32Out160[0] }), .Read1(\Level32Load128[0] ), .Read2(
        \Level32Load160[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_97 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink97[31] , \ScanLink97[30] , 
        \ScanLink97[29] , \ScanLink97[28] , \ScanLink97[27] , \ScanLink97[26] , 
        \ScanLink97[25] , \ScanLink97[24] , \ScanLink97[23] , \ScanLink97[22] , 
        \ScanLink97[21] , \ScanLink97[20] , \ScanLink97[19] , \ScanLink97[18] , 
        \ScanLink97[17] , \ScanLink97[16] , \ScanLink97[15] , \ScanLink97[14] , 
        \ScanLink97[13] , \ScanLink97[12] , \ScanLink97[11] , \ScanLink97[10] , 
        \ScanLink97[9] , \ScanLink97[8] , \ScanLink97[7] , \ScanLink97[6] , 
        \ScanLink97[5] , \ScanLink97[4] , \ScanLink97[3] , \ScanLink97[2] , 
        \ScanLink97[1] , \ScanLink97[0] }), .ScanOut({\ScanLink98[31] , 
        \ScanLink98[30] , \ScanLink98[29] , \ScanLink98[28] , \ScanLink98[27] , 
        \ScanLink98[26] , \ScanLink98[25] , \ScanLink98[24] , \ScanLink98[23] , 
        \ScanLink98[22] , \ScanLink98[21] , \ScanLink98[20] , \ScanLink98[19] , 
        \ScanLink98[18] , \ScanLink98[17] , \ScanLink98[16] , \ScanLink98[15] , 
        \ScanLink98[14] , \ScanLink98[13] , \ScanLink98[12] , \ScanLink98[11] , 
        \ScanLink98[10] , \ScanLink98[9] , \ScanLink98[8] , \ScanLink98[7] , 
        \ScanLink98[6] , \ScanLink98[5] , \ScanLink98[4] , \ScanLink98[3] , 
        \ScanLink98[2] , \ScanLink98[1] , \ScanLink98[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load97[0] ), .Out({
        \Level1Out97[31] , \Level1Out97[30] , \Level1Out97[29] , 
        \Level1Out97[28] , \Level1Out97[27] , \Level1Out97[26] , 
        \Level1Out97[25] , \Level1Out97[24] , \Level1Out97[23] , 
        \Level1Out97[22] , \Level1Out97[21] , \Level1Out97[20] , 
        \Level1Out97[19] , \Level1Out97[18] , \Level1Out97[17] , 
        \Level1Out97[16] , \Level1Out97[15] , \Level1Out97[14] , 
        \Level1Out97[13] , \Level1Out97[12] , \Level1Out97[11] , 
        \Level1Out97[10] , \Level1Out97[9] , \Level1Out97[8] , 
        \Level1Out97[7] , \Level1Out97[6] , \Level1Out97[5] , \Level1Out97[4] , 
        \Level1Out97[3] , \Level1Out97[2] , \Level1Out97[1] , \Level1Out97[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_139 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink139[31] , \ScanLink139[30] , 
        \ScanLink139[29] , \ScanLink139[28] , \ScanLink139[27] , 
        \ScanLink139[26] , \ScanLink139[25] , \ScanLink139[24] , 
        \ScanLink139[23] , \ScanLink139[22] , \ScanLink139[21] , 
        \ScanLink139[20] , \ScanLink139[19] , \ScanLink139[18] , 
        \ScanLink139[17] , \ScanLink139[16] , \ScanLink139[15] , 
        \ScanLink139[14] , \ScanLink139[13] , \ScanLink139[12] , 
        \ScanLink139[11] , \ScanLink139[10] , \ScanLink139[9] , 
        \ScanLink139[8] , \ScanLink139[7] , \ScanLink139[6] , \ScanLink139[5] , 
        \ScanLink139[4] , \ScanLink139[3] , \ScanLink139[2] , \ScanLink139[1] , 
        \ScanLink139[0] }), .ScanOut({\ScanLink140[31] , \ScanLink140[30] , 
        \ScanLink140[29] , \ScanLink140[28] , \ScanLink140[27] , 
        \ScanLink140[26] , \ScanLink140[25] , \ScanLink140[24] , 
        \ScanLink140[23] , \ScanLink140[22] , \ScanLink140[21] , 
        \ScanLink140[20] , \ScanLink140[19] , \ScanLink140[18] , 
        \ScanLink140[17] , \ScanLink140[16] , \ScanLink140[15] , 
        \ScanLink140[14] , \ScanLink140[13] , \ScanLink140[12] , 
        \ScanLink140[11] , \ScanLink140[10] , \ScanLink140[9] , 
        \ScanLink140[8] , \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , 
        \ScanLink140[4] , \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , 
        \ScanLink140[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load139[0] ), .Out({\Level1Out139[31] , \Level1Out139[30] , 
        \Level1Out139[29] , \Level1Out139[28] , \Level1Out139[27] , 
        \Level1Out139[26] , \Level1Out139[25] , \Level1Out139[24] , 
        \Level1Out139[23] , \Level1Out139[22] , \Level1Out139[21] , 
        \Level1Out139[20] , \Level1Out139[19] , \Level1Out139[18] , 
        \Level1Out139[17] , \Level1Out139[16] , \Level1Out139[15] , 
        \Level1Out139[14] , \Level1Out139[13] , \Level1Out139[12] , 
        \Level1Out139[11] , \Level1Out139[10] , \Level1Out139[9] , 
        \Level1Out139[8] , \Level1Out139[7] , \Level1Out139[6] , 
        \Level1Out139[5] , \Level1Out139[4] , \Level1Out139[3] , 
        \Level1Out139[2] , \Level1Out139[1] , \Level1Out139[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_209 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink209[31] , \ScanLink209[30] , 
        \ScanLink209[29] , \ScanLink209[28] , \ScanLink209[27] , 
        \ScanLink209[26] , \ScanLink209[25] , \ScanLink209[24] , 
        \ScanLink209[23] , \ScanLink209[22] , \ScanLink209[21] , 
        \ScanLink209[20] , \ScanLink209[19] , \ScanLink209[18] , 
        \ScanLink209[17] , \ScanLink209[16] , \ScanLink209[15] , 
        \ScanLink209[14] , \ScanLink209[13] , \ScanLink209[12] , 
        \ScanLink209[11] , \ScanLink209[10] , \ScanLink209[9] , 
        \ScanLink209[8] , \ScanLink209[7] , \ScanLink209[6] , \ScanLink209[5] , 
        \ScanLink209[4] , \ScanLink209[3] , \ScanLink209[2] , \ScanLink209[1] , 
        \ScanLink209[0] }), .ScanOut({\ScanLink210[31] , \ScanLink210[30] , 
        \ScanLink210[29] , \ScanLink210[28] , \ScanLink210[27] , 
        \ScanLink210[26] , \ScanLink210[25] , \ScanLink210[24] , 
        \ScanLink210[23] , \ScanLink210[22] , \ScanLink210[21] , 
        \ScanLink210[20] , \ScanLink210[19] , \ScanLink210[18] , 
        \ScanLink210[17] , \ScanLink210[16] , \ScanLink210[15] , 
        \ScanLink210[14] , \ScanLink210[13] , \ScanLink210[12] , 
        \ScanLink210[11] , \ScanLink210[10] , \ScanLink210[9] , 
        \ScanLink210[8] , \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , 
        \ScanLink210[4] , \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , 
        \ScanLink210[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load209[0] ), .Out({\Level1Out209[31] , \Level1Out209[30] , 
        \Level1Out209[29] , \Level1Out209[28] , \Level1Out209[27] , 
        \Level1Out209[26] , \Level1Out209[25] , \Level1Out209[24] , 
        \Level1Out209[23] , \Level1Out209[22] , \Level1Out209[21] , 
        \Level1Out209[20] , \Level1Out209[19] , \Level1Out209[18] , 
        \Level1Out209[17] , \Level1Out209[16] , \Level1Out209[15] , 
        \Level1Out209[14] , \Level1Out209[13] , \Level1Out209[12] , 
        \Level1Out209[11] , \Level1Out209[10] , \Level1Out209[9] , 
        \Level1Out209[8] , \Level1Out209[7] , \Level1Out209[6] , 
        \Level1Out209[5] , \Level1Out209[4] , \Level1Out209[3] , 
        \Level1Out209[2] , \Level1Out209[1] , \Level1Out209[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_192 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink192[31] , \ScanLink192[30] , 
        \ScanLink192[29] , \ScanLink192[28] , \ScanLink192[27] , 
        \ScanLink192[26] , \ScanLink192[25] , \ScanLink192[24] , 
        \ScanLink192[23] , \ScanLink192[22] , \ScanLink192[21] , 
        \ScanLink192[20] , \ScanLink192[19] , \ScanLink192[18] , 
        \ScanLink192[17] , \ScanLink192[16] , \ScanLink192[15] , 
        \ScanLink192[14] , \ScanLink192[13] , \ScanLink192[12] , 
        \ScanLink192[11] , \ScanLink192[10] , \ScanLink192[9] , 
        \ScanLink192[8] , \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , 
        \ScanLink192[4] , \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , 
        \ScanLink192[0] }), .ScanOut({\ScanLink193[31] , \ScanLink193[30] , 
        \ScanLink193[29] , \ScanLink193[28] , \ScanLink193[27] , 
        \ScanLink193[26] , \ScanLink193[25] , \ScanLink193[24] , 
        \ScanLink193[23] , \ScanLink193[22] , \ScanLink193[21] , 
        \ScanLink193[20] , \ScanLink193[19] , \ScanLink193[18] , 
        \ScanLink193[17] , \ScanLink193[16] , \ScanLink193[15] , 
        \ScanLink193[14] , \ScanLink193[13] , \ScanLink193[12] , 
        \ScanLink193[11] , \ScanLink193[10] , \ScanLink193[9] , 
        \ScanLink193[8] , \ScanLink193[7] , \ScanLink193[6] , \ScanLink193[5] , 
        \ScanLink193[4] , \ScanLink193[3] , \ScanLink193[2] , \ScanLink193[1] , 
        \ScanLink193[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load192[0] ), .Out({\Level1Out192[31] , \Level1Out192[30] , 
        \Level1Out192[29] , \Level1Out192[28] , \Level1Out192[27] , 
        \Level1Out192[26] , \Level1Out192[25] , \Level1Out192[24] , 
        \Level1Out192[23] , \Level1Out192[22] , \Level1Out192[21] , 
        \Level1Out192[20] , \Level1Out192[19] , \Level1Out192[18] , 
        \Level1Out192[17] , \Level1Out192[16] , \Level1Out192[15] , 
        \Level1Out192[14] , \Level1Out192[13] , \Level1Out192[12] , 
        \Level1Out192[11] , \Level1Out192[10] , \Level1Out192[9] , 
        \Level1Out192[8] , \Level1Out192[7] , \Level1Out192[6] , 
        \Level1Out192[5] , \Level1Out192[4] , \Level1Out192[3] , 
        \Level1Out192[2] , \Level1Out192[1] , \Level1Out192[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_26_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load26[0] ), .Out({\Level2Out26[31] , \Level2Out26[30] , 
        \Level2Out26[29] , \Level2Out26[28] , \Level2Out26[27] , 
        \Level2Out26[26] , \Level2Out26[25] , \Level2Out26[24] , 
        \Level2Out26[23] , \Level2Out26[22] , \Level2Out26[21] , 
        \Level2Out26[20] , \Level2Out26[19] , \Level2Out26[18] , 
        \Level2Out26[17] , \Level2Out26[16] , \Level2Out26[15] , 
        \Level2Out26[14] , \Level2Out26[13] , \Level2Out26[12] , 
        \Level2Out26[11] , \Level2Out26[10] , \Level2Out26[9] , 
        \Level2Out26[8] , \Level2Out26[7] , \Level2Out26[6] , \Level2Out26[5] , 
        \Level2Out26[4] , \Level2Out26[3] , \Level2Out26[2] , \Level2Out26[1] , 
        \Level2Out26[0] }), .In1({\Level1Out26[31] , \Level1Out26[30] , 
        \Level1Out26[29] , \Level1Out26[28] , \Level1Out26[27] , 
        \Level1Out26[26] , \Level1Out26[25] , \Level1Out26[24] , 
        \Level1Out26[23] , \Level1Out26[22] , \Level1Out26[21] , 
        \Level1Out26[20] , \Level1Out26[19] , \Level1Out26[18] , 
        \Level1Out26[17] , \Level1Out26[16] , \Level1Out26[15] , 
        \Level1Out26[14] , \Level1Out26[13] , \Level1Out26[12] , 
        \Level1Out26[11] , \Level1Out26[10] , \Level1Out26[9] , 
        \Level1Out26[8] , \Level1Out26[7] , \Level1Out26[6] , \Level1Out26[5] , 
        \Level1Out26[4] , \Level1Out26[3] , \Level1Out26[2] , \Level1Out26[1] , 
        \Level1Out26[0] }), .In2({\Level1Out27[31] , \Level1Out27[30] , 
        \Level1Out27[29] , \Level1Out27[28] , \Level1Out27[27] , 
        \Level1Out27[26] , \Level1Out27[25] , \Level1Out27[24] , 
        \Level1Out27[23] , \Level1Out27[22] , \Level1Out27[21] , 
        \Level1Out27[20] , \Level1Out27[19] , \Level1Out27[18] , 
        \Level1Out27[17] , \Level1Out27[16] , \Level1Out27[15] , 
        \Level1Out27[14] , \Level1Out27[13] , \Level1Out27[12] , 
        \Level1Out27[11] , \Level1Out27[10] , \Level1Out27[9] , 
        \Level1Out27[8] , \Level1Out27[7] , \Level1Out27[6] , \Level1Out27[5] , 
        \Level1Out27[4] , \Level1Out27[3] , \Level1Out27[2] , \Level1Out27[1] , 
        \Level1Out27[0] }), .Read1(\Level1Load26[0] ), .Read2(
        \Level1Load27[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_160_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load160[0] ), .Out({\Level2Out160[31] , \Level2Out160[30] , 
        \Level2Out160[29] , \Level2Out160[28] , \Level2Out160[27] , 
        \Level2Out160[26] , \Level2Out160[25] , \Level2Out160[24] , 
        \Level2Out160[23] , \Level2Out160[22] , \Level2Out160[21] , 
        \Level2Out160[20] , \Level2Out160[19] , \Level2Out160[18] , 
        \Level2Out160[17] , \Level2Out160[16] , \Level2Out160[15] , 
        \Level2Out160[14] , \Level2Out160[13] , \Level2Out160[12] , 
        \Level2Out160[11] , \Level2Out160[10] , \Level2Out160[9] , 
        \Level2Out160[8] , \Level2Out160[7] , \Level2Out160[6] , 
        \Level2Out160[5] , \Level2Out160[4] , \Level2Out160[3] , 
        \Level2Out160[2] , \Level2Out160[1] , \Level2Out160[0] }), .In1({
        \Level1Out160[31] , \Level1Out160[30] , \Level1Out160[29] , 
        \Level1Out160[28] , \Level1Out160[27] , \Level1Out160[26] , 
        \Level1Out160[25] , \Level1Out160[24] , \Level1Out160[23] , 
        \Level1Out160[22] , \Level1Out160[21] , \Level1Out160[20] , 
        \Level1Out160[19] , \Level1Out160[18] , \Level1Out160[17] , 
        \Level1Out160[16] , \Level1Out160[15] , \Level1Out160[14] , 
        \Level1Out160[13] , \Level1Out160[12] , \Level1Out160[11] , 
        \Level1Out160[10] , \Level1Out160[9] , \Level1Out160[8] , 
        \Level1Out160[7] , \Level1Out160[6] , \Level1Out160[5] , 
        \Level1Out160[4] , \Level1Out160[3] , \Level1Out160[2] , 
        \Level1Out160[1] , \Level1Out160[0] }), .In2({\Level1Out161[31] , 
        \Level1Out161[30] , \Level1Out161[29] , \Level1Out161[28] , 
        \Level1Out161[27] , \Level1Out161[26] , \Level1Out161[25] , 
        \Level1Out161[24] , \Level1Out161[23] , \Level1Out161[22] , 
        \Level1Out161[21] , \Level1Out161[20] , \Level1Out161[19] , 
        \Level1Out161[18] , \Level1Out161[17] , \Level1Out161[16] , 
        \Level1Out161[15] , \Level1Out161[14] , \Level1Out161[13] , 
        \Level1Out161[12] , \Level1Out161[11] , \Level1Out161[10] , 
        \Level1Out161[9] , \Level1Out161[8] , \Level1Out161[7] , 
        \Level1Out161[6] , \Level1Out161[5] , \Level1Out161[4] , 
        \Level1Out161[3] , \Level1Out161[2] , \Level1Out161[1] , 
        \Level1Out161[0] }), .Read1(\Level1Load160[0] ), .Read2(
        \Level1Load161[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_254_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load254[0] ), .Out({\Level2Out254[31] , \Level2Out254[30] , 
        \Level2Out254[29] , \Level2Out254[28] , \Level2Out254[27] , 
        \Level2Out254[26] , \Level2Out254[25] , \Level2Out254[24] , 
        \Level2Out254[23] , \Level2Out254[22] , \Level2Out254[21] , 
        \Level2Out254[20] , \Level2Out254[19] , \Level2Out254[18] , 
        \Level2Out254[17] , \Level2Out254[16] , \Level2Out254[15] , 
        \Level2Out254[14] , \Level2Out254[13] , \Level2Out254[12] , 
        \Level2Out254[11] , \Level2Out254[10] , \Level2Out254[9] , 
        \Level2Out254[8] , \Level2Out254[7] , \Level2Out254[6] , 
        \Level2Out254[5] , \Level2Out254[4] , \Level2Out254[3] , 
        \Level2Out254[2] , \Level2Out254[1] , \Level2Out254[0] }), .In1({
        \Level1Out254[31] , \Level1Out254[30] , \Level1Out254[29] , 
        \Level1Out254[28] , \Level1Out254[27] , \Level1Out254[26] , 
        \Level1Out254[25] , \Level1Out254[24] , \Level1Out254[23] , 
        \Level1Out254[22] , \Level1Out254[21] , \Level1Out254[20] , 
        \Level1Out254[19] , \Level1Out254[18] , \Level1Out254[17] , 
        \Level1Out254[16] , \Level1Out254[15] , \Level1Out254[14] , 
        \Level1Out254[13] , \Level1Out254[12] , \Level1Out254[11] , 
        \Level1Out254[10] , \Level1Out254[9] , \Level1Out254[8] , 
        \Level1Out254[7] , \Level1Out254[6] , \Level1Out254[5] , 
        \Level1Out254[4] , \Level1Out254[3] , \Level1Out254[2] , 
        \Level1Out254[1] , \Level1Out254[0] }), .In2({\Level1Out255[31] , 
        \Level1Out255[30] , \Level1Out255[29] , \Level1Out255[28] , 
        \Level1Out255[27] , \Level1Out255[26] , \Level1Out255[25] , 
        \Level1Out255[24] , \Level1Out255[23] , \Level1Out255[22] , 
        \Level1Out255[21] , \Level1Out255[20] , \Level1Out255[19] , 
        \Level1Out255[18] , \Level1Out255[17] , \Level1Out255[16] , 
        \Level1Out255[15] , \Level1Out255[14] , \Level1Out255[13] , 
        \Level1Out255[12] , \Level1Out255[11] , \Level1Out255[10] , 
        \Level1Out255[9] , \Level1Out255[8] , \Level1Out255[7] , 
        \Level1Out255[6] , \Level1Out255[5] , \Level1Out255[4] , 
        \Level1Out255[3] , \Level1Out255[2] , \Level1Out255[1] , 
        \Level1Out255[0] }), .Read1(\Level1Load254[0] ), .Read2(
        \Level1Load255[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_156_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load156[0] ), .Out({\Level4Out156[31] , \Level4Out156[30] , 
        \Level4Out156[29] , \Level4Out156[28] , \Level4Out156[27] , 
        \Level4Out156[26] , \Level4Out156[25] , \Level4Out156[24] , 
        \Level4Out156[23] , \Level4Out156[22] , \Level4Out156[21] , 
        \Level4Out156[20] , \Level4Out156[19] , \Level4Out156[18] , 
        \Level4Out156[17] , \Level4Out156[16] , \Level4Out156[15] , 
        \Level4Out156[14] , \Level4Out156[13] , \Level4Out156[12] , 
        \Level4Out156[11] , \Level4Out156[10] , \Level4Out156[9] , 
        \Level4Out156[8] , \Level4Out156[7] , \Level4Out156[6] , 
        \Level4Out156[5] , \Level4Out156[4] , \Level4Out156[3] , 
        \Level4Out156[2] , \Level4Out156[1] , \Level4Out156[0] }), .In1({
        \Level2Out156[31] , \Level2Out156[30] , \Level2Out156[29] , 
        \Level2Out156[28] , \Level2Out156[27] , \Level2Out156[26] , 
        \Level2Out156[25] , \Level2Out156[24] , \Level2Out156[23] , 
        \Level2Out156[22] , \Level2Out156[21] , \Level2Out156[20] , 
        \Level2Out156[19] , \Level2Out156[18] , \Level2Out156[17] , 
        \Level2Out156[16] , \Level2Out156[15] , \Level2Out156[14] , 
        \Level2Out156[13] , \Level2Out156[12] , \Level2Out156[11] , 
        \Level2Out156[10] , \Level2Out156[9] , \Level2Out156[8] , 
        \Level2Out156[7] , \Level2Out156[6] , \Level2Out156[5] , 
        \Level2Out156[4] , \Level2Out156[3] , \Level2Out156[2] , 
        \Level2Out156[1] , \Level2Out156[0] }), .In2({\Level2Out158[31] , 
        \Level2Out158[30] , \Level2Out158[29] , \Level2Out158[28] , 
        \Level2Out158[27] , \Level2Out158[26] , \Level2Out158[25] , 
        \Level2Out158[24] , \Level2Out158[23] , \Level2Out158[22] , 
        \Level2Out158[21] , \Level2Out158[20] , \Level2Out158[19] , 
        \Level2Out158[18] , \Level2Out158[17] , \Level2Out158[16] , 
        \Level2Out158[15] , \Level2Out158[14] , \Level2Out158[13] , 
        \Level2Out158[12] , \Level2Out158[11] , \Level2Out158[10] , 
        \Level2Out158[9] , \Level2Out158[8] , \Level2Out158[7] , 
        \Level2Out158[6] , \Level2Out158[5] , \Level2Out158[4] , 
        \Level2Out158[3] , \Level2Out158[2] , \Level2Out158[1] , 
        \Level2Out158[0] }), .Read1(\Level2Load156[0] ), .Read2(
        \Level2Load158[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_248_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load248[0] ), .Out({\Level4Out248[31] , \Level4Out248[30] , 
        \Level4Out248[29] , \Level4Out248[28] , \Level4Out248[27] , 
        \Level4Out248[26] , \Level4Out248[25] , \Level4Out248[24] , 
        \Level4Out248[23] , \Level4Out248[22] , \Level4Out248[21] , 
        \Level4Out248[20] , \Level4Out248[19] , \Level4Out248[18] , 
        \Level4Out248[17] , \Level4Out248[16] , \Level4Out248[15] , 
        \Level4Out248[14] , \Level4Out248[13] , \Level4Out248[12] , 
        \Level4Out248[11] , \Level4Out248[10] , \Level4Out248[9] , 
        \Level4Out248[8] , \Level4Out248[7] , \Level4Out248[6] , 
        \Level4Out248[5] , \Level4Out248[4] , \Level4Out248[3] , 
        \Level4Out248[2] , \Level4Out248[1] , \Level4Out248[0] }), .In1({
        \Level2Out248[31] , \Level2Out248[30] , \Level2Out248[29] , 
        \Level2Out248[28] , \Level2Out248[27] , \Level2Out248[26] , 
        \Level2Out248[25] , \Level2Out248[24] , \Level2Out248[23] , 
        \Level2Out248[22] , \Level2Out248[21] , \Level2Out248[20] , 
        \Level2Out248[19] , \Level2Out248[18] , \Level2Out248[17] , 
        \Level2Out248[16] , \Level2Out248[15] , \Level2Out248[14] , 
        \Level2Out248[13] , \Level2Out248[12] , \Level2Out248[11] , 
        \Level2Out248[10] , \Level2Out248[9] , \Level2Out248[8] , 
        \Level2Out248[7] , \Level2Out248[6] , \Level2Out248[5] , 
        \Level2Out248[4] , \Level2Out248[3] , \Level2Out248[2] , 
        \Level2Out248[1] , \Level2Out248[0] }), .In2({\Level2Out250[31] , 
        \Level2Out250[30] , \Level2Out250[29] , \Level2Out250[28] , 
        \Level2Out250[27] , \Level2Out250[26] , \Level2Out250[25] , 
        \Level2Out250[24] , \Level2Out250[23] , \Level2Out250[22] , 
        \Level2Out250[21] , \Level2Out250[20] , \Level2Out250[19] , 
        \Level2Out250[18] , \Level2Out250[17] , \Level2Out250[16] , 
        \Level2Out250[15] , \Level2Out250[14] , \Level2Out250[13] , 
        \Level2Out250[12] , \Level2Out250[11] , \Level2Out250[10] , 
        \Level2Out250[9] , \Level2Out250[8] , \Level2Out250[7] , 
        \Level2Out250[6] , \Level2Out250[5] , \Level2Out250[4] , 
        \Level2Out250[3] , \Level2Out250[2] , \Level2Out250[1] , 
        \Level2Out250[0] }), .Read1(\Level2Load248[0] ), .Read2(
        \Level2Load250[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_229 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink229[31] , \ScanLink229[30] , 
        \ScanLink229[29] , \ScanLink229[28] , \ScanLink229[27] , 
        \ScanLink229[26] , \ScanLink229[25] , \ScanLink229[24] , 
        \ScanLink229[23] , \ScanLink229[22] , \ScanLink229[21] , 
        \ScanLink229[20] , \ScanLink229[19] , \ScanLink229[18] , 
        \ScanLink229[17] , \ScanLink229[16] , \ScanLink229[15] , 
        \ScanLink229[14] , \ScanLink229[13] , \ScanLink229[12] , 
        \ScanLink229[11] , \ScanLink229[10] , \ScanLink229[9] , 
        \ScanLink229[8] , \ScanLink229[7] , \ScanLink229[6] , \ScanLink229[5] , 
        \ScanLink229[4] , \ScanLink229[3] , \ScanLink229[2] , \ScanLink229[1] , 
        \ScanLink229[0] }), .ScanOut({\ScanLink230[31] , \ScanLink230[30] , 
        \ScanLink230[29] , \ScanLink230[28] , \ScanLink230[27] , 
        \ScanLink230[26] , \ScanLink230[25] , \ScanLink230[24] , 
        \ScanLink230[23] , \ScanLink230[22] , \ScanLink230[21] , 
        \ScanLink230[20] , \ScanLink230[19] , \ScanLink230[18] , 
        \ScanLink230[17] , \ScanLink230[16] , \ScanLink230[15] , 
        \ScanLink230[14] , \ScanLink230[13] , \ScanLink230[12] , 
        \ScanLink230[11] , \ScanLink230[10] , \ScanLink230[9] , 
        \ScanLink230[8] , \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , 
        \ScanLink230[4] , \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , 
        \ScanLink230[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load229[0] ), .Out({\Level1Out229[31] , \Level1Out229[30] , 
        \Level1Out229[29] , \Level1Out229[28] , \Level1Out229[27] , 
        \Level1Out229[26] , \Level1Out229[25] , \Level1Out229[24] , 
        \Level1Out229[23] , \Level1Out229[22] , \Level1Out229[21] , 
        \Level1Out229[20] , \Level1Out229[19] , \Level1Out229[18] , 
        \Level1Out229[17] , \Level1Out229[16] , \Level1Out229[15] , 
        \Level1Out229[14] , \Level1Out229[13] , \Level1Out229[12] , 
        \Level1Out229[11] , \Level1Out229[10] , \Level1Out229[9] , 
        \Level1Out229[8] , \Level1Out229[7] , \Level1Out229[6] , 
        \Level1Out229[5] , \Level1Out229[4] , \Level1Out229[3] , 
        \Level1Out229[2] , \Level1Out229[1] , \Level1Out229[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_224_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load224[0] ), .Out({\Level16Out224[31] , \Level16Out224[30] , 
        \Level16Out224[29] , \Level16Out224[28] , \Level16Out224[27] , 
        \Level16Out224[26] , \Level16Out224[25] , \Level16Out224[24] , 
        \Level16Out224[23] , \Level16Out224[22] , \Level16Out224[21] , 
        \Level16Out224[20] , \Level16Out224[19] , \Level16Out224[18] , 
        \Level16Out224[17] , \Level16Out224[16] , \Level16Out224[15] , 
        \Level16Out224[14] , \Level16Out224[13] , \Level16Out224[12] , 
        \Level16Out224[11] , \Level16Out224[10] , \Level16Out224[9] , 
        \Level16Out224[8] , \Level16Out224[7] , \Level16Out224[6] , 
        \Level16Out224[5] , \Level16Out224[4] , \Level16Out224[3] , 
        \Level16Out224[2] , \Level16Out224[1] , \Level16Out224[0] }), .In1({
        \Level8Out224[31] , \Level8Out224[30] , \Level8Out224[29] , 
        \Level8Out224[28] , \Level8Out224[27] , \Level8Out224[26] , 
        \Level8Out224[25] , \Level8Out224[24] , \Level8Out224[23] , 
        \Level8Out224[22] , \Level8Out224[21] , \Level8Out224[20] , 
        \Level8Out224[19] , \Level8Out224[18] , \Level8Out224[17] , 
        \Level8Out224[16] , \Level8Out224[15] , \Level8Out224[14] , 
        \Level8Out224[13] , \Level8Out224[12] , \Level8Out224[11] , 
        \Level8Out224[10] , \Level8Out224[9] , \Level8Out224[8] , 
        \Level8Out224[7] , \Level8Out224[6] , \Level8Out224[5] , 
        \Level8Out224[4] , \Level8Out224[3] , \Level8Out224[2] , 
        \Level8Out224[1] , \Level8Out224[0] }), .In2({\Level8Out232[31] , 
        \Level8Out232[30] , \Level8Out232[29] , \Level8Out232[28] , 
        \Level8Out232[27] , \Level8Out232[26] , \Level8Out232[25] , 
        \Level8Out232[24] , \Level8Out232[23] , \Level8Out232[22] , 
        \Level8Out232[21] , \Level8Out232[20] , \Level8Out232[19] , 
        \Level8Out232[18] , \Level8Out232[17] , \Level8Out232[16] , 
        \Level8Out232[15] , \Level8Out232[14] , \Level8Out232[13] , 
        \Level8Out232[12] , \Level8Out232[11] , \Level8Out232[10] , 
        \Level8Out232[9] , \Level8Out232[8] , \Level8Out232[7] , 
        \Level8Out232[6] , \Level8Out232[5] , \Level8Out232[4] , 
        \Level8Out232[3] , \Level8Out232[2] , \Level8Out232[1] , 
        \Level8Out232[0] }), .Read1(\Level8Load224[0] ), .Read2(
        \Level8Load232[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_119 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink119[31] , \ScanLink119[30] , 
        \ScanLink119[29] , \ScanLink119[28] , \ScanLink119[27] , 
        \ScanLink119[26] , \ScanLink119[25] , \ScanLink119[24] , 
        \ScanLink119[23] , \ScanLink119[22] , \ScanLink119[21] , 
        \ScanLink119[20] , \ScanLink119[19] , \ScanLink119[18] , 
        \ScanLink119[17] , \ScanLink119[16] , \ScanLink119[15] , 
        \ScanLink119[14] , \ScanLink119[13] , \ScanLink119[12] , 
        \ScanLink119[11] , \ScanLink119[10] , \ScanLink119[9] , 
        \ScanLink119[8] , \ScanLink119[7] , \ScanLink119[6] , \ScanLink119[5] , 
        \ScanLink119[4] , \ScanLink119[3] , \ScanLink119[2] , \ScanLink119[1] , 
        \ScanLink119[0] }), .ScanOut({\ScanLink120[31] , \ScanLink120[30] , 
        \ScanLink120[29] , \ScanLink120[28] , \ScanLink120[27] , 
        \ScanLink120[26] , \ScanLink120[25] , \ScanLink120[24] , 
        \ScanLink120[23] , \ScanLink120[22] , \ScanLink120[21] , 
        \ScanLink120[20] , \ScanLink120[19] , \ScanLink120[18] , 
        \ScanLink120[17] , \ScanLink120[16] , \ScanLink120[15] , 
        \ScanLink120[14] , \ScanLink120[13] , \ScanLink120[12] , 
        \ScanLink120[11] , \ScanLink120[10] , \ScanLink120[9] , 
        \ScanLink120[8] , \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , 
        \ScanLink120[4] , \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , 
        \ScanLink120[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load119[0] ), .Out({\Level1Out119[31] , \Level1Out119[30] , 
        \Level1Out119[29] , \Level1Out119[28] , \Level1Out119[27] , 
        \Level1Out119[26] , \Level1Out119[25] , \Level1Out119[24] , 
        \Level1Out119[23] , \Level1Out119[22] , \Level1Out119[21] , 
        \Level1Out119[20] , \Level1Out119[19] , \Level1Out119[18] , 
        \Level1Out119[17] , \Level1Out119[16] , \Level1Out119[15] , 
        \Level1Out119[14] , \Level1Out119[13] , \Level1Out119[12] , 
        \Level1Out119[11] , \Level1Out119[10] , \Level1Out119[9] , 
        \Level1Out119[8] , \Level1Out119[7] , \Level1Out119[6] , 
        \Level1Out119[5] , \Level1Out119[4] , \Level1Out119[3] , 
        \Level1Out119[2] , \Level1Out119[1] , \Level1Out119[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_150 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink150[31] , \ScanLink150[30] , 
        \ScanLink150[29] , \ScanLink150[28] , \ScanLink150[27] , 
        \ScanLink150[26] , \ScanLink150[25] , \ScanLink150[24] , 
        \ScanLink150[23] , \ScanLink150[22] , \ScanLink150[21] , 
        \ScanLink150[20] , \ScanLink150[19] , \ScanLink150[18] , 
        \ScanLink150[17] , \ScanLink150[16] , \ScanLink150[15] , 
        \ScanLink150[14] , \ScanLink150[13] , \ScanLink150[12] , 
        \ScanLink150[11] , \ScanLink150[10] , \ScanLink150[9] , 
        \ScanLink150[8] , \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , 
        \ScanLink150[4] , \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , 
        \ScanLink150[0] }), .ScanOut({\ScanLink151[31] , \ScanLink151[30] , 
        \ScanLink151[29] , \ScanLink151[28] , \ScanLink151[27] , 
        \ScanLink151[26] , \ScanLink151[25] , \ScanLink151[24] , 
        \ScanLink151[23] , \ScanLink151[22] , \ScanLink151[21] , 
        \ScanLink151[20] , \ScanLink151[19] , \ScanLink151[18] , 
        \ScanLink151[17] , \ScanLink151[16] , \ScanLink151[15] , 
        \ScanLink151[14] , \ScanLink151[13] , \ScanLink151[12] , 
        \ScanLink151[11] , \ScanLink151[10] , \ScanLink151[9] , 
        \ScanLink151[8] , \ScanLink151[7] , \ScanLink151[6] , \ScanLink151[5] , 
        \ScanLink151[4] , \ScanLink151[3] , \ScanLink151[2] , \ScanLink151[1] , 
        \ScanLink151[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load150[0] ), .Out({\Level1Out150[31] , \Level1Out150[30] , 
        \Level1Out150[29] , \Level1Out150[28] , \Level1Out150[27] , 
        \Level1Out150[26] , \Level1Out150[25] , \Level1Out150[24] , 
        \Level1Out150[23] , \Level1Out150[22] , \Level1Out150[21] , 
        \Level1Out150[20] , \Level1Out150[19] , \Level1Out150[18] , 
        \Level1Out150[17] , \Level1Out150[16] , \Level1Out150[15] , 
        \Level1Out150[14] , \Level1Out150[13] , \Level1Out150[12] , 
        \Level1Out150[11] , \Level1Out150[10] , \Level1Out150[9] , 
        \Level1Out150[8] , \Level1Out150[7] , \Level1Out150[6] , 
        \Level1Out150[5] , \Level1Out150[4] , \Level1Out150[3] , 
        \Level1Out150[2] , \Level1Out150[1] , \Level1Out150[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_177 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink177[31] , \ScanLink177[30] , 
        \ScanLink177[29] , \ScanLink177[28] , \ScanLink177[27] , 
        \ScanLink177[26] , \ScanLink177[25] , \ScanLink177[24] , 
        \ScanLink177[23] , \ScanLink177[22] , \ScanLink177[21] , 
        \ScanLink177[20] , \ScanLink177[19] , \ScanLink177[18] , 
        \ScanLink177[17] , \ScanLink177[16] , \ScanLink177[15] , 
        \ScanLink177[14] , \ScanLink177[13] , \ScanLink177[12] , 
        \ScanLink177[11] , \ScanLink177[10] , \ScanLink177[9] , 
        \ScanLink177[8] , \ScanLink177[7] , \ScanLink177[6] , \ScanLink177[5] , 
        \ScanLink177[4] , \ScanLink177[3] , \ScanLink177[2] , \ScanLink177[1] , 
        \ScanLink177[0] }), .ScanOut({\ScanLink178[31] , \ScanLink178[30] , 
        \ScanLink178[29] , \ScanLink178[28] , \ScanLink178[27] , 
        \ScanLink178[26] , \ScanLink178[25] , \ScanLink178[24] , 
        \ScanLink178[23] , \ScanLink178[22] , \ScanLink178[21] , 
        \ScanLink178[20] , \ScanLink178[19] , \ScanLink178[18] , 
        \ScanLink178[17] , \ScanLink178[16] , \ScanLink178[15] , 
        \ScanLink178[14] , \ScanLink178[13] , \ScanLink178[12] , 
        \ScanLink178[11] , \ScanLink178[10] , \ScanLink178[9] , 
        \ScanLink178[8] , \ScanLink178[7] , \ScanLink178[6] , \ScanLink178[5] , 
        \ScanLink178[4] , \ScanLink178[3] , \ScanLink178[2] , \ScanLink178[1] , 
        \ScanLink178[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load177[0] ), .Out({\Level1Out177[31] , \Level1Out177[30] , 
        \Level1Out177[29] , \Level1Out177[28] , \Level1Out177[27] , 
        \Level1Out177[26] , \Level1Out177[25] , \Level1Out177[24] , 
        \Level1Out177[23] , \Level1Out177[22] , \Level1Out177[21] , 
        \Level1Out177[20] , \Level1Out177[19] , \Level1Out177[18] , 
        \Level1Out177[17] , \Level1Out177[16] , \Level1Out177[15] , 
        \Level1Out177[14] , \Level1Out177[13] , \Level1Out177[12] , 
        \Level1Out177[11] , \Level1Out177[10] , \Level1Out177[9] , 
        \Level1Out177[8] , \Level1Out177[7] , \Level1Out177[6] , 
        \Level1Out177[5] , \Level1Out177[4] , \Level1Out177[3] , 
        \Level1Out177[2] , \Level1Out177[1] , \Level1Out177[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_247 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink247[31] , \ScanLink247[30] , 
        \ScanLink247[29] , \ScanLink247[28] , \ScanLink247[27] , 
        \ScanLink247[26] , \ScanLink247[25] , \ScanLink247[24] , 
        \ScanLink247[23] , \ScanLink247[22] , \ScanLink247[21] , 
        \ScanLink247[20] , \ScanLink247[19] , \ScanLink247[18] , 
        \ScanLink247[17] , \ScanLink247[16] , \ScanLink247[15] , 
        \ScanLink247[14] , \ScanLink247[13] , \ScanLink247[12] , 
        \ScanLink247[11] , \ScanLink247[10] , \ScanLink247[9] , 
        \ScanLink247[8] , \ScanLink247[7] , \ScanLink247[6] , \ScanLink247[5] , 
        \ScanLink247[4] , \ScanLink247[3] , \ScanLink247[2] , \ScanLink247[1] , 
        \ScanLink247[0] }), .ScanOut({\ScanLink248[31] , \ScanLink248[30] , 
        \ScanLink248[29] , \ScanLink248[28] , \ScanLink248[27] , 
        \ScanLink248[26] , \ScanLink248[25] , \ScanLink248[24] , 
        \ScanLink248[23] , \ScanLink248[22] , \ScanLink248[21] , 
        \ScanLink248[20] , \ScanLink248[19] , \ScanLink248[18] , 
        \ScanLink248[17] , \ScanLink248[16] , \ScanLink248[15] , 
        \ScanLink248[14] , \ScanLink248[13] , \ScanLink248[12] , 
        \ScanLink248[11] , \ScanLink248[10] , \ScanLink248[9] , 
        \ScanLink248[8] , \ScanLink248[7] , \ScanLink248[6] , \ScanLink248[5] , 
        \ScanLink248[4] , \ScanLink248[3] , \ScanLink248[2] , \ScanLink248[1] , 
        \ScanLink248[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load247[0] ), .Out({\Level1Out247[31] , \Level1Out247[30] , 
        \Level1Out247[29] , \Level1Out247[28] , \Level1Out247[27] , 
        \Level1Out247[26] , \Level1Out247[25] , \Level1Out247[24] , 
        \Level1Out247[23] , \Level1Out247[22] , \Level1Out247[21] , 
        \Level1Out247[20] , \Level1Out247[19] , \Level1Out247[18] , 
        \Level1Out247[17] , \Level1Out247[16] , \Level1Out247[15] , 
        \Level1Out247[14] , \Level1Out247[13] , \Level1Out247[12] , 
        \Level1Out247[11] , \Level1Out247[10] , \Level1Out247[9] , 
        \Level1Out247[8] , \Level1Out247[7] , \Level1Out247[6] , 
        \Level1Out247[5] , \Level1Out247[4] , \Level1Out247[3] , 
        \Level1Out247[2] , \Level1Out247[1] , \Level1Out247[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_69 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink69[31] , \ScanLink69[30] , 
        \ScanLink69[29] , \ScanLink69[28] , \ScanLink69[27] , \ScanLink69[26] , 
        \ScanLink69[25] , \ScanLink69[24] , \ScanLink69[23] , \ScanLink69[22] , 
        \ScanLink69[21] , \ScanLink69[20] , \ScanLink69[19] , \ScanLink69[18] , 
        \ScanLink69[17] , \ScanLink69[16] , \ScanLink69[15] , \ScanLink69[14] , 
        \ScanLink69[13] , \ScanLink69[12] , \ScanLink69[11] , \ScanLink69[10] , 
        \ScanLink69[9] , \ScanLink69[8] , \ScanLink69[7] , \ScanLink69[6] , 
        \ScanLink69[5] , \ScanLink69[4] , \ScanLink69[3] , \ScanLink69[2] , 
        \ScanLink69[1] , \ScanLink69[0] }), .ScanOut({\ScanLink70[31] , 
        \ScanLink70[30] , \ScanLink70[29] , \ScanLink70[28] , \ScanLink70[27] , 
        \ScanLink70[26] , \ScanLink70[25] , \ScanLink70[24] , \ScanLink70[23] , 
        \ScanLink70[22] , \ScanLink70[21] , \ScanLink70[20] , \ScanLink70[19] , 
        \ScanLink70[18] , \ScanLink70[17] , \ScanLink70[16] , \ScanLink70[15] , 
        \ScanLink70[14] , \ScanLink70[13] , \ScanLink70[12] , \ScanLink70[11] , 
        \ScanLink70[10] , \ScanLink70[9] , \ScanLink70[8] , \ScanLink70[7] , 
        \ScanLink70[6] , \ScanLink70[5] , \ScanLink70[4] , \ScanLink70[3] , 
        \ScanLink70[2] , \ScanLink70[1] , \ScanLink70[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load69[0] ), .Out({
        \Level1Out69[31] , \Level1Out69[30] , \Level1Out69[29] , 
        \Level1Out69[28] , \Level1Out69[27] , \Level1Out69[26] , 
        \Level1Out69[25] , \Level1Out69[24] , \Level1Out69[23] , 
        \Level1Out69[22] , \Level1Out69[21] , \Level1Out69[20] , 
        \Level1Out69[19] , \Level1Out69[18] , \Level1Out69[17] , 
        \Level1Out69[16] , \Level1Out69[15] , \Level1Out69[14] , 
        \Level1Out69[13] , \Level1Out69[12] , \Level1Out69[11] , 
        \Level1Out69[10] , \Level1Out69[9] , \Level1Out69[8] , 
        \Level1Out69[7] , \Level1Out69[6] , \Level1Out69[5] , \Level1Out69[4] , 
        \Level1Out69[3] , \Level1Out69[2] , \Level1Out69[1] , \Level1Out69[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load128[0] ), .Out({\Level16Out128[31] , \Level16Out128[30] , 
        \Level16Out128[29] , \Level16Out128[28] , \Level16Out128[27] , 
        \Level16Out128[26] , \Level16Out128[25] , \Level16Out128[24] , 
        \Level16Out128[23] , \Level16Out128[22] , \Level16Out128[21] , 
        \Level16Out128[20] , \Level16Out128[19] , \Level16Out128[18] , 
        \Level16Out128[17] , \Level16Out128[16] , \Level16Out128[15] , 
        \Level16Out128[14] , \Level16Out128[13] , \Level16Out128[12] , 
        \Level16Out128[11] , \Level16Out128[10] , \Level16Out128[9] , 
        \Level16Out128[8] , \Level16Out128[7] , \Level16Out128[6] , 
        \Level16Out128[5] , \Level16Out128[4] , \Level16Out128[3] , 
        \Level16Out128[2] , \Level16Out128[1] , \Level16Out128[0] }), .In1({
        \Level8Out128[31] , \Level8Out128[30] , \Level8Out128[29] , 
        \Level8Out128[28] , \Level8Out128[27] , \Level8Out128[26] , 
        \Level8Out128[25] , \Level8Out128[24] , \Level8Out128[23] , 
        \Level8Out128[22] , \Level8Out128[21] , \Level8Out128[20] , 
        \Level8Out128[19] , \Level8Out128[18] , \Level8Out128[17] , 
        \Level8Out128[16] , \Level8Out128[15] , \Level8Out128[14] , 
        \Level8Out128[13] , \Level8Out128[12] , \Level8Out128[11] , 
        \Level8Out128[10] , \Level8Out128[9] , \Level8Out128[8] , 
        \Level8Out128[7] , \Level8Out128[6] , \Level8Out128[5] , 
        \Level8Out128[4] , \Level8Out128[3] , \Level8Out128[2] , 
        \Level8Out128[1] , \Level8Out128[0] }), .In2({\Level8Out136[31] , 
        \Level8Out136[30] , \Level8Out136[29] , \Level8Out136[28] , 
        \Level8Out136[27] , \Level8Out136[26] , \Level8Out136[25] , 
        \Level8Out136[24] , \Level8Out136[23] , \Level8Out136[22] , 
        \Level8Out136[21] , \Level8Out136[20] , \Level8Out136[19] , 
        \Level8Out136[18] , \Level8Out136[17] , \Level8Out136[16] , 
        \Level8Out136[15] , \Level8Out136[14] , \Level8Out136[13] , 
        \Level8Out136[12] , \Level8Out136[11] , \Level8Out136[10] , 
        \Level8Out136[9] , \Level8Out136[8] , \Level8Out136[7] , 
        \Level8Out136[6] , \Level8Out136[5] , \Level8Out136[4] , 
        \Level8Out136[3] , \Level8Out136[2] , \Level8Out136[1] , 
        \Level8Out136[0] }), .Read1(\Level8Load128[0] ), .Read2(
        \Level8Load136[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanOut({\ScanLink10[31] , 
        \ScanLink10[30] , \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , 
        \ScanLink10[26] , \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , 
        \ScanLink10[22] , \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , 
        \ScanLink10[18] , \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , 
        \ScanLink10[14] , \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , 
        \ScanLink10[10] , \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , 
        \ScanLink10[6] , \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , 
        \ScanLink10[2] , \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load9[0] ), .Out({
        \Level1Out9[31] , \Level1Out9[30] , \Level1Out9[29] , \Level1Out9[28] , 
        \Level1Out9[27] , \Level1Out9[26] , \Level1Out9[25] , \Level1Out9[24] , 
        \Level1Out9[23] , \Level1Out9[22] , \Level1Out9[21] , \Level1Out9[20] , 
        \Level1Out9[19] , \Level1Out9[18] , \Level1Out9[17] , \Level1Out9[16] , 
        \Level1Out9[15] , \Level1Out9[14] , \Level1Out9[13] , \Level1Out9[12] , 
        \Level1Out9[11] , \Level1Out9[10] , \Level1Out9[9] , \Level1Out9[8] , 
        \Level1Out9[7] , \Level1Out9[6] , \Level1Out9[5] , \Level1Out9[4] , 
        \Level1Out9[3] , \Level1Out9[2] , \Level1Out9[1] , \Level1Out9[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanOut({\ScanLink16[31] , 
        \ScanLink16[30] , \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , 
        \ScanLink16[26] , \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , 
        \ScanLink16[22] , \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , 
        \ScanLink16[18] , \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , 
        \ScanLink16[14] , \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , 
        \ScanLink16[10] , \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , 
        \ScanLink16[6] , \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , 
        \ScanLink16[2] , \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load15[0] ), .Out({
        \Level1Out15[31] , \Level1Out15[30] , \Level1Out15[29] , 
        \Level1Out15[28] , \Level1Out15[27] , \Level1Out15[26] , 
        \Level1Out15[25] , \Level1Out15[24] , \Level1Out15[23] , 
        \Level1Out15[22] , \Level1Out15[21] , \Level1Out15[20] , 
        \Level1Out15[19] , \Level1Out15[18] , \Level1Out15[17] , 
        \Level1Out15[16] , \Level1Out15[15] , \Level1Out15[14] , 
        \Level1Out15[13] , \Level1Out15[12] , \Level1Out15[11] , 
        \Level1Out15[10] , \Level1Out15[9] , \Level1Out15[8] , 
        \Level1Out15[7] , \Level1Out15[6] , \Level1Out15[5] , \Level1Out15[4] , 
        \Level1Out15[3] , \Level1Out15[2] , \Level1Out15[1] , \Level1Out15[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_20 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanOut({\ScanLink21[31] , 
        \ScanLink21[30] , \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , 
        \ScanLink21[26] , \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , 
        \ScanLink21[22] , \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , 
        \ScanLink21[18] , \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , 
        \ScanLink21[14] , \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , 
        \ScanLink21[10] , \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , 
        \ScanLink21[6] , \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , 
        \ScanLink21[2] , \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load20[0] ), .Out({
        \Level1Out20[31] , \Level1Out20[30] , \Level1Out20[29] , 
        \Level1Out20[28] , \Level1Out20[27] , \Level1Out20[26] , 
        \Level1Out20[25] , \Level1Out20[24] , \Level1Out20[23] , 
        \Level1Out20[22] , \Level1Out20[21] , \Level1Out20[20] , 
        \Level1Out20[19] , \Level1Out20[18] , \Level1Out20[17] , 
        \Level1Out20[16] , \Level1Out20[15] , \Level1Out20[14] , 
        \Level1Out20[13] , \Level1Out20[12] , \Level1Out20[11] , 
        \Level1Out20[10] , \Level1Out20[9] , \Level1Out20[8] , 
        \Level1Out20[7] , \Level1Out20[6] , \Level1Out20[5] , \Level1Out20[4] , 
        \Level1Out20[3] , \Level1Out20[2] , \Level1Out20[1] , \Level1Out20[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_102 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink102[31] , \ScanLink102[30] , 
        \ScanLink102[29] , \ScanLink102[28] , \ScanLink102[27] , 
        \ScanLink102[26] , \ScanLink102[25] , \ScanLink102[24] , 
        \ScanLink102[23] , \ScanLink102[22] , \ScanLink102[21] , 
        \ScanLink102[20] , \ScanLink102[19] , \ScanLink102[18] , 
        \ScanLink102[17] , \ScanLink102[16] , \ScanLink102[15] , 
        \ScanLink102[14] , \ScanLink102[13] , \ScanLink102[12] , 
        \ScanLink102[11] , \ScanLink102[10] , \ScanLink102[9] , 
        \ScanLink102[8] , \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , 
        \ScanLink102[4] , \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , 
        \ScanLink102[0] }), .ScanOut({\ScanLink103[31] , \ScanLink103[30] , 
        \ScanLink103[29] , \ScanLink103[28] , \ScanLink103[27] , 
        \ScanLink103[26] , \ScanLink103[25] , \ScanLink103[24] , 
        \ScanLink103[23] , \ScanLink103[22] , \ScanLink103[21] , 
        \ScanLink103[20] , \ScanLink103[19] , \ScanLink103[18] , 
        \ScanLink103[17] , \ScanLink103[16] , \ScanLink103[15] , 
        \ScanLink103[14] , \ScanLink103[13] , \ScanLink103[12] , 
        \ScanLink103[11] , \ScanLink103[10] , \ScanLink103[9] , 
        \ScanLink103[8] , \ScanLink103[7] , \ScanLink103[6] , \ScanLink103[5] , 
        \ScanLink103[4] , \ScanLink103[3] , \ScanLink103[2] , \ScanLink103[1] , 
        \ScanLink103[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load102[0] ), .Out({\Level1Out102[31] , \Level1Out102[30] , 
        \Level1Out102[29] , \Level1Out102[28] , \Level1Out102[27] , 
        \Level1Out102[26] , \Level1Out102[25] , \Level1Out102[24] , 
        \Level1Out102[23] , \Level1Out102[22] , \Level1Out102[21] , 
        \Level1Out102[20] , \Level1Out102[19] , \Level1Out102[18] , 
        \Level1Out102[17] , \Level1Out102[16] , \Level1Out102[15] , 
        \Level1Out102[14] , \Level1Out102[13] , \Level1Out102[12] , 
        \Level1Out102[11] , \Level1Out102[10] , \Level1Out102[9] , 
        \Level1Out102[8] , \Level1Out102[7] , \Level1Out102[6] , 
        \Level1Out102[5] , \Level1Out102[4] , \Level1Out102[3] , 
        \Level1Out102[2] , \Level1Out102[1] , \Level1Out102[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_152_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load152[0] ), .Out({\Level2Out152[31] , \Level2Out152[30] , 
        \Level2Out152[29] , \Level2Out152[28] , \Level2Out152[27] , 
        \Level2Out152[26] , \Level2Out152[25] , \Level2Out152[24] , 
        \Level2Out152[23] , \Level2Out152[22] , \Level2Out152[21] , 
        \Level2Out152[20] , \Level2Out152[19] , \Level2Out152[18] , 
        \Level2Out152[17] , \Level2Out152[16] , \Level2Out152[15] , 
        \Level2Out152[14] , \Level2Out152[13] , \Level2Out152[12] , 
        \Level2Out152[11] , \Level2Out152[10] , \Level2Out152[9] , 
        \Level2Out152[8] , \Level2Out152[7] , \Level2Out152[6] , 
        \Level2Out152[5] , \Level2Out152[4] , \Level2Out152[3] , 
        \Level2Out152[2] , \Level2Out152[1] , \Level2Out152[0] }), .In1({
        \Level1Out152[31] , \Level1Out152[30] , \Level1Out152[29] , 
        \Level1Out152[28] , \Level1Out152[27] , \Level1Out152[26] , 
        \Level1Out152[25] , \Level1Out152[24] , \Level1Out152[23] , 
        \Level1Out152[22] , \Level1Out152[21] , \Level1Out152[20] , 
        \Level1Out152[19] , \Level1Out152[18] , \Level1Out152[17] , 
        \Level1Out152[16] , \Level1Out152[15] , \Level1Out152[14] , 
        \Level1Out152[13] , \Level1Out152[12] , \Level1Out152[11] , 
        \Level1Out152[10] , \Level1Out152[9] , \Level1Out152[8] , 
        \Level1Out152[7] , \Level1Out152[6] , \Level1Out152[5] , 
        \Level1Out152[4] , \Level1Out152[3] , \Level1Out152[2] , 
        \Level1Out152[1] , \Level1Out152[0] }), .In2({\Level1Out153[31] , 
        \Level1Out153[30] , \Level1Out153[29] , \Level1Out153[28] , 
        \Level1Out153[27] , \Level1Out153[26] , \Level1Out153[25] , 
        \Level1Out153[24] , \Level1Out153[23] , \Level1Out153[22] , 
        \Level1Out153[21] , \Level1Out153[20] , \Level1Out153[19] , 
        \Level1Out153[18] , \Level1Out153[17] , \Level1Out153[16] , 
        \Level1Out153[15] , \Level1Out153[14] , \Level1Out153[13] , 
        \Level1Out153[12] , \Level1Out153[11] , \Level1Out153[10] , 
        \Level1Out153[9] , \Level1Out153[8] , \Level1Out153[7] , 
        \Level1Out153[6] , \Level1Out153[5] , \Level1Out153[4] , 
        \Level1Out153[3] , \Level1Out153[2] , \Level1Out153[1] , 
        \Level1Out153[0] }), .Read1(\Level1Load152[0] ), .Read2(
        \Level1Load153[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_125 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink125[31] , \ScanLink125[30] , 
        \ScanLink125[29] , \ScanLink125[28] , \ScanLink125[27] , 
        \ScanLink125[26] , \ScanLink125[25] , \ScanLink125[24] , 
        \ScanLink125[23] , \ScanLink125[22] , \ScanLink125[21] , 
        \ScanLink125[20] , \ScanLink125[19] , \ScanLink125[18] , 
        \ScanLink125[17] , \ScanLink125[16] , \ScanLink125[15] , 
        \ScanLink125[14] , \ScanLink125[13] , \ScanLink125[12] , 
        \ScanLink125[11] , \ScanLink125[10] , \ScanLink125[9] , 
        \ScanLink125[8] , \ScanLink125[7] , \ScanLink125[6] , \ScanLink125[5] , 
        \ScanLink125[4] , \ScanLink125[3] , \ScanLink125[2] , \ScanLink125[1] , 
        \ScanLink125[0] }), .ScanOut({\ScanLink126[31] , \ScanLink126[30] , 
        \ScanLink126[29] , \ScanLink126[28] , \ScanLink126[27] , 
        \ScanLink126[26] , \ScanLink126[25] , \ScanLink126[24] , 
        \ScanLink126[23] , \ScanLink126[22] , \ScanLink126[21] , 
        \ScanLink126[20] , \ScanLink126[19] , \ScanLink126[18] , 
        \ScanLink126[17] , \ScanLink126[16] , \ScanLink126[15] , 
        \ScanLink126[14] , \ScanLink126[13] , \ScanLink126[12] , 
        \ScanLink126[11] , \ScanLink126[10] , \ScanLink126[9] , 
        \ScanLink126[8] , \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , 
        \ScanLink126[4] , \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , 
        \ScanLink126[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load125[0] ), .Out({\Level1Out125[31] , \Level1Out125[30] , 
        \Level1Out125[29] , \Level1Out125[28] , \Level1Out125[27] , 
        \Level1Out125[26] , \Level1Out125[25] , \Level1Out125[24] , 
        \Level1Out125[23] , \Level1Out125[22] , \Level1Out125[21] , 
        \Level1Out125[20] , \Level1Out125[19] , \Level1Out125[18] , 
        \Level1Out125[17] , \Level1Out125[16] , \Level1Out125[15] , 
        \Level1Out125[14] , \Level1Out125[13] , \Level1Out125[12] , 
        \Level1Out125[11] , \Level1Out125[10] , \Level1Out125[9] , 
        \Level1Out125[8] , \Level1Out125[7] , \Level1Out125[6] , 
        \Level1Out125[5] , \Level1Out125[4] , \Level1Out125[3] , 
        \Level1Out125[2] , \Level1Out125[1] , \Level1Out125[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_215 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink215[31] , \ScanLink215[30] , 
        \ScanLink215[29] , \ScanLink215[28] , \ScanLink215[27] , 
        \ScanLink215[26] , \ScanLink215[25] , \ScanLink215[24] , 
        \ScanLink215[23] , \ScanLink215[22] , \ScanLink215[21] , 
        \ScanLink215[20] , \ScanLink215[19] , \ScanLink215[18] , 
        \ScanLink215[17] , \ScanLink215[16] , \ScanLink215[15] , 
        \ScanLink215[14] , \ScanLink215[13] , \ScanLink215[12] , 
        \ScanLink215[11] , \ScanLink215[10] , \ScanLink215[9] , 
        \ScanLink215[8] , \ScanLink215[7] , \ScanLink215[6] , \ScanLink215[5] , 
        \ScanLink215[4] , \ScanLink215[3] , \ScanLink215[2] , \ScanLink215[1] , 
        \ScanLink215[0] }), .ScanOut({\ScanLink216[31] , \ScanLink216[30] , 
        \ScanLink216[29] , \ScanLink216[28] , \ScanLink216[27] , 
        \ScanLink216[26] , \ScanLink216[25] , \ScanLink216[24] , 
        \ScanLink216[23] , \ScanLink216[22] , \ScanLink216[21] , 
        \ScanLink216[20] , \ScanLink216[19] , \ScanLink216[18] , 
        \ScanLink216[17] , \ScanLink216[16] , \ScanLink216[15] , 
        \ScanLink216[14] , \ScanLink216[13] , \ScanLink216[12] , 
        \ScanLink216[11] , \ScanLink216[10] , \ScanLink216[9] , 
        \ScanLink216[8] , \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , 
        \ScanLink216[4] , \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , 
        \ScanLink216[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load215[0] ), .Out({\Level1Out215[31] , \Level1Out215[30] , 
        \Level1Out215[29] , \Level1Out215[28] , \Level1Out215[27] , 
        \Level1Out215[26] , \Level1Out215[25] , \Level1Out215[24] , 
        \Level1Out215[23] , \Level1Out215[22] , \Level1Out215[21] , 
        \Level1Out215[20] , \Level1Out215[19] , \Level1Out215[18] , 
        \Level1Out215[17] , \Level1Out215[16] , \Level1Out215[15] , 
        \Level1Out215[14] , \Level1Out215[13] , \Level1Out215[12] , 
        \Level1Out215[11] , \Level1Out215[10] , \Level1Out215[9] , 
        \Level1Out215[8] , \Level1Out215[7] , \Level1Out215[6] , 
        \Level1Out215[5] , \Level1Out215[4] , \Level1Out215[3] , 
        \Level1Out215[2] , \Level1Out215[1] , \Level1Out215[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_232 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink232[31] , \ScanLink232[30] , 
        \ScanLink232[29] , \ScanLink232[28] , \ScanLink232[27] , 
        \ScanLink232[26] , \ScanLink232[25] , \ScanLink232[24] , 
        \ScanLink232[23] , \ScanLink232[22] , \ScanLink232[21] , 
        \ScanLink232[20] , \ScanLink232[19] , \ScanLink232[18] , 
        \ScanLink232[17] , \ScanLink232[16] , \ScanLink232[15] , 
        \ScanLink232[14] , \ScanLink232[13] , \ScanLink232[12] , 
        \ScanLink232[11] , \ScanLink232[10] , \ScanLink232[9] , 
        \ScanLink232[8] , \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , 
        \ScanLink232[4] , \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , 
        \ScanLink232[0] }), .ScanOut({\ScanLink233[31] , \ScanLink233[30] , 
        \ScanLink233[29] , \ScanLink233[28] , \ScanLink233[27] , 
        \ScanLink233[26] , \ScanLink233[25] , \ScanLink233[24] , 
        \ScanLink233[23] , \ScanLink233[22] , \ScanLink233[21] , 
        \ScanLink233[20] , \ScanLink233[19] , \ScanLink233[18] , 
        \ScanLink233[17] , \ScanLink233[16] , \ScanLink233[15] , 
        \ScanLink233[14] , \ScanLink233[13] , \ScanLink233[12] , 
        \ScanLink233[11] , \ScanLink233[10] , \ScanLink233[9] , 
        \ScanLink233[8] , \ScanLink233[7] , \ScanLink233[6] , \ScanLink233[5] , 
        \ScanLink233[4] , \ScanLink233[3] , \ScanLink233[2] , \ScanLink233[1] , 
        \ScanLink233[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load232[0] ), .Out({\Level1Out232[31] , \Level1Out232[30] , 
        \Level1Out232[29] , \Level1Out232[28] , \Level1Out232[27] , 
        \Level1Out232[26] , \Level1Out232[25] , \Level1Out232[24] , 
        \Level1Out232[23] , \Level1Out232[22] , \Level1Out232[21] , 
        \Level1Out232[20] , \Level1Out232[19] , \Level1Out232[18] , 
        \Level1Out232[17] , \Level1Out232[16] , \Level1Out232[15] , 
        \Level1Out232[14] , \Level1Out232[13] , \Level1Out232[12] , 
        \Level1Out232[11] , \Level1Out232[10] , \Level1Out232[9] , 
        \Level1Out232[8] , \Level1Out232[7] , \Level1Out232[6] , 
        \Level1Out232[5] , \Level1Out232[4] , \Level1Out232[3] , 
        \Level1Out232[2] , \Level1Out232[1] , \Level1Out232[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_14_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load14[0] ), .Out({\Level2Out14[31] , \Level2Out14[30] , 
        \Level2Out14[29] , \Level2Out14[28] , \Level2Out14[27] , 
        \Level2Out14[26] , \Level2Out14[25] , \Level2Out14[24] , 
        \Level2Out14[23] , \Level2Out14[22] , \Level2Out14[21] , 
        \Level2Out14[20] , \Level2Out14[19] , \Level2Out14[18] , 
        \Level2Out14[17] , \Level2Out14[16] , \Level2Out14[15] , 
        \Level2Out14[14] , \Level2Out14[13] , \Level2Out14[12] , 
        \Level2Out14[11] , \Level2Out14[10] , \Level2Out14[9] , 
        \Level2Out14[8] , \Level2Out14[7] , \Level2Out14[6] , \Level2Out14[5] , 
        \Level2Out14[4] , \Level2Out14[3] , \Level2Out14[2] , \Level2Out14[1] , 
        \Level2Out14[0] }), .In1({\Level1Out14[31] , \Level1Out14[30] , 
        \Level1Out14[29] , \Level1Out14[28] , \Level1Out14[27] , 
        \Level1Out14[26] , \Level1Out14[25] , \Level1Out14[24] , 
        \Level1Out14[23] , \Level1Out14[22] , \Level1Out14[21] , 
        \Level1Out14[20] , \Level1Out14[19] , \Level1Out14[18] , 
        \Level1Out14[17] , \Level1Out14[16] , \Level1Out14[15] , 
        \Level1Out14[14] , \Level1Out14[13] , \Level1Out14[12] , 
        \Level1Out14[11] , \Level1Out14[10] , \Level1Out14[9] , 
        \Level1Out14[8] , \Level1Out14[7] , \Level1Out14[6] , \Level1Out14[5] , 
        \Level1Out14[4] , \Level1Out14[3] , \Level1Out14[2] , \Level1Out14[1] , 
        \Level1Out14[0] }), .In2({\Level1Out15[31] , \Level1Out15[30] , 
        \Level1Out15[29] , \Level1Out15[28] , \Level1Out15[27] , 
        \Level1Out15[26] , \Level1Out15[25] , \Level1Out15[24] , 
        \Level1Out15[23] , \Level1Out15[22] , \Level1Out15[21] , 
        \Level1Out15[20] , \Level1Out15[19] , \Level1Out15[18] , 
        \Level1Out15[17] , \Level1Out15[16] , \Level1Out15[15] , 
        \Level1Out15[14] , \Level1Out15[13] , \Level1Out15[12] , 
        \Level1Out15[11] , \Level1Out15[10] , \Level1Out15[9] , 
        \Level1Out15[8] , \Level1Out15[7] , \Level1Out15[6] , \Level1Out15[5] , 
        \Level1Out15[4] , \Level1Out15[3] , \Level1Out15[2] , \Level1Out15[1] , 
        \Level1Out15[0] }), .Read1(\Level1Load14[0] ), .Read2(
        \Level1Load15[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_178_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load178[0] ), .Out({\Level2Out178[31] , \Level2Out178[30] , 
        \Level2Out178[29] , \Level2Out178[28] , \Level2Out178[27] , 
        \Level2Out178[26] , \Level2Out178[25] , \Level2Out178[24] , 
        \Level2Out178[23] , \Level2Out178[22] , \Level2Out178[21] , 
        \Level2Out178[20] , \Level2Out178[19] , \Level2Out178[18] , 
        \Level2Out178[17] , \Level2Out178[16] , \Level2Out178[15] , 
        \Level2Out178[14] , \Level2Out178[13] , \Level2Out178[12] , 
        \Level2Out178[11] , \Level2Out178[10] , \Level2Out178[9] , 
        \Level2Out178[8] , \Level2Out178[7] , \Level2Out178[6] , 
        \Level2Out178[5] , \Level2Out178[4] , \Level2Out178[3] , 
        \Level2Out178[2] , \Level2Out178[1] , \Level2Out178[0] }), .In1({
        \Level1Out178[31] , \Level1Out178[30] , \Level1Out178[29] , 
        \Level1Out178[28] , \Level1Out178[27] , \Level1Out178[26] , 
        \Level1Out178[25] , \Level1Out178[24] , \Level1Out178[23] , 
        \Level1Out178[22] , \Level1Out178[21] , \Level1Out178[20] , 
        \Level1Out178[19] , \Level1Out178[18] , \Level1Out178[17] , 
        \Level1Out178[16] , \Level1Out178[15] , \Level1Out178[14] , 
        \Level1Out178[13] , \Level1Out178[12] , \Level1Out178[11] , 
        \Level1Out178[10] , \Level1Out178[9] , \Level1Out178[8] , 
        \Level1Out178[7] , \Level1Out178[6] , \Level1Out178[5] , 
        \Level1Out178[4] , \Level1Out178[3] , \Level1Out178[2] , 
        \Level1Out178[1] , \Level1Out178[0] }), .In2({\Level1Out179[31] , 
        \Level1Out179[30] , \Level1Out179[29] , \Level1Out179[28] , 
        \Level1Out179[27] , \Level1Out179[26] , \Level1Out179[25] , 
        \Level1Out179[24] , \Level1Out179[23] , \Level1Out179[22] , 
        \Level1Out179[21] , \Level1Out179[20] , \Level1Out179[19] , 
        \Level1Out179[18] , \Level1Out179[17] , \Level1Out179[16] , 
        \Level1Out179[15] , \Level1Out179[14] , \Level1Out179[13] , 
        \Level1Out179[12] , \Level1Out179[11] , \Level1Out179[10] , 
        \Level1Out179[9] , \Level1Out179[8] , \Level1Out179[7] , 
        \Level1Out179[6] , \Level1Out179[5] , \Level1Out179[4] , 
        \Level1Out179[3] , \Level1Out179[2] , \Level1Out179[1] , 
        \Level1Out179[0] }), .Read1(\Level1Load178[0] ), .Read2(
        \Level1Load179[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_164_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load164[0] ), .Out({\Level4Out164[31] , \Level4Out164[30] , 
        \Level4Out164[29] , \Level4Out164[28] , \Level4Out164[27] , 
        \Level4Out164[26] , \Level4Out164[25] , \Level4Out164[24] , 
        \Level4Out164[23] , \Level4Out164[22] , \Level4Out164[21] , 
        \Level4Out164[20] , \Level4Out164[19] , \Level4Out164[18] , 
        \Level4Out164[17] , \Level4Out164[16] , \Level4Out164[15] , 
        \Level4Out164[14] , \Level4Out164[13] , \Level4Out164[12] , 
        \Level4Out164[11] , \Level4Out164[10] , \Level4Out164[9] , 
        \Level4Out164[8] , \Level4Out164[7] , \Level4Out164[6] , 
        \Level4Out164[5] , \Level4Out164[4] , \Level4Out164[3] , 
        \Level4Out164[2] , \Level4Out164[1] , \Level4Out164[0] }), .In1({
        \Level2Out164[31] , \Level2Out164[30] , \Level2Out164[29] , 
        \Level2Out164[28] , \Level2Out164[27] , \Level2Out164[26] , 
        \Level2Out164[25] , \Level2Out164[24] , \Level2Out164[23] , 
        \Level2Out164[22] , \Level2Out164[21] , \Level2Out164[20] , 
        \Level2Out164[19] , \Level2Out164[18] , \Level2Out164[17] , 
        \Level2Out164[16] , \Level2Out164[15] , \Level2Out164[14] , 
        \Level2Out164[13] , \Level2Out164[12] , \Level2Out164[11] , 
        \Level2Out164[10] , \Level2Out164[9] , \Level2Out164[8] , 
        \Level2Out164[7] , \Level2Out164[6] , \Level2Out164[5] , 
        \Level2Out164[4] , \Level2Out164[3] , \Level2Out164[2] , 
        \Level2Out164[1] , \Level2Out164[0] }), .In2({\Level2Out166[31] , 
        \Level2Out166[30] , \Level2Out166[29] , \Level2Out166[28] , 
        \Level2Out166[27] , \Level2Out166[26] , \Level2Out166[25] , 
        \Level2Out166[24] , \Level2Out166[23] , \Level2Out166[22] , 
        \Level2Out166[21] , \Level2Out166[20] , \Level2Out166[19] , 
        \Level2Out166[18] , \Level2Out166[17] , \Level2Out166[16] , 
        \Level2Out166[15] , \Level2Out166[14] , \Level2Out166[13] , 
        \Level2Out166[12] , \Level2Out166[11] , \Level2Out166[10] , 
        \Level2Out166[9] , \Level2Out166[8] , \Level2Out166[7] , 
        \Level2Out166[6] , \Level2Out166[5] , \Level2Out166[4] , 
        \Level2Out166[3] , \Level2Out166[2] , \Level2Out166[1] , 
        \Level2Out166[0] }), .Read1(\Level2Load164[0] ), .Read2(
        \Level2Load166[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_189 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink189[31] , \ScanLink189[30] , 
        \ScanLink189[29] , \ScanLink189[28] , \ScanLink189[27] , 
        \ScanLink189[26] , \ScanLink189[25] , \ScanLink189[24] , 
        \ScanLink189[23] , \ScanLink189[22] , \ScanLink189[21] , 
        \ScanLink189[20] , \ScanLink189[19] , \ScanLink189[18] , 
        \ScanLink189[17] , \ScanLink189[16] , \ScanLink189[15] , 
        \ScanLink189[14] , \ScanLink189[13] , \ScanLink189[12] , 
        \ScanLink189[11] , \ScanLink189[10] , \ScanLink189[9] , 
        \ScanLink189[8] , \ScanLink189[7] , \ScanLink189[6] , \ScanLink189[5] , 
        \ScanLink189[4] , \ScanLink189[3] , \ScanLink189[2] , \ScanLink189[1] , 
        \ScanLink189[0] }), .ScanOut({\ScanLink190[31] , \ScanLink190[30] , 
        \ScanLink190[29] , \ScanLink190[28] , \ScanLink190[27] , 
        \ScanLink190[26] , \ScanLink190[25] , \ScanLink190[24] , 
        \ScanLink190[23] , \ScanLink190[22] , \ScanLink190[21] , 
        \ScanLink190[20] , \ScanLink190[19] , \ScanLink190[18] , 
        \ScanLink190[17] , \ScanLink190[16] , \ScanLink190[15] , 
        \ScanLink190[14] , \ScanLink190[13] , \ScanLink190[12] , 
        \ScanLink190[11] , \ScanLink190[10] , \ScanLink190[9] , 
        \ScanLink190[8] , \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , 
        \ScanLink190[4] , \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , 
        \ScanLink190[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load189[0] ), .Out({\Level1Out189[31] , \Level1Out189[30] , 
        \Level1Out189[29] , \Level1Out189[28] , \Level1Out189[27] , 
        \Level1Out189[26] , \Level1Out189[25] , \Level1Out189[24] , 
        \Level1Out189[23] , \Level1Out189[22] , \Level1Out189[21] , 
        \Level1Out189[20] , \Level1Out189[19] , \Level1Out189[18] , 
        \Level1Out189[17] , \Level1Out189[16] , \Level1Out189[15] , 
        \Level1Out189[14] , \Level1Out189[13] , \Level1Out189[12] , 
        \Level1Out189[11] , \Level1Out189[10] , \Level1Out189[9] , 
        \Level1Out189[8] , \Level1Out189[7] , \Level1Out189[6] , 
        \Level1Out189[5] , \Level1Out189[4] , \Level1Out189[3] , 
        \Level1Out189[2] , \Level1Out189[1] , \Level1Out189[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_82_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load82[0] ), .Out({\Level2Out82[31] , \Level2Out82[30] , 
        \Level2Out82[29] , \Level2Out82[28] , \Level2Out82[27] , 
        \Level2Out82[26] , \Level2Out82[25] , \Level2Out82[24] , 
        \Level2Out82[23] , \Level2Out82[22] , \Level2Out82[21] , 
        \Level2Out82[20] , \Level2Out82[19] , \Level2Out82[18] , 
        \Level2Out82[17] , \Level2Out82[16] , \Level2Out82[15] , 
        \Level2Out82[14] , \Level2Out82[13] , \Level2Out82[12] , 
        \Level2Out82[11] , \Level2Out82[10] , \Level2Out82[9] , 
        \Level2Out82[8] , \Level2Out82[7] , \Level2Out82[6] , \Level2Out82[5] , 
        \Level2Out82[4] , \Level2Out82[3] , \Level2Out82[2] , \Level2Out82[1] , 
        \Level2Out82[0] }), .In1({\Level1Out82[31] , \Level1Out82[30] , 
        \Level1Out82[29] , \Level1Out82[28] , \Level1Out82[27] , 
        \Level1Out82[26] , \Level1Out82[25] , \Level1Out82[24] , 
        \Level1Out82[23] , \Level1Out82[22] , \Level1Out82[21] , 
        \Level1Out82[20] , \Level1Out82[19] , \Level1Out82[18] , 
        \Level1Out82[17] , \Level1Out82[16] , \Level1Out82[15] , 
        \Level1Out82[14] , \Level1Out82[13] , \Level1Out82[12] , 
        \Level1Out82[11] , \Level1Out82[10] , \Level1Out82[9] , 
        \Level1Out82[8] , \Level1Out82[7] , \Level1Out82[6] , \Level1Out82[5] , 
        \Level1Out82[4] , \Level1Out82[3] , \Level1Out82[2] , \Level1Out82[1] , 
        \Level1Out82[0] }), .In2({\Level1Out83[31] , \Level1Out83[30] , 
        \Level1Out83[29] , \Level1Out83[28] , \Level1Out83[27] , 
        \Level1Out83[26] , \Level1Out83[25] , \Level1Out83[24] , 
        \Level1Out83[23] , \Level1Out83[22] , \Level1Out83[21] , 
        \Level1Out83[20] , \Level1Out83[19] , \Level1Out83[18] , 
        \Level1Out83[17] , \Level1Out83[16] , \Level1Out83[15] , 
        \Level1Out83[14] , \Level1Out83[13] , \Level1Out83[12] , 
        \Level1Out83[11] , \Level1Out83[10] , \Level1Out83[9] , 
        \Level1Out83[8] , \Level1Out83[7] , \Level1Out83[6] , \Level1Out83[5] , 
        \Level1Out83[4] , \Level1Out83[3] , \Level1Out83[2] , \Level1Out83[1] , 
        \Level1Out83[0] }), .Read1(\Level1Load82[0] ), .Read2(
        \Level1Load83[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_96_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load96[0] ), .Out({\Level32Out96[31] , \Level32Out96[30] , 
        \Level32Out96[29] , \Level32Out96[28] , \Level32Out96[27] , 
        \Level32Out96[26] , \Level32Out96[25] , \Level32Out96[24] , 
        \Level32Out96[23] , \Level32Out96[22] , \Level32Out96[21] , 
        \Level32Out96[20] , \Level32Out96[19] , \Level32Out96[18] , 
        \Level32Out96[17] , \Level32Out96[16] , \Level32Out96[15] , 
        \Level32Out96[14] , \Level32Out96[13] , \Level32Out96[12] , 
        \Level32Out96[11] , \Level32Out96[10] , \Level32Out96[9] , 
        \Level32Out96[8] , \Level32Out96[7] , \Level32Out96[6] , 
        \Level32Out96[5] , \Level32Out96[4] , \Level32Out96[3] , 
        \Level32Out96[2] , \Level32Out96[1] , \Level32Out96[0] }), .In1({
        \Level16Out96[31] , \Level16Out96[30] , \Level16Out96[29] , 
        \Level16Out96[28] , \Level16Out96[27] , \Level16Out96[26] , 
        \Level16Out96[25] , \Level16Out96[24] , \Level16Out96[23] , 
        \Level16Out96[22] , \Level16Out96[21] , \Level16Out96[20] , 
        \Level16Out96[19] , \Level16Out96[18] , \Level16Out96[17] , 
        \Level16Out96[16] , \Level16Out96[15] , \Level16Out96[14] , 
        \Level16Out96[13] , \Level16Out96[12] , \Level16Out96[11] , 
        \Level16Out96[10] , \Level16Out96[9] , \Level16Out96[8] , 
        \Level16Out96[7] , \Level16Out96[6] , \Level16Out96[5] , 
        \Level16Out96[4] , \Level16Out96[3] , \Level16Out96[2] , 
        \Level16Out96[1] , \Level16Out96[0] }), .In2({\Level16Out112[31] , 
        \Level16Out112[30] , \Level16Out112[29] , \Level16Out112[28] , 
        \Level16Out112[27] , \Level16Out112[26] , \Level16Out112[25] , 
        \Level16Out112[24] , \Level16Out112[23] , \Level16Out112[22] , 
        \Level16Out112[21] , \Level16Out112[20] , \Level16Out112[19] , 
        \Level16Out112[18] , \Level16Out112[17] , \Level16Out112[16] , 
        \Level16Out112[15] , \Level16Out112[14] , \Level16Out112[13] , 
        \Level16Out112[12] , \Level16Out112[11] , \Level16Out112[10] , 
        \Level16Out112[9] , \Level16Out112[8] , \Level16Out112[7] , 
        \Level16Out112[6] , \Level16Out112[5] , \Level16Out112[4] , 
        \Level16Out112[3] , \Level16Out112[2] , \Level16Out112[1] , 
        \Level16Out112[0] }), .Read1(\Level16Load96[0] ), .Read2(
        \Level16Load112[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_32 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanOut({\ScanLink33[31] , 
        \ScanLink33[30] , \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , 
        \ScanLink33[26] , \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , 
        \ScanLink33[22] , \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , 
        \ScanLink33[18] , \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , 
        \ScanLink33[14] , \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , 
        \ScanLink33[10] , \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , 
        \ScanLink33[6] , \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , 
        \ScanLink33[2] , \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load32[0] ), .Out({
        \Level1Out32[31] , \Level1Out32[30] , \Level1Out32[29] , 
        \Level1Out32[28] , \Level1Out32[27] , \Level1Out32[26] , 
        \Level1Out32[25] , \Level1Out32[24] , \Level1Out32[23] , 
        \Level1Out32[22] , \Level1Out32[21] , \Level1Out32[20] , 
        \Level1Out32[19] , \Level1Out32[18] , \Level1Out32[17] , 
        \Level1Out32[16] , \Level1Out32[15] , \Level1Out32[14] , 
        \Level1Out32[13] , \Level1Out32[12] , \Level1Out32[11] , 
        \Level1Out32[10] , \Level1Out32[9] , \Level1Out32[8] , 
        \Level1Out32[7] , \Level1Out32[6] , \Level1Out32[5] , \Level1Out32[4] , 
        \Level1Out32[3] , \Level1Out32[2] , \Level1Out32[1] , \Level1Out32[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_47 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanOut({\ScanLink48[31] , 
        \ScanLink48[30] , \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , 
        \ScanLink48[26] , \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , 
        \ScanLink48[22] , \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , 
        \ScanLink48[18] , \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , 
        \ScanLink48[14] , \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , 
        \ScanLink48[10] , \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , 
        \ScanLink48[6] , \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , 
        \ScanLink48[2] , \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load47[0] ), .Out({
        \Level1Out47[31] , \Level1Out47[30] , \Level1Out47[29] , 
        \Level1Out47[28] , \Level1Out47[27] , \Level1Out47[26] , 
        \Level1Out47[25] , \Level1Out47[24] , \Level1Out47[23] , 
        \Level1Out47[22] , \Level1Out47[21] , \Level1Out47[20] , 
        \Level1Out47[19] , \Level1Out47[18] , \Level1Out47[17] , 
        \Level1Out47[16] , \Level1Out47[15] , \Level1Out47[14] , 
        \Level1Out47[13] , \Level1Out47[12] , \Level1Out47[11] , 
        \Level1Out47[10] , \Level1Out47[9] , \Level1Out47[8] , 
        \Level1Out47[7] , \Level1Out47[6] , \Level1Out47[5] , \Level1Out47[4] , 
        \Level1Out47[3] , \Level1Out47[2] , \Level1Out47[1] , \Level1Out47[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_60 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanOut({\ScanLink61[31] , 
        \ScanLink61[30] , \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , 
        \ScanLink61[26] , \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , 
        \ScanLink61[22] , \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , 
        \ScanLink61[18] , \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , 
        \ScanLink61[14] , \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , 
        \ScanLink61[10] , \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , 
        \ScanLink61[6] , \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , 
        \ScanLink61[2] , \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load60[0] ), .Out({
        \Level1Out60[31] , \Level1Out60[30] , \Level1Out60[29] , 
        \Level1Out60[28] , \Level1Out60[27] , \Level1Out60[26] , 
        \Level1Out60[25] , \Level1Out60[24] , \Level1Out60[23] , 
        \Level1Out60[22] , \Level1Out60[21] , \Level1Out60[20] , 
        \Level1Out60[19] , \Level1Out60[18] , \Level1Out60[17] , 
        \Level1Out60[16] , \Level1Out60[15] , \Level1Out60[14] , 
        \Level1Out60[13] , \Level1Out60[12] , \Level1Out60[11] , 
        \Level1Out60[10] , \Level1Out60[9] , \Level1Out60[8] , 
        \Level1Out60[7] , \Level1Out60[6] , \Level1Out60[5] , \Level1Out60[4] , 
        \Level1Out60[3] , \Level1Out60[2] , \Level1Out60[1] , \Level1Out60[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_110 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink110[31] , \ScanLink110[30] , 
        \ScanLink110[29] , \ScanLink110[28] , \ScanLink110[27] , 
        \ScanLink110[26] , \ScanLink110[25] , \ScanLink110[24] , 
        \ScanLink110[23] , \ScanLink110[22] , \ScanLink110[21] , 
        \ScanLink110[20] , \ScanLink110[19] , \ScanLink110[18] , 
        \ScanLink110[17] , \ScanLink110[16] , \ScanLink110[15] , 
        \ScanLink110[14] , \ScanLink110[13] , \ScanLink110[12] , 
        \ScanLink110[11] , \ScanLink110[10] , \ScanLink110[9] , 
        \ScanLink110[8] , \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , 
        \ScanLink110[4] , \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , 
        \ScanLink110[0] }), .ScanOut({\ScanLink111[31] , \ScanLink111[30] , 
        \ScanLink111[29] , \ScanLink111[28] , \ScanLink111[27] , 
        \ScanLink111[26] , \ScanLink111[25] , \ScanLink111[24] , 
        \ScanLink111[23] , \ScanLink111[22] , \ScanLink111[21] , 
        \ScanLink111[20] , \ScanLink111[19] , \ScanLink111[18] , 
        \ScanLink111[17] , \ScanLink111[16] , \ScanLink111[15] , 
        \ScanLink111[14] , \ScanLink111[13] , \ScanLink111[12] , 
        \ScanLink111[11] , \ScanLink111[10] , \ScanLink111[9] , 
        \ScanLink111[8] , \ScanLink111[7] , \ScanLink111[6] , \ScanLink111[5] , 
        \ScanLink111[4] , \ScanLink111[3] , \ScanLink111[2] , \ScanLink111[1] , 
        \ScanLink111[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load110[0] ), .Out({\Level1Out110[31] , \Level1Out110[30] , 
        \Level1Out110[29] , \Level1Out110[28] , \Level1Out110[27] , 
        \Level1Out110[26] , \Level1Out110[25] , \Level1Out110[24] , 
        \Level1Out110[23] , \Level1Out110[22] , \Level1Out110[21] , 
        \Level1Out110[20] , \Level1Out110[19] , \Level1Out110[18] , 
        \Level1Out110[17] , \Level1Out110[16] , \Level1Out110[15] , 
        \Level1Out110[14] , \Level1Out110[13] , \Level1Out110[12] , 
        \Level1Out110[11] , \Level1Out110[10] , \Level1Out110[9] , 
        \Level1Out110[8] , \Level1Out110[7] , \Level1Out110[6] , 
        \Level1Out110[5] , \Level1Out110[4] , \Level1Out110[3] , 
        \Level1Out110[2] , \Level1Out110[1] , \Level1Out110[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_137 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink137[31] , \ScanLink137[30] , 
        \ScanLink137[29] , \ScanLink137[28] , \ScanLink137[27] , 
        \ScanLink137[26] , \ScanLink137[25] , \ScanLink137[24] , 
        \ScanLink137[23] , \ScanLink137[22] , \ScanLink137[21] , 
        \ScanLink137[20] , \ScanLink137[19] , \ScanLink137[18] , 
        \ScanLink137[17] , \ScanLink137[16] , \ScanLink137[15] , 
        \ScanLink137[14] , \ScanLink137[13] , \ScanLink137[12] , 
        \ScanLink137[11] , \ScanLink137[10] , \ScanLink137[9] , 
        \ScanLink137[8] , \ScanLink137[7] , \ScanLink137[6] , \ScanLink137[5] , 
        \ScanLink137[4] , \ScanLink137[3] , \ScanLink137[2] , \ScanLink137[1] , 
        \ScanLink137[0] }), .ScanOut({\ScanLink138[31] , \ScanLink138[30] , 
        \ScanLink138[29] , \ScanLink138[28] , \ScanLink138[27] , 
        \ScanLink138[26] , \ScanLink138[25] , \ScanLink138[24] , 
        \ScanLink138[23] , \ScanLink138[22] , \ScanLink138[21] , 
        \ScanLink138[20] , \ScanLink138[19] , \ScanLink138[18] , 
        \ScanLink138[17] , \ScanLink138[16] , \ScanLink138[15] , 
        \ScanLink138[14] , \ScanLink138[13] , \ScanLink138[12] , 
        \ScanLink138[11] , \ScanLink138[10] , \ScanLink138[9] , 
        \ScanLink138[8] , \ScanLink138[7] , \ScanLink138[6] , \ScanLink138[5] , 
        \ScanLink138[4] , \ScanLink138[3] , \ScanLink138[2] , \ScanLink138[1] , 
        \ScanLink138[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load137[0] ), .Out({\Level1Out137[31] , \Level1Out137[30] , 
        \Level1Out137[29] , \Level1Out137[28] , \Level1Out137[27] , 
        \Level1Out137[26] , \Level1Out137[25] , \Level1Out137[24] , 
        \Level1Out137[23] , \Level1Out137[22] , \Level1Out137[21] , 
        \Level1Out137[20] , \Level1Out137[19] , \Level1Out137[18] , 
        \Level1Out137[17] , \Level1Out137[16] , \Level1Out137[15] , 
        \Level1Out137[14] , \Level1Out137[13] , \Level1Out137[12] , 
        \Level1Out137[11] , \Level1Out137[10] , \Level1Out137[9] , 
        \Level1Out137[8] , \Level1Out137[7] , \Level1Out137[6] , 
        \Level1Out137[5] , \Level1Out137[4] , \Level1Out137[3] , 
        \Level1Out137[2] , \Level1Out137[1] , \Level1Out137[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_207 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink207[31] , \ScanLink207[30] , 
        \ScanLink207[29] , \ScanLink207[28] , \ScanLink207[27] , 
        \ScanLink207[26] , \ScanLink207[25] , \ScanLink207[24] , 
        \ScanLink207[23] , \ScanLink207[22] , \ScanLink207[21] , 
        \ScanLink207[20] , \ScanLink207[19] , \ScanLink207[18] , 
        \ScanLink207[17] , \ScanLink207[16] , \ScanLink207[15] , 
        \ScanLink207[14] , \ScanLink207[13] , \ScanLink207[12] , 
        \ScanLink207[11] , \ScanLink207[10] , \ScanLink207[9] , 
        \ScanLink207[8] , \ScanLink207[7] , \ScanLink207[6] , \ScanLink207[5] , 
        \ScanLink207[4] , \ScanLink207[3] , \ScanLink207[2] , \ScanLink207[1] , 
        \ScanLink207[0] }), .ScanOut({\ScanLink208[31] , \ScanLink208[30] , 
        \ScanLink208[29] , \ScanLink208[28] , \ScanLink208[27] , 
        \ScanLink208[26] , \ScanLink208[25] , \ScanLink208[24] , 
        \ScanLink208[23] , \ScanLink208[22] , \ScanLink208[21] , 
        \ScanLink208[20] , \ScanLink208[19] , \ScanLink208[18] , 
        \ScanLink208[17] , \ScanLink208[16] , \ScanLink208[15] , 
        \ScanLink208[14] , \ScanLink208[13] , \ScanLink208[12] , 
        \ScanLink208[11] , \ScanLink208[10] , \ScanLink208[9] , 
        \ScanLink208[8] , \ScanLink208[7] , \ScanLink208[6] , \ScanLink208[5] , 
        \ScanLink208[4] , \ScanLink208[3] , \ScanLink208[2] , \ScanLink208[1] , 
        \ScanLink208[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load207[0] ), .Out({\Level1Out207[31] , \Level1Out207[30] , 
        \Level1Out207[29] , \Level1Out207[28] , \Level1Out207[27] , 
        \Level1Out207[26] , \Level1Out207[25] , \Level1Out207[24] , 
        \Level1Out207[23] , \Level1Out207[22] , \Level1Out207[21] , 
        \Level1Out207[20] , \Level1Out207[19] , \Level1Out207[18] , 
        \Level1Out207[17] , \Level1Out207[16] , \Level1Out207[15] , 
        \Level1Out207[14] , \Level1Out207[13] , \Level1Out207[12] , 
        \Level1Out207[11] , \Level1Out207[10] , \Level1Out207[9] , 
        \Level1Out207[8] , \Level1Out207[7] , \Level1Out207[6] , 
        \Level1Out207[5] , \Level1Out207[4] , \Level1Out207[3] , 
        \Level1Out207[2] , \Level1Out207[1] , \Level1Out207[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_220 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink220[31] , \ScanLink220[30] , 
        \ScanLink220[29] , \ScanLink220[28] , \ScanLink220[27] , 
        \ScanLink220[26] , \ScanLink220[25] , \ScanLink220[24] , 
        \ScanLink220[23] , \ScanLink220[22] , \ScanLink220[21] , 
        \ScanLink220[20] , \ScanLink220[19] , \ScanLink220[18] , 
        \ScanLink220[17] , \ScanLink220[16] , \ScanLink220[15] , 
        \ScanLink220[14] , \ScanLink220[13] , \ScanLink220[12] , 
        \ScanLink220[11] , \ScanLink220[10] , \ScanLink220[9] , 
        \ScanLink220[8] , \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , 
        \ScanLink220[4] , \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , 
        \ScanLink220[0] }), .ScanOut({\ScanLink221[31] , \ScanLink221[30] , 
        \ScanLink221[29] , \ScanLink221[28] , \ScanLink221[27] , 
        \ScanLink221[26] , \ScanLink221[25] , \ScanLink221[24] , 
        \ScanLink221[23] , \ScanLink221[22] , \ScanLink221[21] , 
        \ScanLink221[20] , \ScanLink221[19] , \ScanLink221[18] , 
        \ScanLink221[17] , \ScanLink221[16] , \ScanLink221[15] , 
        \ScanLink221[14] , \ScanLink221[13] , \ScanLink221[12] , 
        \ScanLink221[11] , \ScanLink221[10] , \ScanLink221[9] , 
        \ScanLink221[8] , \ScanLink221[7] , \ScanLink221[6] , \ScanLink221[5] , 
        \ScanLink221[4] , \ScanLink221[3] , \ScanLink221[2] , \ScanLink221[1] , 
        \ScanLink221[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load220[0] ), .Out({\Level1Out220[31] , \Level1Out220[30] , 
        \Level1Out220[29] , \Level1Out220[28] , \Level1Out220[27] , 
        \Level1Out220[26] , \Level1Out220[25] , \Level1Out220[24] , 
        \Level1Out220[23] , \Level1Out220[22] , \Level1Out220[21] , 
        \Level1Out220[20] , \Level1Out220[19] , \Level1Out220[18] , 
        \Level1Out220[17] , \Level1Out220[16] , \Level1Out220[15] , 
        \Level1Out220[14] , \Level1Out220[13] , \Level1Out220[12] , 
        \Level1Out220[11] , \Level1Out220[10] , \Level1Out220[9] , 
        \Level1Out220[8] , \Level1Out220[7] , \Level1Out220[6] , 
        \Level1Out220[5] , \Level1Out220[4] , \Level1Out220[3] , 
        \Level1Out220[2] , \Level1Out220[1] , \Level1Out220[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load0[0] ), .Out({\Level4Out0[31] , \Level4Out0[30] , 
        \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , \Level4Out0[26] , 
        \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , \Level4Out0[22] , 
        \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , \Level4Out0[18] , 
        \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , \Level4Out0[14] , 
        \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , \Level4Out0[10] , 
        \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , \Level4Out0[6] , 
        \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , \Level4Out0[2] , 
        \Level4Out0[1] , \Level4Out0[0] }), .In1({\Level2Out0[31] , 
        \Level2Out0[30] , \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , 
        \Level2Out0[26] , \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , 
        \Level2Out0[22] , \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , 
        \Level2Out0[18] , \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , 
        \Level2Out0[14] , \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , 
        \Level2Out0[10] , \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , 
        \Level2Out0[6] , \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , 
        \Level2Out0[2] , \Level2Out0[1] , \Level2Out0[0] }), .In2({
        \Level2Out2[31] , \Level2Out2[30] , \Level2Out2[29] , \Level2Out2[28] , 
        \Level2Out2[27] , \Level2Out2[26] , \Level2Out2[25] , \Level2Out2[24] , 
        \Level2Out2[23] , \Level2Out2[22] , \Level2Out2[21] , \Level2Out2[20] , 
        \Level2Out2[19] , \Level2Out2[18] , \Level2Out2[17] , \Level2Out2[16] , 
        \Level2Out2[15] , \Level2Out2[14] , \Level2Out2[13] , \Level2Out2[12] , 
        \Level2Out2[11] , \Level2Out2[10] , \Level2Out2[9] , \Level2Out2[8] , 
        \Level2Out2[7] , \Level2Out2[6] , \Level2Out2[5] , \Level2Out2[4] , 
        \Level2Out2[3] , \Level2Out2[2] , \Level2Out2[1] , \Level2Out2[0] }), 
        .Read1(\Level2Load0[0] ), .Read2(\Level2Load2[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_159 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink159[31] , \ScanLink159[30] , 
        \ScanLink159[29] , \ScanLink159[28] , \ScanLink159[27] , 
        \ScanLink159[26] , \ScanLink159[25] , \ScanLink159[24] , 
        \ScanLink159[23] , \ScanLink159[22] , \ScanLink159[21] , 
        \ScanLink159[20] , \ScanLink159[19] , \ScanLink159[18] , 
        \ScanLink159[17] , \ScanLink159[16] , \ScanLink159[15] , 
        \ScanLink159[14] , \ScanLink159[13] , \ScanLink159[12] , 
        \ScanLink159[11] , \ScanLink159[10] , \ScanLink159[9] , 
        \ScanLink159[8] , \ScanLink159[7] , \ScanLink159[6] , \ScanLink159[5] , 
        \ScanLink159[4] , \ScanLink159[3] , \ScanLink159[2] , \ScanLink159[1] , 
        \ScanLink159[0] }), .ScanOut({\ScanLink160[31] , \ScanLink160[30] , 
        \ScanLink160[29] , \ScanLink160[28] , \ScanLink160[27] , 
        \ScanLink160[26] , \ScanLink160[25] , \ScanLink160[24] , 
        \ScanLink160[23] , \ScanLink160[22] , \ScanLink160[21] , 
        \ScanLink160[20] , \ScanLink160[19] , \ScanLink160[18] , 
        \ScanLink160[17] , \ScanLink160[16] , \ScanLink160[15] , 
        \ScanLink160[14] , \ScanLink160[13] , \ScanLink160[12] , 
        \ScanLink160[11] , \ScanLink160[10] , \ScanLink160[9] , 
        \ScanLink160[8] , \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , 
        \ScanLink160[4] , \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , 
        \ScanLink160[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load159[0] ), .Out({\Level1Out159[31] , \Level1Out159[30] , 
        \Level1Out159[29] , \Level1Out159[28] , \Level1Out159[27] , 
        \Level1Out159[26] , \Level1Out159[25] , \Level1Out159[24] , 
        \Level1Out159[23] , \Level1Out159[22] , \Level1Out159[21] , 
        \Level1Out159[20] , \Level1Out159[19] , \Level1Out159[18] , 
        \Level1Out159[17] , \Level1Out159[16] , \Level1Out159[15] , 
        \Level1Out159[14] , \Level1Out159[13] , \Level1Out159[12] , 
        \Level1Out159[11] , \Level1Out159[10] , \Level1Out159[9] , 
        \Level1Out159[8] , \Level1Out159[7] , \Level1Out159[6] , 
        \Level1Out159[5] , \Level1Out159[4] , \Level1Out159[3] , 
        \Level1Out159[2] , \Level1Out159[1] , \Level1Out159[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_44_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load44[0] ), .Out({\Level2Out44[31] , \Level2Out44[30] , 
        \Level2Out44[29] , \Level2Out44[28] , \Level2Out44[27] , 
        \Level2Out44[26] , \Level2Out44[25] , \Level2Out44[24] , 
        \Level2Out44[23] , \Level2Out44[22] , \Level2Out44[21] , 
        \Level2Out44[20] , \Level2Out44[19] , \Level2Out44[18] , 
        \Level2Out44[17] , \Level2Out44[16] , \Level2Out44[15] , 
        \Level2Out44[14] , \Level2Out44[13] , \Level2Out44[12] , 
        \Level2Out44[11] , \Level2Out44[10] , \Level2Out44[9] , 
        \Level2Out44[8] , \Level2Out44[7] , \Level2Out44[6] , \Level2Out44[5] , 
        \Level2Out44[4] , \Level2Out44[3] , \Level2Out44[2] , \Level2Out44[1] , 
        \Level2Out44[0] }), .In1({\Level1Out44[31] , \Level1Out44[30] , 
        \Level1Out44[29] , \Level1Out44[28] , \Level1Out44[27] , 
        \Level1Out44[26] , \Level1Out44[25] , \Level1Out44[24] , 
        \Level1Out44[23] , \Level1Out44[22] , \Level1Out44[21] , 
        \Level1Out44[20] , \Level1Out44[19] , \Level1Out44[18] , 
        \Level1Out44[17] , \Level1Out44[16] , \Level1Out44[15] , 
        \Level1Out44[14] , \Level1Out44[13] , \Level1Out44[12] , 
        \Level1Out44[11] , \Level1Out44[10] , \Level1Out44[9] , 
        \Level1Out44[8] , \Level1Out44[7] , \Level1Out44[6] , \Level1Out44[5] , 
        \Level1Out44[4] , \Level1Out44[3] , \Level1Out44[2] , \Level1Out44[1] , 
        \Level1Out44[0] }), .In2({\Level1Out45[31] , \Level1Out45[30] , 
        \Level1Out45[29] , \Level1Out45[28] , \Level1Out45[27] , 
        \Level1Out45[26] , \Level1Out45[25] , \Level1Out45[24] , 
        \Level1Out45[23] , \Level1Out45[22] , \Level1Out45[21] , 
        \Level1Out45[20] , \Level1Out45[19] , \Level1Out45[18] , 
        \Level1Out45[17] , \Level1Out45[16] , \Level1Out45[15] , 
        \Level1Out45[14] , \Level1Out45[13] , \Level1Out45[12] , 
        \Level1Out45[11] , \Level1Out45[10] , \Level1Out45[9] , 
        \Level1Out45[8] , \Level1Out45[7] , \Level1Out45[6] , \Level1Out45[5] , 
        \Level1Out45[4] , \Level1Out45[3] , \Level1Out45[2] , \Level1Out45[1] , 
        \Level1Out45[0] }), .Read1(\Level1Load44[0] ), .Read2(
        \Level1Load45[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load128[0] ), .Out({\Level2Out128[31] , \Level2Out128[30] , 
        \Level2Out128[29] , \Level2Out128[28] , \Level2Out128[27] , 
        \Level2Out128[26] , \Level2Out128[25] , \Level2Out128[24] , 
        \Level2Out128[23] , \Level2Out128[22] , \Level2Out128[21] , 
        \Level2Out128[20] , \Level2Out128[19] , \Level2Out128[18] , 
        \Level2Out128[17] , \Level2Out128[16] , \Level2Out128[15] , 
        \Level2Out128[14] , \Level2Out128[13] , \Level2Out128[12] , 
        \Level2Out128[11] , \Level2Out128[10] , \Level2Out128[9] , 
        \Level2Out128[8] , \Level2Out128[7] , \Level2Out128[6] , 
        \Level2Out128[5] , \Level2Out128[4] , \Level2Out128[3] , 
        \Level2Out128[2] , \Level2Out128[1] , \Level2Out128[0] }), .In1({
        \Level1Out128[31] , \Level1Out128[30] , \Level1Out128[29] , 
        \Level1Out128[28] , \Level1Out128[27] , \Level1Out128[26] , 
        \Level1Out128[25] , \Level1Out128[24] , \Level1Out128[23] , 
        \Level1Out128[22] , \Level1Out128[21] , \Level1Out128[20] , 
        \Level1Out128[19] , \Level1Out128[18] , \Level1Out128[17] , 
        \Level1Out128[16] , \Level1Out128[15] , \Level1Out128[14] , 
        \Level1Out128[13] , \Level1Out128[12] , \Level1Out128[11] , 
        \Level1Out128[10] , \Level1Out128[9] , \Level1Out128[8] , 
        \Level1Out128[7] , \Level1Out128[6] , \Level1Out128[5] , 
        \Level1Out128[4] , \Level1Out128[3] , \Level1Out128[2] , 
        \Level1Out128[1] , \Level1Out128[0] }), .In2({\Level1Out129[31] , 
        \Level1Out129[30] , \Level1Out129[29] , \Level1Out129[28] , 
        \Level1Out129[27] , \Level1Out129[26] , \Level1Out129[25] , 
        \Level1Out129[24] , \Level1Out129[23] , \Level1Out129[22] , 
        \Level1Out129[21] , \Level1Out129[20] , \Level1Out129[19] , 
        \Level1Out129[18] , \Level1Out129[17] , \Level1Out129[16] , 
        \Level1Out129[15] , \Level1Out129[14] , \Level1Out129[13] , 
        \Level1Out129[12] , \Level1Out129[11] , \Level1Out129[10] , 
        \Level1Out129[9] , \Level1Out129[8] , \Level1Out129[7] , 
        \Level1Out129[6] , \Level1Out129[5] , \Level1Out129[4] , 
        \Level1Out129[3] , \Level1Out129[2] , \Level1Out129[1] , 
        \Level1Out129[0] }), .Read1(\Level1Load128[0] ), .Read2(
        \Level1Load129[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_194_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load194[0] ), .Out({\Level2Out194[31] , \Level2Out194[30] , 
        \Level2Out194[29] , \Level2Out194[28] , \Level2Out194[27] , 
        \Level2Out194[26] , \Level2Out194[25] , \Level2Out194[24] , 
        \Level2Out194[23] , \Level2Out194[22] , \Level2Out194[21] , 
        \Level2Out194[20] , \Level2Out194[19] , \Level2Out194[18] , 
        \Level2Out194[17] , \Level2Out194[16] , \Level2Out194[15] , 
        \Level2Out194[14] , \Level2Out194[13] , \Level2Out194[12] , 
        \Level2Out194[11] , \Level2Out194[10] , \Level2Out194[9] , 
        \Level2Out194[8] , \Level2Out194[7] , \Level2Out194[6] , 
        \Level2Out194[5] , \Level2Out194[4] , \Level2Out194[3] , 
        \Level2Out194[2] , \Level2Out194[1] , \Level2Out194[0] }), .In1({
        \Level1Out194[31] , \Level1Out194[30] , \Level1Out194[29] , 
        \Level1Out194[28] , \Level1Out194[27] , \Level1Out194[26] , 
        \Level1Out194[25] , \Level1Out194[24] , \Level1Out194[23] , 
        \Level1Out194[22] , \Level1Out194[21] , \Level1Out194[20] , 
        \Level1Out194[19] , \Level1Out194[18] , \Level1Out194[17] , 
        \Level1Out194[16] , \Level1Out194[15] , \Level1Out194[14] , 
        \Level1Out194[13] , \Level1Out194[12] , \Level1Out194[11] , 
        \Level1Out194[10] , \Level1Out194[9] , \Level1Out194[8] , 
        \Level1Out194[7] , \Level1Out194[6] , \Level1Out194[5] , 
        \Level1Out194[4] , \Level1Out194[3] , \Level1Out194[2] , 
        \Level1Out194[1] , \Level1Out194[0] }), .In2({\Level1Out195[31] , 
        \Level1Out195[30] , \Level1Out195[29] , \Level1Out195[28] , 
        \Level1Out195[27] , \Level1Out195[26] , \Level1Out195[25] , 
        \Level1Out195[24] , \Level1Out195[23] , \Level1Out195[22] , 
        \Level1Out195[21] , \Level1Out195[20] , \Level1Out195[19] , 
        \Level1Out195[18] , \Level1Out195[17] , \Level1Out195[16] , 
        \Level1Out195[15] , \Level1Out195[14] , \Level1Out195[13] , 
        \Level1Out195[12] , \Level1Out195[11] , \Level1Out195[10] , 
        \Level1Out195[9] , \Level1Out195[8] , \Level1Out195[7] , 
        \Level1Out195[6] , \Level1Out195[5] , \Level1Out195[4] , 
        \Level1Out195[3] , \Level1Out195[2] , \Level1Out195[1] , 
        \Level1Out195[0] }), .Read1(\Level1Load194[0] ), .Read2(
        \Level1Load195[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_188_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load188[0] ), .Out({\Level4Out188[31] , \Level4Out188[30] , 
        \Level4Out188[29] , \Level4Out188[28] , \Level4Out188[27] , 
        \Level4Out188[26] , \Level4Out188[25] , \Level4Out188[24] , 
        \Level4Out188[23] , \Level4Out188[22] , \Level4Out188[21] , 
        \Level4Out188[20] , \Level4Out188[19] , \Level4Out188[18] , 
        \Level4Out188[17] , \Level4Out188[16] , \Level4Out188[15] , 
        \Level4Out188[14] , \Level4Out188[13] , \Level4Out188[12] , 
        \Level4Out188[11] , \Level4Out188[10] , \Level4Out188[9] , 
        \Level4Out188[8] , \Level4Out188[7] , \Level4Out188[6] , 
        \Level4Out188[5] , \Level4Out188[4] , \Level4Out188[3] , 
        \Level4Out188[2] , \Level4Out188[1] , \Level4Out188[0] }), .In1({
        \Level2Out188[31] , \Level2Out188[30] , \Level2Out188[29] , 
        \Level2Out188[28] , \Level2Out188[27] , \Level2Out188[26] , 
        \Level2Out188[25] , \Level2Out188[24] , \Level2Out188[23] , 
        \Level2Out188[22] , \Level2Out188[21] , \Level2Out188[20] , 
        \Level2Out188[19] , \Level2Out188[18] , \Level2Out188[17] , 
        \Level2Out188[16] , \Level2Out188[15] , \Level2Out188[14] , 
        \Level2Out188[13] , \Level2Out188[12] , \Level2Out188[11] , 
        \Level2Out188[10] , \Level2Out188[9] , \Level2Out188[8] , 
        \Level2Out188[7] , \Level2Out188[6] , \Level2Out188[5] , 
        \Level2Out188[4] , \Level2Out188[3] , \Level2Out188[2] , 
        \Level2Out188[1] , \Level2Out188[0] }), .In2({\Level2Out190[31] , 
        \Level2Out190[30] , \Level2Out190[29] , \Level2Out190[28] , 
        \Level2Out190[27] , \Level2Out190[26] , \Level2Out190[25] , 
        \Level2Out190[24] , \Level2Out190[23] , \Level2Out190[22] , 
        \Level2Out190[21] , \Level2Out190[20] , \Level2Out190[19] , 
        \Level2Out190[18] , \Level2Out190[17] , \Level2Out190[16] , 
        \Level2Out190[15] , \Level2Out190[14] , \Level2Out190[13] , 
        \Level2Out190[12] , \Level2Out190[11] , \Level2Out190[10] , 
        \Level2Out190[9] , \Level2Out190[8] , \Level2Out190[7] , 
        \Level2Out190[6] , \Level2Out190[5] , \Level2Out190[4] , 
        \Level2Out190[3] , \Level2Out190[2] , \Level2Out190[1] , 
        \Level2Out190[0] }), .Read1(\Level2Load188[0] ), .Read2(
        \Level2Load190[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_240_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load240[0] ), .Out({\Level16Out240[31] , \Level16Out240[30] , 
        \Level16Out240[29] , \Level16Out240[28] , \Level16Out240[27] , 
        \Level16Out240[26] , \Level16Out240[25] , \Level16Out240[24] , 
        \Level16Out240[23] , \Level16Out240[22] , \Level16Out240[21] , 
        \Level16Out240[20] , \Level16Out240[19] , \Level16Out240[18] , 
        \Level16Out240[17] , \Level16Out240[16] , \Level16Out240[15] , 
        \Level16Out240[14] , \Level16Out240[13] , \Level16Out240[12] , 
        \Level16Out240[11] , \Level16Out240[10] , \Level16Out240[9] , 
        \Level16Out240[8] , \Level16Out240[7] , \Level16Out240[6] , 
        \Level16Out240[5] , \Level16Out240[4] , \Level16Out240[3] , 
        \Level16Out240[2] , \Level16Out240[1] , \Level16Out240[0] }), .In1({
        \Level8Out240[31] , \Level8Out240[30] , \Level8Out240[29] , 
        \Level8Out240[28] , \Level8Out240[27] , \Level8Out240[26] , 
        \Level8Out240[25] , \Level8Out240[24] , \Level8Out240[23] , 
        \Level8Out240[22] , \Level8Out240[21] , \Level8Out240[20] , 
        \Level8Out240[19] , \Level8Out240[18] , \Level8Out240[17] , 
        \Level8Out240[16] , \Level8Out240[15] , \Level8Out240[14] , 
        \Level8Out240[13] , \Level8Out240[12] , \Level8Out240[11] , 
        \Level8Out240[10] , \Level8Out240[9] , \Level8Out240[8] , 
        \Level8Out240[7] , \Level8Out240[6] , \Level8Out240[5] , 
        \Level8Out240[4] , \Level8Out240[3] , \Level8Out240[2] , 
        \Level8Out240[1] , \Level8Out240[0] }), .In2({\Level8Out248[31] , 
        \Level8Out248[30] , \Level8Out248[29] , \Level8Out248[28] , 
        \Level8Out248[27] , \Level8Out248[26] , \Level8Out248[25] , 
        \Level8Out248[24] , \Level8Out248[23] , \Level8Out248[22] , 
        \Level8Out248[21] , \Level8Out248[20] , \Level8Out248[19] , 
        \Level8Out248[18] , \Level8Out248[17] , \Level8Out248[16] , 
        \Level8Out248[15] , \Level8Out248[14] , \Level8Out248[13] , 
        \Level8Out248[12] , \Level8Out248[11] , \Level8Out248[10] , 
        \Level8Out248[9] , \Level8Out248[8] , \Level8Out248[7] , 
        \Level8Out248[6] , \Level8Out248[5] , \Level8Out248[4] , 
        \Level8Out248[3] , \Level8Out248[2] , \Level8Out248[1] , 
        \Level8Out248[0] }), .Read1(\Level8Load240[0] ), .Read2(
        \Level8Load248[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_136_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load136[0] ), .Out({\Level8Out136[31] , \Level8Out136[30] , 
        \Level8Out136[29] , \Level8Out136[28] , \Level8Out136[27] , 
        \Level8Out136[26] , \Level8Out136[25] , \Level8Out136[24] , 
        \Level8Out136[23] , \Level8Out136[22] , \Level8Out136[21] , 
        \Level8Out136[20] , \Level8Out136[19] , \Level8Out136[18] , 
        \Level8Out136[17] , \Level8Out136[16] , \Level8Out136[15] , 
        \Level8Out136[14] , \Level8Out136[13] , \Level8Out136[12] , 
        \Level8Out136[11] , \Level8Out136[10] , \Level8Out136[9] , 
        \Level8Out136[8] , \Level8Out136[7] , \Level8Out136[6] , 
        \Level8Out136[5] , \Level8Out136[4] , \Level8Out136[3] , 
        \Level8Out136[2] , \Level8Out136[1] , \Level8Out136[0] }), .In1({
        \Level4Out136[31] , \Level4Out136[30] , \Level4Out136[29] , 
        \Level4Out136[28] , \Level4Out136[27] , \Level4Out136[26] , 
        \Level4Out136[25] , \Level4Out136[24] , \Level4Out136[23] , 
        \Level4Out136[22] , \Level4Out136[21] , \Level4Out136[20] , 
        \Level4Out136[19] , \Level4Out136[18] , \Level4Out136[17] , 
        \Level4Out136[16] , \Level4Out136[15] , \Level4Out136[14] , 
        \Level4Out136[13] , \Level4Out136[12] , \Level4Out136[11] , 
        \Level4Out136[10] , \Level4Out136[9] , \Level4Out136[8] , 
        \Level4Out136[7] , \Level4Out136[6] , \Level4Out136[5] , 
        \Level4Out136[4] , \Level4Out136[3] , \Level4Out136[2] , 
        \Level4Out136[1] , \Level4Out136[0] }), .In2({\Level4Out140[31] , 
        \Level4Out140[30] , \Level4Out140[29] , \Level4Out140[28] , 
        \Level4Out140[27] , \Level4Out140[26] , \Level4Out140[25] , 
        \Level4Out140[24] , \Level4Out140[23] , \Level4Out140[22] , 
        \Level4Out140[21] , \Level4Out140[20] , \Level4Out140[19] , 
        \Level4Out140[18] , \Level4Out140[17] , \Level4Out140[16] , 
        \Level4Out140[15] , \Level4Out140[14] , \Level4Out140[13] , 
        \Level4Out140[12] , \Level4Out140[11] , \Level4Out140[10] , 
        \Level4Out140[9] , \Level4Out140[8] , \Level4Out140[7] , 
        \Level4Out140[6] , \Level4Out140[5] , \Level4Out140[4] , 
        \Level4Out140[3] , \Level4Out140[2] , \Level4Out140[1] , 
        \Level4Out140[0] }), .Read1(\Level4Load136[0] ), .Read2(
        \Level4Load140[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_236_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load236[0] ), .Out({\Level2Out236[31] , \Level2Out236[30] , 
        \Level2Out236[29] , \Level2Out236[28] , \Level2Out236[27] , 
        \Level2Out236[26] , \Level2Out236[25] , \Level2Out236[24] , 
        \Level2Out236[23] , \Level2Out236[22] , \Level2Out236[21] , 
        \Level2Out236[20] , \Level2Out236[19] , \Level2Out236[18] , 
        \Level2Out236[17] , \Level2Out236[16] , \Level2Out236[15] , 
        \Level2Out236[14] , \Level2Out236[13] , \Level2Out236[12] , 
        \Level2Out236[11] , \Level2Out236[10] , \Level2Out236[9] , 
        \Level2Out236[8] , \Level2Out236[7] , \Level2Out236[6] , 
        \Level2Out236[5] , \Level2Out236[4] , \Level2Out236[3] , 
        \Level2Out236[2] , \Level2Out236[1] , \Level2Out236[0] }), .In1({
        \Level1Out236[31] , \Level1Out236[30] , \Level1Out236[29] , 
        \Level1Out236[28] , \Level1Out236[27] , \Level1Out236[26] , 
        \Level1Out236[25] , \Level1Out236[24] , \Level1Out236[23] , 
        \Level1Out236[22] , \Level1Out236[21] , \Level1Out236[20] , 
        \Level1Out236[19] , \Level1Out236[18] , \Level1Out236[17] , 
        \Level1Out236[16] , \Level1Out236[15] , \Level1Out236[14] , 
        \Level1Out236[13] , \Level1Out236[12] , \Level1Out236[11] , 
        \Level1Out236[10] , \Level1Out236[9] , \Level1Out236[8] , 
        \Level1Out236[7] , \Level1Out236[6] , \Level1Out236[5] , 
        \Level1Out236[4] , \Level1Out236[3] , \Level1Out236[2] , 
        \Level1Out236[1] , \Level1Out236[0] }), .In2({\Level1Out237[31] , 
        \Level1Out237[30] , \Level1Out237[29] , \Level1Out237[28] , 
        \Level1Out237[27] , \Level1Out237[26] , \Level1Out237[25] , 
        \Level1Out237[24] , \Level1Out237[23] , \Level1Out237[22] , 
        \Level1Out237[21] , \Level1Out237[20] , \Level1Out237[19] , 
        \Level1Out237[18] , \Level1Out237[17] , \Level1Out237[16] , 
        \Level1Out237[15] , \Level1Out237[14] , \Level1Out237[13] , 
        \Level1Out237[12] , \Level1Out237[11] , \Level1Out237[10] , 
        \Level1Out237[9] , \Level1Out237[8] , \Level1Out237[7] , 
        \Level1Out237[6] , \Level1Out237[5] , \Level1Out237[4] , 
        \Level1Out237[3] , \Level1Out237[2] , \Level1Out237[1] , 
        \Level1Out237[0] }), .Read1(\Level1Load236[0] ), .Read2(
        \Level1Load237[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_102_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load102[0] ), .Out({\Level2Out102[31] , \Level2Out102[30] , 
        \Level2Out102[29] , \Level2Out102[28] , \Level2Out102[27] , 
        \Level2Out102[26] , \Level2Out102[25] , \Level2Out102[24] , 
        \Level2Out102[23] , \Level2Out102[22] , \Level2Out102[21] , 
        \Level2Out102[20] , \Level2Out102[19] , \Level2Out102[18] , 
        \Level2Out102[17] , \Level2Out102[16] , \Level2Out102[15] , 
        \Level2Out102[14] , \Level2Out102[13] , \Level2Out102[12] , 
        \Level2Out102[11] , \Level2Out102[10] , \Level2Out102[9] , 
        \Level2Out102[8] , \Level2Out102[7] , \Level2Out102[6] , 
        \Level2Out102[5] , \Level2Out102[4] , \Level2Out102[3] , 
        \Level2Out102[2] , \Level2Out102[1] , \Level2Out102[0] }), .In1({
        \Level1Out102[31] , \Level1Out102[30] , \Level1Out102[29] , 
        \Level1Out102[28] , \Level1Out102[27] , \Level1Out102[26] , 
        \Level1Out102[25] , \Level1Out102[24] , \Level1Out102[23] , 
        \Level1Out102[22] , \Level1Out102[21] , \Level1Out102[20] , 
        \Level1Out102[19] , \Level1Out102[18] , \Level1Out102[17] , 
        \Level1Out102[16] , \Level1Out102[15] , \Level1Out102[14] , 
        \Level1Out102[13] , \Level1Out102[12] , \Level1Out102[11] , 
        \Level1Out102[10] , \Level1Out102[9] , \Level1Out102[8] , 
        \Level1Out102[7] , \Level1Out102[6] , \Level1Out102[5] , 
        \Level1Out102[4] , \Level1Out102[3] , \Level1Out102[2] , 
        \Level1Out102[1] , \Level1Out102[0] }), .In2({\Level1Out103[31] , 
        \Level1Out103[30] , \Level1Out103[29] , \Level1Out103[28] , 
        \Level1Out103[27] , \Level1Out103[26] , \Level1Out103[25] , 
        \Level1Out103[24] , \Level1Out103[23] , \Level1Out103[22] , 
        \Level1Out103[21] , \Level1Out103[20] , \Level1Out103[19] , 
        \Level1Out103[18] , \Level1Out103[17] , \Level1Out103[16] , 
        \Level1Out103[15] , \Level1Out103[14] , \Level1Out103[13] , 
        \Level1Out103[12] , \Level1Out103[11] , \Level1Out103[10] , 
        \Level1Out103[9] , \Level1Out103[8] , \Level1Out103[7] , 
        \Level1Out103[6] , \Level1Out103[5] , \Level1Out103[4] , 
        \Level1Out103[3] , \Level1Out103[2] , \Level1Out103[1] , 
        \Level1Out103[0] }), .Read1(\Level1Load102[0] ), .Read2(
        \Level1Load103[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_72_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load72[0] ), .Out({\Level4Out72[31] , \Level4Out72[30] , 
        \Level4Out72[29] , \Level4Out72[28] , \Level4Out72[27] , 
        \Level4Out72[26] , \Level4Out72[25] , \Level4Out72[24] , 
        \Level4Out72[23] , \Level4Out72[22] , \Level4Out72[21] , 
        \Level4Out72[20] , \Level4Out72[19] , \Level4Out72[18] , 
        \Level4Out72[17] , \Level4Out72[16] , \Level4Out72[15] , 
        \Level4Out72[14] , \Level4Out72[13] , \Level4Out72[12] , 
        \Level4Out72[11] , \Level4Out72[10] , \Level4Out72[9] , 
        \Level4Out72[8] , \Level4Out72[7] , \Level4Out72[6] , \Level4Out72[5] , 
        \Level4Out72[4] , \Level4Out72[3] , \Level4Out72[2] , \Level4Out72[1] , 
        \Level4Out72[0] }), .In1({\Level2Out72[31] , \Level2Out72[30] , 
        \Level2Out72[29] , \Level2Out72[28] , \Level2Out72[27] , 
        \Level2Out72[26] , \Level2Out72[25] , \Level2Out72[24] , 
        \Level2Out72[23] , \Level2Out72[22] , \Level2Out72[21] , 
        \Level2Out72[20] , \Level2Out72[19] , \Level2Out72[18] , 
        \Level2Out72[17] , \Level2Out72[16] , \Level2Out72[15] , 
        \Level2Out72[14] , \Level2Out72[13] , \Level2Out72[12] , 
        \Level2Out72[11] , \Level2Out72[10] , \Level2Out72[9] , 
        \Level2Out72[8] , \Level2Out72[7] , \Level2Out72[6] , \Level2Out72[5] , 
        \Level2Out72[4] , \Level2Out72[3] , \Level2Out72[2] , \Level2Out72[1] , 
        \Level2Out72[0] }), .In2({\Level2Out74[31] , \Level2Out74[30] , 
        \Level2Out74[29] , \Level2Out74[28] , \Level2Out74[27] , 
        \Level2Out74[26] , \Level2Out74[25] , \Level2Out74[24] , 
        \Level2Out74[23] , \Level2Out74[22] , \Level2Out74[21] , 
        \Level2Out74[20] , \Level2Out74[19] , \Level2Out74[18] , 
        \Level2Out74[17] , \Level2Out74[16] , \Level2Out74[15] , 
        \Level2Out74[14] , \Level2Out74[13] , \Level2Out74[12] , 
        \Level2Out74[11] , \Level2Out74[10] , \Level2Out74[9] , 
        \Level2Out74[8] , \Level2Out74[7] , \Level2Out74[6] , \Level2Out74[5] , 
        \Level2Out74[4] , \Level2Out74[3] , \Level2Out74[2] , \Level2Out74[1] , 
        \Level2Out74[0] }), .Read1(\Level2Load72[0] ), .Read2(
        \Level2Load74[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_200_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load200[0] ), .Out({\Level4Out200[31] , \Level4Out200[30] , 
        \Level4Out200[29] , \Level4Out200[28] , \Level4Out200[27] , 
        \Level4Out200[26] , \Level4Out200[25] , \Level4Out200[24] , 
        \Level4Out200[23] , \Level4Out200[22] , \Level4Out200[21] , 
        \Level4Out200[20] , \Level4Out200[19] , \Level4Out200[18] , 
        \Level4Out200[17] , \Level4Out200[16] , \Level4Out200[15] , 
        \Level4Out200[14] , \Level4Out200[13] , \Level4Out200[12] , 
        \Level4Out200[11] , \Level4Out200[10] , \Level4Out200[9] , 
        \Level4Out200[8] , \Level4Out200[7] , \Level4Out200[6] , 
        \Level4Out200[5] , \Level4Out200[4] , \Level4Out200[3] , 
        \Level4Out200[2] , \Level4Out200[1] , \Level4Out200[0] }), .In1({
        \Level2Out200[31] , \Level2Out200[30] , \Level2Out200[29] , 
        \Level2Out200[28] , \Level2Out200[27] , \Level2Out200[26] , 
        \Level2Out200[25] , \Level2Out200[24] , \Level2Out200[23] , 
        \Level2Out200[22] , \Level2Out200[21] , \Level2Out200[20] , 
        \Level2Out200[19] , \Level2Out200[18] , \Level2Out200[17] , 
        \Level2Out200[16] , \Level2Out200[15] , \Level2Out200[14] , 
        \Level2Out200[13] , \Level2Out200[12] , \Level2Out200[11] , 
        \Level2Out200[10] , \Level2Out200[9] , \Level2Out200[8] , 
        \Level2Out200[7] , \Level2Out200[6] , \Level2Out200[5] , 
        \Level2Out200[4] , \Level2Out200[3] , \Level2Out200[2] , 
        \Level2Out200[1] , \Level2Out200[0] }), .In2({\Level2Out202[31] , 
        \Level2Out202[30] , \Level2Out202[29] , \Level2Out202[28] , 
        \Level2Out202[27] , \Level2Out202[26] , \Level2Out202[25] , 
        \Level2Out202[24] , \Level2Out202[23] , \Level2Out202[22] , 
        \Level2Out202[21] , \Level2Out202[20] , \Level2Out202[19] , 
        \Level2Out202[18] , \Level2Out202[17] , \Level2Out202[16] , 
        \Level2Out202[15] , \Level2Out202[14] , \Level2Out202[13] , 
        \Level2Out202[12] , \Level2Out202[11] , \Level2Out202[10] , 
        \Level2Out202[9] , \Level2Out202[8] , \Level2Out202[7] , 
        \Level2Out202[6] , \Level2Out202[5] , \Level2Out202[4] , 
        \Level2Out202[3] , \Level2Out202[2] , \Level2Out202[1] , 
        \Level2Out202[0] }), .Read1(\Level2Load200[0] ), .Read2(
        \Level2Load202[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_104_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load104[0] ), .Out({\Level8Out104[31] , \Level8Out104[30] , 
        \Level8Out104[29] , \Level8Out104[28] , \Level8Out104[27] , 
        \Level8Out104[26] , \Level8Out104[25] , \Level8Out104[24] , 
        \Level8Out104[23] , \Level8Out104[22] , \Level8Out104[21] , 
        \Level8Out104[20] , \Level8Out104[19] , \Level8Out104[18] , 
        \Level8Out104[17] , \Level8Out104[16] , \Level8Out104[15] , 
        \Level8Out104[14] , \Level8Out104[13] , \Level8Out104[12] , 
        \Level8Out104[11] , \Level8Out104[10] , \Level8Out104[9] , 
        \Level8Out104[8] , \Level8Out104[7] , \Level8Out104[6] , 
        \Level8Out104[5] , \Level8Out104[4] , \Level8Out104[3] , 
        \Level8Out104[2] , \Level8Out104[1] , \Level8Out104[0] }), .In1({
        \Level4Out104[31] , \Level4Out104[30] , \Level4Out104[29] , 
        \Level4Out104[28] , \Level4Out104[27] , \Level4Out104[26] , 
        \Level4Out104[25] , \Level4Out104[24] , \Level4Out104[23] , 
        \Level4Out104[22] , \Level4Out104[21] , \Level4Out104[20] , 
        \Level4Out104[19] , \Level4Out104[18] , \Level4Out104[17] , 
        \Level4Out104[16] , \Level4Out104[15] , \Level4Out104[14] , 
        \Level4Out104[13] , \Level4Out104[12] , \Level4Out104[11] , 
        \Level4Out104[10] , \Level4Out104[9] , \Level4Out104[8] , 
        \Level4Out104[7] , \Level4Out104[6] , \Level4Out104[5] , 
        \Level4Out104[4] , \Level4Out104[3] , \Level4Out104[2] , 
        \Level4Out104[1] , \Level4Out104[0] }), .In2({\Level4Out108[31] , 
        \Level4Out108[30] , \Level4Out108[29] , \Level4Out108[28] , 
        \Level4Out108[27] , \Level4Out108[26] , \Level4Out108[25] , 
        \Level4Out108[24] , \Level4Out108[23] , \Level4Out108[22] , 
        \Level4Out108[21] , \Level4Out108[20] , \Level4Out108[19] , 
        \Level4Out108[18] , \Level4Out108[17] , \Level4Out108[16] , 
        \Level4Out108[15] , \Level4Out108[14] , \Level4Out108[13] , 
        \Level4Out108[12] , \Level4Out108[11] , \Level4Out108[10] , 
        \Level4Out108[9] , \Level4Out108[8] , \Level4Out108[7] , 
        \Level4Out108[6] , \Level4Out108[5] , \Level4Out108[4] , 
        \Level4Out108[3] , \Level4Out108[2] , \Level4Out108[1] , 
        \Level4Out108[0] }), .Read1(\Level4Load104[0] ), .Read2(
        \Level4Load108[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_255 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink255[31] , \ScanLink255[30] , 
        \ScanLink255[29] , \ScanLink255[28] , \ScanLink255[27] , 
        \ScanLink255[26] , \ScanLink255[25] , \ScanLink255[24] , 
        \ScanLink255[23] , \ScanLink255[22] , \ScanLink255[21] , 
        \ScanLink255[20] , \ScanLink255[19] , \ScanLink255[18] , 
        \ScanLink255[17] , \ScanLink255[16] , \ScanLink255[15] , 
        \ScanLink255[14] , \ScanLink255[13] , \ScanLink255[12] , 
        \ScanLink255[11] , \ScanLink255[10] , \ScanLink255[9] , 
        \ScanLink255[8] , \ScanLink255[7] , \ScanLink255[6] , \ScanLink255[5] , 
        \ScanLink255[4] , \ScanLink255[3] , \ScanLink255[2] , \ScanLink255[1] , 
        \ScanLink255[0] }), .ScanOut({\ScanLink256[31] , \ScanLink256[30] , 
        \ScanLink256[29] , \ScanLink256[28] , \ScanLink256[27] , 
        \ScanLink256[26] , \ScanLink256[25] , \ScanLink256[24] , 
        \ScanLink256[23] , \ScanLink256[22] , \ScanLink256[21] , 
        \ScanLink256[20] , \ScanLink256[19] , \ScanLink256[18] , 
        \ScanLink256[17] , \ScanLink256[16] , \ScanLink256[15] , 
        \ScanLink256[14] , \ScanLink256[13] , \ScanLink256[12] , 
        \ScanLink256[11] , \ScanLink256[10] , \ScanLink256[9] , 
        \ScanLink256[8] , \ScanLink256[7] , \ScanLink256[6] , \ScanLink256[5] , 
        \ScanLink256[4] , \ScanLink256[3] , \ScanLink256[2] , \ScanLink256[1] , 
        \ScanLink256[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load255[0] ), .Out({\Level1Out255[31] , \Level1Out255[30] , 
        \Level1Out255[29] , \Level1Out255[28] , \Level1Out255[27] , 
        \Level1Out255[26] , \Level1Out255[25] , \Level1Out255[24] , 
        \Level1Out255[23] , \Level1Out255[22] , \Level1Out255[21] , 
        \Level1Out255[20] , \Level1Out255[19] , \Level1Out255[18] , 
        \Level1Out255[17] , \Level1Out255[16] , \Level1Out255[15] , 
        \Level1Out255[14] , \Level1Out255[13] , \Level1Out255[12] , 
        \Level1Out255[11] , \Level1Out255[10] , \Level1Out255[9] , 
        \Level1Out255[8] , \Level1Out255[7] , \Level1Out255[6] , 
        \Level1Out255[5] , \Level1Out255[4] , \Level1Out255[3] , 
        \Level1Out255[2] , \Level1Out255[1] , \Level1Out255[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load40[0] ), .Out({\Level4Out40[31] , \Level4Out40[30] , 
        \Level4Out40[29] , \Level4Out40[28] , \Level4Out40[27] , 
        \Level4Out40[26] , \Level4Out40[25] , \Level4Out40[24] , 
        \Level4Out40[23] , \Level4Out40[22] , \Level4Out40[21] , 
        \Level4Out40[20] , \Level4Out40[19] , \Level4Out40[18] , 
        \Level4Out40[17] , \Level4Out40[16] , \Level4Out40[15] , 
        \Level4Out40[14] , \Level4Out40[13] , \Level4Out40[12] , 
        \Level4Out40[11] , \Level4Out40[10] , \Level4Out40[9] , 
        \Level4Out40[8] , \Level4Out40[7] , \Level4Out40[6] , \Level4Out40[5] , 
        \Level4Out40[4] , \Level4Out40[3] , \Level4Out40[2] , \Level4Out40[1] , 
        \Level4Out40[0] }), .In1({\Level2Out40[31] , \Level2Out40[30] , 
        \Level2Out40[29] , \Level2Out40[28] , \Level2Out40[27] , 
        \Level2Out40[26] , \Level2Out40[25] , \Level2Out40[24] , 
        \Level2Out40[23] , \Level2Out40[22] , \Level2Out40[21] , 
        \Level2Out40[20] , \Level2Out40[19] , \Level2Out40[18] , 
        \Level2Out40[17] , \Level2Out40[16] , \Level2Out40[15] , 
        \Level2Out40[14] , \Level2Out40[13] , \Level2Out40[12] , 
        \Level2Out40[11] , \Level2Out40[10] , \Level2Out40[9] , 
        \Level2Out40[8] , \Level2Out40[7] , \Level2Out40[6] , \Level2Out40[5] , 
        \Level2Out40[4] , \Level2Out40[3] , \Level2Out40[2] , \Level2Out40[1] , 
        \Level2Out40[0] }), .In2({\Level2Out42[31] , \Level2Out42[30] , 
        \Level2Out42[29] , \Level2Out42[28] , \Level2Out42[27] , 
        \Level2Out42[26] , \Level2Out42[25] , \Level2Out42[24] , 
        \Level2Out42[23] , \Level2Out42[22] , \Level2Out42[21] , 
        \Level2Out42[20] , \Level2Out42[19] , \Level2Out42[18] , 
        \Level2Out42[17] , \Level2Out42[16] , \Level2Out42[15] , 
        \Level2Out42[14] , \Level2Out42[13] , \Level2Out42[12] , 
        \Level2Out42[11] , \Level2Out42[10] , \Level2Out42[9] , 
        \Level2Out42[8] , \Level2Out42[7] , \Level2Out42[6] , \Level2Out42[5] , 
        \Level2Out42[4] , \Level2Out42[3] , \Level2Out42[2] , \Level2Out42[1] , 
        \Level2Out42[0] }), .Read1(\Level2Load40[0] ), .Read2(
        \Level2Load42[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_130_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load130[0] ), .Out({\Level2Out130[31] , \Level2Out130[30] , 
        \Level2Out130[29] , \Level2Out130[28] , \Level2Out130[27] , 
        \Level2Out130[26] , \Level2Out130[25] , \Level2Out130[24] , 
        \Level2Out130[23] , \Level2Out130[22] , \Level2Out130[21] , 
        \Level2Out130[20] , \Level2Out130[19] , \Level2Out130[18] , 
        \Level2Out130[17] , \Level2Out130[16] , \Level2Out130[15] , 
        \Level2Out130[14] , \Level2Out130[13] , \Level2Out130[12] , 
        \Level2Out130[11] , \Level2Out130[10] , \Level2Out130[9] , 
        \Level2Out130[8] , \Level2Out130[7] , \Level2Out130[6] , 
        \Level2Out130[5] , \Level2Out130[4] , \Level2Out130[3] , 
        \Level2Out130[2] , \Level2Out130[1] , \Level2Out130[0] }), .In1({
        \Level1Out130[31] , \Level1Out130[30] , \Level1Out130[29] , 
        \Level1Out130[28] , \Level1Out130[27] , \Level1Out130[26] , 
        \Level1Out130[25] , \Level1Out130[24] , \Level1Out130[23] , 
        \Level1Out130[22] , \Level1Out130[21] , \Level1Out130[20] , 
        \Level1Out130[19] , \Level1Out130[18] , \Level1Out130[17] , 
        \Level1Out130[16] , \Level1Out130[15] , \Level1Out130[14] , 
        \Level1Out130[13] , \Level1Out130[12] , \Level1Out130[11] , 
        \Level1Out130[10] , \Level1Out130[9] , \Level1Out130[8] , 
        \Level1Out130[7] , \Level1Out130[6] , \Level1Out130[5] , 
        \Level1Out130[4] , \Level1Out130[3] , \Level1Out130[2] , 
        \Level1Out130[1] , \Level1Out130[0] }), .In2({\Level1Out131[31] , 
        \Level1Out131[30] , \Level1Out131[29] , \Level1Out131[28] , 
        \Level1Out131[27] , \Level1Out131[26] , \Level1Out131[25] , 
        \Level1Out131[24] , \Level1Out131[23] , \Level1Out131[22] , 
        \Level1Out131[21] , \Level1Out131[20] , \Level1Out131[19] , 
        \Level1Out131[18] , \Level1Out131[17] , \Level1Out131[16] , 
        \Level1Out131[15] , \Level1Out131[14] , \Level1Out131[13] , 
        \Level1Out131[12] , \Level1Out131[11] , \Level1Out131[10] , 
        \Level1Out131[9] , \Level1Out131[8] , \Level1Out131[7] , 
        \Level1Out131[6] , \Level1Out131[5] , \Level1Out131[4] , 
        \Level1Out131[3] , \Level1Out131[2] , \Level1Out131[1] , 
        \Level1Out131[0] }), .Read1(\Level1Load130[0] ), .Read2(
        \Level1Load131[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load192[0] ), .Out({\Level8Out192[31] , \Level8Out192[30] , 
        \Level8Out192[29] , \Level8Out192[28] , \Level8Out192[27] , 
        \Level8Out192[26] , \Level8Out192[25] , \Level8Out192[24] , 
        \Level8Out192[23] , \Level8Out192[22] , \Level8Out192[21] , 
        \Level8Out192[20] , \Level8Out192[19] , \Level8Out192[18] , 
        \Level8Out192[17] , \Level8Out192[16] , \Level8Out192[15] , 
        \Level8Out192[14] , \Level8Out192[13] , \Level8Out192[12] , 
        \Level8Out192[11] , \Level8Out192[10] , \Level8Out192[9] , 
        \Level8Out192[8] , \Level8Out192[7] , \Level8Out192[6] , 
        \Level8Out192[5] , \Level8Out192[4] , \Level8Out192[3] , 
        \Level8Out192[2] , \Level8Out192[1] , \Level8Out192[0] }), .In1({
        \Level4Out192[31] , \Level4Out192[30] , \Level4Out192[29] , 
        \Level4Out192[28] , \Level4Out192[27] , \Level4Out192[26] , 
        \Level4Out192[25] , \Level4Out192[24] , \Level4Out192[23] , 
        \Level4Out192[22] , \Level4Out192[21] , \Level4Out192[20] , 
        \Level4Out192[19] , \Level4Out192[18] , \Level4Out192[17] , 
        \Level4Out192[16] , \Level4Out192[15] , \Level4Out192[14] , 
        \Level4Out192[13] , \Level4Out192[12] , \Level4Out192[11] , 
        \Level4Out192[10] , \Level4Out192[9] , \Level4Out192[8] , 
        \Level4Out192[7] , \Level4Out192[6] , \Level4Out192[5] , 
        \Level4Out192[4] , \Level4Out192[3] , \Level4Out192[2] , 
        \Level4Out192[1] , \Level4Out192[0] }), .In2({\Level4Out196[31] , 
        \Level4Out196[30] , \Level4Out196[29] , \Level4Out196[28] , 
        \Level4Out196[27] , \Level4Out196[26] , \Level4Out196[25] , 
        \Level4Out196[24] , \Level4Out196[23] , \Level4Out196[22] , 
        \Level4Out196[21] , \Level4Out196[20] , \Level4Out196[19] , 
        \Level4Out196[18] , \Level4Out196[17] , \Level4Out196[16] , 
        \Level4Out196[15] , \Level4Out196[14] , \Level4Out196[13] , 
        \Level4Out196[12] , \Level4Out196[11] , \Level4Out196[10] , 
        \Level4Out196[9] , \Level4Out196[8] , \Level4Out196[7] , 
        \Level4Out196[6] , \Level4Out196[5] , \Level4Out196[4] , 
        \Level4Out196[3] , \Level4Out196[2] , \Level4Out196[1] , 
        \Level4Out196[0] }), .Read1(\Level4Load192[0] ), .Read2(
        \Level4Load196[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_142 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink142[31] , \ScanLink142[30] , 
        \ScanLink142[29] , \ScanLink142[28] , \ScanLink142[27] , 
        \ScanLink142[26] , \ScanLink142[25] , \ScanLink142[24] , 
        \ScanLink142[23] , \ScanLink142[22] , \ScanLink142[21] , 
        \ScanLink142[20] , \ScanLink142[19] , \ScanLink142[18] , 
        \ScanLink142[17] , \ScanLink142[16] , \ScanLink142[15] , 
        \ScanLink142[14] , \ScanLink142[13] , \ScanLink142[12] , 
        \ScanLink142[11] , \ScanLink142[10] , \ScanLink142[9] , 
        \ScanLink142[8] , \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , 
        \ScanLink142[4] , \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , 
        \ScanLink142[0] }), .ScanOut({\ScanLink143[31] , \ScanLink143[30] , 
        \ScanLink143[29] , \ScanLink143[28] , \ScanLink143[27] , 
        \ScanLink143[26] , \ScanLink143[25] , \ScanLink143[24] , 
        \ScanLink143[23] , \ScanLink143[22] , \ScanLink143[21] , 
        \ScanLink143[20] , \ScanLink143[19] , \ScanLink143[18] , 
        \ScanLink143[17] , \ScanLink143[16] , \ScanLink143[15] , 
        \ScanLink143[14] , \ScanLink143[13] , \ScanLink143[12] , 
        \ScanLink143[11] , \ScanLink143[10] , \ScanLink143[9] , 
        \ScanLink143[8] , \ScanLink143[7] , \ScanLink143[6] , \ScanLink143[5] , 
        \ScanLink143[4] , \ScanLink143[3] , \ScanLink143[2] , \ScanLink143[1] , 
        \ScanLink143[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load142[0] ), .Out({\Level1Out142[31] , \Level1Out142[30] , 
        \Level1Out142[29] , \Level1Out142[28] , \Level1Out142[27] , 
        \Level1Out142[26] , \Level1Out142[25] , \Level1Out142[24] , 
        \Level1Out142[23] , \Level1Out142[22] , \Level1Out142[21] , 
        \Level1Out142[20] , \Level1Out142[19] , \Level1Out142[18] , 
        \Level1Out142[17] , \Level1Out142[16] , \Level1Out142[15] , 
        \Level1Out142[14] , \Level1Out142[13] , \Level1Out142[12] , 
        \Level1Out142[11] , \Level1Out142[10] , \Level1Out142[9] , 
        \Level1Out142[8] , \Level1Out142[7] , \Level1Out142[6] , 
        \Level1Out142[5] , \Level1Out142[4] , \Level1Out142[3] , 
        \Level1Out142[2] , \Level1Out142[1] , \Level1Out142[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_165 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink165[31] , \ScanLink165[30] , 
        \ScanLink165[29] , \ScanLink165[28] , \ScanLink165[27] , 
        \ScanLink165[26] , \ScanLink165[25] , \ScanLink165[24] , 
        \ScanLink165[23] , \ScanLink165[22] , \ScanLink165[21] , 
        \ScanLink165[20] , \ScanLink165[19] , \ScanLink165[18] , 
        \ScanLink165[17] , \ScanLink165[16] , \ScanLink165[15] , 
        \ScanLink165[14] , \ScanLink165[13] , \ScanLink165[12] , 
        \ScanLink165[11] , \ScanLink165[10] , \ScanLink165[9] , 
        \ScanLink165[8] , \ScanLink165[7] , \ScanLink165[6] , \ScanLink165[5] , 
        \ScanLink165[4] , \ScanLink165[3] , \ScanLink165[2] , \ScanLink165[1] , 
        \ScanLink165[0] }), .ScanOut({\ScanLink166[31] , \ScanLink166[30] , 
        \ScanLink166[29] , \ScanLink166[28] , \ScanLink166[27] , 
        \ScanLink166[26] , \ScanLink166[25] , \ScanLink166[24] , 
        \ScanLink166[23] , \ScanLink166[22] , \ScanLink166[21] , 
        \ScanLink166[20] , \ScanLink166[19] , \ScanLink166[18] , 
        \ScanLink166[17] , \ScanLink166[16] , \ScanLink166[15] , 
        \ScanLink166[14] , \ScanLink166[13] , \ScanLink166[12] , 
        \ScanLink166[11] , \ScanLink166[10] , \ScanLink166[9] , 
        \ScanLink166[8] , \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , 
        \ScanLink166[4] , \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , 
        \ScanLink166[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load165[0] ), .Out({\Level1Out165[31] , \Level1Out165[30] , 
        \Level1Out165[29] , \Level1Out165[28] , \Level1Out165[27] , 
        \Level1Out165[26] , \Level1Out165[25] , \Level1Out165[24] , 
        \Level1Out165[23] , \Level1Out165[22] , \Level1Out165[21] , 
        \Level1Out165[20] , \Level1Out165[19] , \Level1Out165[18] , 
        \Level1Out165[17] , \Level1Out165[16] , \Level1Out165[15] , 
        \Level1Out165[14] , \Level1Out165[13] , \Level1Out165[12] , 
        \Level1Out165[11] , \Level1Out165[10] , \Level1Out165[9] , 
        \Level1Out165[8] , \Level1Out165[7] , \Level1Out165[6] , 
        \Level1Out165[5] , \Level1Out165[4] , \Level1Out165[3] , 
        \Level1Out165[2] , \Level1Out165[1] , \Level1Out165[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_204_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load204[0] ), .Out({\Level2Out204[31] , \Level2Out204[30] , 
        \Level2Out204[29] , \Level2Out204[28] , \Level2Out204[27] , 
        \Level2Out204[26] , \Level2Out204[25] , \Level2Out204[24] , 
        \Level2Out204[23] , \Level2Out204[22] , \Level2Out204[21] , 
        \Level2Out204[20] , \Level2Out204[19] , \Level2Out204[18] , 
        \Level2Out204[17] , \Level2Out204[16] , \Level2Out204[15] , 
        \Level2Out204[14] , \Level2Out204[13] , \Level2Out204[12] , 
        \Level2Out204[11] , \Level2Out204[10] , \Level2Out204[9] , 
        \Level2Out204[8] , \Level2Out204[7] , \Level2Out204[6] , 
        \Level2Out204[5] , \Level2Out204[4] , \Level2Out204[3] , 
        \Level2Out204[2] , \Level2Out204[1] , \Level2Out204[0] }), .In1({
        \Level1Out204[31] , \Level1Out204[30] , \Level1Out204[29] , 
        \Level1Out204[28] , \Level1Out204[27] , \Level1Out204[26] , 
        \Level1Out204[25] , \Level1Out204[24] , \Level1Out204[23] , 
        \Level1Out204[22] , \Level1Out204[21] , \Level1Out204[20] , 
        \Level1Out204[19] , \Level1Out204[18] , \Level1Out204[17] , 
        \Level1Out204[16] , \Level1Out204[15] , \Level1Out204[14] , 
        \Level1Out204[13] , \Level1Out204[12] , \Level1Out204[11] , 
        \Level1Out204[10] , \Level1Out204[9] , \Level1Out204[8] , 
        \Level1Out204[7] , \Level1Out204[6] , \Level1Out204[5] , 
        \Level1Out204[4] , \Level1Out204[3] , \Level1Out204[2] , 
        \Level1Out204[1] , \Level1Out204[0] }), .In2({\Level1Out205[31] , 
        \Level1Out205[30] , \Level1Out205[29] , \Level1Out205[28] , 
        \Level1Out205[27] , \Level1Out205[26] , \Level1Out205[25] , 
        \Level1Out205[24] , \Level1Out205[23] , \Level1Out205[22] , 
        \Level1Out205[21] , \Level1Out205[20] , \Level1Out205[19] , 
        \Level1Out205[18] , \Level1Out205[17] , \Level1Out205[16] , 
        \Level1Out205[15] , \Level1Out205[14] , \Level1Out205[13] , 
        \Level1Out205[12] , \Level1Out205[11] , \Level1Out205[10] , 
        \Level1Out205[9] , \Level1Out205[8] , \Level1Out205[7] , 
        \Level1Out205[6] , \Level1Out205[5] , \Level1Out205[4] , 
        \Level1Out205[3] , \Level1Out205[2] , \Level1Out205[1] , 
        \Level1Out205[0] }), .Read1(\Level1Load204[0] ), .Read2(
        \Level1Load205[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_232_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load232[0] ), .Out({\Level4Out232[31] , \Level4Out232[30] , 
        \Level4Out232[29] , \Level4Out232[28] , \Level4Out232[27] , 
        \Level4Out232[26] , \Level4Out232[25] , \Level4Out232[24] , 
        \Level4Out232[23] , \Level4Out232[22] , \Level4Out232[21] , 
        \Level4Out232[20] , \Level4Out232[19] , \Level4Out232[18] , 
        \Level4Out232[17] , \Level4Out232[16] , \Level4Out232[15] , 
        \Level4Out232[14] , \Level4Out232[13] , \Level4Out232[12] , 
        \Level4Out232[11] , \Level4Out232[10] , \Level4Out232[9] , 
        \Level4Out232[8] , \Level4Out232[7] , \Level4Out232[6] , 
        \Level4Out232[5] , \Level4Out232[4] , \Level4Out232[3] , 
        \Level4Out232[2] , \Level4Out232[1] , \Level4Out232[0] }), .In1({
        \Level2Out232[31] , \Level2Out232[30] , \Level2Out232[29] , 
        \Level2Out232[28] , \Level2Out232[27] , \Level2Out232[26] , 
        \Level2Out232[25] , \Level2Out232[24] , \Level2Out232[23] , 
        \Level2Out232[22] , \Level2Out232[21] , \Level2Out232[20] , 
        \Level2Out232[19] , \Level2Out232[18] , \Level2Out232[17] , 
        \Level2Out232[16] , \Level2Out232[15] , \Level2Out232[14] , 
        \Level2Out232[13] , \Level2Out232[12] , \Level2Out232[11] , 
        \Level2Out232[10] , \Level2Out232[9] , \Level2Out232[8] , 
        \Level2Out232[7] , \Level2Out232[6] , \Level2Out232[5] , 
        \Level2Out232[4] , \Level2Out232[3] , \Level2Out232[2] , 
        \Level2Out232[1] , \Level2Out232[0] }), .In2({\Level2Out234[31] , 
        \Level2Out234[30] , \Level2Out234[29] , \Level2Out234[28] , 
        \Level2Out234[27] , \Level2Out234[26] , \Level2Out234[25] , 
        \Level2Out234[24] , \Level2Out234[23] , \Level2Out234[22] , 
        \Level2Out234[21] , \Level2Out234[20] , \Level2Out234[19] , 
        \Level2Out234[18] , \Level2Out234[17] , \Level2Out234[16] , 
        \Level2Out234[15] , \Level2Out234[14] , \Level2Out234[13] , 
        \Level2Out234[12] , \Level2Out234[11] , \Level2Out234[10] , 
        \Level2Out234[9] , \Level2Out234[8] , \Level2Out234[7] , 
        \Level2Out234[6] , \Level2Out234[5] , \Level2Out234[4] , 
        \Level2Out234[3] , \Level2Out234[2] , \Level2Out234[1] , 
        \Level2Out234[0] }), .Read1(\Level2Load232[0] ), .Read2(
        \Level2Load234[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_76_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load76[0] ), .Out({\Level2Out76[31] , \Level2Out76[30] , 
        \Level2Out76[29] , \Level2Out76[28] , \Level2Out76[27] , 
        \Level2Out76[26] , \Level2Out76[25] , \Level2Out76[24] , 
        \Level2Out76[23] , \Level2Out76[22] , \Level2Out76[21] , 
        \Level2Out76[20] , \Level2Out76[19] , \Level2Out76[18] , 
        \Level2Out76[17] , \Level2Out76[16] , \Level2Out76[15] , 
        \Level2Out76[14] , \Level2Out76[13] , \Level2Out76[12] , 
        \Level2Out76[11] , \Level2Out76[10] , \Level2Out76[9] , 
        \Level2Out76[8] , \Level2Out76[7] , \Level2Out76[6] , \Level2Out76[5] , 
        \Level2Out76[4] , \Level2Out76[3] , \Level2Out76[2] , \Level2Out76[1] , 
        \Level2Out76[0] }), .In1({\Level1Out76[31] , \Level1Out76[30] , 
        \Level1Out76[29] , \Level1Out76[28] , \Level1Out76[27] , 
        \Level1Out76[26] , \Level1Out76[25] , \Level1Out76[24] , 
        \Level1Out76[23] , \Level1Out76[22] , \Level1Out76[21] , 
        \Level1Out76[20] , \Level1Out76[19] , \Level1Out76[18] , 
        \Level1Out76[17] , \Level1Out76[16] , \Level1Out76[15] , 
        \Level1Out76[14] , \Level1Out76[13] , \Level1Out76[12] , 
        \Level1Out76[11] , \Level1Out76[10] , \Level1Out76[9] , 
        \Level1Out76[8] , \Level1Out76[7] , \Level1Out76[6] , \Level1Out76[5] , 
        \Level1Out76[4] , \Level1Out76[3] , \Level1Out76[2] , \Level1Out76[1] , 
        \Level1Out76[0] }), .In2({\Level1Out77[31] , \Level1Out77[30] , 
        \Level1Out77[29] , \Level1Out77[28] , \Level1Out77[27] , 
        \Level1Out77[26] , \Level1Out77[25] , \Level1Out77[24] , 
        \Level1Out77[23] , \Level1Out77[22] , \Level1Out77[21] , 
        \Level1Out77[20] , \Level1Out77[19] , \Level1Out77[18] , 
        \Level1Out77[17] , \Level1Out77[16] , \Level1Out77[15] , 
        \Level1Out77[14] , \Level1Out77[13] , \Level1Out77[12] , 
        \Level1Out77[11] , \Level1Out77[10] , \Level1Out77[9] , 
        \Level1Out77[8] , \Level1Out77[7] , \Level1Out77[6] , \Level1Out77[5] , 
        \Level1Out77[4] , \Level1Out77[3] , \Level1Out77[2] , \Level1Out77[1] , 
        \Level1Out77[0] }), .Read1(\Level1Load76[0] ), .Read2(
        \Level1Load77[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanOut({\ScanLink3[31] , 
        \ScanLink3[30] , \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , 
        \ScanLink3[26] , \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , 
        \ScanLink3[22] , \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , 
        \ScanLink3[18] , \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , 
        \ScanLink3[14] , \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , 
        \ScanLink3[10] , \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , 
        \ScanLink3[6] , \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , 
        \ScanLink3[2] , \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load2[0] ), .Out({
        \Level1Out2[31] , \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , 
        \Level1Out2[27] , \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , 
        \Level1Out2[23] , \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , 
        \Level1Out2[19] , \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , 
        \Level1Out2[15] , \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , 
        \Level1Out2[11] , \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , 
        \Level1Out2[7] , \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , 
        \Level1Out2[3] , \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_22 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanOut({\ScanLink23[31] , 
        \ScanLink23[30] , \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , 
        \ScanLink23[26] , \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , 
        \ScanLink23[22] , \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , 
        \ScanLink23[18] , \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , 
        \ScanLink23[14] , \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , 
        \ScanLink23[10] , \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , 
        \ScanLink23[6] , \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , 
        \ScanLink23[2] , \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load22[0] ), .Out({
        \Level1Out22[31] , \Level1Out22[30] , \Level1Out22[29] , 
        \Level1Out22[28] , \Level1Out22[27] , \Level1Out22[26] , 
        \Level1Out22[25] , \Level1Out22[24] , \Level1Out22[23] , 
        \Level1Out22[22] , \Level1Out22[21] , \Level1Out22[20] , 
        \Level1Out22[19] , \Level1Out22[18] , \Level1Out22[17] , 
        \Level1Out22[16] , \Level1Out22[15] , \Level1Out22[14] , 
        \Level1Out22[13] , \Level1Out22[12] , \Level1Out22[11] , 
        \Level1Out22[10] , \Level1Out22[9] , \Level1Out22[8] , 
        \Level1Out22[7] , \Level1Out22[6] , \Level1Out22[5] , \Level1Out22[4] , 
        \Level1Out22[3] , \Level1Out22[2] , \Level1Out22[1] , \Level1Out22[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_29 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanOut({\ScanLink30[31] , 
        \ScanLink30[30] , \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , 
        \ScanLink30[26] , \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , 
        \ScanLink30[22] , \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , 
        \ScanLink30[18] , \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , 
        \ScanLink30[14] , \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , 
        \ScanLink30[10] , \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , 
        \ScanLink30[6] , \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , 
        \ScanLink30[2] , \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load29[0] ), .Out({
        \Level1Out29[31] , \Level1Out29[30] , \Level1Out29[29] , 
        \Level1Out29[28] , \Level1Out29[27] , \Level1Out29[26] , 
        \Level1Out29[25] , \Level1Out29[24] , \Level1Out29[23] , 
        \Level1Out29[22] , \Level1Out29[21] , \Level1Out29[20] , 
        \Level1Out29[19] , \Level1Out29[18] , \Level1Out29[17] , 
        \Level1Out29[16] , \Level1Out29[15] , \Level1Out29[14] , 
        \Level1Out29[13] , \Level1Out29[12] , \Level1Out29[11] , 
        \Level1Out29[10] , \Level1Out29[9] , \Level1Out29[8] , 
        \Level1Out29[7] , \Level1Out29[6] , \Level1Out29[5] , \Level1Out29[4] , 
        \Level1Out29[3] , \Level1Out29[2] , \Level1Out29[1] , \Level1Out29[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_85 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink85[31] , \ScanLink85[30] , 
        \ScanLink85[29] , \ScanLink85[28] , \ScanLink85[27] , \ScanLink85[26] , 
        \ScanLink85[25] , \ScanLink85[24] , \ScanLink85[23] , \ScanLink85[22] , 
        \ScanLink85[21] , \ScanLink85[20] , \ScanLink85[19] , \ScanLink85[18] , 
        \ScanLink85[17] , \ScanLink85[16] , \ScanLink85[15] , \ScanLink85[14] , 
        \ScanLink85[13] , \ScanLink85[12] , \ScanLink85[11] , \ScanLink85[10] , 
        \ScanLink85[9] , \ScanLink85[8] , \ScanLink85[7] , \ScanLink85[6] , 
        \ScanLink85[5] , \ScanLink85[4] , \ScanLink85[3] , \ScanLink85[2] , 
        \ScanLink85[1] , \ScanLink85[0] }), .ScanOut({\ScanLink86[31] , 
        \ScanLink86[30] , \ScanLink86[29] , \ScanLink86[28] , \ScanLink86[27] , 
        \ScanLink86[26] , \ScanLink86[25] , \ScanLink86[24] , \ScanLink86[23] , 
        \ScanLink86[22] , \ScanLink86[21] , \ScanLink86[20] , \ScanLink86[19] , 
        \ScanLink86[18] , \ScanLink86[17] , \ScanLink86[16] , \ScanLink86[15] , 
        \ScanLink86[14] , \ScanLink86[13] , \ScanLink86[12] , \ScanLink86[11] , 
        \ScanLink86[10] , \ScanLink86[9] , \ScanLink86[8] , \ScanLink86[7] , 
        \ScanLink86[6] , \ScanLink86[5] , \ScanLink86[4] , \ScanLink86[3] , 
        \ScanLink86[2] , \ScanLink86[1] , \ScanLink86[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load85[0] ), .Out({
        \Level1Out85[31] , \Level1Out85[30] , \Level1Out85[29] , 
        \Level1Out85[28] , \Level1Out85[27] , \Level1Out85[26] , 
        \Level1Out85[25] , \Level1Out85[24] , \Level1Out85[23] , 
        \Level1Out85[22] , \Level1Out85[21] , \Level1Out85[20] , 
        \Level1Out85[19] , \Level1Out85[18] , \Level1Out85[17] , 
        \Level1Out85[16] , \Level1Out85[15] , \Level1Out85[14] , 
        \Level1Out85[13] , \Level1Out85[12] , \Level1Out85[11] , 
        \Level1Out85[10] , \Level1Out85[9] , \Level1Out85[8] , 
        \Level1Out85[7] , \Level1Out85[6] , \Level1Out85[5] , \Level1Out85[4] , 
        \Level1Out85[3] , \Level1Out85[2] , \Level1Out85[1] , \Level1Out85[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_180 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink180[31] , \ScanLink180[30] , 
        \ScanLink180[29] , \ScanLink180[28] , \ScanLink180[27] , 
        \ScanLink180[26] , \ScanLink180[25] , \ScanLink180[24] , 
        \ScanLink180[23] , \ScanLink180[22] , \ScanLink180[21] , 
        \ScanLink180[20] , \ScanLink180[19] , \ScanLink180[18] , 
        \ScanLink180[17] , \ScanLink180[16] , \ScanLink180[15] , 
        \ScanLink180[14] , \ScanLink180[13] , \ScanLink180[12] , 
        \ScanLink180[11] , \ScanLink180[10] , \ScanLink180[9] , 
        \ScanLink180[8] , \ScanLink180[7] , \ScanLink180[6] , \ScanLink180[5] , 
        \ScanLink180[4] , \ScanLink180[3] , \ScanLink180[2] , \ScanLink180[1] , 
        \ScanLink180[0] }), .ScanOut({\ScanLink181[31] , \ScanLink181[30] , 
        \ScanLink181[29] , \ScanLink181[28] , \ScanLink181[27] , 
        \ScanLink181[26] , \ScanLink181[25] , \ScanLink181[24] , 
        \ScanLink181[23] , \ScanLink181[22] , \ScanLink181[21] , 
        \ScanLink181[20] , \ScanLink181[19] , \ScanLink181[18] , 
        \ScanLink181[17] , \ScanLink181[16] , \ScanLink181[15] , 
        \ScanLink181[14] , \ScanLink181[13] , \ScanLink181[12] , 
        \ScanLink181[11] , \ScanLink181[10] , \ScanLink181[9] , 
        \ScanLink181[8] , \ScanLink181[7] , \ScanLink181[6] , \ScanLink181[5] , 
        \ScanLink181[4] , \ScanLink181[3] , \ScanLink181[2] , \ScanLink181[1] , 
        \ScanLink181[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load180[0] ), .Out({\Level1Out180[31] , \Level1Out180[30] , 
        \Level1Out180[29] , \Level1Out180[28] , \Level1Out180[27] , 
        \Level1Out180[26] , \Level1Out180[25] , \Level1Out180[24] , 
        \Level1Out180[23] , \Level1Out180[22] , \Level1Out180[21] , 
        \Level1Out180[20] , \Level1Out180[19] , \Level1Out180[18] , 
        \Level1Out180[17] , \Level1Out180[16] , \Level1Out180[15] , 
        \Level1Out180[14] , \Level1Out180[13] , \Level1Out180[12] , 
        \Level1Out180[11] , \Level1Out180[10] , \Level1Out180[9] , 
        \Level1Out180[8] , \Level1Out180[7] , \Level1Out180[6] , 
        \Level1Out180[5] , \Level1Out180[4] , \Level1Out180[3] , 
        \Level1Out180[2] , \Level1Out180[1] , \Level1Out180[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load4[0] ), .Out({\Level2Out4[31] , \Level2Out4[30] , 
        \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , \Level2Out4[26] , 
        \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , \Level2Out4[22] , 
        \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , \Level2Out4[18] , 
        \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , \Level2Out4[14] , 
        \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , \Level2Out4[10] , 
        \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , \Level2Out4[6] , 
        \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , \Level2Out4[2] , 
        \Level2Out4[1] , \Level2Out4[0] }), .In1({\Level1Out4[31] , 
        \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , \Level1Out4[27] , 
        \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , \Level1Out4[23] , 
        \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , \Level1Out4[19] , 
        \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , \Level1Out4[15] , 
        \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , \Level1Out4[11] , 
        \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , \Level1Out4[7] , 
        \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , \Level1Out4[3] , 
        \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] }), .In2({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] }), 
        .Read1(\Level1Load4[0] ), .Read2(\Level1Load5[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_100 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink100[31] , \ScanLink100[30] , 
        \ScanLink100[29] , \ScanLink100[28] , \ScanLink100[27] , 
        \ScanLink100[26] , \ScanLink100[25] , \ScanLink100[24] , 
        \ScanLink100[23] , \ScanLink100[22] , \ScanLink100[21] , 
        \ScanLink100[20] , \ScanLink100[19] , \ScanLink100[18] , 
        \ScanLink100[17] , \ScanLink100[16] , \ScanLink100[15] , 
        \ScanLink100[14] , \ScanLink100[13] , \ScanLink100[12] , 
        \ScanLink100[11] , \ScanLink100[10] , \ScanLink100[9] , 
        \ScanLink100[8] , \ScanLink100[7] , \ScanLink100[6] , \ScanLink100[5] , 
        \ScanLink100[4] , \ScanLink100[3] , \ScanLink100[2] , \ScanLink100[1] , 
        \ScanLink100[0] }), .ScanOut({\ScanLink101[31] , \ScanLink101[30] , 
        \ScanLink101[29] , \ScanLink101[28] , \ScanLink101[27] , 
        \ScanLink101[26] , \ScanLink101[25] , \ScanLink101[24] , 
        \ScanLink101[23] , \ScanLink101[22] , \ScanLink101[21] , 
        \ScanLink101[20] , \ScanLink101[19] , \ScanLink101[18] , 
        \ScanLink101[17] , \ScanLink101[16] , \ScanLink101[15] , 
        \ScanLink101[14] , \ScanLink101[13] , \ScanLink101[12] , 
        \ScanLink101[11] , \ScanLink101[10] , \ScanLink101[9] , 
        \ScanLink101[8] , \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , 
        \ScanLink101[4] , \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , 
        \ScanLink101[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load100[0] ), .Out({\Level1Out100[31] , \Level1Out100[30] , 
        \Level1Out100[29] , \Level1Out100[28] , \Level1Out100[27] , 
        \Level1Out100[26] , \Level1Out100[25] , \Level1Out100[24] , 
        \Level1Out100[23] , \Level1Out100[22] , \Level1Out100[21] , 
        \Level1Out100[20] , \Level1Out100[19] , \Level1Out100[18] , 
        \Level1Out100[17] , \Level1Out100[16] , \Level1Out100[15] , 
        \Level1Out100[14] , \Level1Out100[13] , \Level1Out100[12] , 
        \Level1Out100[11] , \Level1Out100[10] , \Level1Out100[9] , 
        \Level1Out100[8] , \Level1Out100[7] , \Level1Out100[6] , 
        \Level1Out100[5] , \Level1Out100[4] , \Level1Out100[3] , 
        \Level1Out100[2] , \Level1Out100[1] , \Level1Out100[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_127 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink127[31] , \ScanLink127[30] , 
        \ScanLink127[29] , \ScanLink127[28] , \ScanLink127[27] , 
        \ScanLink127[26] , \ScanLink127[25] , \ScanLink127[24] , 
        \ScanLink127[23] , \ScanLink127[22] , \ScanLink127[21] , 
        \ScanLink127[20] , \ScanLink127[19] , \ScanLink127[18] , 
        \ScanLink127[17] , \ScanLink127[16] , \ScanLink127[15] , 
        \ScanLink127[14] , \ScanLink127[13] , \ScanLink127[12] , 
        \ScanLink127[11] , \ScanLink127[10] , \ScanLink127[9] , 
        \ScanLink127[8] , \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , 
        \ScanLink127[4] , \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , 
        \ScanLink127[0] }), .ScanOut({\ScanLink128[31] , \ScanLink128[30] , 
        \ScanLink128[29] , \ScanLink128[28] , \ScanLink128[27] , 
        \ScanLink128[26] , \ScanLink128[25] , \ScanLink128[24] , 
        \ScanLink128[23] , \ScanLink128[22] , \ScanLink128[21] , 
        \ScanLink128[20] , \ScanLink128[19] , \ScanLink128[18] , 
        \ScanLink128[17] , \ScanLink128[16] , \ScanLink128[15] , 
        \ScanLink128[14] , \ScanLink128[13] , \ScanLink128[12] , 
        \ScanLink128[11] , \ScanLink128[10] , \ScanLink128[9] , 
        \ScanLink128[8] , \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , 
        \ScanLink128[4] , \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , 
        \ScanLink128[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load127[0] ), .Out({\Level1Out127[31] , \Level1Out127[30] , 
        \Level1Out127[29] , \Level1Out127[28] , \Level1Out127[27] , 
        \Level1Out127[26] , \Level1Out127[25] , \Level1Out127[24] , 
        \Level1Out127[23] , \Level1Out127[22] , \Level1Out127[21] , 
        \Level1Out127[20] , \Level1Out127[19] , \Level1Out127[18] , 
        \Level1Out127[17] , \Level1Out127[16] , \Level1Out127[15] , 
        \Level1Out127[14] , \Level1Out127[13] , \Level1Out127[12] , 
        \Level1Out127[11] , \Level1Out127[10] , \Level1Out127[9] , 
        \Level1Out127[8] , \Level1Out127[7] , \Level1Out127[6] , 
        \Level1Out127[5] , \Level1Out127[4] , \Level1Out127[3] , 
        \Level1Out127[2] , \Level1Out127[1] , \Level1Out127[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_217 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink217[31] , \ScanLink217[30] , 
        \ScanLink217[29] , \ScanLink217[28] , \ScanLink217[27] , 
        \ScanLink217[26] , \ScanLink217[25] , \ScanLink217[24] , 
        \ScanLink217[23] , \ScanLink217[22] , \ScanLink217[21] , 
        \ScanLink217[20] , \ScanLink217[19] , \ScanLink217[18] , 
        \ScanLink217[17] , \ScanLink217[16] , \ScanLink217[15] , 
        \ScanLink217[14] , \ScanLink217[13] , \ScanLink217[12] , 
        \ScanLink217[11] , \ScanLink217[10] , \ScanLink217[9] , 
        \ScanLink217[8] , \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , 
        \ScanLink217[4] , \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , 
        \ScanLink217[0] }), .ScanOut({\ScanLink218[31] , \ScanLink218[30] , 
        \ScanLink218[29] , \ScanLink218[28] , \ScanLink218[27] , 
        \ScanLink218[26] , \ScanLink218[25] , \ScanLink218[24] , 
        \ScanLink218[23] , \ScanLink218[22] , \ScanLink218[21] , 
        \ScanLink218[20] , \ScanLink218[19] , \ScanLink218[18] , 
        \ScanLink218[17] , \ScanLink218[16] , \ScanLink218[15] , 
        \ScanLink218[14] , \ScanLink218[13] , \ScanLink218[12] , 
        \ScanLink218[11] , \ScanLink218[10] , \ScanLink218[9] , 
        \ScanLink218[8] , \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , 
        \ScanLink218[4] , \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , 
        \ScanLink218[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load217[0] ), .Out({\Level1Out217[31] , \Level1Out217[30] , 
        \Level1Out217[29] , \Level1Out217[28] , \Level1Out217[27] , 
        \Level1Out217[26] , \Level1Out217[25] , \Level1Out217[24] , 
        \Level1Out217[23] , \Level1Out217[22] , \Level1Out217[21] , 
        \Level1Out217[20] , \Level1Out217[19] , \Level1Out217[18] , 
        \Level1Out217[17] , \Level1Out217[16] , \Level1Out217[15] , 
        \Level1Out217[14] , \Level1Out217[13] , \Level1Out217[12] , 
        \Level1Out217[11] , \Level1Out217[10] , \Level1Out217[9] , 
        \Level1Out217[8] , \Level1Out217[7] , \Level1Out217[6] , 
        \Level1Out217[5] , \Level1Out217[4] , \Level1Out217[3] , 
        \Level1Out217[2] , \Level1Out217[1] , \Level1Out217[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_112_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load112[0] ), .Out({\Level8Out112[31] , \Level8Out112[30] , 
        \Level8Out112[29] , \Level8Out112[28] , \Level8Out112[27] , 
        \Level8Out112[26] , \Level8Out112[25] , \Level8Out112[24] , 
        \Level8Out112[23] , \Level8Out112[22] , \Level8Out112[21] , 
        \Level8Out112[20] , \Level8Out112[19] , \Level8Out112[18] , 
        \Level8Out112[17] , \Level8Out112[16] , \Level8Out112[15] , 
        \Level8Out112[14] , \Level8Out112[13] , \Level8Out112[12] , 
        \Level8Out112[11] , \Level8Out112[10] , \Level8Out112[9] , 
        \Level8Out112[8] , \Level8Out112[7] , \Level8Out112[6] , 
        \Level8Out112[5] , \Level8Out112[4] , \Level8Out112[3] , 
        \Level8Out112[2] , \Level8Out112[1] , \Level8Out112[0] }), .In1({
        \Level4Out112[31] , \Level4Out112[30] , \Level4Out112[29] , 
        \Level4Out112[28] , \Level4Out112[27] , \Level4Out112[26] , 
        \Level4Out112[25] , \Level4Out112[24] , \Level4Out112[23] , 
        \Level4Out112[22] , \Level4Out112[21] , \Level4Out112[20] , 
        \Level4Out112[19] , \Level4Out112[18] , \Level4Out112[17] , 
        \Level4Out112[16] , \Level4Out112[15] , \Level4Out112[14] , 
        \Level4Out112[13] , \Level4Out112[12] , \Level4Out112[11] , 
        \Level4Out112[10] , \Level4Out112[9] , \Level4Out112[8] , 
        \Level4Out112[7] , \Level4Out112[6] , \Level4Out112[5] , 
        \Level4Out112[4] , \Level4Out112[3] , \Level4Out112[2] , 
        \Level4Out112[1] , \Level4Out112[0] }), .In2({\Level4Out116[31] , 
        \Level4Out116[30] , \Level4Out116[29] , \Level4Out116[28] , 
        \Level4Out116[27] , \Level4Out116[26] , \Level4Out116[25] , 
        \Level4Out116[24] , \Level4Out116[23] , \Level4Out116[22] , 
        \Level4Out116[21] , \Level4Out116[20] , \Level4Out116[19] , 
        \Level4Out116[18] , \Level4Out116[17] , \Level4Out116[16] , 
        \Level4Out116[15] , \Level4Out116[14] , \Level4Out116[13] , 
        \Level4Out116[12] , \Level4Out116[11] , \Level4Out116[10] , 
        \Level4Out116[9] , \Level4Out116[8] , \Level4Out116[7] , 
        \Level4Out116[6] , \Level4Out116[5] , \Level4Out116[4] , 
        \Level4Out116[3] , \Level4Out116[2] , \Level4Out116[1] , 
        \Level4Out116[0] }), .Read1(\Level4Load112[0] ), .Read2(
        \Level4Load116[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_60_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load60[0] ), .Out({\Level2Out60[31] , \Level2Out60[30] , 
        \Level2Out60[29] , \Level2Out60[28] , \Level2Out60[27] , 
        \Level2Out60[26] , \Level2Out60[25] , \Level2Out60[24] , 
        \Level2Out60[23] , \Level2Out60[22] , \Level2Out60[21] , 
        \Level2Out60[20] , \Level2Out60[19] , \Level2Out60[18] , 
        \Level2Out60[17] , \Level2Out60[16] , \Level2Out60[15] , 
        \Level2Out60[14] , \Level2Out60[13] , \Level2Out60[12] , 
        \Level2Out60[11] , \Level2Out60[10] , \Level2Out60[9] , 
        \Level2Out60[8] , \Level2Out60[7] , \Level2Out60[6] , \Level2Out60[5] , 
        \Level2Out60[4] , \Level2Out60[3] , \Level2Out60[2] , \Level2Out60[1] , 
        \Level2Out60[0] }), .In1({\Level1Out60[31] , \Level1Out60[30] , 
        \Level1Out60[29] , \Level1Out60[28] , \Level1Out60[27] , 
        \Level1Out60[26] , \Level1Out60[25] , \Level1Out60[24] , 
        \Level1Out60[23] , \Level1Out60[22] , \Level1Out60[21] , 
        \Level1Out60[20] , \Level1Out60[19] , \Level1Out60[18] , 
        \Level1Out60[17] , \Level1Out60[16] , \Level1Out60[15] , 
        \Level1Out60[14] , \Level1Out60[13] , \Level1Out60[12] , 
        \Level1Out60[11] , \Level1Out60[10] , \Level1Out60[9] , 
        \Level1Out60[8] , \Level1Out60[7] , \Level1Out60[6] , \Level1Out60[5] , 
        \Level1Out60[4] , \Level1Out60[3] , \Level1Out60[2] , \Level1Out60[1] , 
        \Level1Out60[0] }), .In2({\Level1Out61[31] , \Level1Out61[30] , 
        \Level1Out61[29] , \Level1Out61[28] , \Level1Out61[27] , 
        \Level1Out61[26] , \Level1Out61[25] , \Level1Out61[24] , 
        \Level1Out61[23] , \Level1Out61[22] , \Level1Out61[21] , 
        \Level1Out61[20] , \Level1Out61[19] , \Level1Out61[18] , 
        \Level1Out61[17] , \Level1Out61[16] , \Level1Out61[15] , 
        \Level1Out61[14] , \Level1Out61[13] , \Level1Out61[12] , 
        \Level1Out61[11] , \Level1Out61[10] , \Level1Out61[9] , 
        \Level1Out61[8] , \Level1Out61[7] , \Level1Out61[6] , \Level1Out61[5] , 
        \Level1Out61[4] , \Level1Out61[3] , \Level1Out61[2] , \Level1Out61[1] , 
        \Level1Out61[0] }), .Read1(\Level1Load60[0] ), .Read2(
        \Level1Load61[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_212_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load212[0] ), .Out({\Level2Out212[31] , \Level2Out212[30] , 
        \Level2Out212[29] , \Level2Out212[28] , \Level2Out212[27] , 
        \Level2Out212[26] , \Level2Out212[25] , \Level2Out212[24] , 
        \Level2Out212[23] , \Level2Out212[22] , \Level2Out212[21] , 
        \Level2Out212[20] , \Level2Out212[19] , \Level2Out212[18] , 
        \Level2Out212[17] , \Level2Out212[16] , \Level2Out212[15] , 
        \Level2Out212[14] , \Level2Out212[13] , \Level2Out212[12] , 
        \Level2Out212[11] , \Level2Out212[10] , \Level2Out212[9] , 
        \Level2Out212[8] , \Level2Out212[7] , \Level2Out212[6] , 
        \Level2Out212[5] , \Level2Out212[4] , \Level2Out212[3] , 
        \Level2Out212[2] , \Level2Out212[1] , \Level2Out212[0] }), .In1({
        \Level1Out212[31] , \Level1Out212[30] , \Level1Out212[29] , 
        \Level1Out212[28] , \Level1Out212[27] , \Level1Out212[26] , 
        \Level1Out212[25] , \Level1Out212[24] , \Level1Out212[23] , 
        \Level1Out212[22] , \Level1Out212[21] , \Level1Out212[20] , 
        \Level1Out212[19] , \Level1Out212[18] , \Level1Out212[17] , 
        \Level1Out212[16] , \Level1Out212[15] , \Level1Out212[14] , 
        \Level1Out212[13] , \Level1Out212[12] , \Level1Out212[11] , 
        \Level1Out212[10] , \Level1Out212[9] , \Level1Out212[8] , 
        \Level1Out212[7] , \Level1Out212[6] , \Level1Out212[5] , 
        \Level1Out212[4] , \Level1Out212[3] , \Level1Out212[2] , 
        \Level1Out212[1] , \Level1Out212[0] }), .In2({\Level1Out213[31] , 
        \Level1Out213[30] , \Level1Out213[29] , \Level1Out213[28] , 
        \Level1Out213[27] , \Level1Out213[26] , \Level1Out213[25] , 
        \Level1Out213[24] , \Level1Out213[23] , \Level1Out213[22] , 
        \Level1Out213[21] , \Level1Out213[20] , \Level1Out213[19] , 
        \Level1Out213[18] , \Level1Out213[17] , \Level1Out213[16] , 
        \Level1Out213[15] , \Level1Out213[14] , \Level1Out213[13] , 
        \Level1Out213[12] , \Level1Out213[11] , \Level1Out213[10] , 
        \Level1Out213[9] , \Level1Out213[8] , \Level1Out213[7] , 
        \Level1Out213[6] , \Level1Out213[5] , \Level1Out213[4] , 
        \Level1Out213[3] , \Level1Out213[2] , \Level1Out213[1] , 
        \Level1Out213[0] }), .Read1(\Level1Load212[0] ), .Read2(
        \Level1Load213[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_230 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink230[31] , \ScanLink230[30] , 
        \ScanLink230[29] , \ScanLink230[28] , \ScanLink230[27] , 
        \ScanLink230[26] , \ScanLink230[25] , \ScanLink230[24] , 
        \ScanLink230[23] , \ScanLink230[22] , \ScanLink230[21] , 
        \ScanLink230[20] , \ScanLink230[19] , \ScanLink230[18] , 
        \ScanLink230[17] , \ScanLink230[16] , \ScanLink230[15] , 
        \ScanLink230[14] , \ScanLink230[13] , \ScanLink230[12] , 
        \ScanLink230[11] , \ScanLink230[10] , \ScanLink230[9] , 
        \ScanLink230[8] , \ScanLink230[7] , \ScanLink230[6] , \ScanLink230[5] , 
        \ScanLink230[4] , \ScanLink230[3] , \ScanLink230[2] , \ScanLink230[1] , 
        \ScanLink230[0] }), .ScanOut({\ScanLink231[31] , \ScanLink231[30] , 
        \ScanLink231[29] , \ScanLink231[28] , \ScanLink231[27] , 
        \ScanLink231[26] , \ScanLink231[25] , \ScanLink231[24] , 
        \ScanLink231[23] , \ScanLink231[22] , \ScanLink231[21] , 
        \ScanLink231[20] , \ScanLink231[19] , \ScanLink231[18] , 
        \ScanLink231[17] , \ScanLink231[16] , \ScanLink231[15] , 
        \ScanLink231[14] , \ScanLink231[13] , \ScanLink231[12] , 
        \ScanLink231[11] , \ScanLink231[10] , \ScanLink231[9] , 
        \ScanLink231[8] , \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , 
        \ScanLink231[4] , \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , 
        \ScanLink231[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load230[0] ), .Out({\Level1Out230[31] , \Level1Out230[30] , 
        \Level1Out230[29] , \Level1Out230[28] , \Level1Out230[27] , 
        \Level1Out230[26] , \Level1Out230[25] , \Level1Out230[24] , 
        \Level1Out230[23] , \Level1Out230[22] , \Level1Out230[21] , 
        \Level1Out230[20] , \Level1Out230[19] , \Level1Out230[18] , 
        \Level1Out230[17] , \Level1Out230[16] , \Level1Out230[15] , 
        \Level1Out230[14] , \Level1Out230[13] , \Level1Out230[12] , 
        \Level1Out230[11] , \Level1Out230[10] , \Level1Out230[9] , 
        \Level1Out230[8] , \Level1Out230[7] , \Level1Out230[6] , 
        \Level1Out230[5] , \Level1Out230[4] , \Level1Out230[3] , 
        \Level1Out230[2] , \Level1Out230[1] , \Level1Out230[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_126_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load126[0] ), .Out({\Level2Out126[31] , \Level2Out126[30] , 
        \Level2Out126[29] , \Level2Out126[28] , \Level2Out126[27] , 
        \Level2Out126[26] , \Level2Out126[25] , \Level2Out126[24] , 
        \Level2Out126[23] , \Level2Out126[22] , \Level2Out126[21] , 
        \Level2Out126[20] , \Level2Out126[19] , \Level2Out126[18] , 
        \Level2Out126[17] , \Level2Out126[16] , \Level2Out126[15] , 
        \Level2Out126[14] , \Level2Out126[13] , \Level2Out126[12] , 
        \Level2Out126[11] , \Level2Out126[10] , \Level2Out126[9] , 
        \Level2Out126[8] , \Level2Out126[7] , \Level2Out126[6] , 
        \Level2Out126[5] , \Level2Out126[4] , \Level2Out126[3] , 
        \Level2Out126[2] , \Level2Out126[1] , \Level2Out126[0] }), .In1({
        \Level1Out126[31] , \Level1Out126[30] , \Level1Out126[29] , 
        \Level1Out126[28] , \Level1Out126[27] , \Level1Out126[26] , 
        \Level1Out126[25] , \Level1Out126[24] , \Level1Out126[23] , 
        \Level1Out126[22] , \Level1Out126[21] , \Level1Out126[20] , 
        \Level1Out126[19] , \Level1Out126[18] , \Level1Out126[17] , 
        \Level1Out126[16] , \Level1Out126[15] , \Level1Out126[14] , 
        \Level1Out126[13] , \Level1Out126[12] , \Level1Out126[11] , 
        \Level1Out126[10] , \Level1Out126[9] , \Level1Out126[8] , 
        \Level1Out126[7] , \Level1Out126[6] , \Level1Out126[5] , 
        \Level1Out126[4] , \Level1Out126[3] , \Level1Out126[2] , 
        \Level1Out126[1] , \Level1Out126[0] }), .In2({\Level1Out127[31] , 
        \Level1Out127[30] , \Level1Out127[29] , \Level1Out127[28] , 
        \Level1Out127[27] , \Level1Out127[26] , \Level1Out127[25] , 
        \Level1Out127[24] , \Level1Out127[23] , \Level1Out127[22] , 
        \Level1Out127[21] , \Level1Out127[20] , \Level1Out127[19] , 
        \Level1Out127[18] , \Level1Out127[17] , \Level1Out127[16] , 
        \Level1Out127[15] , \Level1Out127[14] , \Level1Out127[13] , 
        \Level1Out127[12] , \Level1Out127[11] , \Level1Out127[10] , 
        \Level1Out127[9] , \Level1Out127[8] , \Level1Out127[7] , 
        \Level1Out127[6] , \Level1Out127[5] , \Level1Out127[4] , 
        \Level1Out127[3] , \Level1Out127[2] , \Level1Out127[1] , 
        \Level1Out127[0] }), .Read1(\Level1Load126[0] ), .Read2(
        \Level1Load127[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_238_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load238[0] ), .Out({\Level2Out238[31] , \Level2Out238[30] , 
        \Level2Out238[29] , \Level2Out238[28] , \Level2Out238[27] , 
        \Level2Out238[26] , \Level2Out238[25] , \Level2Out238[24] , 
        \Level2Out238[23] , \Level2Out238[22] , \Level2Out238[21] , 
        \Level2Out238[20] , \Level2Out238[19] , \Level2Out238[18] , 
        \Level2Out238[17] , \Level2Out238[16] , \Level2Out238[15] , 
        \Level2Out238[14] , \Level2Out238[13] , \Level2Out238[12] , 
        \Level2Out238[11] , \Level2Out238[10] , \Level2Out238[9] , 
        \Level2Out238[8] , \Level2Out238[7] , \Level2Out238[6] , 
        \Level2Out238[5] , \Level2Out238[4] , \Level2Out238[3] , 
        \Level2Out238[2] , \Level2Out238[1] , \Level2Out238[0] }), .In1({
        \Level1Out238[31] , \Level1Out238[30] , \Level1Out238[29] , 
        \Level1Out238[28] , \Level1Out238[27] , \Level1Out238[26] , 
        \Level1Out238[25] , \Level1Out238[24] , \Level1Out238[23] , 
        \Level1Out238[22] , \Level1Out238[21] , \Level1Out238[20] , 
        \Level1Out238[19] , \Level1Out238[18] , \Level1Out238[17] , 
        \Level1Out238[16] , \Level1Out238[15] , \Level1Out238[14] , 
        \Level1Out238[13] , \Level1Out238[12] , \Level1Out238[11] , 
        \Level1Out238[10] , \Level1Out238[9] , \Level1Out238[8] , 
        \Level1Out238[7] , \Level1Out238[6] , \Level1Out238[5] , 
        \Level1Out238[4] , \Level1Out238[3] , \Level1Out238[2] , 
        \Level1Out238[1] , \Level1Out238[0] }), .In2({\Level1Out239[31] , 
        \Level1Out239[30] , \Level1Out239[29] , \Level1Out239[28] , 
        \Level1Out239[27] , \Level1Out239[26] , \Level1Out239[25] , 
        \Level1Out239[24] , \Level1Out239[23] , \Level1Out239[22] , 
        \Level1Out239[21] , \Level1Out239[20] , \Level1Out239[19] , 
        \Level1Out239[18] , \Level1Out239[17] , \Level1Out239[16] , 
        \Level1Out239[15] , \Level1Out239[14] , \Level1Out239[13] , 
        \Level1Out239[12] , \Level1Out239[11] , \Level1Out239[10] , 
        \Level1Out239[9] , \Level1Out239[8] , \Level1Out239[7] , 
        \Level1Out239[6] , \Level1Out239[5] , \Level1Out239[4] , 
        \Level1Out239[3] , \Level1Out239[2] , \Level1Out239[1] , 
        \Level1Out239[0] }), .Read1(\Level1Load238[0] ), .Read2(
        \Level1Load239[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_224_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load224[0] ), .Out({\Level4Out224[31] , \Level4Out224[30] , 
        \Level4Out224[29] , \Level4Out224[28] , \Level4Out224[27] , 
        \Level4Out224[26] , \Level4Out224[25] , \Level4Out224[24] , 
        \Level4Out224[23] , \Level4Out224[22] , \Level4Out224[21] , 
        \Level4Out224[20] , \Level4Out224[19] , \Level4Out224[18] , 
        \Level4Out224[17] , \Level4Out224[16] , \Level4Out224[15] , 
        \Level4Out224[14] , \Level4Out224[13] , \Level4Out224[12] , 
        \Level4Out224[11] , \Level4Out224[10] , \Level4Out224[9] , 
        \Level4Out224[8] , \Level4Out224[7] , \Level4Out224[6] , 
        \Level4Out224[5] , \Level4Out224[4] , \Level4Out224[3] , 
        \Level4Out224[2] , \Level4Out224[1] , \Level4Out224[0] }), .In1({
        \Level2Out224[31] , \Level2Out224[30] , \Level2Out224[29] , 
        \Level2Out224[28] , \Level2Out224[27] , \Level2Out224[26] , 
        \Level2Out224[25] , \Level2Out224[24] , \Level2Out224[23] , 
        \Level2Out224[22] , \Level2Out224[21] , \Level2Out224[20] , 
        \Level2Out224[19] , \Level2Out224[18] , \Level2Out224[17] , 
        \Level2Out224[16] , \Level2Out224[15] , \Level2Out224[14] , 
        \Level2Out224[13] , \Level2Out224[12] , \Level2Out224[11] , 
        \Level2Out224[10] , \Level2Out224[9] , \Level2Out224[8] , 
        \Level2Out224[7] , \Level2Out224[6] , \Level2Out224[5] , 
        \Level2Out224[4] , \Level2Out224[3] , \Level2Out224[2] , 
        \Level2Out224[1] , \Level2Out224[0] }), .In2({\Level2Out226[31] , 
        \Level2Out226[30] , \Level2Out226[29] , \Level2Out226[28] , 
        \Level2Out226[27] , \Level2Out226[26] , \Level2Out226[25] , 
        \Level2Out226[24] , \Level2Out226[23] , \Level2Out226[22] , 
        \Level2Out226[21] , \Level2Out226[20] , \Level2Out226[19] , 
        \Level2Out226[18] , \Level2Out226[17] , \Level2Out226[16] , 
        \Level2Out226[15] , \Level2Out226[14] , \Level2Out226[13] , 
        \Level2Out226[12] , \Level2Out226[11] , \Level2Out226[10] , 
        \Level2Out226[9] , \Level2Out226[8] , \Level2Out226[7] , 
        \Level2Out226[6] , \Level2Out226[5] , \Level2Out226[4] , 
        \Level2Out226[3] , \Level2Out226[2] , \Level2Out226[1] , 
        \Level2Out226[0] }), .Read1(\Level2Load224[0] ), .Read2(
        \Level2Load226[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_184_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load184[0] ), .Out({\Level8Out184[31] , \Level8Out184[30] , 
        \Level8Out184[29] , \Level8Out184[28] , \Level8Out184[27] , 
        \Level8Out184[26] , \Level8Out184[25] , \Level8Out184[24] , 
        \Level8Out184[23] , \Level8Out184[22] , \Level8Out184[21] , 
        \Level8Out184[20] , \Level8Out184[19] , \Level8Out184[18] , 
        \Level8Out184[17] , \Level8Out184[16] , \Level8Out184[15] , 
        \Level8Out184[14] , \Level8Out184[13] , \Level8Out184[12] , 
        \Level8Out184[11] , \Level8Out184[10] , \Level8Out184[9] , 
        \Level8Out184[8] , \Level8Out184[7] , \Level8Out184[6] , 
        \Level8Out184[5] , \Level8Out184[4] , \Level8Out184[3] , 
        \Level8Out184[2] , \Level8Out184[1] , \Level8Out184[0] }), .In1({
        \Level4Out184[31] , \Level4Out184[30] , \Level4Out184[29] , 
        \Level4Out184[28] , \Level4Out184[27] , \Level4Out184[26] , 
        \Level4Out184[25] , \Level4Out184[24] , \Level4Out184[23] , 
        \Level4Out184[22] , \Level4Out184[21] , \Level4Out184[20] , 
        \Level4Out184[19] , \Level4Out184[18] , \Level4Out184[17] , 
        \Level4Out184[16] , \Level4Out184[15] , \Level4Out184[14] , 
        \Level4Out184[13] , \Level4Out184[12] , \Level4Out184[11] , 
        \Level4Out184[10] , \Level4Out184[9] , \Level4Out184[8] , 
        \Level4Out184[7] , \Level4Out184[6] , \Level4Out184[5] , 
        \Level4Out184[4] , \Level4Out184[3] , \Level4Out184[2] , 
        \Level4Out184[1] , \Level4Out184[0] }), .In2({\Level4Out188[31] , 
        \Level4Out188[30] , \Level4Out188[29] , \Level4Out188[28] , 
        \Level4Out188[27] , \Level4Out188[26] , \Level4Out188[25] , 
        \Level4Out188[24] , \Level4Out188[23] , \Level4Out188[22] , 
        \Level4Out188[21] , \Level4Out188[20] , \Level4Out188[19] , 
        \Level4Out188[18] , \Level4Out188[17] , \Level4Out188[16] , 
        \Level4Out188[15] , \Level4Out188[14] , \Level4Out188[13] , 
        \Level4Out188[12] , \Level4Out188[11] , \Level4Out188[10] , 
        \Level4Out188[9] , \Level4Out188[8] , \Level4Out188[7] , 
        \Level4Out188[6] , \Level4Out188[5] , \Level4Out188[4] , 
        \Level4Out188[3] , \Level4Out188[2] , \Level4Out188[1] , 
        \Level4Out188[0] }), .Read1(\Level4Load184[0] ), .Read2(
        \Level4Load188[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load56[0] ), .Out({\Level4Out56[31] , \Level4Out56[30] , 
        \Level4Out56[29] , \Level4Out56[28] , \Level4Out56[27] , 
        \Level4Out56[26] , \Level4Out56[25] , \Level4Out56[24] , 
        \Level4Out56[23] , \Level4Out56[22] , \Level4Out56[21] , 
        \Level4Out56[20] , \Level4Out56[19] , \Level4Out56[18] , 
        \Level4Out56[17] , \Level4Out56[16] , \Level4Out56[15] , 
        \Level4Out56[14] , \Level4Out56[13] , \Level4Out56[12] , 
        \Level4Out56[11] , \Level4Out56[10] , \Level4Out56[9] , 
        \Level4Out56[8] , \Level4Out56[7] , \Level4Out56[6] , \Level4Out56[5] , 
        \Level4Out56[4] , \Level4Out56[3] , \Level4Out56[2] , \Level4Out56[1] , 
        \Level4Out56[0] }), .In1({\Level2Out56[31] , \Level2Out56[30] , 
        \Level2Out56[29] , \Level2Out56[28] , \Level2Out56[27] , 
        \Level2Out56[26] , \Level2Out56[25] , \Level2Out56[24] , 
        \Level2Out56[23] , \Level2Out56[22] , \Level2Out56[21] , 
        \Level2Out56[20] , \Level2Out56[19] , \Level2Out56[18] , 
        \Level2Out56[17] , \Level2Out56[16] , \Level2Out56[15] , 
        \Level2Out56[14] , \Level2Out56[13] , \Level2Out56[12] , 
        \Level2Out56[11] , \Level2Out56[10] , \Level2Out56[9] , 
        \Level2Out56[8] , \Level2Out56[7] , \Level2Out56[6] , \Level2Out56[5] , 
        \Level2Out56[4] , \Level2Out56[3] , \Level2Out56[2] , \Level2Out56[1] , 
        \Level2Out56[0] }), .In2({\Level2Out58[31] , \Level2Out58[30] , 
        \Level2Out58[29] , \Level2Out58[28] , \Level2Out58[27] , 
        \Level2Out58[26] , \Level2Out58[25] , \Level2Out58[24] , 
        \Level2Out58[23] , \Level2Out58[22] , \Level2Out58[21] , 
        \Level2Out58[20] , \Level2Out58[19] , \Level2Out58[18] , 
        \Level2Out58[17] , \Level2Out58[16] , \Level2Out58[15] , 
        \Level2Out58[14] , \Level2Out58[13] , \Level2Out58[12] , 
        \Level2Out58[11] , \Level2Out58[10] , \Level2Out58[9] , 
        \Level2Out58[8] , \Level2Out58[7] , \Level2Out58[6] , \Level2Out58[5] , 
        \Level2Out58[4] , \Level2Out58[3] , \Level2Out58[2] , \Level2Out58[1] , 
        \Level2Out58[0] }), .Read1(\Level2Load56[0] ), .Read2(
        \Level2Load58[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanOut({\ScanLink4[31] , 
        \ScanLink4[30] , \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , 
        \ScanLink4[26] , \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , 
        \ScanLink4[22] , \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , 
        \ScanLink4[18] , \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , 
        \ScanLink4[14] , \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , 
        \ScanLink4[10] , \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , 
        \ScanLink4[6] , \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , 
        \ScanLink4[2] , \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load3[0] ), .Out({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanOut({\ScanLink5[31] , 
        \ScanLink5[30] , \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , 
        \ScanLink5[26] , \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , 
        \ScanLink5[22] , \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , 
        \ScanLink5[18] , \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , 
        \ScanLink5[14] , \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , 
        \ScanLink5[10] , \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , 
        \ScanLink5[6] , \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , 
        \ScanLink5[2] , \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load4[0] ), .Out({
        \Level1Out4[31] , \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , 
        \Level1Out4[27] , \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , 
        \Level1Out4[23] , \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , 
        \Level1Out4[19] , \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , 
        \Level1Out4[15] , \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , 
        \Level1Out4[11] , \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , 
        \Level1Out4[7] , \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , 
        \Level1Out4[3] , \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanOut({\ScanLink6[31] , 
        \ScanLink6[30] , \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , 
        \ScanLink6[26] , \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , 
        \ScanLink6[22] , \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , 
        \ScanLink6[18] , \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , 
        \ScanLink6[14] , \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , 
        \ScanLink6[10] , \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , 
        \ScanLink6[6] , \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , 
        \ScanLink6[2] , \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load5[0] ), .Out({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanOut({\ScanLink11[31] , 
        \ScanLink11[30] , \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , 
        \ScanLink11[26] , \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , 
        \ScanLink11[22] , \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , 
        \ScanLink11[18] , \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , 
        \ScanLink11[14] , \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , 
        \ScanLink11[10] , \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , 
        \ScanLink11[6] , \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , 
        \ScanLink11[2] , \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load10[0] ), .Out({
        \Level1Out10[31] , \Level1Out10[30] , \Level1Out10[29] , 
        \Level1Out10[28] , \Level1Out10[27] , \Level1Out10[26] , 
        \Level1Out10[25] , \Level1Out10[24] , \Level1Out10[23] , 
        \Level1Out10[22] , \Level1Out10[21] , \Level1Out10[20] , 
        \Level1Out10[19] , \Level1Out10[18] , \Level1Out10[17] , 
        \Level1Out10[16] , \Level1Out10[15] , \Level1Out10[14] , 
        \Level1Out10[13] , \Level1Out10[12] , \Level1Out10[11] , 
        \Level1Out10[10] , \Level1Out10[9] , \Level1Out10[8] , 
        \Level1Out10[7] , \Level1Out10[6] , \Level1Out10[5] , \Level1Out10[4] , 
        \Level1Out10[3] , \Level1Out10[2] , \Level1Out10[1] , \Level1Out10[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_17 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanOut({\ScanLink18[31] , 
        \ScanLink18[30] , \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , 
        \ScanLink18[26] , \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , 
        \ScanLink18[22] , \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , 
        \ScanLink18[18] , \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , 
        \ScanLink18[14] , \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , 
        \ScanLink18[10] , \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , 
        \ScanLink18[6] , \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , 
        \ScanLink18[2] , \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load17[0] ), .Out({
        \Level1Out17[31] , \Level1Out17[30] , \Level1Out17[29] , 
        \Level1Out17[28] , \Level1Out17[27] , \Level1Out17[26] , 
        \Level1Out17[25] , \Level1Out17[24] , \Level1Out17[23] , 
        \Level1Out17[22] , \Level1Out17[21] , \Level1Out17[20] , 
        \Level1Out17[19] , \Level1Out17[18] , \Level1Out17[17] , 
        \Level1Out17[16] , \Level1Out17[15] , \Level1Out17[14] , 
        \Level1Out17[13] , \Level1Out17[12] , \Level1Out17[11] , 
        \Level1Out17[10] , \Level1Out17[9] , \Level1Out17[8] , 
        \Level1Out17[7] , \Level1Out17[6] , \Level1Out17[5] , \Level1Out17[4] , 
        \Level1Out17[3] , \Level1Out17[2] , \Level1Out17[1] , \Level1Out17[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_30 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanOut({\ScanLink31[31] , 
        \ScanLink31[30] , \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , 
        \ScanLink31[26] , \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , 
        \ScanLink31[22] , \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , 
        \ScanLink31[18] , \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , 
        \ScanLink31[14] , \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , 
        \ScanLink31[10] , \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , 
        \ScanLink31[6] , \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , 
        \ScanLink31[2] , \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load30[0] ), .Out({
        \Level1Out30[31] , \Level1Out30[30] , \Level1Out30[29] , 
        \Level1Out30[28] , \Level1Out30[27] , \Level1Out30[26] , 
        \Level1Out30[25] , \Level1Out30[24] , \Level1Out30[23] , 
        \Level1Out30[22] , \Level1Out30[21] , \Level1Out30[20] , 
        \Level1Out30[19] , \Level1Out30[18] , \Level1Out30[17] , 
        \Level1Out30[16] , \Level1Out30[15] , \Level1Out30[14] , 
        \Level1Out30[13] , \Level1Out30[12] , \Level1Out30[11] , 
        \Level1Out30[10] , \Level1Out30[9] , \Level1Out30[8] , 
        \Level1Out30[7] , \Level1Out30[6] , \Level1Out30[5] , \Level1Out30[4] , 
        \Level1Out30[3] , \Level1Out30[2] , \Level1Out30[1] , \Level1Out30[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_39 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanOut({\ScanLink40[31] , 
        \ScanLink40[30] , \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , 
        \ScanLink40[26] , \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , 
        \ScanLink40[22] , \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , 
        \ScanLink40[18] , \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , 
        \ScanLink40[14] , \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , 
        \ScanLink40[10] , \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , 
        \ScanLink40[6] , \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , 
        \ScanLink40[2] , \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load39[0] ), .Out({
        \Level1Out39[31] , \Level1Out39[30] , \Level1Out39[29] , 
        \Level1Out39[28] , \Level1Out39[27] , \Level1Out39[26] , 
        \Level1Out39[25] , \Level1Out39[24] , \Level1Out39[23] , 
        \Level1Out39[22] , \Level1Out39[21] , \Level1Out39[20] , 
        \Level1Out39[19] , \Level1Out39[18] , \Level1Out39[17] , 
        \Level1Out39[16] , \Level1Out39[15] , \Level1Out39[14] , 
        \Level1Out39[13] , \Level1Out39[12] , \Level1Out39[11] , 
        \Level1Out39[10] , \Level1Out39[9] , \Level1Out39[8] , 
        \Level1Out39[7] , \Level1Out39[6] , \Level1Out39[5] , \Level1Out39[4] , 
        \Level1Out39[3] , \Level1Out39[2] , \Level1Out39[1] , \Level1Out39[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_57 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanOut({\ScanLink58[31] , 
        \ScanLink58[30] , \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , 
        \ScanLink58[26] , \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , 
        \ScanLink58[22] , \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , 
        \ScanLink58[18] , \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , 
        \ScanLink58[14] , \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , 
        \ScanLink58[10] , \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , 
        \ScanLink58[6] , \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , 
        \ScanLink58[2] , \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load57[0] ), .Out({
        \Level1Out57[31] , \Level1Out57[30] , \Level1Out57[29] , 
        \Level1Out57[28] , \Level1Out57[27] , \Level1Out57[26] , 
        \Level1Out57[25] , \Level1Out57[24] , \Level1Out57[23] , 
        \Level1Out57[22] , \Level1Out57[21] , \Level1Out57[20] , 
        \Level1Out57[19] , \Level1Out57[18] , \Level1Out57[17] , 
        \Level1Out57[16] , \Level1Out57[15] , \Level1Out57[14] , 
        \Level1Out57[13] , \Level1Out57[12] , \Level1Out57[11] , 
        \Level1Out57[10] , \Level1Out57[9] , \Level1Out57[8] , 
        \Level1Out57[7] , \Level1Out57[6] , \Level1Out57[5] , \Level1Out57[4] , 
        \Level1Out57[3] , \Level1Out57[2] , \Level1Out57[1] , \Level1Out57[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_149 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink149[31] , \ScanLink149[30] , 
        \ScanLink149[29] , \ScanLink149[28] , \ScanLink149[27] , 
        \ScanLink149[26] , \ScanLink149[25] , \ScanLink149[24] , 
        \ScanLink149[23] , \ScanLink149[22] , \ScanLink149[21] , 
        \ScanLink149[20] , \ScanLink149[19] , \ScanLink149[18] , 
        \ScanLink149[17] , \ScanLink149[16] , \ScanLink149[15] , 
        \ScanLink149[14] , \ScanLink149[13] , \ScanLink149[12] , 
        \ScanLink149[11] , \ScanLink149[10] , \ScanLink149[9] , 
        \ScanLink149[8] , \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , 
        \ScanLink149[4] , \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , 
        \ScanLink149[0] }), .ScanOut({\ScanLink150[31] , \ScanLink150[30] , 
        \ScanLink150[29] , \ScanLink150[28] , \ScanLink150[27] , 
        \ScanLink150[26] , \ScanLink150[25] , \ScanLink150[24] , 
        \ScanLink150[23] , \ScanLink150[22] , \ScanLink150[21] , 
        \ScanLink150[20] , \ScanLink150[19] , \ScanLink150[18] , 
        \ScanLink150[17] , \ScanLink150[16] , \ScanLink150[15] , 
        \ScanLink150[14] , \ScanLink150[13] , \ScanLink150[12] , 
        \ScanLink150[11] , \ScanLink150[10] , \ScanLink150[9] , 
        \ScanLink150[8] , \ScanLink150[7] , \ScanLink150[6] , \ScanLink150[5] , 
        \ScanLink150[4] , \ScanLink150[3] , \ScanLink150[2] , \ScanLink150[1] , 
        \ScanLink150[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load149[0] ), .Out({\Level1Out149[31] , \Level1Out149[30] , 
        \Level1Out149[29] , \Level1Out149[28] , \Level1Out149[27] , 
        \Level1Out149[26] , \Level1Out149[25] , \Level1Out149[24] , 
        \Level1Out149[23] , \Level1Out149[22] , \Level1Out149[21] , 
        \Level1Out149[20] , \Level1Out149[19] , \Level1Out149[18] , 
        \Level1Out149[17] , \Level1Out149[16] , \Level1Out149[15] , 
        \Level1Out149[14] , \Level1Out149[13] , \Level1Out149[12] , 
        \Level1Out149[11] , \Level1Out149[10] , \Level1Out149[9] , 
        \Level1Out149[8] , \Level1Out149[7] , \Level1Out149[6] , 
        \Level1Out149[5] , \Level1Out149[4] , \Level1Out149[3] , 
        \Level1Out149[2] , \Level1Out149[1] , \Level1Out149[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_144_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load144[0] ), .Out({\Level16Out144[31] , \Level16Out144[30] , 
        \Level16Out144[29] , \Level16Out144[28] , \Level16Out144[27] , 
        \Level16Out144[26] , \Level16Out144[25] , \Level16Out144[24] , 
        \Level16Out144[23] , \Level16Out144[22] , \Level16Out144[21] , 
        \Level16Out144[20] , \Level16Out144[19] , \Level16Out144[18] , 
        \Level16Out144[17] , \Level16Out144[16] , \Level16Out144[15] , 
        \Level16Out144[14] , \Level16Out144[13] , \Level16Out144[12] , 
        \Level16Out144[11] , \Level16Out144[10] , \Level16Out144[9] , 
        \Level16Out144[8] , \Level16Out144[7] , \Level16Out144[6] , 
        \Level16Out144[5] , \Level16Out144[4] , \Level16Out144[3] , 
        \Level16Out144[2] , \Level16Out144[1] , \Level16Out144[0] }), .In1({
        \Level8Out144[31] , \Level8Out144[30] , \Level8Out144[29] , 
        \Level8Out144[28] , \Level8Out144[27] , \Level8Out144[26] , 
        \Level8Out144[25] , \Level8Out144[24] , \Level8Out144[23] , 
        \Level8Out144[22] , \Level8Out144[21] , \Level8Out144[20] , 
        \Level8Out144[19] , \Level8Out144[18] , \Level8Out144[17] , 
        \Level8Out144[16] , \Level8Out144[15] , \Level8Out144[14] , 
        \Level8Out144[13] , \Level8Out144[12] , \Level8Out144[11] , 
        \Level8Out144[10] , \Level8Out144[9] , \Level8Out144[8] , 
        \Level8Out144[7] , \Level8Out144[6] , \Level8Out144[5] , 
        \Level8Out144[4] , \Level8Out144[3] , \Level8Out144[2] , 
        \Level8Out144[1] , \Level8Out144[0] }), .In2({\Level8Out152[31] , 
        \Level8Out152[30] , \Level8Out152[29] , \Level8Out152[28] , 
        \Level8Out152[27] , \Level8Out152[26] , \Level8Out152[25] , 
        \Level8Out152[24] , \Level8Out152[23] , \Level8Out152[22] , 
        \Level8Out152[21] , \Level8Out152[20] , \Level8Out152[19] , 
        \Level8Out152[18] , \Level8Out152[17] , \Level8Out152[16] , 
        \Level8Out152[15] , \Level8Out152[14] , \Level8Out152[13] , 
        \Level8Out152[12] , \Level8Out152[11] , \Level8Out152[10] , 
        \Level8Out152[9] , \Level8Out152[8] , \Level8Out152[7] , 
        \Level8Out152[6] , \Level8Out152[5] , \Level8Out152[4] , 
        \Level8Out152[3] , \Level8Out152[2] , \Level8Out152[1] , 
        \Level8Out152[0] }), .Read1(\Level8Load144[0] ), .Read2(
        \Level8Load152[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_70 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink70[31] , \ScanLink70[30] , 
        \ScanLink70[29] , \ScanLink70[28] , \ScanLink70[27] , \ScanLink70[26] , 
        \ScanLink70[25] , \ScanLink70[24] , \ScanLink70[23] , \ScanLink70[22] , 
        \ScanLink70[21] , \ScanLink70[20] , \ScanLink70[19] , \ScanLink70[18] , 
        \ScanLink70[17] , \ScanLink70[16] , \ScanLink70[15] , \ScanLink70[14] , 
        \ScanLink70[13] , \ScanLink70[12] , \ScanLink70[11] , \ScanLink70[10] , 
        \ScanLink70[9] , \ScanLink70[8] , \ScanLink70[7] , \ScanLink70[6] , 
        \ScanLink70[5] , \ScanLink70[4] , \ScanLink70[3] , \ScanLink70[2] , 
        \ScanLink70[1] , \ScanLink70[0] }), .ScanOut({\ScanLink71[31] , 
        \ScanLink71[30] , \ScanLink71[29] , \ScanLink71[28] , \ScanLink71[27] , 
        \ScanLink71[26] , \ScanLink71[25] , \ScanLink71[24] , \ScanLink71[23] , 
        \ScanLink71[22] , \ScanLink71[21] , \ScanLink71[20] , \ScanLink71[19] , 
        \ScanLink71[18] , \ScanLink71[17] , \ScanLink71[16] , \ScanLink71[15] , 
        \ScanLink71[14] , \ScanLink71[13] , \ScanLink71[12] , \ScanLink71[11] , 
        \ScanLink71[10] , \ScanLink71[9] , \ScanLink71[8] , \ScanLink71[7] , 
        \ScanLink71[6] , \ScanLink71[5] , \ScanLink71[4] , \ScanLink71[3] , 
        \ScanLink71[2] , \ScanLink71[1] , \ScanLink71[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load70[0] ), .Out({
        \Level1Out70[31] , \Level1Out70[30] , \Level1Out70[29] , 
        \Level1Out70[28] , \Level1Out70[27] , \Level1Out70[26] , 
        \Level1Out70[25] , \Level1Out70[24] , \Level1Out70[23] , 
        \Level1Out70[22] , \Level1Out70[21] , \Level1Out70[20] , 
        \Level1Out70[19] , \Level1Out70[18] , \Level1Out70[17] , 
        \Level1Out70[16] , \Level1Out70[15] , \Level1Out70[14] , 
        \Level1Out70[13] , \Level1Out70[12] , \Level1Out70[11] , 
        \Level1Out70[10] , \Level1Out70[9] , \Level1Out70[8] , 
        \Level1Out70[7] , \Level1Out70[6] , \Level1Out70[5] , \Level1Out70[4] , 
        \Level1Out70[3] , \Level1Out70[2] , \Level1Out70[1] , \Level1Out70[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_95 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink95[31] , \ScanLink95[30] , 
        \ScanLink95[29] , \ScanLink95[28] , \ScanLink95[27] , \ScanLink95[26] , 
        \ScanLink95[25] , \ScanLink95[24] , \ScanLink95[23] , \ScanLink95[22] , 
        \ScanLink95[21] , \ScanLink95[20] , \ScanLink95[19] , \ScanLink95[18] , 
        \ScanLink95[17] , \ScanLink95[16] , \ScanLink95[15] , \ScanLink95[14] , 
        \ScanLink95[13] , \ScanLink95[12] , \ScanLink95[11] , \ScanLink95[10] , 
        \ScanLink95[9] , \ScanLink95[8] , \ScanLink95[7] , \ScanLink95[6] , 
        \ScanLink95[5] , \ScanLink95[4] , \ScanLink95[3] , \ScanLink95[2] , 
        \ScanLink95[1] , \ScanLink95[0] }), .ScanOut({\ScanLink96[31] , 
        \ScanLink96[30] , \ScanLink96[29] , \ScanLink96[28] , \ScanLink96[27] , 
        \ScanLink96[26] , \ScanLink96[25] , \ScanLink96[24] , \ScanLink96[23] , 
        \ScanLink96[22] , \ScanLink96[21] , \ScanLink96[20] , \ScanLink96[19] , 
        \ScanLink96[18] , \ScanLink96[17] , \ScanLink96[16] , \ScanLink96[15] , 
        \ScanLink96[14] , \ScanLink96[13] , \ScanLink96[12] , \ScanLink96[11] , 
        \ScanLink96[10] , \ScanLink96[9] , \ScanLink96[8] , \ScanLink96[7] , 
        \ScanLink96[6] , \ScanLink96[5] , \ScanLink96[4] , \ScanLink96[3] , 
        \ScanLink96[2] , \ScanLink96[1] , \ScanLink96[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load95[0] ), .Out({
        \Level1Out95[31] , \Level1Out95[30] , \Level1Out95[29] , 
        \Level1Out95[28] , \Level1Out95[27] , \Level1Out95[26] , 
        \Level1Out95[25] , \Level1Out95[24] , \Level1Out95[23] , 
        \Level1Out95[22] , \Level1Out95[21] , \Level1Out95[20] , 
        \Level1Out95[19] , \Level1Out95[18] , \Level1Out95[17] , 
        \Level1Out95[16] , \Level1Out95[15] , \Level1Out95[14] , 
        \Level1Out95[13] , \Level1Out95[12] , \Level1Out95[11] , 
        \Level1Out95[10] , \Level1Out95[9] , \Level1Out95[8] , 
        \Level1Out95[7] , \Level1Out95[6] , \Level1Out95[5] , \Level1Out95[4] , 
        \Level1Out95[3] , \Level1Out95[2] , \Level1Out95[1] , \Level1Out95[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_152 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink152[31] , \ScanLink152[30] , 
        \ScanLink152[29] , \ScanLink152[28] , \ScanLink152[27] , 
        \ScanLink152[26] , \ScanLink152[25] , \ScanLink152[24] , 
        \ScanLink152[23] , \ScanLink152[22] , \ScanLink152[21] , 
        \ScanLink152[20] , \ScanLink152[19] , \ScanLink152[18] , 
        \ScanLink152[17] , \ScanLink152[16] , \ScanLink152[15] , 
        \ScanLink152[14] , \ScanLink152[13] , \ScanLink152[12] , 
        \ScanLink152[11] , \ScanLink152[10] , \ScanLink152[9] , 
        \ScanLink152[8] , \ScanLink152[7] , \ScanLink152[6] , \ScanLink152[5] , 
        \ScanLink152[4] , \ScanLink152[3] , \ScanLink152[2] , \ScanLink152[1] , 
        \ScanLink152[0] }), .ScanOut({\ScanLink153[31] , \ScanLink153[30] , 
        \ScanLink153[29] , \ScanLink153[28] , \ScanLink153[27] , 
        \ScanLink153[26] , \ScanLink153[25] , \ScanLink153[24] , 
        \ScanLink153[23] , \ScanLink153[22] , \ScanLink153[21] , 
        \ScanLink153[20] , \ScanLink153[19] , \ScanLink153[18] , 
        \ScanLink153[17] , \ScanLink153[16] , \ScanLink153[15] , 
        \ScanLink153[14] , \ScanLink153[13] , \ScanLink153[12] , 
        \ScanLink153[11] , \ScanLink153[10] , \ScanLink153[9] , 
        \ScanLink153[8] , \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , 
        \ScanLink153[4] , \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , 
        \ScanLink153[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load152[0] ), .Out({\Level1Out152[31] , \Level1Out152[30] , 
        \Level1Out152[29] , \Level1Out152[28] , \Level1Out152[27] , 
        \Level1Out152[26] , \Level1Out152[25] , \Level1Out152[24] , 
        \Level1Out152[23] , \Level1Out152[22] , \Level1Out152[21] , 
        \Level1Out152[20] , \Level1Out152[19] , \Level1Out152[18] , 
        \Level1Out152[17] , \Level1Out152[16] , \Level1Out152[15] , 
        \Level1Out152[14] , \Level1Out152[13] , \Level1Out152[12] , 
        \Level1Out152[11] , \Level1Out152[10] , \Level1Out152[9] , 
        \Level1Out152[8] , \Level1Out152[7] , \Level1Out152[6] , 
        \Level1Out152[5] , \Level1Out152[4] , \Level1Out152[3] , 
        \Level1Out152[2] , \Level1Out152[1] , \Level1Out152[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_175 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink175[31] , \ScanLink175[30] , 
        \ScanLink175[29] , \ScanLink175[28] , \ScanLink175[27] , 
        \ScanLink175[26] , \ScanLink175[25] , \ScanLink175[24] , 
        \ScanLink175[23] , \ScanLink175[22] , \ScanLink175[21] , 
        \ScanLink175[20] , \ScanLink175[19] , \ScanLink175[18] , 
        \ScanLink175[17] , \ScanLink175[16] , \ScanLink175[15] , 
        \ScanLink175[14] , \ScanLink175[13] , \ScanLink175[12] , 
        \ScanLink175[11] , \ScanLink175[10] , \ScanLink175[9] , 
        \ScanLink175[8] , \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , 
        \ScanLink175[4] , \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , 
        \ScanLink175[0] }), .ScanOut({\ScanLink176[31] , \ScanLink176[30] , 
        \ScanLink176[29] , \ScanLink176[28] , \ScanLink176[27] , 
        \ScanLink176[26] , \ScanLink176[25] , \ScanLink176[24] , 
        \ScanLink176[23] , \ScanLink176[22] , \ScanLink176[21] , 
        \ScanLink176[20] , \ScanLink176[19] , \ScanLink176[18] , 
        \ScanLink176[17] , \ScanLink176[16] , \ScanLink176[15] , 
        \ScanLink176[14] , \ScanLink176[13] , \ScanLink176[12] , 
        \ScanLink176[11] , \ScanLink176[10] , \ScanLink176[9] , 
        \ScanLink176[8] , \ScanLink176[7] , \ScanLink176[6] , \ScanLink176[5] , 
        \ScanLink176[4] , \ScanLink176[3] , \ScanLink176[2] , \ScanLink176[1] , 
        \ScanLink176[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load175[0] ), .Out({\Level1Out175[31] , \Level1Out175[30] , 
        \Level1Out175[29] , \Level1Out175[28] , \Level1Out175[27] , 
        \Level1Out175[26] , \Level1Out175[25] , \Level1Out175[24] , 
        \Level1Out175[23] , \Level1Out175[22] , \Level1Out175[21] , 
        \Level1Out175[20] , \Level1Out175[19] , \Level1Out175[18] , 
        \Level1Out175[17] , \Level1Out175[16] , \Level1Out175[15] , 
        \Level1Out175[14] , \Level1Out175[13] , \Level1Out175[12] , 
        \Level1Out175[11] , \Level1Out175[10] , \Level1Out175[9] , 
        \Level1Out175[8] , \Level1Out175[7] , \Level1Out175[6] , 
        \Level1Out175[5] , \Level1Out175[4] , \Level1Out175[3] , 
        \Level1Out175[2] , \Level1Out175[1] , \Level1Out175[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_245 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink245[31] , \ScanLink245[30] , 
        \ScanLink245[29] , \ScanLink245[28] , \ScanLink245[27] , 
        \ScanLink245[26] , \ScanLink245[25] , \ScanLink245[24] , 
        \ScanLink245[23] , \ScanLink245[22] , \ScanLink245[21] , 
        \ScanLink245[20] , \ScanLink245[19] , \ScanLink245[18] , 
        \ScanLink245[17] , \ScanLink245[16] , \ScanLink245[15] , 
        \ScanLink245[14] , \ScanLink245[13] , \ScanLink245[12] , 
        \ScanLink245[11] , \ScanLink245[10] , \ScanLink245[9] , 
        \ScanLink245[8] , \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , 
        \ScanLink245[4] , \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , 
        \ScanLink245[0] }), .ScanOut({\ScanLink246[31] , \ScanLink246[30] , 
        \ScanLink246[29] , \ScanLink246[28] , \ScanLink246[27] , 
        \ScanLink246[26] , \ScanLink246[25] , \ScanLink246[24] , 
        \ScanLink246[23] , \ScanLink246[22] , \ScanLink246[21] , 
        \ScanLink246[20] , \ScanLink246[19] , \ScanLink246[18] , 
        \ScanLink246[17] , \ScanLink246[16] , \ScanLink246[15] , 
        \ScanLink246[14] , \ScanLink246[13] , \ScanLink246[12] , 
        \ScanLink246[11] , \ScanLink246[10] , \ScanLink246[9] , 
        \ScanLink246[8] , \ScanLink246[7] , \ScanLink246[6] , \ScanLink246[5] , 
        \ScanLink246[4] , \ScanLink246[3] , \ScanLink246[2] , \ScanLink246[1] , 
        \ScanLink246[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load245[0] ), .Out({\Level1Out245[31] , \Level1Out245[30] , 
        \Level1Out245[29] , \Level1Out245[28] , \Level1Out245[27] , 
        \Level1Out245[26] , \Level1Out245[25] , \Level1Out245[24] , 
        \Level1Out245[23] , \Level1Out245[22] , \Level1Out245[21] , 
        \Level1Out245[20] , \Level1Out245[19] , \Level1Out245[18] , 
        \Level1Out245[17] , \Level1Out245[16] , \Level1Out245[15] , 
        \Level1Out245[14] , \Level1Out245[13] , \Level1Out245[12] , 
        \Level1Out245[11] , \Level1Out245[10] , \Level1Out245[9] , 
        \Level1Out245[8] , \Level1Out245[7] , \Level1Out245[6] , 
        \Level1Out245[5] , \Level1Out245[4] , \Level1Out245[3] , 
        \Level1Out245[2] , \Level1Out245[1] , \Level1Out245[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_182_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load182[0] ), .Out({\Level2Out182[31] , \Level2Out182[30] , 
        \Level2Out182[29] , \Level2Out182[28] , \Level2Out182[27] , 
        \Level2Out182[26] , \Level2Out182[25] , \Level2Out182[24] , 
        \Level2Out182[23] , \Level2Out182[22] , \Level2Out182[21] , 
        \Level2Out182[20] , \Level2Out182[19] , \Level2Out182[18] , 
        \Level2Out182[17] , \Level2Out182[16] , \Level2Out182[15] , 
        \Level2Out182[14] , \Level2Out182[13] , \Level2Out182[12] , 
        \Level2Out182[11] , \Level2Out182[10] , \Level2Out182[9] , 
        \Level2Out182[8] , \Level2Out182[7] , \Level2Out182[6] , 
        \Level2Out182[5] , \Level2Out182[4] , \Level2Out182[3] , 
        \Level2Out182[2] , \Level2Out182[1] , \Level2Out182[0] }), .In1({
        \Level1Out182[31] , \Level1Out182[30] , \Level1Out182[29] , 
        \Level1Out182[28] , \Level1Out182[27] , \Level1Out182[26] , 
        \Level1Out182[25] , \Level1Out182[24] , \Level1Out182[23] , 
        \Level1Out182[22] , \Level1Out182[21] , \Level1Out182[20] , 
        \Level1Out182[19] , \Level1Out182[18] , \Level1Out182[17] , 
        \Level1Out182[16] , \Level1Out182[15] , \Level1Out182[14] , 
        \Level1Out182[13] , \Level1Out182[12] , \Level1Out182[11] , 
        \Level1Out182[10] , \Level1Out182[9] , \Level1Out182[8] , 
        \Level1Out182[7] , \Level1Out182[6] , \Level1Out182[5] , 
        \Level1Out182[4] , \Level1Out182[3] , \Level1Out182[2] , 
        \Level1Out182[1] , \Level1Out182[0] }), .In2({\Level1Out183[31] , 
        \Level1Out183[30] , \Level1Out183[29] , \Level1Out183[28] , 
        \Level1Out183[27] , \Level1Out183[26] , \Level1Out183[25] , 
        \Level1Out183[24] , \Level1Out183[23] , \Level1Out183[22] , 
        \Level1Out183[21] , \Level1Out183[20] , \Level1Out183[19] , 
        \Level1Out183[18] , \Level1Out183[17] , \Level1Out183[16] , 
        \Level1Out183[15] , \Level1Out183[14] , \Level1Out183[13] , 
        \Level1Out183[12] , \Level1Out183[11] , \Level1Out183[10] , 
        \Level1Out183[9] , \Level1Out183[8] , \Level1Out183[7] , 
        \Level1Out183[6] , \Level1Out183[5] , \Level1Out183[4] , 
        \Level1Out183[3] , \Level1Out183[2] , \Level1Out183[1] , 
        \Level1Out183[0] }), .Read1(\Level1Load182[0] ), .Read2(
        \Level1Load183[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_120_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load120[0] ), .Out({\Level8Out120[31] , \Level8Out120[30] , 
        \Level8Out120[29] , \Level8Out120[28] , \Level8Out120[27] , 
        \Level8Out120[26] , \Level8Out120[25] , \Level8Out120[24] , 
        \Level8Out120[23] , \Level8Out120[22] , \Level8Out120[21] , 
        \Level8Out120[20] , \Level8Out120[19] , \Level8Out120[18] , 
        \Level8Out120[17] , \Level8Out120[16] , \Level8Out120[15] , 
        \Level8Out120[14] , \Level8Out120[13] , \Level8Out120[12] , 
        \Level8Out120[11] , \Level8Out120[10] , \Level8Out120[9] , 
        \Level8Out120[8] , \Level8Out120[7] , \Level8Out120[6] , 
        \Level8Out120[5] , \Level8Out120[4] , \Level8Out120[3] , 
        \Level8Out120[2] , \Level8Out120[1] , \Level8Out120[0] }), .In1({
        \Level4Out120[31] , \Level4Out120[30] , \Level4Out120[29] , 
        \Level4Out120[28] , \Level4Out120[27] , \Level4Out120[26] , 
        \Level4Out120[25] , \Level4Out120[24] , \Level4Out120[23] , 
        \Level4Out120[22] , \Level4Out120[21] , \Level4Out120[20] , 
        \Level4Out120[19] , \Level4Out120[18] , \Level4Out120[17] , 
        \Level4Out120[16] , \Level4Out120[15] , \Level4Out120[14] , 
        \Level4Out120[13] , \Level4Out120[12] , \Level4Out120[11] , 
        \Level4Out120[10] , \Level4Out120[9] , \Level4Out120[8] , 
        \Level4Out120[7] , \Level4Out120[6] , \Level4Out120[5] , 
        \Level4Out120[4] , \Level4Out120[3] , \Level4Out120[2] , 
        \Level4Out120[1] , \Level4Out120[0] }), .In2({\Level4Out124[31] , 
        \Level4Out124[30] , \Level4Out124[29] , \Level4Out124[28] , 
        \Level4Out124[27] , \Level4Out124[26] , \Level4Out124[25] , 
        \Level4Out124[24] , \Level4Out124[23] , \Level4Out124[22] , 
        \Level4Out124[21] , \Level4Out124[20] , \Level4Out124[19] , 
        \Level4Out124[18] , \Level4Out124[17] , \Level4Out124[16] , 
        \Level4Out124[15] , \Level4Out124[14] , \Level4Out124[13] , 
        \Level4Out124[12] , \Level4Out124[11] , \Level4Out124[10] , 
        \Level4Out124[9] , \Level4Out124[8] , \Level4Out124[7] , 
        \Level4Out124[6] , \Level4Out124[5] , \Level4Out124[4] , 
        \Level4Out124[3] , \Level4Out124[2] , \Level4Out124[1] , 
        \Level4Out124[0] }), .Read1(\Level4Load120[0] ), .Read2(
        \Level4Load124[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_190 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink190[31] , \ScanLink190[30] , 
        \ScanLink190[29] , \ScanLink190[28] , \ScanLink190[27] , 
        \ScanLink190[26] , \ScanLink190[25] , \ScanLink190[24] , 
        \ScanLink190[23] , \ScanLink190[22] , \ScanLink190[21] , 
        \ScanLink190[20] , \ScanLink190[19] , \ScanLink190[18] , 
        \ScanLink190[17] , \ScanLink190[16] , \ScanLink190[15] , 
        \ScanLink190[14] , \ScanLink190[13] , \ScanLink190[12] , 
        \ScanLink190[11] , \ScanLink190[10] , \ScanLink190[9] , 
        \ScanLink190[8] , \ScanLink190[7] , \ScanLink190[6] , \ScanLink190[5] , 
        \ScanLink190[4] , \ScanLink190[3] , \ScanLink190[2] , \ScanLink190[1] , 
        \ScanLink190[0] }), .ScanOut({\ScanLink191[31] , \ScanLink191[30] , 
        \ScanLink191[29] , \ScanLink191[28] , \ScanLink191[27] , 
        \ScanLink191[26] , \ScanLink191[25] , \ScanLink191[24] , 
        \ScanLink191[23] , \ScanLink191[22] , \ScanLink191[21] , 
        \ScanLink191[20] , \ScanLink191[19] , \ScanLink191[18] , 
        \ScanLink191[17] , \ScanLink191[16] , \ScanLink191[15] , 
        \ScanLink191[14] , \ScanLink191[13] , \ScanLink191[12] , 
        \ScanLink191[11] , \ScanLink191[10] , \ScanLink191[9] , 
        \ScanLink191[8] , \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , 
        \ScanLink191[4] , \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , 
        \ScanLink191[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load190[0] ), .Out({\Level1Out190[31] , \Level1Out190[30] , 
        \Level1Out190[29] , \Level1Out190[28] , \Level1Out190[27] , 
        \Level1Out190[26] , \Level1Out190[25] , \Level1Out190[24] , 
        \Level1Out190[23] , \Level1Out190[22] , \Level1Out190[21] , 
        \Level1Out190[20] , \Level1Out190[19] , \Level1Out190[18] , 
        \Level1Out190[17] , \Level1Out190[16] , \Level1Out190[15] , 
        \Level1Out190[14] , \Level1Out190[13] , \Level1Out190[12] , 
        \Level1Out190[11] , \Level1Out190[10] , \Level1Out190[9] , 
        \Level1Out190[8] , \Level1Out190[7] , \Level1Out190[6] , 
        \Level1Out190[5] , \Level1Out190[4] , \Level1Out190[3] , 
        \Level1Out190[2] , \Level1Out190[1] , \Level1Out190[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_114_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load114[0] ), .Out({\Level2Out114[31] , \Level2Out114[30] , 
        \Level2Out114[29] , \Level2Out114[28] , \Level2Out114[27] , 
        \Level2Out114[26] , \Level2Out114[25] , \Level2Out114[24] , 
        \Level2Out114[23] , \Level2Out114[22] , \Level2Out114[21] , 
        \Level2Out114[20] , \Level2Out114[19] , \Level2Out114[18] , 
        \Level2Out114[17] , \Level2Out114[16] , \Level2Out114[15] , 
        \Level2Out114[14] , \Level2Out114[13] , \Level2Out114[12] , 
        \Level2Out114[11] , \Level2Out114[10] , \Level2Out114[9] , 
        \Level2Out114[8] , \Level2Out114[7] , \Level2Out114[6] , 
        \Level2Out114[5] , \Level2Out114[4] , \Level2Out114[3] , 
        \Level2Out114[2] , \Level2Out114[1] , \Level2Out114[0] }), .In1({
        \Level1Out114[31] , \Level1Out114[30] , \Level1Out114[29] , 
        \Level1Out114[28] , \Level1Out114[27] , \Level1Out114[26] , 
        \Level1Out114[25] , \Level1Out114[24] , \Level1Out114[23] , 
        \Level1Out114[22] , \Level1Out114[21] , \Level1Out114[20] , 
        \Level1Out114[19] , \Level1Out114[18] , \Level1Out114[17] , 
        \Level1Out114[16] , \Level1Out114[15] , \Level1Out114[14] , 
        \Level1Out114[13] , \Level1Out114[12] , \Level1Out114[11] , 
        \Level1Out114[10] , \Level1Out114[9] , \Level1Out114[8] , 
        \Level1Out114[7] , \Level1Out114[6] , \Level1Out114[5] , 
        \Level1Out114[4] , \Level1Out114[3] , \Level1Out114[2] , 
        \Level1Out114[1] , \Level1Out114[0] }), .In2({\Level1Out115[31] , 
        \Level1Out115[30] , \Level1Out115[29] , \Level1Out115[28] , 
        \Level1Out115[27] , \Level1Out115[26] , \Level1Out115[25] , 
        \Level1Out115[24] , \Level1Out115[23] , \Level1Out115[22] , 
        \Level1Out115[21] , \Level1Out115[20] , \Level1Out115[19] , 
        \Level1Out115[18] , \Level1Out115[17] , \Level1Out115[16] , 
        \Level1Out115[15] , \Level1Out115[14] , \Level1Out115[13] , 
        \Level1Out115[12] , \Level1Out115[11] , \Level1Out115[10] , 
        \Level1Out115[9] , \Level1Out115[8] , \Level1Out115[7] , 
        \Level1Out115[6] , \Level1Out115[5] , \Level1Out115[4] , 
        \Level1Out115[3] , \Level1Out115[2] , \Level1Out115[1] , 
        \Level1Out115[0] }), .Read1(\Level1Load114[0] ), .Read2(
        \Level1Load115[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level128Load0[0] ), .Out({\Level128Out0[31] , \Level128Out0[30] , 
        \Level128Out0[29] , \Level128Out0[28] , \Level128Out0[27] , 
        \Level128Out0[26] , \Level128Out0[25] , \Level128Out0[24] , 
        \Level128Out0[23] , \Level128Out0[22] , \Level128Out0[21] , 
        \Level128Out0[20] , \Level128Out0[19] , \Level128Out0[18] , 
        \Level128Out0[17] , \Level128Out0[16] , \Level128Out0[15] , 
        \Level128Out0[14] , \Level128Out0[13] , \Level128Out0[12] , 
        \Level128Out0[11] , \Level128Out0[10] , \Level128Out0[9] , 
        \Level128Out0[8] , \Level128Out0[7] , \Level128Out0[6] , 
        \Level128Out0[5] , \Level128Out0[4] , \Level128Out0[3] , 
        \Level128Out0[2] , \Level128Out0[1] , \Level128Out0[0] }), .In1({
        \Level64Out0[31] , \Level64Out0[30] , \Level64Out0[29] , 
        \Level64Out0[28] , \Level64Out0[27] , \Level64Out0[26] , 
        \Level64Out0[25] , \Level64Out0[24] , \Level64Out0[23] , 
        \Level64Out0[22] , \Level64Out0[21] , \Level64Out0[20] , 
        \Level64Out0[19] , \Level64Out0[18] , \Level64Out0[17] , 
        \Level64Out0[16] , \Level64Out0[15] , \Level64Out0[14] , 
        \Level64Out0[13] , \Level64Out0[12] , \Level64Out0[11] , 
        \Level64Out0[10] , \Level64Out0[9] , \Level64Out0[8] , 
        \Level64Out0[7] , \Level64Out0[6] , \Level64Out0[5] , \Level64Out0[4] , 
        \Level64Out0[3] , \Level64Out0[2] , \Level64Out0[1] , \Level64Out0[0] 
        }), .In2({\Level64Out64[31] , \Level64Out64[30] , \Level64Out64[29] , 
        \Level64Out64[28] , \Level64Out64[27] , \Level64Out64[26] , 
        \Level64Out64[25] , \Level64Out64[24] , \Level64Out64[23] , 
        \Level64Out64[22] , \Level64Out64[21] , \Level64Out64[20] , 
        \Level64Out64[19] , \Level64Out64[18] , \Level64Out64[17] , 
        \Level64Out64[16] , \Level64Out64[15] , \Level64Out64[14] , 
        \Level64Out64[13] , \Level64Out64[12] , \Level64Out64[11] , 
        \Level64Out64[10] , \Level64Out64[9] , \Level64Out64[8] , 
        \Level64Out64[7] , \Level64Out64[6] , \Level64Out64[5] , 
        \Level64Out64[4] , \Level64Out64[3] , \Level64Out64[2] , 
        \Level64Out64[1] , \Level64Out64[0] }), .Read1(\Level64Load0[0] ), 
        .Read2(\Level64Load64[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load64[0] ), .Out({\Level4Out64[31] , \Level4Out64[30] , 
        \Level4Out64[29] , \Level4Out64[28] , \Level4Out64[27] , 
        \Level4Out64[26] , \Level4Out64[25] , \Level4Out64[24] , 
        \Level4Out64[23] , \Level4Out64[22] , \Level4Out64[21] , 
        \Level4Out64[20] , \Level4Out64[19] , \Level4Out64[18] , 
        \Level4Out64[17] , \Level4Out64[16] , \Level4Out64[15] , 
        \Level4Out64[14] , \Level4Out64[13] , \Level4Out64[12] , 
        \Level4Out64[11] , \Level4Out64[10] , \Level4Out64[9] , 
        \Level4Out64[8] , \Level4Out64[7] , \Level4Out64[6] , \Level4Out64[5] , 
        \Level4Out64[4] , \Level4Out64[3] , \Level4Out64[2] , \Level4Out64[1] , 
        \Level4Out64[0] }), .In1({\Level2Out64[31] , \Level2Out64[30] , 
        \Level2Out64[29] , \Level2Out64[28] , \Level2Out64[27] , 
        \Level2Out64[26] , \Level2Out64[25] , \Level2Out64[24] , 
        \Level2Out64[23] , \Level2Out64[22] , \Level2Out64[21] , 
        \Level2Out64[20] , \Level2Out64[19] , \Level2Out64[18] , 
        \Level2Out64[17] , \Level2Out64[16] , \Level2Out64[15] , 
        \Level2Out64[14] , \Level2Out64[13] , \Level2Out64[12] , 
        \Level2Out64[11] , \Level2Out64[10] , \Level2Out64[9] , 
        \Level2Out64[8] , \Level2Out64[7] , \Level2Out64[6] , \Level2Out64[5] , 
        \Level2Out64[4] , \Level2Out64[3] , \Level2Out64[2] , \Level2Out64[1] , 
        \Level2Out64[0] }), .In2({\Level2Out66[31] , \Level2Out66[30] , 
        \Level2Out66[29] , \Level2Out66[28] , \Level2Out66[27] , 
        \Level2Out66[26] , \Level2Out66[25] , \Level2Out66[24] , 
        \Level2Out66[23] , \Level2Out66[22] , \Level2Out66[21] , 
        \Level2Out66[20] , \Level2Out66[19] , \Level2Out66[18] , 
        \Level2Out66[17] , \Level2Out66[16] , \Level2Out66[15] , 
        \Level2Out66[14] , \Level2Out66[13] , \Level2Out66[12] , 
        \Level2Out66[11] , \Level2Out66[10] , \Level2Out66[9] , 
        \Level2Out66[8] , \Level2Out66[7] , \Level2Out66[6] , \Level2Out66[5] , 
        \Level2Out66[4] , \Level2Out66[3] , \Level2Out66[2] , \Level2Out66[1] , 
        \Level2Out66[0] }), .Read1(\Level2Load64[0] ), .Read2(
        \Level2Load66[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_108_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load108[0] ), .Out({\Level4Out108[31] , \Level4Out108[30] , 
        \Level4Out108[29] , \Level4Out108[28] , \Level4Out108[27] , 
        \Level4Out108[26] , \Level4Out108[25] , \Level4Out108[24] , 
        \Level4Out108[23] , \Level4Out108[22] , \Level4Out108[21] , 
        \Level4Out108[20] , \Level4Out108[19] , \Level4Out108[18] , 
        \Level4Out108[17] , \Level4Out108[16] , \Level4Out108[15] , 
        \Level4Out108[14] , \Level4Out108[13] , \Level4Out108[12] , 
        \Level4Out108[11] , \Level4Out108[10] , \Level4Out108[9] , 
        \Level4Out108[8] , \Level4Out108[7] , \Level4Out108[6] , 
        \Level4Out108[5] , \Level4Out108[4] , \Level4Out108[3] , 
        \Level4Out108[2] , \Level4Out108[1] , \Level4Out108[0] }), .In1({
        \Level2Out108[31] , \Level2Out108[30] , \Level2Out108[29] , 
        \Level2Out108[28] , \Level2Out108[27] , \Level2Out108[26] , 
        \Level2Out108[25] , \Level2Out108[24] , \Level2Out108[23] , 
        \Level2Out108[22] , \Level2Out108[21] , \Level2Out108[20] , 
        \Level2Out108[19] , \Level2Out108[18] , \Level2Out108[17] , 
        \Level2Out108[16] , \Level2Out108[15] , \Level2Out108[14] , 
        \Level2Out108[13] , \Level2Out108[12] , \Level2Out108[11] , 
        \Level2Out108[10] , \Level2Out108[9] , \Level2Out108[8] , 
        \Level2Out108[7] , \Level2Out108[6] , \Level2Out108[5] , 
        \Level2Out108[4] , \Level2Out108[3] , \Level2Out108[2] , 
        \Level2Out108[1] , \Level2Out108[0] }), .In2({\Level2Out110[31] , 
        \Level2Out110[30] , \Level2Out110[29] , \Level2Out110[28] , 
        \Level2Out110[27] , \Level2Out110[26] , \Level2Out110[25] , 
        \Level2Out110[24] , \Level2Out110[23] , \Level2Out110[22] , 
        \Level2Out110[21] , \Level2Out110[20] , \Level2Out110[19] , 
        \Level2Out110[18] , \Level2Out110[17] , \Level2Out110[16] , 
        \Level2Out110[15] , \Level2Out110[14] , \Level2Out110[13] , 
        \Level2Out110[12] , \Level2Out110[11] , \Level2Out110[10] , 
        \Level2Out110[9] , \Level2Out110[8] , \Level2Out110[7] , 
        \Level2Out110[6] , \Level2Out110[5] , \Level2Out110[4] , 
        \Level2Out110[3] , \Level2Out110[2] , \Level2Out110[1] , 
        \Level2Out110[0] }), .Read1(\Level2Load108[0] ), .Read2(
        \Level2Load110[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_216_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load216[0] ), .Out({\Level4Out216[31] , \Level4Out216[30] , 
        \Level4Out216[29] , \Level4Out216[28] , \Level4Out216[27] , 
        \Level4Out216[26] , \Level4Out216[25] , \Level4Out216[24] , 
        \Level4Out216[23] , \Level4Out216[22] , \Level4Out216[21] , 
        \Level4Out216[20] , \Level4Out216[19] , \Level4Out216[18] , 
        \Level4Out216[17] , \Level4Out216[16] , \Level4Out216[15] , 
        \Level4Out216[14] , \Level4Out216[13] , \Level4Out216[12] , 
        \Level4Out216[11] , \Level4Out216[10] , \Level4Out216[9] , 
        \Level4Out216[8] , \Level4Out216[7] , \Level4Out216[6] , 
        \Level4Out216[5] , \Level4Out216[4] , \Level4Out216[3] , 
        \Level4Out216[2] , \Level4Out216[1] , \Level4Out216[0] }), .In1({
        \Level2Out216[31] , \Level2Out216[30] , \Level2Out216[29] , 
        \Level2Out216[28] , \Level2Out216[27] , \Level2Out216[26] , 
        \Level2Out216[25] , \Level2Out216[24] , \Level2Out216[23] , 
        \Level2Out216[22] , \Level2Out216[21] , \Level2Out216[20] , 
        \Level2Out216[19] , \Level2Out216[18] , \Level2Out216[17] , 
        \Level2Out216[16] , \Level2Out216[15] , \Level2Out216[14] , 
        \Level2Out216[13] , \Level2Out216[12] , \Level2Out216[11] , 
        \Level2Out216[10] , \Level2Out216[9] , \Level2Out216[8] , 
        \Level2Out216[7] , \Level2Out216[6] , \Level2Out216[5] , 
        \Level2Out216[4] , \Level2Out216[3] , \Level2Out216[2] , 
        \Level2Out216[1] , \Level2Out216[0] }), .In2({\Level2Out218[31] , 
        \Level2Out218[30] , \Level2Out218[29] , \Level2Out218[28] , 
        \Level2Out218[27] , \Level2Out218[26] , \Level2Out218[25] , 
        \Level2Out218[24] , \Level2Out218[23] , \Level2Out218[22] , 
        \Level2Out218[21] , \Level2Out218[20] , \Level2Out218[19] , 
        \Level2Out218[18] , \Level2Out218[17] , \Level2Out218[16] , 
        \Level2Out218[15] , \Level2Out218[14] , \Level2Out218[13] , 
        \Level2Out218[12] , \Level2Out218[11] , \Level2Out218[10] , 
        \Level2Out218[9] , \Level2Out218[8] , \Level2Out218[7] , 
        \Level2Out218[6] , \Level2Out218[5] , \Level2Out218[4] , 
        \Level2Out218[3] , \Level2Out218[2] , \Level2Out218[1] , 
        \Level2Out218[0] }), .Read1(\Level2Load216[0] ), .Read2(
        \Level2Load218[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_78_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load78[0] ), .Out({\Level2Out78[31] , \Level2Out78[30] , 
        \Level2Out78[29] , \Level2Out78[28] , \Level2Out78[27] , 
        \Level2Out78[26] , \Level2Out78[25] , \Level2Out78[24] , 
        \Level2Out78[23] , \Level2Out78[22] , \Level2Out78[21] , 
        \Level2Out78[20] , \Level2Out78[19] , \Level2Out78[18] , 
        \Level2Out78[17] , \Level2Out78[16] , \Level2Out78[15] , 
        \Level2Out78[14] , \Level2Out78[13] , \Level2Out78[12] , 
        \Level2Out78[11] , \Level2Out78[10] , \Level2Out78[9] , 
        \Level2Out78[8] , \Level2Out78[7] , \Level2Out78[6] , \Level2Out78[5] , 
        \Level2Out78[4] , \Level2Out78[3] , \Level2Out78[2] , \Level2Out78[1] , 
        \Level2Out78[0] }), .In1({\Level1Out78[31] , \Level1Out78[30] , 
        \Level1Out78[29] , \Level1Out78[28] , \Level1Out78[27] , 
        \Level1Out78[26] , \Level1Out78[25] , \Level1Out78[24] , 
        \Level1Out78[23] , \Level1Out78[22] , \Level1Out78[21] , 
        \Level1Out78[20] , \Level1Out78[19] , \Level1Out78[18] , 
        \Level1Out78[17] , \Level1Out78[16] , \Level1Out78[15] , 
        \Level1Out78[14] , \Level1Out78[13] , \Level1Out78[12] , 
        \Level1Out78[11] , \Level1Out78[10] , \Level1Out78[9] , 
        \Level1Out78[8] , \Level1Out78[7] , \Level1Out78[6] , \Level1Out78[5] , 
        \Level1Out78[4] , \Level1Out78[3] , \Level1Out78[2] , \Level1Out78[1] , 
        \Level1Out78[0] }), .In2({\Level1Out79[31] , \Level1Out79[30] , 
        \Level1Out79[29] , \Level1Out79[28] , \Level1Out79[27] , 
        \Level1Out79[26] , \Level1Out79[25] , \Level1Out79[24] , 
        \Level1Out79[23] , \Level1Out79[22] , \Level1Out79[21] , 
        \Level1Out79[20] , \Level1Out79[19] , \Level1Out79[18] , 
        \Level1Out79[17] , \Level1Out79[16] , \Level1Out79[15] , 
        \Level1Out79[14] , \Level1Out79[13] , \Level1Out79[12] , 
        \Level1Out79[11] , \Level1Out79[10] , \Level1Out79[9] , 
        \Level1Out79[8] , \Level1Out79[7] , \Level1Out79[6] , \Level1Out79[5] , 
        \Level1Out79[4] , \Level1Out79[3] , \Level1Out79[2] , \Level1Out79[1] , 
        \Level1Out79[0] }), .Read1(\Level1Load78[0] ), .Read2(
        \Level1Load79[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_45 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanOut({\ScanLink46[31] , 
        \ScanLink46[30] , \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , 
        \ScanLink46[26] , \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , 
        \ScanLink46[22] , \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , 
        \ScanLink46[18] , \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , 
        \ScanLink46[14] , \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , 
        \ScanLink46[10] , \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , 
        \ScanLink46[6] , \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , 
        \ScanLink46[2] , \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load45[0] ), .Out({
        \Level1Out45[31] , \Level1Out45[30] , \Level1Out45[29] , 
        \Level1Out45[28] , \Level1Out45[27] , \Level1Out45[26] , 
        \Level1Out45[25] , \Level1Out45[24] , \Level1Out45[23] , 
        \Level1Out45[22] , \Level1Out45[21] , \Level1Out45[20] , 
        \Level1Out45[19] , \Level1Out45[18] , \Level1Out45[17] , 
        \Level1Out45[16] , \Level1Out45[15] , \Level1Out45[14] , 
        \Level1Out45[13] , \Level1Out45[12] , \Level1Out45[11] , 
        \Level1Out45[10] , \Level1Out45[9] , \Level1Out45[8] , 
        \Level1Out45[7] , \Level1Out45[6] , \Level1Out45[5] , \Level1Out45[4] , 
        \Level1Out45[3] , \Level1Out45[2] , \Level1Out45[1] , \Level1Out45[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_87 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink87[31] , \ScanLink87[30] , 
        \ScanLink87[29] , \ScanLink87[28] , \ScanLink87[27] , \ScanLink87[26] , 
        \ScanLink87[25] , \ScanLink87[24] , \ScanLink87[23] , \ScanLink87[22] , 
        \ScanLink87[21] , \ScanLink87[20] , \ScanLink87[19] , \ScanLink87[18] , 
        \ScanLink87[17] , \ScanLink87[16] , \ScanLink87[15] , \ScanLink87[14] , 
        \ScanLink87[13] , \ScanLink87[12] , \ScanLink87[11] , \ScanLink87[10] , 
        \ScanLink87[9] , \ScanLink87[8] , \ScanLink87[7] , \ScanLink87[6] , 
        \ScanLink87[5] , \ScanLink87[4] , \ScanLink87[3] , \ScanLink87[2] , 
        \ScanLink87[1] , \ScanLink87[0] }), .ScanOut({\ScanLink88[31] , 
        \ScanLink88[30] , \ScanLink88[29] , \ScanLink88[28] , \ScanLink88[27] , 
        \ScanLink88[26] , \ScanLink88[25] , \ScanLink88[24] , \ScanLink88[23] , 
        \ScanLink88[22] , \ScanLink88[21] , \ScanLink88[20] , \ScanLink88[19] , 
        \ScanLink88[18] , \ScanLink88[17] , \ScanLink88[16] , \ScanLink88[15] , 
        \ScanLink88[14] , \ScanLink88[13] , \ScanLink88[12] , \ScanLink88[11] , 
        \ScanLink88[10] , \ScanLink88[9] , \ScanLink88[8] , \ScanLink88[7] , 
        \ScanLink88[6] , \ScanLink88[5] , \ScanLink88[4] , \ScanLink88[3] , 
        \ScanLink88[2] , \ScanLink88[1] , \ScanLink88[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load87[0] ), .Out({
        \Level1Out87[31] , \Level1Out87[30] , \Level1Out87[29] , 
        \Level1Out87[28] , \Level1Out87[27] , \Level1Out87[26] , 
        \Level1Out87[25] , \Level1Out87[24] , \Level1Out87[23] , 
        \Level1Out87[22] , \Level1Out87[21] , \Level1Out87[20] , 
        \Level1Out87[19] , \Level1Out87[18] , \Level1Out87[17] , 
        \Level1Out87[16] , \Level1Out87[15] , \Level1Out87[14] , 
        \Level1Out87[13] , \Level1Out87[12] , \Level1Out87[11] , 
        \Level1Out87[10] , \Level1Out87[9] , \Level1Out87[8] , 
        \Level1Out87[7] , \Level1Out87[6] , \Level1Out87[5] , \Level1Out87[4] , 
        \Level1Out87[3] , \Level1Out87[2] , \Level1Out87[1] , \Level1Out87[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_109 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink109[31] , \ScanLink109[30] , 
        \ScanLink109[29] , \ScanLink109[28] , \ScanLink109[27] , 
        \ScanLink109[26] , \ScanLink109[25] , \ScanLink109[24] , 
        \ScanLink109[23] , \ScanLink109[22] , \ScanLink109[21] , 
        \ScanLink109[20] , \ScanLink109[19] , \ScanLink109[18] , 
        \ScanLink109[17] , \ScanLink109[16] , \ScanLink109[15] , 
        \ScanLink109[14] , \ScanLink109[13] , \ScanLink109[12] , 
        \ScanLink109[11] , \ScanLink109[10] , \ScanLink109[9] , 
        \ScanLink109[8] , \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , 
        \ScanLink109[4] , \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , 
        \ScanLink109[0] }), .ScanOut({\ScanLink110[31] , \ScanLink110[30] , 
        \ScanLink110[29] , \ScanLink110[28] , \ScanLink110[27] , 
        \ScanLink110[26] , \ScanLink110[25] , \ScanLink110[24] , 
        \ScanLink110[23] , \ScanLink110[22] , \ScanLink110[21] , 
        \ScanLink110[20] , \ScanLink110[19] , \ScanLink110[18] , 
        \ScanLink110[17] , \ScanLink110[16] , \ScanLink110[15] , 
        \ScanLink110[14] , \ScanLink110[13] , \ScanLink110[12] , 
        \ScanLink110[11] , \ScanLink110[10] , \ScanLink110[9] , 
        \ScanLink110[8] , \ScanLink110[7] , \ScanLink110[6] , \ScanLink110[5] , 
        \ScanLink110[4] , \ScanLink110[3] , \ScanLink110[2] , \ScanLink110[1] , 
        \ScanLink110[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load109[0] ), .Out({\Level1Out109[31] , \Level1Out109[30] , 
        \Level1Out109[29] , \Level1Out109[28] , \Level1Out109[27] , 
        \Level1Out109[26] , \Level1Out109[25] , \Level1Out109[24] , 
        \Level1Out109[23] , \Level1Out109[22] , \Level1Out109[21] , 
        \Level1Out109[20] , \Level1Out109[19] , \Level1Out109[18] , 
        \Level1Out109[17] , \Level1Out109[16] , \Level1Out109[15] , 
        \Level1Out109[14] , \Level1Out109[13] , \Level1Out109[12] , 
        \Level1Out109[11] , \Level1Out109[10] , \Level1Out109[9] , 
        \Level1Out109[8] , \Level1Out109[7] , \Level1Out109[6] , 
        \Level1Out109[5] , \Level1Out109[4] , \Level1Out109[3] , 
        \Level1Out109[2] , \Level1Out109[1] , \Level1Out109[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_182 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink182[31] , \ScanLink182[30] , 
        \ScanLink182[29] , \ScanLink182[28] , \ScanLink182[27] , 
        \ScanLink182[26] , \ScanLink182[25] , \ScanLink182[24] , 
        \ScanLink182[23] , \ScanLink182[22] , \ScanLink182[21] , 
        \ScanLink182[20] , \ScanLink182[19] , \ScanLink182[18] , 
        \ScanLink182[17] , \ScanLink182[16] , \ScanLink182[15] , 
        \ScanLink182[14] , \ScanLink182[13] , \ScanLink182[12] , 
        \ScanLink182[11] , \ScanLink182[10] , \ScanLink182[9] , 
        \ScanLink182[8] , \ScanLink182[7] , \ScanLink182[6] , \ScanLink182[5] , 
        \ScanLink182[4] , \ScanLink182[3] , \ScanLink182[2] , \ScanLink182[1] , 
        \ScanLink182[0] }), .ScanOut({\ScanLink183[31] , \ScanLink183[30] , 
        \ScanLink183[29] , \ScanLink183[28] , \ScanLink183[27] , 
        \ScanLink183[26] , \ScanLink183[25] , \ScanLink183[24] , 
        \ScanLink183[23] , \ScanLink183[22] , \ScanLink183[21] , 
        \ScanLink183[20] , \ScanLink183[19] , \ScanLink183[18] , 
        \ScanLink183[17] , \ScanLink183[16] , \ScanLink183[15] , 
        \ScanLink183[14] , \ScanLink183[13] , \ScanLink183[12] , 
        \ScanLink183[11] , \ScanLink183[10] , \ScanLink183[9] , 
        \ScanLink183[8] , \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , 
        \ScanLink183[4] , \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , 
        \ScanLink183[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load182[0] ), .Out({\Level1Out182[31] , \Level1Out182[30] , 
        \Level1Out182[29] , \Level1Out182[28] , \Level1Out182[27] , 
        \Level1Out182[26] , \Level1Out182[25] , \Level1Out182[24] , 
        \Level1Out182[23] , \Level1Out182[22] , \Level1Out182[21] , 
        \Level1Out182[20] , \Level1Out182[19] , \Level1Out182[18] , 
        \Level1Out182[17] , \Level1Out182[16] , \Level1Out182[15] , 
        \Level1Out182[14] , \Level1Out182[13] , \Level1Out182[12] , 
        \Level1Out182[11] , \Level1Out182[10] , \Level1Out182[9] , 
        \Level1Out182[8] , \Level1Out182[7] , \Level1Out182[6] , 
        \Level1Out182[5] , \Level1Out182[4] , \Level1Out182[3] , 
        \Level1Out182[2] , \Level1Out182[1] , \Level1Out182[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_52_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load52[0] ), .Out({\Level2Out52[31] , \Level2Out52[30] , 
        \Level2Out52[29] , \Level2Out52[28] , \Level2Out52[27] , 
        \Level2Out52[26] , \Level2Out52[25] , \Level2Out52[24] , 
        \Level2Out52[23] , \Level2Out52[22] , \Level2Out52[21] , 
        \Level2Out52[20] , \Level2Out52[19] , \Level2Out52[18] , 
        \Level2Out52[17] , \Level2Out52[16] , \Level2Out52[15] , 
        \Level2Out52[14] , \Level2Out52[13] , \Level2Out52[12] , 
        \Level2Out52[11] , \Level2Out52[10] , \Level2Out52[9] , 
        \Level2Out52[8] , \Level2Out52[7] , \Level2Out52[6] , \Level2Out52[5] , 
        \Level2Out52[4] , \Level2Out52[3] , \Level2Out52[2] , \Level2Out52[1] , 
        \Level2Out52[0] }), .In1({\Level1Out52[31] , \Level1Out52[30] , 
        \Level1Out52[29] , \Level1Out52[28] , \Level1Out52[27] , 
        \Level1Out52[26] , \Level1Out52[25] , \Level1Out52[24] , 
        \Level1Out52[23] , \Level1Out52[22] , \Level1Out52[21] , 
        \Level1Out52[20] , \Level1Out52[19] , \Level1Out52[18] , 
        \Level1Out52[17] , \Level1Out52[16] , \Level1Out52[15] , 
        \Level1Out52[14] , \Level1Out52[13] , \Level1Out52[12] , 
        \Level1Out52[11] , \Level1Out52[10] , \Level1Out52[9] , 
        \Level1Out52[8] , \Level1Out52[7] , \Level1Out52[6] , \Level1Out52[5] , 
        \Level1Out52[4] , \Level1Out52[3] , \Level1Out52[2] , \Level1Out52[1] , 
        \Level1Out52[0] }), .In2({\Level1Out53[31] , \Level1Out53[30] , 
        \Level1Out53[29] , \Level1Out53[28] , \Level1Out53[27] , 
        \Level1Out53[26] , \Level1Out53[25] , \Level1Out53[24] , 
        \Level1Out53[23] , \Level1Out53[22] , \Level1Out53[21] , 
        \Level1Out53[20] , \Level1Out53[19] , \Level1Out53[18] , 
        \Level1Out53[17] , \Level1Out53[16] , \Level1Out53[15] , 
        \Level1Out53[14] , \Level1Out53[13] , \Level1Out53[12] , 
        \Level1Out53[11] , \Level1Out53[10] , \Level1Out53[9] , 
        \Level1Out53[8] , \Level1Out53[7] , \Level1Out53[6] , \Level1Out53[5] , 
        \Level1Out53[4] , \Level1Out53[3] , \Level1Out53[2] , \Level1Out53[1] , 
        \Level1Out53[0] }), .Read1(\Level1Load52[0] ), .Read2(
        \Level1Load53[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_220_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load220[0] ), .Out({\Level2Out220[31] , \Level2Out220[30] , 
        \Level2Out220[29] , \Level2Out220[28] , \Level2Out220[27] , 
        \Level2Out220[26] , \Level2Out220[25] , \Level2Out220[24] , 
        \Level2Out220[23] , \Level2Out220[22] , \Level2Out220[21] , 
        \Level2Out220[20] , \Level2Out220[19] , \Level2Out220[18] , 
        \Level2Out220[17] , \Level2Out220[16] , \Level2Out220[15] , 
        \Level2Out220[14] , \Level2Out220[13] , \Level2Out220[12] , 
        \Level2Out220[11] , \Level2Out220[10] , \Level2Out220[9] , 
        \Level2Out220[8] , \Level2Out220[7] , \Level2Out220[6] , 
        \Level2Out220[5] , \Level2Out220[4] , \Level2Out220[3] , 
        \Level2Out220[2] , \Level2Out220[1] , \Level2Out220[0] }), .In1({
        \Level1Out220[31] , \Level1Out220[30] , \Level1Out220[29] , 
        \Level1Out220[28] , \Level1Out220[27] , \Level1Out220[26] , 
        \Level1Out220[25] , \Level1Out220[24] , \Level1Out220[23] , 
        \Level1Out220[22] , \Level1Out220[21] , \Level1Out220[20] , 
        \Level1Out220[19] , \Level1Out220[18] , \Level1Out220[17] , 
        \Level1Out220[16] , \Level1Out220[15] , \Level1Out220[14] , 
        \Level1Out220[13] , \Level1Out220[12] , \Level1Out220[11] , 
        \Level1Out220[10] , \Level1Out220[9] , \Level1Out220[8] , 
        \Level1Out220[7] , \Level1Out220[6] , \Level1Out220[5] , 
        \Level1Out220[4] , \Level1Out220[3] , \Level1Out220[2] , 
        \Level1Out220[1] , \Level1Out220[0] }), .In2({\Level1Out221[31] , 
        \Level1Out221[30] , \Level1Out221[29] , \Level1Out221[28] , 
        \Level1Out221[27] , \Level1Out221[26] , \Level1Out221[25] , 
        \Level1Out221[24] , \Level1Out221[23] , \Level1Out221[22] , 
        \Level1Out221[21] , \Level1Out221[20] , \Level1Out221[19] , 
        \Level1Out221[18] , \Level1Out221[17] , \Level1Out221[16] , 
        \Level1Out221[15] , \Level1Out221[14] , \Level1Out221[13] , 
        \Level1Out221[12] , \Level1Out221[11] , \Level1Out221[10] , 
        \Level1Out221[9] , \Level1Out221[8] , \Level1Out221[7] , 
        \Level1Out221[6] , \Level1Out221[5] , \Level1Out221[4] , 
        \Level1Out221[3] , \Level1Out221[2] , \Level1Out221[1] , 
        \Level1Out221[0] }), .Read1(\Level1Load220[0] ), .Read2(
        \Level1Load221[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_239 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink239[31] , \ScanLink239[30] , 
        \ScanLink239[29] , \ScanLink239[28] , \ScanLink239[27] , 
        \ScanLink239[26] , \ScanLink239[25] , \ScanLink239[24] , 
        \ScanLink239[23] , \ScanLink239[22] , \ScanLink239[21] , 
        \ScanLink239[20] , \ScanLink239[19] , \ScanLink239[18] , 
        \ScanLink239[17] , \ScanLink239[16] , \ScanLink239[15] , 
        \ScanLink239[14] , \ScanLink239[13] , \ScanLink239[12] , 
        \ScanLink239[11] , \ScanLink239[10] , \ScanLink239[9] , 
        \ScanLink239[8] , \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , 
        \ScanLink239[4] , \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , 
        \ScanLink239[0] }), .ScanOut({\ScanLink240[31] , \ScanLink240[30] , 
        \ScanLink240[29] , \ScanLink240[28] , \ScanLink240[27] , 
        \ScanLink240[26] , \ScanLink240[25] , \ScanLink240[24] , 
        \ScanLink240[23] , \ScanLink240[22] , \ScanLink240[21] , 
        \ScanLink240[20] , \ScanLink240[19] , \ScanLink240[18] , 
        \ScanLink240[17] , \ScanLink240[16] , \ScanLink240[15] , 
        \ScanLink240[14] , \ScanLink240[13] , \ScanLink240[12] , 
        \ScanLink240[11] , \ScanLink240[10] , \ScanLink240[9] , 
        \ScanLink240[8] , \ScanLink240[7] , \ScanLink240[6] , \ScanLink240[5] , 
        \ScanLink240[4] , \ScanLink240[3] , \ScanLink240[2] , \ScanLink240[1] , 
        \ScanLink240[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load239[0] ), .Out({\Level1Out239[31] , \Level1Out239[30] , 
        \Level1Out239[29] , \Level1Out239[28] , \Level1Out239[27] , 
        \Level1Out239[26] , \Level1Out239[25] , \Level1Out239[24] , 
        \Level1Out239[23] , \Level1Out239[22] , \Level1Out239[21] , 
        \Level1Out239[20] , \Level1Out239[19] , \Level1Out239[18] , 
        \Level1Out239[17] , \Level1Out239[16] , \Level1Out239[15] , 
        \Level1Out239[14] , \Level1Out239[13] , \Level1Out239[12] , 
        \Level1Out239[11] , \Level1Out239[10] , \Level1Out239[9] , 
        \Level1Out239[8] , \Level1Out239[7] , \Level1Out239[6] , 
        \Level1Out239[5] , \Level1Out239[4] , \Level1Out239[3] , 
        \Level1Out239[2] , \Level1Out239[1] , \Level1Out239[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load64[0] ), .Out({\Level16Out64[31] , \Level16Out64[30] , 
        \Level16Out64[29] , \Level16Out64[28] , \Level16Out64[27] , 
        \Level16Out64[26] , \Level16Out64[25] , \Level16Out64[24] , 
        \Level16Out64[23] , \Level16Out64[22] , \Level16Out64[21] , 
        \Level16Out64[20] , \Level16Out64[19] , \Level16Out64[18] , 
        \Level16Out64[17] , \Level16Out64[16] , \Level16Out64[15] , 
        \Level16Out64[14] , \Level16Out64[13] , \Level16Out64[12] , 
        \Level16Out64[11] , \Level16Out64[10] , \Level16Out64[9] , 
        \Level16Out64[8] , \Level16Out64[7] , \Level16Out64[6] , 
        \Level16Out64[5] , \Level16Out64[4] , \Level16Out64[3] , 
        \Level16Out64[2] , \Level16Out64[1] , \Level16Out64[0] }), .In1({
        \Level8Out64[31] , \Level8Out64[30] , \Level8Out64[29] , 
        \Level8Out64[28] , \Level8Out64[27] , \Level8Out64[26] , 
        \Level8Out64[25] , \Level8Out64[24] , \Level8Out64[23] , 
        \Level8Out64[22] , \Level8Out64[21] , \Level8Out64[20] , 
        \Level8Out64[19] , \Level8Out64[18] , \Level8Out64[17] , 
        \Level8Out64[16] , \Level8Out64[15] , \Level8Out64[14] , 
        \Level8Out64[13] , \Level8Out64[12] , \Level8Out64[11] , 
        \Level8Out64[10] , \Level8Out64[9] , \Level8Out64[8] , 
        \Level8Out64[7] , \Level8Out64[6] , \Level8Out64[5] , \Level8Out64[4] , 
        \Level8Out64[3] , \Level8Out64[2] , \Level8Out64[1] , \Level8Out64[0] 
        }), .In2({\Level8Out72[31] , \Level8Out72[30] , \Level8Out72[29] , 
        \Level8Out72[28] , \Level8Out72[27] , \Level8Out72[26] , 
        \Level8Out72[25] , \Level8Out72[24] , \Level8Out72[23] , 
        \Level8Out72[22] , \Level8Out72[21] , \Level8Out72[20] , 
        \Level8Out72[19] , \Level8Out72[18] , \Level8Out72[17] , 
        \Level8Out72[16] , \Level8Out72[15] , \Level8Out72[14] , 
        \Level8Out72[13] , \Level8Out72[12] , \Level8Out72[11] , 
        \Level8Out72[10] , \Level8Out72[9] , \Level8Out72[8] , 
        \Level8Out72[7] , \Level8Out72[6] , \Level8Out72[5] , \Level8Out72[4] , 
        \Level8Out72[3] , \Level8Out72[2] , \Level8Out72[1] , \Level8Out72[0] 
        }), .Read1(\Level8Load64[0] ), .Read2(\Level8Load72[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_140 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink140[31] , \ScanLink140[30] , 
        \ScanLink140[29] , \ScanLink140[28] , \ScanLink140[27] , 
        \ScanLink140[26] , \ScanLink140[25] , \ScanLink140[24] , 
        \ScanLink140[23] , \ScanLink140[22] , \ScanLink140[21] , 
        \ScanLink140[20] , \ScanLink140[19] , \ScanLink140[18] , 
        \ScanLink140[17] , \ScanLink140[16] , \ScanLink140[15] , 
        \ScanLink140[14] , \ScanLink140[13] , \ScanLink140[12] , 
        \ScanLink140[11] , \ScanLink140[10] , \ScanLink140[9] , 
        \ScanLink140[8] , \ScanLink140[7] , \ScanLink140[6] , \ScanLink140[5] , 
        \ScanLink140[4] , \ScanLink140[3] , \ScanLink140[2] , \ScanLink140[1] , 
        \ScanLink140[0] }), .ScanOut({\ScanLink141[31] , \ScanLink141[30] , 
        \ScanLink141[29] , \ScanLink141[28] , \ScanLink141[27] , 
        \ScanLink141[26] , \ScanLink141[25] , \ScanLink141[24] , 
        \ScanLink141[23] , \ScanLink141[22] , \ScanLink141[21] , 
        \ScanLink141[20] , \ScanLink141[19] , \ScanLink141[18] , 
        \ScanLink141[17] , \ScanLink141[16] , \ScanLink141[15] , 
        \ScanLink141[14] , \ScanLink141[13] , \ScanLink141[12] , 
        \ScanLink141[11] , \ScanLink141[10] , \ScanLink141[9] , 
        \ScanLink141[8] , \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , 
        \ScanLink141[4] , \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , 
        \ScanLink141[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load140[0] ), .Out({\Level1Out140[31] , \Level1Out140[30] , 
        \Level1Out140[29] , \Level1Out140[28] , \Level1Out140[27] , 
        \Level1Out140[26] , \Level1Out140[25] , \Level1Out140[24] , 
        \Level1Out140[23] , \Level1Out140[22] , \Level1Out140[21] , 
        \Level1Out140[20] , \Level1Out140[19] , \Level1Out140[18] , 
        \Level1Out140[17] , \Level1Out140[16] , \Level1Out140[15] , 
        \Level1Out140[14] , \Level1Out140[13] , \Level1Out140[12] , 
        \Level1Out140[11] , \Level1Out140[10] , \Level1Out140[9] , 
        \Level1Out140[8] , \Level1Out140[7] , \Level1Out140[6] , 
        \Level1Out140[5] , \Level1Out140[4] , \Level1Out140[3] , 
        \Level1Out140[2] , \Level1Out140[1] , \Level1Out140[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_167 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink167[31] , \ScanLink167[30] , 
        \ScanLink167[29] , \ScanLink167[28] , \ScanLink167[27] , 
        \ScanLink167[26] , \ScanLink167[25] , \ScanLink167[24] , 
        \ScanLink167[23] , \ScanLink167[22] , \ScanLink167[21] , 
        \ScanLink167[20] , \ScanLink167[19] , \ScanLink167[18] , 
        \ScanLink167[17] , \ScanLink167[16] , \ScanLink167[15] , 
        \ScanLink167[14] , \ScanLink167[13] , \ScanLink167[12] , 
        \ScanLink167[11] , \ScanLink167[10] , \ScanLink167[9] , 
        \ScanLink167[8] , \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , 
        \ScanLink167[4] , \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , 
        \ScanLink167[0] }), .ScanOut({\ScanLink168[31] , \ScanLink168[30] , 
        \ScanLink168[29] , \ScanLink168[28] , \ScanLink168[27] , 
        \ScanLink168[26] , \ScanLink168[25] , \ScanLink168[24] , 
        \ScanLink168[23] , \ScanLink168[22] , \ScanLink168[21] , 
        \ScanLink168[20] , \ScanLink168[19] , \ScanLink168[18] , 
        \ScanLink168[17] , \ScanLink168[16] , \ScanLink168[15] , 
        \ScanLink168[14] , \ScanLink168[13] , \ScanLink168[12] , 
        \ScanLink168[11] , \ScanLink168[10] , \ScanLink168[9] , 
        \ScanLink168[8] , \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , 
        \ScanLink168[4] , \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , 
        \ScanLink168[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load167[0] ), .Out({\Level1Out167[31] , \Level1Out167[30] , 
        \Level1Out167[29] , \Level1Out167[28] , \Level1Out167[27] , 
        \Level1Out167[26] , \Level1Out167[25] , \Level1Out167[24] , 
        \Level1Out167[23] , \Level1Out167[22] , \Level1Out167[21] , 
        \Level1Out167[20] , \Level1Out167[19] , \Level1Out167[18] , 
        \Level1Out167[17] , \Level1Out167[16] , \Level1Out167[15] , 
        \Level1Out167[14] , \Level1Out167[13] , \Level1Out167[12] , 
        \Level1Out167[11] , \Level1Out167[10] , \Level1Out167[9] , 
        \Level1Out167[8] , \Level1Out167[7] , \Level1Out167[6] , 
        \Level1Out167[5] , \Level1Out167[4] , \Level1Out167[3] , 
        \Level1Out167[2] , \Level1Out167[1] , \Level1Out167[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_28_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load28[0] ), .Out({\Level2Out28[31] , \Level2Out28[30] , 
        \Level2Out28[29] , \Level2Out28[28] , \Level2Out28[27] , 
        \Level2Out28[26] , \Level2Out28[25] , \Level2Out28[24] , 
        \Level2Out28[23] , \Level2Out28[22] , \Level2Out28[21] , 
        \Level2Out28[20] , \Level2Out28[19] , \Level2Out28[18] , 
        \Level2Out28[17] , \Level2Out28[16] , \Level2Out28[15] , 
        \Level2Out28[14] , \Level2Out28[13] , \Level2Out28[12] , 
        \Level2Out28[11] , \Level2Out28[10] , \Level2Out28[9] , 
        \Level2Out28[8] , \Level2Out28[7] , \Level2Out28[6] , \Level2Out28[5] , 
        \Level2Out28[4] , \Level2Out28[3] , \Level2Out28[2] , \Level2Out28[1] , 
        \Level2Out28[0] }), .In1({\Level1Out28[31] , \Level1Out28[30] , 
        \Level1Out28[29] , \Level1Out28[28] , \Level1Out28[27] , 
        \Level1Out28[26] , \Level1Out28[25] , \Level1Out28[24] , 
        \Level1Out28[23] , \Level1Out28[22] , \Level1Out28[21] , 
        \Level1Out28[20] , \Level1Out28[19] , \Level1Out28[18] , 
        \Level1Out28[17] , \Level1Out28[16] , \Level1Out28[15] , 
        \Level1Out28[14] , \Level1Out28[13] , \Level1Out28[12] , 
        \Level1Out28[11] , \Level1Out28[10] , \Level1Out28[9] , 
        \Level1Out28[8] , \Level1Out28[7] , \Level1Out28[6] , \Level1Out28[5] , 
        \Level1Out28[4] , \Level1Out28[3] , \Level1Out28[2] , \Level1Out28[1] , 
        \Level1Out28[0] }), .In2({\Level1Out29[31] , \Level1Out29[30] , 
        \Level1Out29[29] , \Level1Out29[28] , \Level1Out29[27] , 
        \Level1Out29[26] , \Level1Out29[25] , \Level1Out29[24] , 
        \Level1Out29[23] , \Level1Out29[22] , \Level1Out29[21] , 
        \Level1Out29[20] , \Level1Out29[19] , \Level1Out29[18] , 
        \Level1Out29[17] , \Level1Out29[16] , \Level1Out29[15] , 
        \Level1Out29[14] , \Level1Out29[13] , \Level1Out29[12] , 
        \Level1Out29[11] , \Level1Out29[10] , \Level1Out29[9] , 
        \Level1Out29[8] , \Level1Out29[7] , \Level1Out29[6] , \Level1Out29[5] , 
        \Level1Out29[4] , \Level1Out29[3] , \Level1Out29[2] , \Level1Out29[1] , 
        \Level1Out29[0] }), .Read1(\Level1Load28[0] ), .Read2(
        \Level1Load29[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_172_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load172[0] ), .Out({\Level4Out172[31] , \Level4Out172[30] , 
        \Level4Out172[29] , \Level4Out172[28] , \Level4Out172[27] , 
        \Level4Out172[26] , \Level4Out172[25] , \Level4Out172[24] , 
        \Level4Out172[23] , \Level4Out172[22] , \Level4Out172[21] , 
        \Level4Out172[20] , \Level4Out172[19] , \Level4Out172[18] , 
        \Level4Out172[17] , \Level4Out172[16] , \Level4Out172[15] , 
        \Level4Out172[14] , \Level4Out172[13] , \Level4Out172[12] , 
        \Level4Out172[11] , \Level4Out172[10] , \Level4Out172[9] , 
        \Level4Out172[8] , \Level4Out172[7] , \Level4Out172[6] , 
        \Level4Out172[5] , \Level4Out172[4] , \Level4Out172[3] , 
        \Level4Out172[2] , \Level4Out172[1] , \Level4Out172[0] }), .In1({
        \Level2Out172[31] , \Level2Out172[30] , \Level2Out172[29] , 
        \Level2Out172[28] , \Level2Out172[27] , \Level2Out172[26] , 
        \Level2Out172[25] , \Level2Out172[24] , \Level2Out172[23] , 
        \Level2Out172[22] , \Level2Out172[21] , \Level2Out172[20] , 
        \Level2Out172[19] , \Level2Out172[18] , \Level2Out172[17] , 
        \Level2Out172[16] , \Level2Out172[15] , \Level2Out172[14] , 
        \Level2Out172[13] , \Level2Out172[12] , \Level2Out172[11] , 
        \Level2Out172[10] , \Level2Out172[9] , \Level2Out172[8] , 
        \Level2Out172[7] , \Level2Out172[6] , \Level2Out172[5] , 
        \Level2Out172[4] , \Level2Out172[3] , \Level2Out172[2] , 
        \Level2Out172[1] , \Level2Out172[0] }), .In2({\Level2Out174[31] , 
        \Level2Out174[30] , \Level2Out174[29] , \Level2Out174[28] , 
        \Level2Out174[27] , \Level2Out174[26] , \Level2Out174[25] , 
        \Level2Out174[24] , \Level2Out174[23] , \Level2Out174[22] , 
        \Level2Out174[21] , \Level2Out174[20] , \Level2Out174[19] , 
        \Level2Out174[18] , \Level2Out174[17] , \Level2Out174[16] , 
        \Level2Out174[15] , \Level2Out174[14] , \Level2Out174[13] , 
        \Level2Out174[12] , \Level2Out174[11] , \Level2Out174[10] , 
        \Level2Out174[9] , \Level2Out174[8] , \Level2Out174[7] , 
        \Level2Out174[6] , \Level2Out174[5] , \Level2Out174[4] , 
        \Level2Out174[3] , \Level2Out174[2] , \Level2Out174[1] , 
        \Level2Out174[0] }), .Read1(\Level2Load172[0] ), .Read2(
        \Level2Load174[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_144_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load144[0] ), .Out({\Level2Out144[31] , \Level2Out144[30] , 
        \Level2Out144[29] , \Level2Out144[28] , \Level2Out144[27] , 
        \Level2Out144[26] , \Level2Out144[25] , \Level2Out144[24] , 
        \Level2Out144[23] , \Level2Out144[22] , \Level2Out144[21] , 
        \Level2Out144[20] , \Level2Out144[19] , \Level2Out144[18] , 
        \Level2Out144[17] , \Level2Out144[16] , \Level2Out144[15] , 
        \Level2Out144[14] , \Level2Out144[13] , \Level2Out144[12] , 
        \Level2Out144[11] , \Level2Out144[10] , \Level2Out144[9] , 
        \Level2Out144[8] , \Level2Out144[7] , \Level2Out144[6] , 
        \Level2Out144[5] , \Level2Out144[4] , \Level2Out144[3] , 
        \Level2Out144[2] , \Level2Out144[1] , \Level2Out144[0] }), .In1({
        \Level1Out144[31] , \Level1Out144[30] , \Level1Out144[29] , 
        \Level1Out144[28] , \Level1Out144[27] , \Level1Out144[26] , 
        \Level1Out144[25] , \Level1Out144[24] , \Level1Out144[23] , 
        \Level1Out144[22] , \Level1Out144[21] , \Level1Out144[20] , 
        \Level1Out144[19] , \Level1Out144[18] , \Level1Out144[17] , 
        \Level1Out144[16] , \Level1Out144[15] , \Level1Out144[14] , 
        \Level1Out144[13] , \Level1Out144[12] , \Level1Out144[11] , 
        \Level1Out144[10] , \Level1Out144[9] , \Level1Out144[8] , 
        \Level1Out144[7] , \Level1Out144[6] , \Level1Out144[5] , 
        \Level1Out144[4] , \Level1Out144[3] , \Level1Out144[2] , 
        \Level1Out144[1] , \Level1Out144[0] }), .In2({\Level1Out145[31] , 
        \Level1Out145[30] , \Level1Out145[29] , \Level1Out145[28] , 
        \Level1Out145[27] , \Level1Out145[26] , \Level1Out145[25] , 
        \Level1Out145[24] , \Level1Out145[23] , \Level1Out145[22] , 
        \Level1Out145[21] , \Level1Out145[20] , \Level1Out145[19] , 
        \Level1Out145[18] , \Level1Out145[17] , \Level1Out145[16] , 
        \Level1Out145[15] , \Level1Out145[14] , \Level1Out145[13] , 
        \Level1Out145[12] , \Level1Out145[11] , \Level1Out145[10] , 
        \Level1Out145[9] , \Level1Out145[8] , \Level1Out145[7] , 
        \Level1Out145[6] , \Level1Out145[5] , \Level1Out145[4] , 
        \Level1Out145[3] , \Level1Out145[2] , \Level1Out145[1] , 
        \Level1Out145[0] }), .Read1(\Level1Load144[0] ), .Read2(
        \Level1Load145[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_88_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load88[0] ), .Out({\Level4Out88[31] , \Level4Out88[30] , 
        \Level4Out88[29] , \Level4Out88[28] , \Level4Out88[27] , 
        \Level4Out88[26] , \Level4Out88[25] , \Level4Out88[24] , 
        \Level4Out88[23] , \Level4Out88[22] , \Level4Out88[21] , 
        \Level4Out88[20] , \Level4Out88[19] , \Level4Out88[18] , 
        \Level4Out88[17] , \Level4Out88[16] , \Level4Out88[15] , 
        \Level4Out88[14] , \Level4Out88[13] , \Level4Out88[12] , 
        \Level4Out88[11] , \Level4Out88[10] , \Level4Out88[9] , 
        \Level4Out88[8] , \Level4Out88[7] , \Level4Out88[6] , \Level4Out88[5] , 
        \Level4Out88[4] , \Level4Out88[3] , \Level4Out88[2] , \Level4Out88[1] , 
        \Level4Out88[0] }), .In1({\Level2Out88[31] , \Level2Out88[30] , 
        \Level2Out88[29] , \Level2Out88[28] , \Level2Out88[27] , 
        \Level2Out88[26] , \Level2Out88[25] , \Level2Out88[24] , 
        \Level2Out88[23] , \Level2Out88[22] , \Level2Out88[21] , 
        \Level2Out88[20] , \Level2Out88[19] , \Level2Out88[18] , 
        \Level2Out88[17] , \Level2Out88[16] , \Level2Out88[15] , 
        \Level2Out88[14] , \Level2Out88[13] , \Level2Out88[12] , 
        \Level2Out88[11] , \Level2Out88[10] , \Level2Out88[9] , 
        \Level2Out88[8] , \Level2Out88[7] , \Level2Out88[6] , \Level2Out88[5] , 
        \Level2Out88[4] , \Level2Out88[3] , \Level2Out88[2] , \Level2Out88[1] , 
        \Level2Out88[0] }), .In2({\Level2Out90[31] , \Level2Out90[30] , 
        \Level2Out90[29] , \Level2Out90[28] , \Level2Out90[27] , 
        \Level2Out90[26] , \Level2Out90[25] , \Level2Out90[24] , 
        \Level2Out90[23] , \Level2Out90[22] , \Level2Out90[21] , 
        \Level2Out90[20] , \Level2Out90[19] , \Level2Out90[18] , 
        \Level2Out90[17] , \Level2Out90[16] , \Level2Out90[15] , 
        \Level2Out90[14] , \Level2Out90[13] , \Level2Out90[12] , 
        \Level2Out90[11] , \Level2Out90[10] , \Level2Out90[9] , 
        \Level2Out90[8] , \Level2Out90[7] , \Level2Out90[6] , \Level2Out90[5] , 
        \Level2Out90[4] , \Level2Out90[3] , \Level2Out90[2] , \Level2Out90[1] , 
        \Level2Out90[0] }), .Read1(\Level2Load88[0] ), .Read2(
        \Level2Load90[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_62 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanOut({\ScanLink63[31] , 
        \ScanLink63[30] , \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , 
        \ScanLink63[26] , \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , 
        \ScanLink63[22] , \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , 
        \ScanLink63[18] , \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , 
        \ScanLink63[14] , \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , 
        \ScanLink63[10] , \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , 
        \ScanLink63[6] , \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , 
        \ScanLink63[2] , \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load62[0] ), .Out({
        \Level1Out62[31] , \Level1Out62[30] , \Level1Out62[29] , 
        \Level1Out62[28] , \Level1Out62[27] , \Level1Out62[26] , 
        \Level1Out62[25] , \Level1Out62[24] , \Level1Out62[23] , 
        \Level1Out62[22] , \Level1Out62[21] , \Level1Out62[20] , 
        \Level1Out62[19] , \Level1Out62[18] , \Level1Out62[17] , 
        \Level1Out62[16] , \Level1Out62[15] , \Level1Out62[14] , 
        \Level1Out62[13] , \Level1Out62[12] , \Level1Out62[11] , 
        \Level1Out62[10] , \Level1Out62[9] , \Level1Out62[8] , 
        \Level1Out62[7] , \Level1Out62[6] , \Level1Out62[5] , \Level1Out62[4] , 
        \Level1Out62[3] , \Level1Out62[2] , \Level1Out62[1] , \Level1Out62[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_94_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load94[0] ), .Out({\Level2Out94[31] , \Level2Out94[30] , 
        \Level2Out94[29] , \Level2Out94[28] , \Level2Out94[27] , 
        \Level2Out94[26] , \Level2Out94[25] , \Level2Out94[24] , 
        \Level2Out94[23] , \Level2Out94[22] , \Level2Out94[21] , 
        \Level2Out94[20] , \Level2Out94[19] , \Level2Out94[18] , 
        \Level2Out94[17] , \Level2Out94[16] , \Level2Out94[15] , 
        \Level2Out94[14] , \Level2Out94[13] , \Level2Out94[12] , 
        \Level2Out94[11] , \Level2Out94[10] , \Level2Out94[9] , 
        \Level2Out94[8] , \Level2Out94[7] , \Level2Out94[6] , \Level2Out94[5] , 
        \Level2Out94[4] , \Level2Out94[3] , \Level2Out94[2] , \Level2Out94[1] , 
        \Level2Out94[0] }), .In1({\Level1Out94[31] , \Level1Out94[30] , 
        \Level1Out94[29] , \Level1Out94[28] , \Level1Out94[27] , 
        \Level1Out94[26] , \Level1Out94[25] , \Level1Out94[24] , 
        \Level1Out94[23] , \Level1Out94[22] , \Level1Out94[21] , 
        \Level1Out94[20] , \Level1Out94[19] , \Level1Out94[18] , 
        \Level1Out94[17] , \Level1Out94[16] , \Level1Out94[15] , 
        \Level1Out94[14] , \Level1Out94[13] , \Level1Out94[12] , 
        \Level1Out94[11] , \Level1Out94[10] , \Level1Out94[9] , 
        \Level1Out94[8] , \Level1Out94[7] , \Level1Out94[6] , \Level1Out94[5] , 
        \Level1Out94[4] , \Level1Out94[3] , \Level1Out94[2] , \Level1Out94[1] , 
        \Level1Out94[0] }), .In2({\Level1Out95[31] , \Level1Out95[30] , 
        \Level1Out95[29] , \Level1Out95[28] , \Level1Out95[27] , 
        \Level1Out95[26] , \Level1Out95[25] , \Level1Out95[24] , 
        \Level1Out95[23] , \Level1Out95[22] , \Level1Out95[21] , 
        \Level1Out95[20] , \Level1Out95[19] , \Level1Out95[18] , 
        \Level1Out95[17] , \Level1Out95[16] , \Level1Out95[15] , 
        \Level1Out95[14] , \Level1Out95[13] , \Level1Out95[12] , 
        \Level1Out95[11] , \Level1Out95[10] , \Level1Out95[9] , 
        \Level1Out95[8] , \Level1Out95[7] , \Level1Out95[6] , \Level1Out95[5] , 
        \Level1Out95[4] , \Level1Out95[3] , \Level1Out95[2] , \Level1Out95[1] , 
        \Level1Out95[0] }), .Read1(\Level1Load94[0] ), .Read2(
        \Level1Load95[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load16[0] ), .Out({\Level16Out16[31] , \Level16Out16[30] , 
        \Level16Out16[29] , \Level16Out16[28] , \Level16Out16[27] , 
        \Level16Out16[26] , \Level16Out16[25] , \Level16Out16[24] , 
        \Level16Out16[23] , \Level16Out16[22] , \Level16Out16[21] , 
        \Level16Out16[20] , \Level16Out16[19] , \Level16Out16[18] , 
        \Level16Out16[17] , \Level16Out16[16] , \Level16Out16[15] , 
        \Level16Out16[14] , \Level16Out16[13] , \Level16Out16[12] , 
        \Level16Out16[11] , \Level16Out16[10] , \Level16Out16[9] , 
        \Level16Out16[8] , \Level16Out16[7] , \Level16Out16[6] , 
        \Level16Out16[5] , \Level16Out16[4] , \Level16Out16[3] , 
        \Level16Out16[2] , \Level16Out16[1] , \Level16Out16[0] }), .In1({
        \Level8Out16[31] , \Level8Out16[30] , \Level8Out16[29] , 
        \Level8Out16[28] , \Level8Out16[27] , \Level8Out16[26] , 
        \Level8Out16[25] , \Level8Out16[24] , \Level8Out16[23] , 
        \Level8Out16[22] , \Level8Out16[21] , \Level8Out16[20] , 
        \Level8Out16[19] , \Level8Out16[18] , \Level8Out16[17] , 
        \Level8Out16[16] , \Level8Out16[15] , \Level8Out16[14] , 
        \Level8Out16[13] , \Level8Out16[12] , \Level8Out16[11] , 
        \Level8Out16[10] , \Level8Out16[9] , \Level8Out16[8] , 
        \Level8Out16[7] , \Level8Out16[6] , \Level8Out16[5] , \Level8Out16[4] , 
        \Level8Out16[3] , \Level8Out16[2] , \Level8Out16[1] , \Level8Out16[0] 
        }), .In2({\Level8Out24[31] , \Level8Out24[30] , \Level8Out24[29] , 
        \Level8Out24[28] , \Level8Out24[27] , \Level8Out24[26] , 
        \Level8Out24[25] , \Level8Out24[24] , \Level8Out24[23] , 
        \Level8Out24[22] , \Level8Out24[21] , \Level8Out24[20] , 
        \Level8Out24[19] , \Level8Out24[18] , \Level8Out24[17] , 
        \Level8Out24[16] , \Level8Out24[15] , \Level8Out24[14] , 
        \Level8Out24[13] , \Level8Out24[12] , \Level8Out24[11] , 
        \Level8Out24[10] , \Level8Out24[9] , \Level8Out24[8] , 
        \Level8Out24[7] , \Level8Out24[6] , \Level8Out24[5] , \Level8Out24[4] , 
        \Level8Out24[3] , \Level8Out24[2] , \Level8Out24[1] , \Level8Out24[0] 
        }), .Read1(\Level8Load16[0] ), .Read2(\Level8Load24[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level64Load0[0] ), .Out({\Level64Out0[31] , \Level64Out0[30] , 
        \Level64Out0[29] , \Level64Out0[28] , \Level64Out0[27] , 
        \Level64Out0[26] , \Level64Out0[25] , \Level64Out0[24] , 
        \Level64Out0[23] , \Level64Out0[22] , \Level64Out0[21] , 
        \Level64Out0[20] , \Level64Out0[19] , \Level64Out0[18] , 
        \Level64Out0[17] , \Level64Out0[16] , \Level64Out0[15] , 
        \Level64Out0[14] , \Level64Out0[13] , \Level64Out0[12] , 
        \Level64Out0[11] , \Level64Out0[10] , \Level64Out0[9] , 
        \Level64Out0[8] , \Level64Out0[7] , \Level64Out0[6] , \Level64Out0[5] , 
        \Level64Out0[4] , \Level64Out0[3] , \Level64Out0[2] , \Level64Out0[1] , 
        \Level64Out0[0] }), .In1({\Level32Out0[31] , \Level32Out0[30] , 
        \Level32Out0[29] , \Level32Out0[28] , \Level32Out0[27] , 
        \Level32Out0[26] , \Level32Out0[25] , \Level32Out0[24] , 
        \Level32Out0[23] , \Level32Out0[22] , \Level32Out0[21] , 
        \Level32Out0[20] , \Level32Out0[19] , \Level32Out0[18] , 
        \Level32Out0[17] , \Level32Out0[16] , \Level32Out0[15] , 
        \Level32Out0[14] , \Level32Out0[13] , \Level32Out0[12] , 
        \Level32Out0[11] , \Level32Out0[10] , \Level32Out0[9] , 
        \Level32Out0[8] , \Level32Out0[7] , \Level32Out0[6] , \Level32Out0[5] , 
        \Level32Out0[4] , \Level32Out0[3] , \Level32Out0[2] , \Level32Out0[1] , 
        \Level32Out0[0] }), .In2({\Level32Out32[31] , \Level32Out32[30] , 
        \Level32Out32[29] , \Level32Out32[28] , \Level32Out32[27] , 
        \Level32Out32[26] , \Level32Out32[25] , \Level32Out32[24] , 
        \Level32Out32[23] , \Level32Out32[22] , \Level32Out32[21] , 
        \Level32Out32[20] , \Level32Out32[19] , \Level32Out32[18] , 
        \Level32Out32[17] , \Level32Out32[16] , \Level32Out32[15] , 
        \Level32Out32[14] , \Level32Out32[13] , \Level32Out32[12] , 
        \Level32Out32[11] , \Level32Out32[10] , \Level32Out32[9] , 
        \Level32Out32[8] , \Level32Out32[7] , \Level32Out32[6] , 
        \Level32Out32[5] , \Level32Out32[4] , \Level32Out32[3] , 
        \Level32Out32[2] , \Level32Out32[1] , \Level32Out32[0] }), .Read1(
        \Level32Load0[0] ), .Read2(\Level32Load32[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_79 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink79[31] , \ScanLink79[30] , 
        \ScanLink79[29] , \ScanLink79[28] , \ScanLink79[27] , \ScanLink79[26] , 
        \ScanLink79[25] , \ScanLink79[24] , \ScanLink79[23] , \ScanLink79[22] , 
        \ScanLink79[21] , \ScanLink79[20] , \ScanLink79[19] , \ScanLink79[18] , 
        \ScanLink79[17] , \ScanLink79[16] , \ScanLink79[15] , \ScanLink79[14] , 
        \ScanLink79[13] , \ScanLink79[12] , \ScanLink79[11] , \ScanLink79[10] , 
        \ScanLink79[9] , \ScanLink79[8] , \ScanLink79[7] , \ScanLink79[6] , 
        \ScanLink79[5] , \ScanLink79[4] , \ScanLink79[3] , \ScanLink79[2] , 
        \ScanLink79[1] , \ScanLink79[0] }), .ScanOut({\ScanLink80[31] , 
        \ScanLink80[30] , \ScanLink80[29] , \ScanLink80[28] , \ScanLink80[27] , 
        \ScanLink80[26] , \ScanLink80[25] , \ScanLink80[24] , \ScanLink80[23] , 
        \ScanLink80[22] , \ScanLink80[21] , \ScanLink80[20] , \ScanLink80[19] , 
        \ScanLink80[18] , \ScanLink80[17] , \ScanLink80[16] , \ScanLink80[15] , 
        \ScanLink80[14] , \ScanLink80[13] , \ScanLink80[12] , \ScanLink80[11] , 
        \ScanLink80[10] , \ScanLink80[9] , \ScanLink80[8] , \ScanLink80[7] , 
        \ScanLink80[6] , \ScanLink80[5] , \ScanLink80[4] , \ScanLink80[3] , 
        \ScanLink80[2] , \ScanLink80[1] , \ScanLink80[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load79[0] ), .Out({
        \Level1Out79[31] , \Level1Out79[30] , \Level1Out79[29] , 
        \Level1Out79[28] , \Level1Out79[27] , \Level1Out79[26] , 
        \Level1Out79[25] , \Level1Out79[24] , \Level1Out79[23] , 
        \Level1Out79[22] , \Level1Out79[21] , \Level1Out79[20] , 
        \Level1Out79[19] , \Level1Out79[18] , \Level1Out79[17] , 
        \Level1Out79[16] , \Level1Out79[15] , \Level1Out79[14] , 
        \Level1Out79[13] , \Level1Out79[12] , \Level1Out79[11] , 
        \Level1Out79[10] , \Level1Out79[9] , \Level1Out79[8] , 
        \Level1Out79[7] , \Level1Out79[6] , \Level1Out79[5] , \Level1Out79[4] , 
        \Level1Out79[3] , \Level1Out79[2] , \Level1Out79[1] , \Level1Out79[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_112 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink112[31] , \ScanLink112[30] , 
        \ScanLink112[29] , \ScanLink112[28] , \ScanLink112[27] , 
        \ScanLink112[26] , \ScanLink112[25] , \ScanLink112[24] , 
        \ScanLink112[23] , \ScanLink112[22] , \ScanLink112[21] , 
        \ScanLink112[20] , \ScanLink112[19] , \ScanLink112[18] , 
        \ScanLink112[17] , \ScanLink112[16] , \ScanLink112[15] , 
        \ScanLink112[14] , \ScanLink112[13] , \ScanLink112[12] , 
        \ScanLink112[11] , \ScanLink112[10] , \ScanLink112[9] , 
        \ScanLink112[8] , \ScanLink112[7] , \ScanLink112[6] , \ScanLink112[5] , 
        \ScanLink112[4] , \ScanLink112[3] , \ScanLink112[2] , \ScanLink112[1] , 
        \ScanLink112[0] }), .ScanOut({\ScanLink113[31] , \ScanLink113[30] , 
        \ScanLink113[29] , \ScanLink113[28] , \ScanLink113[27] , 
        \ScanLink113[26] , \ScanLink113[25] , \ScanLink113[24] , 
        \ScanLink113[23] , \ScanLink113[22] , \ScanLink113[21] , 
        \ScanLink113[20] , \ScanLink113[19] , \ScanLink113[18] , 
        \ScanLink113[17] , \ScanLink113[16] , \ScanLink113[15] , 
        \ScanLink113[14] , \ScanLink113[13] , \ScanLink113[12] , 
        \ScanLink113[11] , \ScanLink113[10] , \ScanLink113[9] , 
        \ScanLink113[8] , \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , 
        \ScanLink113[4] , \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , 
        \ScanLink113[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load112[0] ), .Out({\Level1Out112[31] , \Level1Out112[30] , 
        \Level1Out112[29] , \Level1Out112[28] , \Level1Out112[27] , 
        \Level1Out112[26] , \Level1Out112[25] , \Level1Out112[24] , 
        \Level1Out112[23] , \Level1Out112[22] , \Level1Out112[21] , 
        \Level1Out112[20] , \Level1Out112[19] , \Level1Out112[18] , 
        \Level1Out112[17] , \Level1Out112[16] , \Level1Out112[15] , 
        \Level1Out112[14] , \Level1Out112[13] , \Level1Out112[12] , 
        \Level1Out112[11] , \Level1Out112[10] , \Level1Out112[9] , 
        \Level1Out112[8] , \Level1Out112[7] , \Level1Out112[6] , 
        \Level1Out112[5] , \Level1Out112[4] , \Level1Out112[3] , 
        \Level1Out112[2] , \Level1Out112[1] , \Level1Out112[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_135 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink135[31] , \ScanLink135[30] , 
        \ScanLink135[29] , \ScanLink135[28] , \ScanLink135[27] , 
        \ScanLink135[26] , \ScanLink135[25] , \ScanLink135[24] , 
        \ScanLink135[23] , \ScanLink135[22] , \ScanLink135[21] , 
        \ScanLink135[20] , \ScanLink135[19] , \ScanLink135[18] , 
        \ScanLink135[17] , \ScanLink135[16] , \ScanLink135[15] , 
        \ScanLink135[14] , \ScanLink135[13] , \ScanLink135[12] , 
        \ScanLink135[11] , \ScanLink135[10] , \ScanLink135[9] , 
        \ScanLink135[8] , \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , 
        \ScanLink135[4] , \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , 
        \ScanLink135[0] }), .ScanOut({\ScanLink136[31] , \ScanLink136[30] , 
        \ScanLink136[29] , \ScanLink136[28] , \ScanLink136[27] , 
        \ScanLink136[26] , \ScanLink136[25] , \ScanLink136[24] , 
        \ScanLink136[23] , \ScanLink136[22] , \ScanLink136[21] , 
        \ScanLink136[20] , \ScanLink136[19] , \ScanLink136[18] , 
        \ScanLink136[17] , \ScanLink136[16] , \ScanLink136[15] , 
        \ScanLink136[14] , \ScanLink136[13] , \ScanLink136[12] , 
        \ScanLink136[11] , \ScanLink136[10] , \ScanLink136[9] , 
        \ScanLink136[8] , \ScanLink136[7] , \ScanLink136[6] , \ScanLink136[5] , 
        \ScanLink136[4] , \ScanLink136[3] , \ScanLink136[2] , \ScanLink136[1] , 
        \ScanLink136[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load135[0] ), .Out({\Level1Out135[31] , \Level1Out135[30] , 
        \Level1Out135[29] , \Level1Out135[28] , \Level1Out135[27] , 
        \Level1Out135[26] , \Level1Out135[25] , \Level1Out135[24] , 
        \Level1Out135[23] , \Level1Out135[22] , \Level1Out135[21] , 
        \Level1Out135[20] , \Level1Out135[19] , \Level1Out135[18] , 
        \Level1Out135[17] , \Level1Out135[16] , \Level1Out135[15] , 
        \Level1Out135[14] , \Level1Out135[13] , \Level1Out135[12] , 
        \Level1Out135[11] , \Level1Out135[10] , \Level1Out135[9] , 
        \Level1Out135[8] , \Level1Out135[7] , \Level1Out135[6] , 
        \Level1Out135[5] , \Level1Out135[4] , \Level1Out135[3] , 
        \Level1Out135[2] , \Level1Out135[1] , \Level1Out135[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_205 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink205[31] , \ScanLink205[30] , 
        \ScanLink205[29] , \ScanLink205[28] , \ScanLink205[27] , 
        \ScanLink205[26] , \ScanLink205[25] , \ScanLink205[24] , 
        \ScanLink205[23] , \ScanLink205[22] , \ScanLink205[21] , 
        \ScanLink205[20] , \ScanLink205[19] , \ScanLink205[18] , 
        \ScanLink205[17] , \ScanLink205[16] , \ScanLink205[15] , 
        \ScanLink205[14] , \ScanLink205[13] , \ScanLink205[12] , 
        \ScanLink205[11] , \ScanLink205[10] , \ScanLink205[9] , 
        \ScanLink205[8] , \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , 
        \ScanLink205[4] , \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , 
        \ScanLink205[0] }), .ScanOut({\ScanLink206[31] , \ScanLink206[30] , 
        \ScanLink206[29] , \ScanLink206[28] , \ScanLink206[27] , 
        \ScanLink206[26] , \ScanLink206[25] , \ScanLink206[24] , 
        \ScanLink206[23] , \ScanLink206[22] , \ScanLink206[21] , 
        \ScanLink206[20] , \ScanLink206[19] , \ScanLink206[18] , 
        \ScanLink206[17] , \ScanLink206[16] , \ScanLink206[15] , 
        \ScanLink206[14] , \ScanLink206[13] , \ScanLink206[12] , 
        \ScanLink206[11] , \ScanLink206[10] , \ScanLink206[9] , 
        \ScanLink206[8] , \ScanLink206[7] , \ScanLink206[6] , \ScanLink206[5] , 
        \ScanLink206[4] , \ScanLink206[3] , \ScanLink206[2] , \ScanLink206[1] , 
        \ScanLink206[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load205[0] ), .Out({\Level1Out205[31] , \Level1Out205[30] , 
        \Level1Out205[29] , \Level1Out205[28] , \Level1Out205[27] , 
        \Level1Out205[26] , \Level1Out205[25] , \Level1Out205[24] , 
        \Level1Out205[23] , \Level1Out205[22] , \Level1Out205[21] , 
        \Level1Out205[20] , \Level1Out205[19] , \Level1Out205[18] , 
        \Level1Out205[17] , \Level1Out205[16] , \Level1Out205[15] , 
        \Level1Out205[14] , \Level1Out205[13] , \Level1Out205[12] , 
        \Level1Out205[11] , \Level1Out205[10] , \Level1Out205[9] , 
        \Level1Out205[8] , \Level1Out205[7] , \Level1Out205[6] , 
        \Level1Out205[5] , \Level1Out205[4] , \Level1Out205[3] , 
        \Level1Out205[2] , \Level1Out205[1] , \Level1Out205[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_30_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load30[0] ), .Out({\Level2Out30[31] , \Level2Out30[30] , 
        \Level2Out30[29] , \Level2Out30[28] , \Level2Out30[27] , 
        \Level2Out30[26] , \Level2Out30[25] , \Level2Out30[24] , 
        \Level2Out30[23] , \Level2Out30[22] , \Level2Out30[21] , 
        \Level2Out30[20] , \Level2Out30[19] , \Level2Out30[18] , 
        \Level2Out30[17] , \Level2Out30[16] , \Level2Out30[15] , 
        \Level2Out30[14] , \Level2Out30[13] , \Level2Out30[12] , 
        \Level2Out30[11] , \Level2Out30[10] , \Level2Out30[9] , 
        \Level2Out30[8] , \Level2Out30[7] , \Level2Out30[6] , \Level2Out30[5] , 
        \Level2Out30[4] , \Level2Out30[3] , \Level2Out30[2] , \Level2Out30[1] , 
        \Level2Out30[0] }), .In1({\Level1Out30[31] , \Level1Out30[30] , 
        \Level1Out30[29] , \Level1Out30[28] , \Level1Out30[27] , 
        \Level1Out30[26] , \Level1Out30[25] , \Level1Out30[24] , 
        \Level1Out30[23] , \Level1Out30[22] , \Level1Out30[21] , 
        \Level1Out30[20] , \Level1Out30[19] , \Level1Out30[18] , 
        \Level1Out30[17] , \Level1Out30[16] , \Level1Out30[15] , 
        \Level1Out30[14] , \Level1Out30[13] , \Level1Out30[12] , 
        \Level1Out30[11] , \Level1Out30[10] , \Level1Out30[9] , 
        \Level1Out30[8] , \Level1Out30[7] , \Level1Out30[6] , \Level1Out30[5] , 
        \Level1Out30[4] , \Level1Out30[3] , \Level1Out30[2] , \Level1Out30[1] , 
        \Level1Out30[0] }), .In2({\Level1Out31[31] , \Level1Out31[30] , 
        \Level1Out31[29] , \Level1Out31[28] , \Level1Out31[27] , 
        \Level1Out31[26] , \Level1Out31[25] , \Level1Out31[24] , 
        \Level1Out31[23] , \Level1Out31[22] , \Level1Out31[21] , 
        \Level1Out31[20] , \Level1Out31[19] , \Level1Out31[18] , 
        \Level1Out31[17] , \Level1Out31[16] , \Level1Out31[15] , 
        \Level1Out31[14] , \Level1Out31[13] , \Level1Out31[12] , 
        \Level1Out31[11] , \Level1Out31[10] , \Level1Out31[9] , 
        \Level1Out31[8] , \Level1Out31[7] , \Level1Out31[6] , \Level1Out31[5] , 
        \Level1Out31[4] , \Level1Out31[3] , \Level1Out31[2] , \Level1Out31[1] , 
        \Level1Out31[0] }), .Read1(\Level1Load30[0] ), .Read2(
        \Level1Load31[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_176_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load176[0] ), .Out({\Level2Out176[31] , \Level2Out176[30] , 
        \Level2Out176[29] , \Level2Out176[28] , \Level2Out176[27] , 
        \Level2Out176[26] , \Level2Out176[25] , \Level2Out176[24] , 
        \Level2Out176[23] , \Level2Out176[22] , \Level2Out176[21] , 
        \Level2Out176[20] , \Level2Out176[19] , \Level2Out176[18] , 
        \Level2Out176[17] , \Level2Out176[16] , \Level2Out176[15] , 
        \Level2Out176[14] , \Level2Out176[13] , \Level2Out176[12] , 
        \Level2Out176[11] , \Level2Out176[10] , \Level2Out176[9] , 
        \Level2Out176[8] , \Level2Out176[7] , \Level2Out176[6] , 
        \Level2Out176[5] , \Level2Out176[4] , \Level2Out176[3] , 
        \Level2Out176[2] , \Level2Out176[1] , \Level2Out176[0] }), .In1({
        \Level1Out176[31] , \Level1Out176[30] , \Level1Out176[29] , 
        \Level1Out176[28] , \Level1Out176[27] , \Level1Out176[26] , 
        \Level1Out176[25] , \Level1Out176[24] , \Level1Out176[23] , 
        \Level1Out176[22] , \Level1Out176[21] , \Level1Out176[20] , 
        \Level1Out176[19] , \Level1Out176[18] , \Level1Out176[17] , 
        \Level1Out176[16] , \Level1Out176[15] , \Level1Out176[14] , 
        \Level1Out176[13] , \Level1Out176[12] , \Level1Out176[11] , 
        \Level1Out176[10] , \Level1Out176[9] , \Level1Out176[8] , 
        \Level1Out176[7] , \Level1Out176[6] , \Level1Out176[5] , 
        \Level1Out176[4] , \Level1Out176[3] , \Level1Out176[2] , 
        \Level1Out176[1] , \Level1Out176[0] }), .In2({\Level1Out177[31] , 
        \Level1Out177[30] , \Level1Out177[29] , \Level1Out177[28] , 
        \Level1Out177[27] , \Level1Out177[26] , \Level1Out177[25] , 
        \Level1Out177[24] , \Level1Out177[23] , \Level1Out177[22] , 
        \Level1Out177[21] , \Level1Out177[20] , \Level1Out177[19] , 
        \Level1Out177[18] , \Level1Out177[17] , \Level1Out177[16] , 
        \Level1Out177[15] , \Level1Out177[14] , \Level1Out177[13] , 
        \Level1Out177[12] , \Level1Out177[11] , \Level1Out177[10] , 
        \Level1Out177[9] , \Level1Out177[8] , \Level1Out177[7] , 
        \Level1Out177[6] , \Level1Out177[5] , \Level1Out177[4] , 
        \Level1Out177[3] , \Level1Out177[2] , \Level1Out177[1] , 
        \Level1Out177[0] }), .Read1(\Level1Load176[0] ), .Read2(
        \Level1Load177[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_242_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load242[0] ), .Out({\Level2Out242[31] , \Level2Out242[30] , 
        \Level2Out242[29] , \Level2Out242[28] , \Level2Out242[27] , 
        \Level2Out242[26] , \Level2Out242[25] , \Level2Out242[24] , 
        \Level2Out242[23] , \Level2Out242[22] , \Level2Out242[21] , 
        \Level2Out242[20] , \Level2Out242[19] , \Level2Out242[18] , 
        \Level2Out242[17] , \Level2Out242[16] , \Level2Out242[15] , 
        \Level2Out242[14] , \Level2Out242[13] , \Level2Out242[12] , 
        \Level2Out242[11] , \Level2Out242[10] , \Level2Out242[9] , 
        \Level2Out242[8] , \Level2Out242[7] , \Level2Out242[6] , 
        \Level2Out242[5] , \Level2Out242[4] , \Level2Out242[3] , 
        \Level2Out242[2] , \Level2Out242[1] , \Level2Out242[0] }), .In1({
        \Level1Out242[31] , \Level1Out242[30] , \Level1Out242[29] , 
        \Level1Out242[28] , \Level1Out242[27] , \Level1Out242[26] , 
        \Level1Out242[25] , \Level1Out242[24] , \Level1Out242[23] , 
        \Level1Out242[22] , \Level1Out242[21] , \Level1Out242[20] , 
        \Level1Out242[19] , \Level1Out242[18] , \Level1Out242[17] , 
        \Level1Out242[16] , \Level1Out242[15] , \Level1Out242[14] , 
        \Level1Out242[13] , \Level1Out242[12] , \Level1Out242[11] , 
        \Level1Out242[10] , \Level1Out242[9] , \Level1Out242[8] , 
        \Level1Out242[7] , \Level1Out242[6] , \Level1Out242[5] , 
        \Level1Out242[4] , \Level1Out242[3] , \Level1Out242[2] , 
        \Level1Out242[1] , \Level1Out242[0] }), .In2({\Level1Out243[31] , 
        \Level1Out243[30] , \Level1Out243[29] , \Level1Out243[28] , 
        \Level1Out243[27] , \Level1Out243[26] , \Level1Out243[25] , 
        \Level1Out243[24] , \Level1Out243[23] , \Level1Out243[22] , 
        \Level1Out243[21] , \Level1Out243[20] , \Level1Out243[19] , 
        \Level1Out243[18] , \Level1Out243[17] , \Level1Out243[16] , 
        \Level1Out243[15] , \Level1Out243[14] , \Level1Out243[13] , 
        \Level1Out243[12] , \Level1Out243[11] , \Level1Out243[10] , 
        \Level1Out243[9] , \Level1Out243[8] , \Level1Out243[7] , 
        \Level1Out243[6] , \Level1Out243[5] , \Level1Out243[4] , 
        \Level1Out243[3] , \Level1Out243[2] , \Level1Out243[1] , 
        \Level1Out243[0] }), .Read1(\Level1Load242[0] ), .Read2(
        \Level1Load243[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_140_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load140[0] ), .Out({\Level4Out140[31] , \Level4Out140[30] , 
        \Level4Out140[29] , \Level4Out140[28] , \Level4Out140[27] , 
        \Level4Out140[26] , \Level4Out140[25] , \Level4Out140[24] , 
        \Level4Out140[23] , \Level4Out140[22] , \Level4Out140[21] , 
        \Level4Out140[20] , \Level4Out140[19] , \Level4Out140[18] , 
        \Level4Out140[17] , \Level4Out140[16] , \Level4Out140[15] , 
        \Level4Out140[14] , \Level4Out140[13] , \Level4Out140[12] , 
        \Level4Out140[11] , \Level4Out140[10] , \Level4Out140[9] , 
        \Level4Out140[8] , \Level4Out140[7] , \Level4Out140[6] , 
        \Level4Out140[5] , \Level4Out140[4] , \Level4Out140[3] , 
        \Level4Out140[2] , \Level4Out140[1] , \Level4Out140[0] }), .In1({
        \Level2Out140[31] , \Level2Out140[30] , \Level2Out140[29] , 
        \Level2Out140[28] , \Level2Out140[27] , \Level2Out140[26] , 
        \Level2Out140[25] , \Level2Out140[24] , \Level2Out140[23] , 
        \Level2Out140[22] , \Level2Out140[21] , \Level2Out140[20] , 
        \Level2Out140[19] , \Level2Out140[18] , \Level2Out140[17] , 
        \Level2Out140[16] , \Level2Out140[15] , \Level2Out140[14] , 
        \Level2Out140[13] , \Level2Out140[12] , \Level2Out140[11] , 
        \Level2Out140[10] , \Level2Out140[9] , \Level2Out140[8] , 
        \Level2Out140[7] , \Level2Out140[6] , \Level2Out140[5] , 
        \Level2Out140[4] , \Level2Out140[3] , \Level2Out140[2] , 
        \Level2Out140[1] , \Level2Out140[0] }), .In2({\Level2Out142[31] , 
        \Level2Out142[30] , \Level2Out142[29] , \Level2Out142[28] , 
        \Level2Out142[27] , \Level2Out142[26] , \Level2Out142[25] , 
        \Level2Out142[24] , \Level2Out142[23] , \Level2Out142[22] , 
        \Level2Out142[21] , \Level2Out142[20] , \Level2Out142[19] , 
        \Level2Out142[18] , \Level2Out142[17] , \Level2Out142[16] , 
        \Level2Out142[15] , \Level2Out142[14] , \Level2Out142[13] , 
        \Level2Out142[12] , \Level2Out142[11] , \Level2Out142[10] , 
        \Level2Out142[9] , \Level2Out142[8] , \Level2Out142[7] , 
        \Level2Out142[6] , \Level2Out142[5] , \Level2Out142[4] , 
        \Level2Out142[3] , \Level2Out142[2] , \Level2Out142[1] , 
        \Level2Out142[0] }), .Read1(\Level2Load140[0] ), .Read2(
        \Level2Load142[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_168_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load168[0] ), .Out({\Level8Out168[31] , \Level8Out168[30] , 
        \Level8Out168[29] , \Level8Out168[28] , \Level8Out168[27] , 
        \Level8Out168[26] , \Level8Out168[25] , \Level8Out168[24] , 
        \Level8Out168[23] , \Level8Out168[22] , \Level8Out168[21] , 
        \Level8Out168[20] , \Level8Out168[19] , \Level8Out168[18] , 
        \Level8Out168[17] , \Level8Out168[16] , \Level8Out168[15] , 
        \Level8Out168[14] , \Level8Out168[13] , \Level8Out168[12] , 
        \Level8Out168[11] , \Level8Out168[10] , \Level8Out168[9] , 
        \Level8Out168[8] , \Level8Out168[7] , \Level8Out168[6] , 
        \Level8Out168[5] , \Level8Out168[4] , \Level8Out168[3] , 
        \Level8Out168[2] , \Level8Out168[1] , \Level8Out168[0] }), .In1({
        \Level4Out168[31] , \Level4Out168[30] , \Level4Out168[29] , 
        \Level4Out168[28] , \Level4Out168[27] , \Level4Out168[26] , 
        \Level4Out168[25] , \Level4Out168[24] , \Level4Out168[23] , 
        \Level4Out168[22] , \Level4Out168[21] , \Level4Out168[20] , 
        \Level4Out168[19] , \Level4Out168[18] , \Level4Out168[17] , 
        \Level4Out168[16] , \Level4Out168[15] , \Level4Out168[14] , 
        \Level4Out168[13] , \Level4Out168[12] , \Level4Out168[11] , 
        \Level4Out168[10] , \Level4Out168[9] , \Level4Out168[8] , 
        \Level4Out168[7] , \Level4Out168[6] , \Level4Out168[5] , 
        \Level4Out168[4] , \Level4Out168[3] , \Level4Out168[2] , 
        \Level4Out168[1] , \Level4Out168[0] }), .In2({\Level4Out172[31] , 
        \Level4Out172[30] , \Level4Out172[29] , \Level4Out172[28] , 
        \Level4Out172[27] , \Level4Out172[26] , \Level4Out172[25] , 
        \Level4Out172[24] , \Level4Out172[23] , \Level4Out172[22] , 
        \Level4Out172[21] , \Level4Out172[20] , \Level4Out172[19] , 
        \Level4Out172[18] , \Level4Out172[17] , \Level4Out172[16] , 
        \Level4Out172[15] , \Level4Out172[14] , \Level4Out172[13] , 
        \Level4Out172[12] , \Level4Out172[11] , \Level4Out172[10] , 
        \Level4Out172[9] , \Level4Out172[8] , \Level4Out172[7] , 
        \Level4Out172[6] , \Level4Out172[5] , \Level4Out172[4] , 
        \Level4Out172[3] , \Level4Out172[2] , \Level4Out172[1] , 
        \Level4Out172[0] }), .Read1(\Level4Load168[0] ), .Read2(
        \Level4Load172[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_222 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink222[31] , \ScanLink222[30] , 
        \ScanLink222[29] , \ScanLink222[28] , \ScanLink222[27] , 
        \ScanLink222[26] , \ScanLink222[25] , \ScanLink222[24] , 
        \ScanLink222[23] , \ScanLink222[22] , \ScanLink222[21] , 
        \ScanLink222[20] , \ScanLink222[19] , \ScanLink222[18] , 
        \ScanLink222[17] , \ScanLink222[16] , \ScanLink222[15] , 
        \ScanLink222[14] , \ScanLink222[13] , \ScanLink222[12] , 
        \ScanLink222[11] , \ScanLink222[10] , \ScanLink222[9] , 
        \ScanLink222[8] , \ScanLink222[7] , \ScanLink222[6] , \ScanLink222[5] , 
        \ScanLink222[4] , \ScanLink222[3] , \ScanLink222[2] , \ScanLink222[1] , 
        \ScanLink222[0] }), .ScanOut({\ScanLink223[31] , \ScanLink223[30] , 
        \ScanLink223[29] , \ScanLink223[28] , \ScanLink223[27] , 
        \ScanLink223[26] , \ScanLink223[25] , \ScanLink223[24] , 
        \ScanLink223[23] , \ScanLink223[22] , \ScanLink223[21] , 
        \ScanLink223[20] , \ScanLink223[19] , \ScanLink223[18] , 
        \ScanLink223[17] , \ScanLink223[16] , \ScanLink223[15] , 
        \ScanLink223[14] , \ScanLink223[13] , \ScanLink223[12] , 
        \ScanLink223[11] , \ScanLink223[10] , \ScanLink223[9] , 
        \ScanLink223[8] , \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , 
        \ScanLink223[4] , \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , 
        \ScanLink223[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load222[0] ), .Out({\Level1Out222[31] , \Level1Out222[30] , 
        \Level1Out222[29] , \Level1Out222[28] , \Level1Out222[27] , 
        \Level1Out222[26] , \Level1Out222[25] , \Level1Out222[24] , 
        \Level1Out222[23] , \Level1Out222[22] , \Level1Out222[21] , 
        \Level1Out222[20] , \Level1Out222[19] , \Level1Out222[18] , 
        \Level1Out222[17] , \Level1Out222[16] , \Level1Out222[15] , 
        \Level1Out222[14] , \Level1Out222[13] , \Level1Out222[12] , 
        \Level1Out222[11] , \Level1Out222[10] , \Level1Out222[9] , 
        \Level1Out222[8] , \Level1Out222[7] , \Level1Out222[6] , 
        \Level1Out222[5] , \Level1Out222[4] , \Level1Out222[3] , 
        \Level1Out222[2] , \Level1Out222[1] , \Level1Out222[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_199 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink199[31] , \ScanLink199[30] , 
        \ScanLink199[29] , \ScanLink199[28] , \ScanLink199[27] , 
        \ScanLink199[26] , \ScanLink199[25] , \ScanLink199[24] , 
        \ScanLink199[23] , \ScanLink199[22] , \ScanLink199[21] , 
        \ScanLink199[20] , \ScanLink199[19] , \ScanLink199[18] , 
        \ScanLink199[17] , \ScanLink199[16] , \ScanLink199[15] , 
        \ScanLink199[14] , \ScanLink199[13] , \ScanLink199[12] , 
        \ScanLink199[11] , \ScanLink199[10] , \ScanLink199[9] , 
        \ScanLink199[8] , \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , 
        \ScanLink199[4] , \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , 
        \ScanLink199[0] }), .ScanOut({\ScanLink200[31] , \ScanLink200[30] , 
        \ScanLink200[29] , \ScanLink200[28] , \ScanLink200[27] , 
        \ScanLink200[26] , \ScanLink200[25] , \ScanLink200[24] , 
        \ScanLink200[23] , \ScanLink200[22] , \ScanLink200[21] , 
        \ScanLink200[20] , \ScanLink200[19] , \ScanLink200[18] , 
        \ScanLink200[17] , \ScanLink200[16] , \ScanLink200[15] , 
        \ScanLink200[14] , \ScanLink200[13] , \ScanLink200[12] , 
        \ScanLink200[11] , \ScanLink200[10] , \ScanLink200[9] , 
        \ScanLink200[8] , \ScanLink200[7] , \ScanLink200[6] , \ScanLink200[5] , 
        \ScanLink200[4] , \ScanLink200[3] , \ScanLink200[2] , \ScanLink200[1] , 
        \ScanLink200[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load199[0] ), .Out({\Level1Out199[31] , \Level1Out199[30] , 
        \Level1Out199[29] , \Level1Out199[28] , \Level1Out199[27] , 
        \Level1Out199[26] , \Level1Out199[25] , \Level1Out199[24] , 
        \Level1Out199[23] , \Level1Out199[22] , \Level1Out199[21] , 
        \Level1Out199[20] , \Level1Out199[19] , \Level1Out199[18] , 
        \Level1Out199[17] , \Level1Out199[16] , \Level1Out199[15] , 
        \Level1Out199[14] , \Level1Out199[13] , \Level1Out199[12] , 
        \Level1Out199[11] , \Level1Out199[10] , \Level1Out199[9] , 
        \Level1Out199[8] , \Level1Out199[7] , \Level1Out199[6] , 
        \Level1Out199[5] , \Level1Out199[4] , \Level1Out199[3] , 
        \Level1Out199[2] , \Level1Out199[1] , \Level1Out199[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_115 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink115[31] , \ScanLink115[30] , 
        \ScanLink115[29] , \ScanLink115[28] , \ScanLink115[27] , 
        \ScanLink115[26] , \ScanLink115[25] , \ScanLink115[24] , 
        \ScanLink115[23] , \ScanLink115[22] , \ScanLink115[21] , 
        \ScanLink115[20] , \ScanLink115[19] , \ScanLink115[18] , 
        \ScanLink115[17] , \ScanLink115[16] , \ScanLink115[15] , 
        \ScanLink115[14] , \ScanLink115[13] , \ScanLink115[12] , 
        \ScanLink115[11] , \ScanLink115[10] , \ScanLink115[9] , 
        \ScanLink115[8] , \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , 
        \ScanLink115[4] , \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , 
        \ScanLink115[0] }), .ScanOut({\ScanLink116[31] , \ScanLink116[30] , 
        \ScanLink116[29] , \ScanLink116[28] , \ScanLink116[27] , 
        \ScanLink116[26] , \ScanLink116[25] , \ScanLink116[24] , 
        \ScanLink116[23] , \ScanLink116[22] , \ScanLink116[21] , 
        \ScanLink116[20] , \ScanLink116[19] , \ScanLink116[18] , 
        \ScanLink116[17] , \ScanLink116[16] , \ScanLink116[15] , 
        \ScanLink116[14] , \ScanLink116[13] , \ScanLink116[12] , 
        \ScanLink116[11] , \ScanLink116[10] , \ScanLink116[9] , 
        \ScanLink116[8] , \ScanLink116[7] , \ScanLink116[6] , \ScanLink116[5] , 
        \ScanLink116[4] , \ScanLink116[3] , \ScanLink116[2] , \ScanLink116[1] , 
        \ScanLink116[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load115[0] ), .Out({\Level1Out115[31] , \Level1Out115[30] , 
        \Level1Out115[29] , \Level1Out115[28] , \Level1Out115[27] , 
        \Level1Out115[26] , \Level1Out115[25] , \Level1Out115[24] , 
        \Level1Out115[23] , \Level1Out115[22] , \Level1Out115[21] , 
        \Level1Out115[20] , \Level1Out115[19] , \Level1Out115[18] , 
        \Level1Out115[17] , \Level1Out115[16] , \Level1Out115[15] , 
        \Level1Out115[14] , \Level1Out115[13] , \Level1Out115[12] , 
        \Level1Out115[11] , \Level1Out115[10] , \Level1Out115[9] , 
        \Level1Out115[8] , \Level1Out115[7] , \Level1Out115[6] , 
        \Level1Out115[5] , \Level1Out115[4] , \Level1Out115[3] , 
        \Level1Out115[2] , \Level1Out115[1] , \Level1Out115[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_225 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink225[31] , \ScanLink225[30] , 
        \ScanLink225[29] , \ScanLink225[28] , \ScanLink225[27] , 
        \ScanLink225[26] , \ScanLink225[25] , \ScanLink225[24] , 
        \ScanLink225[23] , \ScanLink225[22] , \ScanLink225[21] , 
        \ScanLink225[20] , \ScanLink225[19] , \ScanLink225[18] , 
        \ScanLink225[17] , \ScanLink225[16] , \ScanLink225[15] , 
        \ScanLink225[14] , \ScanLink225[13] , \ScanLink225[12] , 
        \ScanLink225[11] , \ScanLink225[10] , \ScanLink225[9] , 
        \ScanLink225[8] , \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , 
        \ScanLink225[4] , \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , 
        \ScanLink225[0] }), .ScanOut({\ScanLink226[31] , \ScanLink226[30] , 
        \ScanLink226[29] , \ScanLink226[28] , \ScanLink226[27] , 
        \ScanLink226[26] , \ScanLink226[25] , \ScanLink226[24] , 
        \ScanLink226[23] , \ScanLink226[22] , \ScanLink226[21] , 
        \ScanLink226[20] , \ScanLink226[19] , \ScanLink226[18] , 
        \ScanLink226[17] , \ScanLink226[16] , \ScanLink226[15] , 
        \ScanLink226[14] , \ScanLink226[13] , \ScanLink226[12] , 
        \ScanLink226[11] , \ScanLink226[10] , \ScanLink226[9] , 
        \ScanLink226[8] , \ScanLink226[7] , \ScanLink226[6] , \ScanLink226[5] , 
        \ScanLink226[4] , \ScanLink226[3] , \ScanLink226[2] , \ScanLink226[1] , 
        \ScanLink226[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load225[0] ), .Out({\Level1Out225[31] , \Level1Out225[30] , 
        \Level1Out225[29] , \Level1Out225[28] , \Level1Out225[27] , 
        \Level1Out225[26] , \Level1Out225[25] , \Level1Out225[24] , 
        \Level1Out225[23] , \Level1Out225[22] , \Level1Out225[21] , 
        \Level1Out225[20] , \Level1Out225[19] , \Level1Out225[18] , 
        \Level1Out225[17] , \Level1Out225[16] , \Level1Out225[15] , 
        \Level1Out225[14] , \Level1Out225[13] , \Level1Out225[12] , 
        \Level1Out225[11] , \Level1Out225[10] , \Level1Out225[9] , 
        \Level1Out225[8] , \Level1Out225[7] , \Level1Out225[6] , 
        \Level1Out225[5] , \Level1Out225[4] , \Level1Out225[3] , 
        \Level1Out225[2] , \Level1Out225[1] , \Level1Out225[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load24[0] ), .Out({\Level2Out24[31] , \Level2Out24[30] , 
        \Level2Out24[29] , \Level2Out24[28] , \Level2Out24[27] , 
        \Level2Out24[26] , \Level2Out24[25] , \Level2Out24[24] , 
        \Level2Out24[23] , \Level2Out24[22] , \Level2Out24[21] , 
        \Level2Out24[20] , \Level2Out24[19] , \Level2Out24[18] , 
        \Level2Out24[17] , \Level2Out24[16] , \Level2Out24[15] , 
        \Level2Out24[14] , \Level2Out24[13] , \Level2Out24[12] , 
        \Level2Out24[11] , \Level2Out24[10] , \Level2Out24[9] , 
        \Level2Out24[8] , \Level2Out24[7] , \Level2Out24[6] , \Level2Out24[5] , 
        \Level2Out24[4] , \Level2Out24[3] , \Level2Out24[2] , \Level2Out24[1] , 
        \Level2Out24[0] }), .In1({\Level1Out24[31] , \Level1Out24[30] , 
        \Level1Out24[29] , \Level1Out24[28] , \Level1Out24[27] , 
        \Level1Out24[26] , \Level1Out24[25] , \Level1Out24[24] , 
        \Level1Out24[23] , \Level1Out24[22] , \Level1Out24[21] , 
        \Level1Out24[20] , \Level1Out24[19] , \Level1Out24[18] , 
        \Level1Out24[17] , \Level1Out24[16] , \Level1Out24[15] , 
        \Level1Out24[14] , \Level1Out24[13] , \Level1Out24[12] , 
        \Level1Out24[11] , \Level1Out24[10] , \Level1Out24[9] , 
        \Level1Out24[8] , \Level1Out24[7] , \Level1Out24[6] , \Level1Out24[5] , 
        \Level1Out24[4] , \Level1Out24[3] , \Level1Out24[2] , \Level1Out24[1] , 
        \Level1Out24[0] }), .In2({\Level1Out25[31] , \Level1Out25[30] , 
        \Level1Out25[29] , \Level1Out25[28] , \Level1Out25[27] , 
        \Level1Out25[26] , \Level1Out25[25] , \Level1Out25[24] , 
        \Level1Out25[23] , \Level1Out25[22] , \Level1Out25[21] , 
        \Level1Out25[20] , \Level1Out25[19] , \Level1Out25[18] , 
        \Level1Out25[17] , \Level1Out25[16] , \Level1Out25[15] , 
        \Level1Out25[14] , \Level1Out25[13] , \Level1Out25[12] , 
        \Level1Out25[11] , \Level1Out25[10] , \Level1Out25[9] , 
        \Level1Out25[8] , \Level1Out25[7] , \Level1Out25[6] , \Level1Out25[5] , 
        \Level1Out25[4] , \Level1Out25[3] , \Level1Out25[2] , \Level1Out25[1] , 
        \Level1Out25[0] }), .Read1(\Level1Load24[0] ), .Read2(
        \Level1Load25[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_148_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load148[0] ), .Out({\Level2Out148[31] , \Level2Out148[30] , 
        \Level2Out148[29] , \Level2Out148[28] , \Level2Out148[27] , 
        \Level2Out148[26] , \Level2Out148[25] , \Level2Out148[24] , 
        \Level2Out148[23] , \Level2Out148[22] , \Level2Out148[21] , 
        \Level2Out148[20] , \Level2Out148[19] , \Level2Out148[18] , 
        \Level2Out148[17] , \Level2Out148[16] , \Level2Out148[15] , 
        \Level2Out148[14] , \Level2Out148[13] , \Level2Out148[12] , 
        \Level2Out148[11] , \Level2Out148[10] , \Level2Out148[9] , 
        \Level2Out148[8] , \Level2Out148[7] , \Level2Out148[6] , 
        \Level2Out148[5] , \Level2Out148[4] , \Level2Out148[3] , 
        \Level2Out148[2] , \Level2Out148[1] , \Level2Out148[0] }), .In1({
        \Level1Out148[31] , \Level1Out148[30] , \Level1Out148[29] , 
        \Level1Out148[28] , \Level1Out148[27] , \Level1Out148[26] , 
        \Level1Out148[25] , \Level1Out148[24] , \Level1Out148[23] , 
        \Level1Out148[22] , \Level1Out148[21] , \Level1Out148[20] , 
        \Level1Out148[19] , \Level1Out148[18] , \Level1Out148[17] , 
        \Level1Out148[16] , \Level1Out148[15] , \Level1Out148[14] , 
        \Level1Out148[13] , \Level1Out148[12] , \Level1Out148[11] , 
        \Level1Out148[10] , \Level1Out148[9] , \Level1Out148[8] , 
        \Level1Out148[7] , \Level1Out148[6] , \Level1Out148[5] , 
        \Level1Out148[4] , \Level1Out148[3] , \Level1Out148[2] , 
        \Level1Out148[1] , \Level1Out148[0] }), .In2({\Level1Out149[31] , 
        \Level1Out149[30] , \Level1Out149[29] , \Level1Out149[28] , 
        \Level1Out149[27] , \Level1Out149[26] , \Level1Out149[25] , 
        \Level1Out149[24] , \Level1Out149[23] , \Level1Out149[22] , 
        \Level1Out149[21] , \Level1Out149[20] , \Level1Out149[19] , 
        \Level1Out149[18] , \Level1Out149[17] , \Level1Out149[16] , 
        \Level1Out149[15] , \Level1Out149[14] , \Level1Out149[13] , 
        \Level1Out149[12] , \Level1Out149[11] , \Level1Out149[10] , 
        \Level1Out149[9] , \Level1Out149[8] , \Level1Out149[7] , 
        \Level1Out149[6] , \Level1Out149[5] , \Level1Out149[4] , 
        \Level1Out149[3] , \Level1Out149[2] , \Level1Out149[1] , 
        \Level1Out149[0] }), .Read1(\Level1Load148[0] ), .Read2(
        \Level1Load149[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_132 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink132[31] , \ScanLink132[30] , 
        \ScanLink132[29] , \ScanLink132[28] , \ScanLink132[27] , 
        \ScanLink132[26] , \ScanLink132[25] , \ScanLink132[24] , 
        \ScanLink132[23] , \ScanLink132[22] , \ScanLink132[21] , 
        \ScanLink132[20] , \ScanLink132[19] , \ScanLink132[18] , 
        \ScanLink132[17] , \ScanLink132[16] , \ScanLink132[15] , 
        \ScanLink132[14] , \ScanLink132[13] , \ScanLink132[12] , 
        \ScanLink132[11] , \ScanLink132[10] , \ScanLink132[9] , 
        \ScanLink132[8] , \ScanLink132[7] , \ScanLink132[6] , \ScanLink132[5] , 
        \ScanLink132[4] , \ScanLink132[3] , \ScanLink132[2] , \ScanLink132[1] , 
        \ScanLink132[0] }), .ScanOut({\ScanLink133[31] , \ScanLink133[30] , 
        \ScanLink133[29] , \ScanLink133[28] , \ScanLink133[27] , 
        \ScanLink133[26] , \ScanLink133[25] , \ScanLink133[24] , 
        \ScanLink133[23] , \ScanLink133[22] , \ScanLink133[21] , 
        \ScanLink133[20] , \ScanLink133[19] , \ScanLink133[18] , 
        \ScanLink133[17] , \ScanLink133[16] , \ScanLink133[15] , 
        \ScanLink133[14] , \ScanLink133[13] , \ScanLink133[12] , 
        \ScanLink133[11] , \ScanLink133[10] , \ScanLink133[9] , 
        \ScanLink133[8] , \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , 
        \ScanLink133[4] , \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , 
        \ScanLink133[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load132[0] ), .Out({\Level1Out132[31] , \Level1Out132[30] , 
        \Level1Out132[29] , \Level1Out132[28] , \Level1Out132[27] , 
        \Level1Out132[26] , \Level1Out132[25] , \Level1Out132[24] , 
        \Level1Out132[23] , \Level1Out132[22] , \Level1Out132[21] , 
        \Level1Out132[20] , \Level1Out132[19] , \Level1Out132[18] , 
        \Level1Out132[17] , \Level1Out132[16] , \Level1Out132[15] , 
        \Level1Out132[14] , \Level1Out132[13] , \Level1Out132[12] , 
        \Level1Out132[11] , \Level1Out132[10] , \Level1Out132[9] , 
        \Level1Out132[8] , \Level1Out132[7] , \Level1Out132[6] , 
        \Level1Out132[5] , \Level1Out132[4] , \Level1Out132[3] , 
        \Level1Out132[2] , \Level1Out132[1] , \Level1Out132[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_162_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load162[0] ), .Out({\Level2Out162[31] , \Level2Out162[30] , 
        \Level2Out162[29] , \Level2Out162[28] , \Level2Out162[27] , 
        \Level2Out162[26] , \Level2Out162[25] , \Level2Out162[24] , 
        \Level2Out162[23] , \Level2Out162[22] , \Level2Out162[21] , 
        \Level2Out162[20] , \Level2Out162[19] , \Level2Out162[18] , 
        \Level2Out162[17] , \Level2Out162[16] , \Level2Out162[15] , 
        \Level2Out162[14] , \Level2Out162[13] , \Level2Out162[12] , 
        \Level2Out162[11] , \Level2Out162[10] , \Level2Out162[9] , 
        \Level2Out162[8] , \Level2Out162[7] , \Level2Out162[6] , 
        \Level2Out162[5] , \Level2Out162[4] , \Level2Out162[3] , 
        \Level2Out162[2] , \Level2Out162[1] , \Level2Out162[0] }), .In1({
        \Level1Out162[31] , \Level1Out162[30] , \Level1Out162[29] , 
        \Level1Out162[28] , \Level1Out162[27] , \Level1Out162[26] , 
        \Level1Out162[25] , \Level1Out162[24] , \Level1Out162[23] , 
        \Level1Out162[22] , \Level1Out162[21] , \Level1Out162[20] , 
        \Level1Out162[19] , \Level1Out162[18] , \Level1Out162[17] , 
        \Level1Out162[16] , \Level1Out162[15] , \Level1Out162[14] , 
        \Level1Out162[13] , \Level1Out162[12] , \Level1Out162[11] , 
        \Level1Out162[10] , \Level1Out162[9] , \Level1Out162[8] , 
        \Level1Out162[7] , \Level1Out162[6] , \Level1Out162[5] , 
        \Level1Out162[4] , \Level1Out162[3] , \Level1Out162[2] , 
        \Level1Out162[1] , \Level1Out162[0] }), .In2({\Level1Out163[31] , 
        \Level1Out163[30] , \Level1Out163[29] , \Level1Out163[28] , 
        \Level1Out163[27] , \Level1Out163[26] , \Level1Out163[25] , 
        \Level1Out163[24] , \Level1Out163[23] , \Level1Out163[22] , 
        \Level1Out163[21] , \Level1Out163[20] , \Level1Out163[19] , 
        \Level1Out163[18] , \Level1Out163[17] , \Level1Out163[16] , 
        \Level1Out163[15] , \Level1Out163[14] , \Level1Out163[13] , 
        \Level1Out163[12] , \Level1Out163[11] , \Level1Out163[10] , 
        \Level1Out163[9] , \Level1Out163[8] , \Level1Out163[7] , 
        \Level1Out163[6] , \Level1Out163[5] , \Level1Out163[4] , 
        \Level1Out163[3] , \Level1Out163[2] , \Level1Out163[1] , 
        \Level1Out163[0] }), .Read1(\Level1Load162[0] ), .Read2(
        \Level1Load163[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_202 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink202[31] , \ScanLink202[30] , 
        \ScanLink202[29] , \ScanLink202[28] , \ScanLink202[27] , 
        \ScanLink202[26] , \ScanLink202[25] , \ScanLink202[24] , 
        \ScanLink202[23] , \ScanLink202[22] , \ScanLink202[21] , 
        \ScanLink202[20] , \ScanLink202[19] , \ScanLink202[18] , 
        \ScanLink202[17] , \ScanLink202[16] , \ScanLink202[15] , 
        \ScanLink202[14] , \ScanLink202[13] , \ScanLink202[12] , 
        \ScanLink202[11] , \ScanLink202[10] , \ScanLink202[9] , 
        \ScanLink202[8] , \ScanLink202[7] , \ScanLink202[6] , \ScanLink202[5] , 
        \ScanLink202[4] , \ScanLink202[3] , \ScanLink202[2] , \ScanLink202[1] , 
        \ScanLink202[0] }), .ScanOut({\ScanLink203[31] , \ScanLink203[30] , 
        \ScanLink203[29] , \ScanLink203[28] , \ScanLink203[27] , 
        \ScanLink203[26] , \ScanLink203[25] , \ScanLink203[24] , 
        \ScanLink203[23] , \ScanLink203[22] , \ScanLink203[21] , 
        \ScanLink203[20] , \ScanLink203[19] , \ScanLink203[18] , 
        \ScanLink203[17] , \ScanLink203[16] , \ScanLink203[15] , 
        \ScanLink203[14] , \ScanLink203[13] , \ScanLink203[12] , 
        \ScanLink203[11] , \ScanLink203[10] , \ScanLink203[9] , 
        \ScanLink203[8] , \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , 
        \ScanLink203[4] , \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , 
        \ScanLink203[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load202[0] ), .Out({\Level1Out202[31] , \Level1Out202[30] , 
        \Level1Out202[29] , \Level1Out202[28] , \Level1Out202[27] , 
        \Level1Out202[26] , \Level1Out202[25] , \Level1Out202[24] , 
        \Level1Out202[23] , \Level1Out202[22] , \Level1Out202[21] , 
        \Level1Out202[20] , \Level1Out202[19] , \Level1Out202[18] , 
        \Level1Out202[17] , \Level1Out202[16] , \Level1Out202[15] , 
        \Level1Out202[14] , \Level1Out202[13] , \Level1Out202[12] , 
        \Level1Out202[11] , \Level1Out202[10] , \Level1Out202[9] , 
        \Level1Out202[8] , \Level1Out202[7] , \Level1Out202[6] , 
        \Level1Out202[5] , \Level1Out202[4] , \Level1Out202[3] , 
        \Level1Out202[2] , \Level1Out202[1] , \Level1Out202[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_12_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load12[0] ), .Out({\Level4Out12[31] , \Level4Out12[30] , 
        \Level4Out12[29] , \Level4Out12[28] , \Level4Out12[27] , 
        \Level4Out12[26] , \Level4Out12[25] , \Level4Out12[24] , 
        \Level4Out12[23] , \Level4Out12[22] , \Level4Out12[21] , 
        \Level4Out12[20] , \Level4Out12[19] , \Level4Out12[18] , 
        \Level4Out12[17] , \Level4Out12[16] , \Level4Out12[15] , 
        \Level4Out12[14] , \Level4Out12[13] , \Level4Out12[12] , 
        \Level4Out12[11] , \Level4Out12[10] , \Level4Out12[9] , 
        \Level4Out12[8] , \Level4Out12[7] , \Level4Out12[6] , \Level4Out12[5] , 
        \Level4Out12[4] , \Level4Out12[3] , \Level4Out12[2] , \Level4Out12[1] , 
        \Level4Out12[0] }), .In1({\Level2Out12[31] , \Level2Out12[30] , 
        \Level2Out12[29] , \Level2Out12[28] , \Level2Out12[27] , 
        \Level2Out12[26] , \Level2Out12[25] , \Level2Out12[24] , 
        \Level2Out12[23] , \Level2Out12[22] , \Level2Out12[21] , 
        \Level2Out12[20] , \Level2Out12[19] , \Level2Out12[18] , 
        \Level2Out12[17] , \Level2Out12[16] , \Level2Out12[15] , 
        \Level2Out12[14] , \Level2Out12[13] , \Level2Out12[12] , 
        \Level2Out12[11] , \Level2Out12[10] , \Level2Out12[9] , 
        \Level2Out12[8] , \Level2Out12[7] , \Level2Out12[6] , \Level2Out12[5] , 
        \Level2Out12[4] , \Level2Out12[3] , \Level2Out12[2] , \Level2Out12[1] , 
        \Level2Out12[0] }), .In2({\Level2Out14[31] , \Level2Out14[30] , 
        \Level2Out14[29] , \Level2Out14[28] , \Level2Out14[27] , 
        \Level2Out14[26] , \Level2Out14[25] , \Level2Out14[24] , 
        \Level2Out14[23] , \Level2Out14[22] , \Level2Out14[21] , 
        \Level2Out14[20] , \Level2Out14[19] , \Level2Out14[18] , 
        \Level2Out14[17] , \Level2Out14[16] , \Level2Out14[15] , 
        \Level2Out14[14] , \Level2Out14[13] , \Level2Out14[12] , 
        \Level2Out14[11] , \Level2Out14[10] , \Level2Out14[9] , 
        \Level2Out14[8] , \Level2Out14[7] , \Level2Out14[6] , \Level2Out14[5] , 
        \Level2Out14[4] , \Level2Out14[3] , \Level2Out14[2] , \Level2Out14[1] , 
        \Level2Out14[0] }), .Read1(\Level2Load12[0] ), .Read2(
        \Level2Load14[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_19 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanOut({\ScanLink20[31] , 
        \ScanLink20[30] , \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , 
        \ScanLink20[26] , \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , 
        \ScanLink20[22] , \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , 
        \ScanLink20[18] , \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , 
        \ScanLink20[14] , \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , 
        \ScanLink20[10] , \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , 
        \ScanLink20[6] , \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , 
        \ScanLink20[2] , \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load19[0] ), .Out({
        \Level1Out19[31] , \Level1Out19[30] , \Level1Out19[29] , 
        \Level1Out19[28] , \Level1Out19[27] , \Level1Out19[26] , 
        \Level1Out19[25] , \Level1Out19[24] , \Level1Out19[23] , 
        \Level1Out19[22] , \Level1Out19[21] , \Level1Out19[20] , 
        \Level1Out19[19] , \Level1Out19[18] , \Level1Out19[17] , 
        \Level1Out19[16] , \Level1Out19[15] , \Level1Out19[14] , 
        \Level1Out19[13] , \Level1Out19[12] , \Level1Out19[11] , 
        \Level1Out19[10] , \Level1Out19[9] , \Level1Out19[8] , 
        \Level1Out19[7] , \Level1Out19[6] , \Level1Out19[5] , \Level1Out19[4] , 
        \Level1Out19[3] , \Level1Out19[2] , \Level1Out19[1] , \Level1Out19[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_37 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanOut({\ScanLink38[31] , 
        \ScanLink38[30] , \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , 
        \ScanLink38[26] , \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , 
        \ScanLink38[22] , \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , 
        \ScanLink38[18] , \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , 
        \ScanLink38[14] , \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , 
        \ScanLink38[10] , \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , 
        \ScanLink38[6] , \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , 
        \ScanLink38[2] , \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load37[0] ), .Out({
        \Level1Out37[31] , \Level1Out37[30] , \Level1Out37[29] , 
        \Level1Out37[28] , \Level1Out37[27] , \Level1Out37[26] , 
        \Level1Out37[25] , \Level1Out37[24] , \Level1Out37[23] , 
        \Level1Out37[22] , \Level1Out37[21] , \Level1Out37[20] , 
        \Level1Out37[19] , \Level1Out37[18] , \Level1Out37[17] , 
        \Level1Out37[16] , \Level1Out37[15] , \Level1Out37[14] , 
        \Level1Out37[13] , \Level1Out37[12] , \Level1Out37[11] , 
        \Level1Out37[10] , \Level1Out37[9] , \Level1Out37[8] , 
        \Level1Out37[7] , \Level1Out37[6] , \Level1Out37[5] , \Level1Out37[4] , 
        \Level1Out37[3] , \Level1Out37[2] , \Level1Out37[1] , \Level1Out37[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_42 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanOut({\ScanLink43[31] , 
        \ScanLink43[30] , \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , 
        \ScanLink43[26] , \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , 
        \ScanLink43[22] , \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , 
        \ScanLink43[18] , \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , 
        \ScanLink43[14] , \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , 
        \ScanLink43[10] , \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , 
        \ScanLink43[6] , \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , 
        \ScanLink43[2] , \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load42[0] ), .Out({
        \Level1Out42[31] , \Level1Out42[30] , \Level1Out42[29] , 
        \Level1Out42[28] , \Level1Out42[27] , \Level1Out42[26] , 
        \Level1Out42[25] , \Level1Out42[24] , \Level1Out42[23] , 
        \Level1Out42[22] , \Level1Out42[21] , \Level1Out42[20] , 
        \Level1Out42[19] , \Level1Out42[18] , \Level1Out42[17] , 
        \Level1Out42[16] , \Level1Out42[15] , \Level1Out42[14] , 
        \Level1Out42[13] , \Level1Out42[12] , \Level1Out42[11] , 
        \Level1Out42[10] , \Level1Out42[9] , \Level1Out42[8] , 
        \Level1Out42[7] , \Level1Out42[6] , \Level1Out42[5] , \Level1Out42[4] , 
        \Level1Out42[3] , \Level1Out42[2] , \Level1Out42[1] , \Level1Out42[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_59 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanOut({\ScanLink60[31] , 
        \ScanLink60[30] , \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , 
        \ScanLink60[26] , \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , 
        \ScanLink60[22] , \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , 
        \ScanLink60[18] , \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , 
        \ScanLink60[14] , \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , 
        \ScanLink60[10] , \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , 
        \ScanLink60[6] , \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , 
        \ScanLink60[2] , \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load59[0] ), .Out({
        \Level1Out59[31] , \Level1Out59[30] , \Level1Out59[29] , 
        \Level1Out59[28] , \Level1Out59[27] , \Level1Out59[26] , 
        \Level1Out59[25] , \Level1Out59[24] , \Level1Out59[23] , 
        \Level1Out59[22] , \Level1Out59[21] , \Level1Out59[20] , 
        \Level1Out59[19] , \Level1Out59[18] , \Level1Out59[17] , 
        \Level1Out59[16] , \Level1Out59[15] , \Level1Out59[14] , 
        \Level1Out59[13] , \Level1Out59[12] , \Level1Out59[11] , 
        \Level1Out59[10] , \Level1Out59[9] , \Level1Out59[8] , 
        \Level1Out59[7] , \Level1Out59[6] , \Level1Out59[5] , \Level1Out59[4] , 
        \Level1Out59[3] , \Level1Out59[2] , \Level1Out59[1] , \Level1Out59[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_98_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load98[0] ), .Out({\Level2Out98[31] , \Level2Out98[30] , 
        \Level2Out98[29] , \Level2Out98[28] , \Level2Out98[27] , 
        \Level2Out98[26] , \Level2Out98[25] , \Level2Out98[24] , 
        \Level2Out98[23] , \Level2Out98[22] , \Level2Out98[21] , 
        \Level2Out98[20] , \Level2Out98[19] , \Level2Out98[18] , 
        \Level2Out98[17] , \Level2Out98[16] , \Level2Out98[15] , 
        \Level2Out98[14] , \Level2Out98[13] , \Level2Out98[12] , 
        \Level2Out98[11] , \Level2Out98[10] , \Level2Out98[9] , 
        \Level2Out98[8] , \Level2Out98[7] , \Level2Out98[6] , \Level2Out98[5] , 
        \Level2Out98[4] , \Level2Out98[3] , \Level2Out98[2] , \Level2Out98[1] , 
        \Level2Out98[0] }), .In1({\Level1Out98[31] , \Level1Out98[30] , 
        \Level1Out98[29] , \Level1Out98[28] , \Level1Out98[27] , 
        \Level1Out98[26] , \Level1Out98[25] , \Level1Out98[24] , 
        \Level1Out98[23] , \Level1Out98[22] , \Level1Out98[21] , 
        \Level1Out98[20] , \Level1Out98[19] , \Level1Out98[18] , 
        \Level1Out98[17] , \Level1Out98[16] , \Level1Out98[15] , 
        \Level1Out98[14] , \Level1Out98[13] , \Level1Out98[12] , 
        \Level1Out98[11] , \Level1Out98[10] , \Level1Out98[9] , 
        \Level1Out98[8] , \Level1Out98[7] , \Level1Out98[6] , \Level1Out98[5] , 
        \Level1Out98[4] , \Level1Out98[3] , \Level1Out98[2] , \Level1Out98[1] , 
        \Level1Out98[0] }), .In2({\Level1Out99[31] , \Level1Out99[30] , 
        \Level1Out99[29] , \Level1Out99[28] , \Level1Out99[27] , 
        \Level1Out99[26] , \Level1Out99[25] , \Level1Out99[24] , 
        \Level1Out99[23] , \Level1Out99[22] , \Level1Out99[21] , 
        \Level1Out99[20] , \Level1Out99[19] , \Level1Out99[18] , 
        \Level1Out99[17] , \Level1Out99[16] , \Level1Out99[15] , 
        \Level1Out99[14] , \Level1Out99[13] , \Level1Out99[12] , 
        \Level1Out99[11] , \Level1Out99[10] , \Level1Out99[9] , 
        \Level1Out99[8] , \Level1Out99[7] , \Level1Out99[6] , \Level1Out99[5] , 
        \Level1Out99[4] , \Level1Out99[3] , \Level1Out99[2] , \Level1Out99[1] , 
        \Level1Out99[0] }), .Read1(\Level1Load98[0] ), .Read2(
        \Level1Load99[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_84_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load84[0] ), .Out({\Level4Out84[31] , \Level4Out84[30] , 
        \Level4Out84[29] , \Level4Out84[28] , \Level4Out84[27] , 
        \Level4Out84[26] , \Level4Out84[25] , \Level4Out84[24] , 
        \Level4Out84[23] , \Level4Out84[22] , \Level4Out84[21] , 
        \Level4Out84[20] , \Level4Out84[19] , \Level4Out84[18] , 
        \Level4Out84[17] , \Level4Out84[16] , \Level4Out84[15] , 
        \Level4Out84[14] , \Level4Out84[13] , \Level4Out84[12] , 
        \Level4Out84[11] , \Level4Out84[10] , \Level4Out84[9] , 
        \Level4Out84[8] , \Level4Out84[7] , \Level4Out84[6] , \Level4Out84[5] , 
        \Level4Out84[4] , \Level4Out84[3] , \Level4Out84[2] , \Level4Out84[1] , 
        \Level4Out84[0] }), .In1({\Level2Out84[31] , \Level2Out84[30] , 
        \Level2Out84[29] , \Level2Out84[28] , \Level2Out84[27] , 
        \Level2Out84[26] , \Level2Out84[25] , \Level2Out84[24] , 
        \Level2Out84[23] , \Level2Out84[22] , \Level2Out84[21] , 
        \Level2Out84[20] , \Level2Out84[19] , \Level2Out84[18] , 
        \Level2Out84[17] , \Level2Out84[16] , \Level2Out84[15] , 
        \Level2Out84[14] , \Level2Out84[13] , \Level2Out84[12] , 
        \Level2Out84[11] , \Level2Out84[10] , \Level2Out84[9] , 
        \Level2Out84[8] , \Level2Out84[7] , \Level2Out84[6] , \Level2Out84[5] , 
        \Level2Out84[4] , \Level2Out84[3] , \Level2Out84[2] , \Level2Out84[1] , 
        \Level2Out84[0] }), .In2({\Level2Out86[31] , \Level2Out86[30] , 
        \Level2Out86[29] , \Level2Out86[28] , \Level2Out86[27] , 
        \Level2Out86[26] , \Level2Out86[25] , \Level2Out86[24] , 
        \Level2Out86[23] , \Level2Out86[22] , \Level2Out86[21] , 
        \Level2Out86[20] , \Level2Out86[19] , \Level2Out86[18] , 
        \Level2Out86[17] , \Level2Out86[16] , \Level2Out86[15] , 
        \Level2Out86[14] , \Level2Out86[13] , \Level2Out86[12] , 
        \Level2Out86[11] , \Level2Out86[10] , \Level2Out86[9] , 
        \Level2Out86[8] , \Level2Out86[7] , \Level2Out86[6] , \Level2Out86[5] , 
        \Level2Out86[4] , \Level2Out86[3] , \Level2Out86[2] , \Level2Out86[1] , 
        \Level2Out86[0] }), .Read1(\Level2Load84[0] ), .Read2(
        \Level2Load86[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_248_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load248[0] ), .Out({\Level8Out248[31] , \Level8Out248[30] , 
        \Level8Out248[29] , \Level8Out248[28] , \Level8Out248[27] , 
        \Level8Out248[26] , \Level8Out248[25] , \Level8Out248[24] , 
        \Level8Out248[23] , \Level8Out248[22] , \Level8Out248[21] , 
        \Level8Out248[20] , \Level8Out248[19] , \Level8Out248[18] , 
        \Level8Out248[17] , \Level8Out248[16] , \Level8Out248[15] , 
        \Level8Out248[14] , \Level8Out248[13] , \Level8Out248[12] , 
        \Level8Out248[11] , \Level8Out248[10] , \Level8Out248[9] , 
        \Level8Out248[8] , \Level8Out248[7] , \Level8Out248[6] , 
        \Level8Out248[5] , \Level8Out248[4] , \Level8Out248[3] , 
        \Level8Out248[2] , \Level8Out248[1] , \Level8Out248[0] }), .In1({
        \Level4Out248[31] , \Level4Out248[30] , \Level4Out248[29] , 
        \Level4Out248[28] , \Level4Out248[27] , \Level4Out248[26] , 
        \Level4Out248[25] , \Level4Out248[24] , \Level4Out248[23] , 
        \Level4Out248[22] , \Level4Out248[21] , \Level4Out248[20] , 
        \Level4Out248[19] , \Level4Out248[18] , \Level4Out248[17] , 
        \Level4Out248[16] , \Level4Out248[15] , \Level4Out248[14] , 
        \Level4Out248[13] , \Level4Out248[12] , \Level4Out248[11] , 
        \Level4Out248[10] , \Level4Out248[9] , \Level4Out248[8] , 
        \Level4Out248[7] , \Level4Out248[6] , \Level4Out248[5] , 
        \Level4Out248[4] , \Level4Out248[3] , \Level4Out248[2] , 
        \Level4Out248[1] , \Level4Out248[0] }), .In2({\Level4Out252[31] , 
        \Level4Out252[30] , \Level4Out252[29] , \Level4Out252[28] , 
        \Level4Out252[27] , \Level4Out252[26] , \Level4Out252[25] , 
        \Level4Out252[24] , \Level4Out252[23] , \Level4Out252[22] , 
        \Level4Out252[21] , \Level4Out252[20] , \Level4Out252[19] , 
        \Level4Out252[18] , \Level4Out252[17] , \Level4Out252[16] , 
        \Level4Out252[15] , \Level4Out252[14] , \Level4Out252[13] , 
        \Level4Out252[12] , \Level4Out252[11] , \Level4Out252[10] , 
        \Level4Out252[9] , \Level4Out252[8] , \Level4Out252[7] , 
        \Level4Out252[6] , \Level4Out252[5] , \Level4Out252[4] , 
        \Level4Out252[3] , \Level4Out252[2] , \Level4Out252[1] , 
        \Level4Out252[0] }), .Read1(\Level4Load248[0] ), .Read2(
        \Level4Load252[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load0[0] ), .Out({\Level16Out0[31] , \Level16Out0[30] , 
        \Level16Out0[29] , \Level16Out0[28] , \Level16Out0[27] , 
        \Level16Out0[26] , \Level16Out0[25] , \Level16Out0[24] , 
        \Level16Out0[23] , \Level16Out0[22] , \Level16Out0[21] , 
        \Level16Out0[20] , \Level16Out0[19] , \Level16Out0[18] , 
        \Level16Out0[17] , \Level16Out0[16] , \Level16Out0[15] , 
        \Level16Out0[14] , \Level16Out0[13] , \Level16Out0[12] , 
        \Level16Out0[11] , \Level16Out0[10] , \Level16Out0[9] , 
        \Level16Out0[8] , \Level16Out0[7] , \Level16Out0[6] , \Level16Out0[5] , 
        \Level16Out0[4] , \Level16Out0[3] , \Level16Out0[2] , \Level16Out0[1] , 
        \Level16Out0[0] }), .In1({\Level8Out0[31] , \Level8Out0[30] , 
        \Level8Out0[29] , \Level8Out0[28] , \Level8Out0[27] , \Level8Out0[26] , 
        \Level8Out0[25] , \Level8Out0[24] , \Level8Out0[23] , \Level8Out0[22] , 
        \Level8Out0[21] , \Level8Out0[20] , \Level8Out0[19] , \Level8Out0[18] , 
        \Level8Out0[17] , \Level8Out0[16] , \Level8Out0[15] , \Level8Out0[14] , 
        \Level8Out0[13] , \Level8Out0[12] , \Level8Out0[11] , \Level8Out0[10] , 
        \Level8Out0[9] , \Level8Out0[8] , \Level8Out0[7] , \Level8Out0[6] , 
        \Level8Out0[5] , \Level8Out0[4] , \Level8Out0[3] , \Level8Out0[2] , 
        \Level8Out0[1] , \Level8Out0[0] }), .In2({\Level8Out8[31] , 
        \Level8Out8[30] , \Level8Out8[29] , \Level8Out8[28] , \Level8Out8[27] , 
        \Level8Out8[26] , \Level8Out8[25] , \Level8Out8[24] , \Level8Out8[23] , 
        \Level8Out8[22] , \Level8Out8[21] , \Level8Out8[20] , \Level8Out8[19] , 
        \Level8Out8[18] , \Level8Out8[17] , \Level8Out8[16] , \Level8Out8[15] , 
        \Level8Out8[14] , \Level8Out8[13] , \Level8Out8[12] , \Level8Out8[11] , 
        \Level8Out8[10] , \Level8Out8[9] , \Level8Out8[8] , \Level8Out8[7] , 
        \Level8Out8[6] , \Level8Out8[5] , \Level8Out8[4] , \Level8Out8[3] , 
        \Level8Out8[2] , \Level8Out8[1] , \Level8Out8[0] }), .Read1(
        \Level8Load0[0] ), .Read2(\Level8Load8[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_65 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink65[31] , \ScanLink65[30] , 
        \ScanLink65[29] , \ScanLink65[28] , \ScanLink65[27] , \ScanLink65[26] , 
        \ScanLink65[25] , \ScanLink65[24] , \ScanLink65[23] , \ScanLink65[22] , 
        \ScanLink65[21] , \ScanLink65[20] , \ScanLink65[19] , \ScanLink65[18] , 
        \ScanLink65[17] , \ScanLink65[16] , \ScanLink65[15] , \ScanLink65[14] , 
        \ScanLink65[13] , \ScanLink65[12] , \ScanLink65[11] , \ScanLink65[10] , 
        \ScanLink65[9] , \ScanLink65[8] , \ScanLink65[7] , \ScanLink65[6] , 
        \ScanLink65[5] , \ScanLink65[4] , \ScanLink65[3] , \ScanLink65[2] , 
        \ScanLink65[1] , \ScanLink65[0] }), .ScanOut({\ScanLink66[31] , 
        \ScanLink66[30] , \ScanLink66[29] , \ScanLink66[28] , \ScanLink66[27] , 
        \ScanLink66[26] , \ScanLink66[25] , \ScanLink66[24] , \ScanLink66[23] , 
        \ScanLink66[22] , \ScanLink66[21] , \ScanLink66[20] , \ScanLink66[19] , 
        \ScanLink66[18] , \ScanLink66[17] , \ScanLink66[16] , \ScanLink66[15] , 
        \ScanLink66[14] , \ScanLink66[13] , \ScanLink66[12] , \ScanLink66[11] , 
        \ScanLink66[10] , \ScanLink66[9] , \ScanLink66[8] , \ScanLink66[7] , 
        \ScanLink66[6] , \ScanLink66[5] , \ScanLink66[4] , \ScanLink66[3] , 
        \ScanLink66[2] , \ScanLink66[1] , \ScanLink66[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load65[0] ), .Out({
        \Level1Out65[31] , \Level1Out65[30] , \Level1Out65[29] , 
        \Level1Out65[28] , \Level1Out65[27] , \Level1Out65[26] , 
        \Level1Out65[25] , \Level1Out65[24] , \Level1Out65[23] , 
        \Level1Out65[22] , \Level1Out65[21] , \Level1Out65[20] , 
        \Level1Out65[19] , \Level1Out65[18] , \Level1Out65[17] , 
        \Level1Out65[16] , \Level1Out65[15] , \Level1Out65[14] , 
        \Level1Out65[13] , \Level1Out65[12] , \Level1Out65[11] , 
        \Level1Out65[10] , \Level1Out65[9] , \Level1Out65[8] , 
        \Level1Out65[7] , \Level1Out65[6] , \Level1Out65[5] , \Level1Out65[4] , 
        \Level1Out65[3] , \Level1Out65[2] , \Level1Out65[1] , \Level1Out65[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_147 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink147[31] , \ScanLink147[30] , 
        \ScanLink147[29] , \ScanLink147[28] , \ScanLink147[27] , 
        \ScanLink147[26] , \ScanLink147[25] , \ScanLink147[24] , 
        \ScanLink147[23] , \ScanLink147[22] , \ScanLink147[21] , 
        \ScanLink147[20] , \ScanLink147[19] , \ScanLink147[18] , 
        \ScanLink147[17] , \ScanLink147[16] , \ScanLink147[15] , 
        \ScanLink147[14] , \ScanLink147[13] , \ScanLink147[12] , 
        \ScanLink147[11] , \ScanLink147[10] , \ScanLink147[9] , 
        \ScanLink147[8] , \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , 
        \ScanLink147[4] , \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , 
        \ScanLink147[0] }), .ScanOut({\ScanLink148[31] , \ScanLink148[30] , 
        \ScanLink148[29] , \ScanLink148[28] , \ScanLink148[27] , 
        \ScanLink148[26] , \ScanLink148[25] , \ScanLink148[24] , 
        \ScanLink148[23] , \ScanLink148[22] , \ScanLink148[21] , 
        \ScanLink148[20] , \ScanLink148[19] , \ScanLink148[18] , 
        \ScanLink148[17] , \ScanLink148[16] , \ScanLink148[15] , 
        \ScanLink148[14] , \ScanLink148[13] , \ScanLink148[12] , 
        \ScanLink148[11] , \ScanLink148[10] , \ScanLink148[9] , 
        \ScanLink148[8] , \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , 
        \ScanLink148[4] , \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , 
        \ScanLink148[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load147[0] ), .Out({\Level1Out147[31] , \Level1Out147[30] , 
        \Level1Out147[29] , \Level1Out147[28] , \Level1Out147[27] , 
        \Level1Out147[26] , \Level1Out147[25] , \Level1Out147[24] , 
        \Level1Out147[23] , \Level1Out147[22] , \Level1Out147[21] , 
        \Level1Out147[20] , \Level1Out147[19] , \Level1Out147[18] , 
        \Level1Out147[17] , \Level1Out147[16] , \Level1Out147[15] , 
        \Level1Out147[14] , \Level1Out147[13] , \Level1Out147[12] , 
        \Level1Out147[11] , \Level1Out147[10] , \Level1Out147[9] , 
        \Level1Out147[8] , \Level1Out147[7] , \Level1Out147[6] , 
        \Level1Out147[5] , \Level1Out147[4] , \Level1Out147[3] , 
        \Level1Out147[2] , \Level1Out147[1] , \Level1Out147[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_160 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink160[31] , \ScanLink160[30] , 
        \ScanLink160[29] , \ScanLink160[28] , \ScanLink160[27] , 
        \ScanLink160[26] , \ScanLink160[25] , \ScanLink160[24] , 
        \ScanLink160[23] , \ScanLink160[22] , \ScanLink160[21] , 
        \ScanLink160[20] , \ScanLink160[19] , \ScanLink160[18] , 
        \ScanLink160[17] , \ScanLink160[16] , \ScanLink160[15] , 
        \ScanLink160[14] , \ScanLink160[13] , \ScanLink160[12] , 
        \ScanLink160[11] , \ScanLink160[10] , \ScanLink160[9] , 
        \ScanLink160[8] , \ScanLink160[7] , \ScanLink160[6] , \ScanLink160[5] , 
        \ScanLink160[4] , \ScanLink160[3] , \ScanLink160[2] , \ScanLink160[1] , 
        \ScanLink160[0] }), .ScanOut({\ScanLink161[31] , \ScanLink161[30] , 
        \ScanLink161[29] , \ScanLink161[28] , \ScanLink161[27] , 
        \ScanLink161[26] , \ScanLink161[25] , \ScanLink161[24] , 
        \ScanLink161[23] , \ScanLink161[22] , \ScanLink161[21] , 
        \ScanLink161[20] , \ScanLink161[19] , \ScanLink161[18] , 
        \ScanLink161[17] , \ScanLink161[16] , \ScanLink161[15] , 
        \ScanLink161[14] , \ScanLink161[13] , \ScanLink161[12] , 
        \ScanLink161[11] , \ScanLink161[10] , \ScanLink161[9] , 
        \ScanLink161[8] , \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , 
        \ScanLink161[4] , \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , 
        \ScanLink161[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load160[0] ), .Out({\Level1Out160[31] , \Level1Out160[30] , 
        \Level1Out160[29] , \Level1Out160[28] , \Level1Out160[27] , 
        \Level1Out160[26] , \Level1Out160[25] , \Level1Out160[24] , 
        \Level1Out160[23] , \Level1Out160[22] , \Level1Out160[21] , 
        \Level1Out160[20] , \Level1Out160[19] , \Level1Out160[18] , 
        \Level1Out160[17] , \Level1Out160[16] , \Level1Out160[15] , 
        \Level1Out160[14] , \Level1Out160[13] , \Level1Out160[12] , 
        \Level1Out160[11] , \Level1Out160[10] , \Level1Out160[9] , 
        \Level1Out160[8] , \Level1Out160[7] , \Level1Out160[6] , 
        \Level1Out160[5] , \Level1Out160[4] , \Level1Out160[3] , 
        \Level1Out160[2] , \Level1Out160[1] , \Level1Out160[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level64Load64[0] ), .Out({\Level64Out64[31] , \Level64Out64[30] , 
        \Level64Out64[29] , \Level64Out64[28] , \Level64Out64[27] , 
        \Level64Out64[26] , \Level64Out64[25] , \Level64Out64[24] , 
        \Level64Out64[23] , \Level64Out64[22] , \Level64Out64[21] , 
        \Level64Out64[20] , \Level64Out64[19] , \Level64Out64[18] , 
        \Level64Out64[17] , \Level64Out64[16] , \Level64Out64[15] , 
        \Level64Out64[14] , \Level64Out64[13] , \Level64Out64[12] , 
        \Level64Out64[11] , \Level64Out64[10] , \Level64Out64[9] , 
        \Level64Out64[8] , \Level64Out64[7] , \Level64Out64[6] , 
        \Level64Out64[5] , \Level64Out64[4] , \Level64Out64[3] , 
        \Level64Out64[2] , \Level64Out64[1] , \Level64Out64[0] }), .In1({
        \Level32Out64[31] , \Level32Out64[30] , \Level32Out64[29] , 
        \Level32Out64[28] , \Level32Out64[27] , \Level32Out64[26] , 
        \Level32Out64[25] , \Level32Out64[24] , \Level32Out64[23] , 
        \Level32Out64[22] , \Level32Out64[21] , \Level32Out64[20] , 
        \Level32Out64[19] , \Level32Out64[18] , \Level32Out64[17] , 
        \Level32Out64[16] , \Level32Out64[15] , \Level32Out64[14] , 
        \Level32Out64[13] , \Level32Out64[12] , \Level32Out64[11] , 
        \Level32Out64[10] , \Level32Out64[9] , \Level32Out64[8] , 
        \Level32Out64[7] , \Level32Out64[6] , \Level32Out64[5] , 
        \Level32Out64[4] , \Level32Out64[3] , \Level32Out64[2] , 
        \Level32Out64[1] , \Level32Out64[0] }), .In2({\Level32Out96[31] , 
        \Level32Out96[30] , \Level32Out96[29] , \Level32Out96[28] , 
        \Level32Out96[27] , \Level32Out96[26] , \Level32Out96[25] , 
        \Level32Out96[24] , \Level32Out96[23] , \Level32Out96[22] , 
        \Level32Out96[21] , \Level32Out96[20] , \Level32Out96[19] , 
        \Level32Out96[18] , \Level32Out96[17] , \Level32Out96[16] , 
        \Level32Out96[15] , \Level32Out96[14] , \Level32Out96[13] , 
        \Level32Out96[12] , \Level32Out96[11] , \Level32Out96[10] , 
        \Level32Out96[9] , \Level32Out96[8] , \Level32Out96[7] , 
        \Level32Out96[6] , \Level32Out96[5] , \Level32Out96[4] , 
        \Level32Out96[3] , \Level32Out96[2] , \Level32Out96[1] , 
        \Level32Out96[0] }), .Read1(\Level32Load64[0] ), .Read2(
        \Level32Load96[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_250 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink250[31] , \ScanLink250[30] , 
        \ScanLink250[29] , \ScanLink250[28] , \ScanLink250[27] , 
        \ScanLink250[26] , \ScanLink250[25] , \ScanLink250[24] , 
        \ScanLink250[23] , \ScanLink250[22] , \ScanLink250[21] , 
        \ScanLink250[20] , \ScanLink250[19] , \ScanLink250[18] , 
        \ScanLink250[17] , \ScanLink250[16] , \ScanLink250[15] , 
        \ScanLink250[14] , \ScanLink250[13] , \ScanLink250[12] , 
        \ScanLink250[11] , \ScanLink250[10] , \ScanLink250[9] , 
        \ScanLink250[8] , \ScanLink250[7] , \ScanLink250[6] , \ScanLink250[5] , 
        \ScanLink250[4] , \ScanLink250[3] , \ScanLink250[2] , \ScanLink250[1] , 
        \ScanLink250[0] }), .ScanOut({\ScanLink251[31] , \ScanLink251[30] , 
        \ScanLink251[29] , \ScanLink251[28] , \ScanLink251[27] , 
        \ScanLink251[26] , \ScanLink251[25] , \ScanLink251[24] , 
        \ScanLink251[23] , \ScanLink251[22] , \ScanLink251[21] , 
        \ScanLink251[20] , \ScanLink251[19] , \ScanLink251[18] , 
        \ScanLink251[17] , \ScanLink251[16] , \ScanLink251[15] , 
        \ScanLink251[14] , \ScanLink251[13] , \ScanLink251[12] , 
        \ScanLink251[11] , \ScanLink251[10] , \ScanLink251[9] , 
        \ScanLink251[8] , \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , 
        \ScanLink251[4] , \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , 
        \ScanLink251[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load250[0] ), .Out({\Level1Out250[31] , \Level1Out250[30] , 
        \Level1Out250[29] , \Level1Out250[28] , \Level1Out250[27] , 
        \Level1Out250[26] , \Level1Out250[25] , \Level1Out250[24] , 
        \Level1Out250[23] , \Level1Out250[22] , \Level1Out250[21] , 
        \Level1Out250[20] , \Level1Out250[19] , \Level1Out250[18] , 
        \Level1Out250[17] , \Level1Out250[16] , \Level1Out250[15] , 
        \Level1Out250[14] , \Level1Out250[13] , \Level1Out250[12] , 
        \Level1Out250[11] , \Level1Out250[10] , \Level1Out250[9] , 
        \Level1Out250[8] , \Level1Out250[7] , \Level1Out250[6] , 
        \Level1Out250[5] , \Level1Out250[4] , \Level1Out250[3] , 
        \Level1Out250[2] , \Level1Out250[1] , \Level1Out250[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_112_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load112[0] ), .Out({\Level16Out112[31] , \Level16Out112[30] , 
        \Level16Out112[29] , \Level16Out112[28] , \Level16Out112[27] , 
        \Level16Out112[26] , \Level16Out112[25] , \Level16Out112[24] , 
        \Level16Out112[23] , \Level16Out112[22] , \Level16Out112[21] , 
        \Level16Out112[20] , \Level16Out112[19] , \Level16Out112[18] , 
        \Level16Out112[17] , \Level16Out112[16] , \Level16Out112[15] , 
        \Level16Out112[14] , \Level16Out112[13] , \Level16Out112[12] , 
        \Level16Out112[11] , \Level16Out112[10] , \Level16Out112[9] , 
        \Level16Out112[8] , \Level16Out112[7] , \Level16Out112[6] , 
        \Level16Out112[5] , \Level16Out112[4] , \Level16Out112[3] , 
        \Level16Out112[2] , \Level16Out112[1] , \Level16Out112[0] }), .In1({
        \Level8Out112[31] , \Level8Out112[30] , \Level8Out112[29] , 
        \Level8Out112[28] , \Level8Out112[27] , \Level8Out112[26] , 
        \Level8Out112[25] , \Level8Out112[24] , \Level8Out112[23] , 
        \Level8Out112[22] , \Level8Out112[21] , \Level8Out112[20] , 
        \Level8Out112[19] , \Level8Out112[18] , \Level8Out112[17] , 
        \Level8Out112[16] , \Level8Out112[15] , \Level8Out112[14] , 
        \Level8Out112[13] , \Level8Out112[12] , \Level8Out112[11] , 
        \Level8Out112[10] , \Level8Out112[9] , \Level8Out112[8] , 
        \Level8Out112[7] , \Level8Out112[6] , \Level8Out112[5] , 
        \Level8Out112[4] , \Level8Out112[3] , \Level8Out112[2] , 
        \Level8Out112[1] , \Level8Out112[0] }), .In2({\Level8Out120[31] , 
        \Level8Out120[30] , \Level8Out120[29] , \Level8Out120[28] , 
        \Level8Out120[27] , \Level8Out120[26] , \Level8Out120[25] , 
        \Level8Out120[24] , \Level8Out120[23] , \Level8Out120[22] , 
        \Level8Out120[21] , \Level8Out120[20] , \Level8Out120[19] , 
        \Level8Out120[18] , \Level8Out120[17] , \Level8Out120[16] , 
        \Level8Out120[15] , \Level8Out120[14] , \Level8Out120[13] , 
        \Level8Out120[12] , \Level8Out120[11] , \Level8Out120[10] , 
        \Level8Out120[9] , \Level8Out120[8] , \Level8Out120[7] , 
        \Level8Out120[6] , \Level8Out120[5] , \Level8Out120[4] , 
        \Level8Out120[3] , \Level8Out120[2] , \Level8Out120[1] , 
        \Level8Out120[0] }), .Read1(\Level8Load112[0] ), .Read2(
        \Level8Load120[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_80 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink80[31] , \ScanLink80[30] , 
        \ScanLink80[29] , \ScanLink80[28] , \ScanLink80[27] , \ScanLink80[26] , 
        \ScanLink80[25] , \ScanLink80[24] , \ScanLink80[23] , \ScanLink80[22] , 
        \ScanLink80[21] , \ScanLink80[20] , \ScanLink80[19] , \ScanLink80[18] , 
        \ScanLink80[17] , \ScanLink80[16] , \ScanLink80[15] , \ScanLink80[14] , 
        \ScanLink80[13] , \ScanLink80[12] , \ScanLink80[11] , \ScanLink80[10] , 
        \ScanLink80[9] , \ScanLink80[8] , \ScanLink80[7] , \ScanLink80[6] , 
        \ScanLink80[5] , \ScanLink80[4] , \ScanLink80[3] , \ScanLink80[2] , 
        \ScanLink80[1] , \ScanLink80[0] }), .ScanOut({\ScanLink81[31] , 
        \ScanLink81[30] , \ScanLink81[29] , \ScanLink81[28] , \ScanLink81[27] , 
        \ScanLink81[26] , \ScanLink81[25] , \ScanLink81[24] , \ScanLink81[23] , 
        \ScanLink81[22] , \ScanLink81[21] , \ScanLink81[20] , \ScanLink81[19] , 
        \ScanLink81[18] , \ScanLink81[17] , \ScanLink81[16] , \ScanLink81[15] , 
        \ScanLink81[14] , \ScanLink81[13] , \ScanLink81[12] , \ScanLink81[11] , 
        \ScanLink81[10] , \ScanLink81[9] , \ScanLink81[8] , \ScanLink81[7] , 
        \ScanLink81[6] , \ScanLink81[5] , \ScanLink81[4] , \ScanLink81[3] , 
        \ScanLink81[2] , \ScanLink81[1] , \ScanLink81[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load80[0] ), .Out({
        \Level1Out80[31] , \Level1Out80[30] , \Level1Out80[29] , 
        \Level1Out80[28] , \Level1Out80[27] , \Level1Out80[26] , 
        \Level1Out80[25] , \Level1Out80[24] , \Level1Out80[23] , 
        \Level1Out80[22] , \Level1Out80[21] , \Level1Out80[20] , 
        \Level1Out80[19] , \Level1Out80[18] , \Level1Out80[17] , 
        \Level1Out80[16] , \Level1Out80[15] , \Level1Out80[14] , 
        \Level1Out80[13] , \Level1Out80[12] , \Level1Out80[11] , 
        \Level1Out80[10] , \Level1Out80[9] , \Level1Out80[8] , 
        \Level1Out80[7] , \Level1Out80[6] , \Level1Out80[5] , \Level1Out80[4] , 
        \Level1Out80[3] , \Level1Out80[2] , \Level1Out80[1] , \Level1Out80[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_129 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink129[31] , \ScanLink129[30] , 
        \ScanLink129[29] , \ScanLink129[28] , \ScanLink129[27] , 
        \ScanLink129[26] , \ScanLink129[25] , \ScanLink129[24] , 
        \ScanLink129[23] , \ScanLink129[22] , \ScanLink129[21] , 
        \ScanLink129[20] , \ScanLink129[19] , \ScanLink129[18] , 
        \ScanLink129[17] , \ScanLink129[16] , \ScanLink129[15] , 
        \ScanLink129[14] , \ScanLink129[13] , \ScanLink129[12] , 
        \ScanLink129[11] , \ScanLink129[10] , \ScanLink129[9] , 
        \ScanLink129[8] , \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , 
        \ScanLink129[4] , \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , 
        \ScanLink129[0] }), .ScanOut({\ScanLink130[31] , \ScanLink130[30] , 
        \ScanLink130[29] , \ScanLink130[28] , \ScanLink130[27] , 
        \ScanLink130[26] , \ScanLink130[25] , \ScanLink130[24] , 
        \ScanLink130[23] , \ScanLink130[22] , \ScanLink130[21] , 
        \ScanLink130[20] , \ScanLink130[19] , \ScanLink130[18] , 
        \ScanLink130[17] , \ScanLink130[16] , \ScanLink130[15] , 
        \ScanLink130[14] , \ScanLink130[13] , \ScanLink130[12] , 
        \ScanLink130[11] , \ScanLink130[10] , \ScanLink130[9] , 
        \ScanLink130[8] , \ScanLink130[7] , \ScanLink130[6] , \ScanLink130[5] , 
        \ScanLink130[4] , \ScanLink130[3] , \ScanLink130[2] , \ScanLink130[1] , 
        \ScanLink130[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load129[0] ), .Out({\Level1Out129[31] , \Level1Out129[30] , 
        \Level1Out129[29] , \Level1Out129[28] , \Level1Out129[27] , 
        \Level1Out129[26] , \Level1Out129[25] , \Level1Out129[24] , 
        \Level1Out129[23] , \Level1Out129[22] , \Level1Out129[21] , 
        \Level1Out129[20] , \Level1Out129[19] , \Level1Out129[18] , 
        \Level1Out129[17] , \Level1Out129[16] , \Level1Out129[15] , 
        \Level1Out129[14] , \Level1Out129[13] , \Level1Out129[12] , 
        \Level1Out129[11] , \Level1Out129[10] , \Level1Out129[9] , 
        \Level1Out129[8] , \Level1Out129[7] , \Level1Out129[6] , 
        \Level1Out129[5] , \Level1Out129[4] , \Level1Out129[3] , 
        \Level1Out129[2] , \Level1Out129[1] , \Level1Out129[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_185 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink185[31] , \ScanLink185[30] , 
        \ScanLink185[29] , \ScanLink185[28] , \ScanLink185[27] , 
        \ScanLink185[26] , \ScanLink185[25] , \ScanLink185[24] , 
        \ScanLink185[23] , \ScanLink185[22] , \ScanLink185[21] , 
        \ScanLink185[20] , \ScanLink185[19] , \ScanLink185[18] , 
        \ScanLink185[17] , \ScanLink185[16] , \ScanLink185[15] , 
        \ScanLink185[14] , \ScanLink185[13] , \ScanLink185[12] , 
        \ScanLink185[11] , \ScanLink185[10] , \ScanLink185[9] , 
        \ScanLink185[8] , \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , 
        \ScanLink185[4] , \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , 
        \ScanLink185[0] }), .ScanOut({\ScanLink186[31] , \ScanLink186[30] , 
        \ScanLink186[29] , \ScanLink186[28] , \ScanLink186[27] , 
        \ScanLink186[26] , \ScanLink186[25] , \ScanLink186[24] , 
        \ScanLink186[23] , \ScanLink186[22] , \ScanLink186[21] , 
        \ScanLink186[20] , \ScanLink186[19] , \ScanLink186[18] , 
        \ScanLink186[17] , \ScanLink186[16] , \ScanLink186[15] , 
        \ScanLink186[14] , \ScanLink186[13] , \ScanLink186[12] , 
        \ScanLink186[11] , \ScanLink186[10] , \ScanLink186[9] , 
        \ScanLink186[8] , \ScanLink186[7] , \ScanLink186[6] , \ScanLink186[5] , 
        \ScanLink186[4] , \ScanLink186[3] , \ScanLink186[2] , \ScanLink186[1] , 
        \ScanLink186[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load185[0] ), .Out({\Level1Out185[31] , \Level1Out185[30] , 
        \Level1Out185[29] , \Level1Out185[28] , \Level1Out185[27] , 
        \Level1Out185[26] , \Level1Out185[25] , \Level1Out185[24] , 
        \Level1Out185[23] , \Level1Out185[22] , \Level1Out185[21] , 
        \Level1Out185[20] , \Level1Out185[19] , \Level1Out185[18] , 
        \Level1Out185[17] , \Level1Out185[16] , \Level1Out185[15] , 
        \Level1Out185[14] , \Level1Out185[13] , \Level1Out185[12] , 
        \Level1Out185[11] , \Level1Out185[10] , \Level1Out185[9] , 
        \Level1Out185[8] , \Level1Out185[7] , \Level1Out185[6] , 
        \Level1Out185[5] , \Level1Out185[4] , \Level1Out185[3] , 
        \Level1Out185[2] , \Level1Out185[1] , \Level1Out185[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load16[0] ), .Out({\Level2Out16[31] , \Level2Out16[30] , 
        \Level2Out16[29] , \Level2Out16[28] , \Level2Out16[27] , 
        \Level2Out16[26] , \Level2Out16[25] , \Level2Out16[24] , 
        \Level2Out16[23] , \Level2Out16[22] , \Level2Out16[21] , 
        \Level2Out16[20] , \Level2Out16[19] , \Level2Out16[18] , 
        \Level2Out16[17] , \Level2Out16[16] , \Level2Out16[15] , 
        \Level2Out16[14] , \Level2Out16[13] , \Level2Out16[12] , 
        \Level2Out16[11] , \Level2Out16[10] , \Level2Out16[9] , 
        \Level2Out16[8] , \Level2Out16[7] , \Level2Out16[6] , \Level2Out16[5] , 
        \Level2Out16[4] , \Level2Out16[3] , \Level2Out16[2] , \Level2Out16[1] , 
        \Level2Out16[0] }), .In1({\Level1Out16[31] , \Level1Out16[30] , 
        \Level1Out16[29] , \Level1Out16[28] , \Level1Out16[27] , 
        \Level1Out16[26] , \Level1Out16[25] , \Level1Out16[24] , 
        \Level1Out16[23] , \Level1Out16[22] , \Level1Out16[21] , 
        \Level1Out16[20] , \Level1Out16[19] , \Level1Out16[18] , 
        \Level1Out16[17] , \Level1Out16[16] , \Level1Out16[15] , 
        \Level1Out16[14] , \Level1Out16[13] , \Level1Out16[12] , 
        \Level1Out16[11] , \Level1Out16[10] , \Level1Out16[9] , 
        \Level1Out16[8] , \Level1Out16[7] , \Level1Out16[6] , \Level1Out16[5] , 
        \Level1Out16[4] , \Level1Out16[3] , \Level1Out16[2] , \Level1Out16[1] , 
        \Level1Out16[0] }), .In2({\Level1Out17[31] , \Level1Out17[30] , 
        \Level1Out17[29] , \Level1Out17[28] , \Level1Out17[27] , 
        \Level1Out17[26] , \Level1Out17[25] , \Level1Out17[24] , 
        \Level1Out17[23] , \Level1Out17[22] , \Level1Out17[21] , 
        \Level1Out17[20] , \Level1Out17[19] , \Level1Out17[18] , 
        \Level1Out17[17] , \Level1Out17[16] , \Level1Out17[15] , 
        \Level1Out17[14] , \Level1Out17[13] , \Level1Out17[12] , 
        \Level1Out17[11] , \Level1Out17[10] , \Level1Out17[9] , 
        \Level1Out17[8] , \Level1Out17[7] , \Level1Out17[6] , \Level1Out17[5] , 
        \Level1Out17[4] , \Level1Out17[3] , \Level1Out17[2] , \Level1Out17[1] , 
        \Level1Out17[0] }), .Read1(\Level1Load16[0] ), .Read2(
        \Level1Load17[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_150_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load150[0] ), .Out({\Level2Out150[31] , \Level2Out150[30] , 
        \Level2Out150[29] , \Level2Out150[28] , \Level2Out150[27] , 
        \Level2Out150[26] , \Level2Out150[25] , \Level2Out150[24] , 
        \Level2Out150[23] , \Level2Out150[22] , \Level2Out150[21] , 
        \Level2Out150[20] , \Level2Out150[19] , \Level2Out150[18] , 
        \Level2Out150[17] , \Level2Out150[16] , \Level2Out150[15] , 
        \Level2Out150[14] , \Level2Out150[13] , \Level2Out150[12] , 
        \Level2Out150[11] , \Level2Out150[10] , \Level2Out150[9] , 
        \Level2Out150[8] , \Level2Out150[7] , \Level2Out150[6] , 
        \Level2Out150[5] , \Level2Out150[4] , \Level2Out150[3] , 
        \Level2Out150[2] , \Level2Out150[1] , \Level2Out150[0] }), .In1({
        \Level1Out150[31] , \Level1Out150[30] , \Level1Out150[29] , 
        \Level1Out150[28] , \Level1Out150[27] , \Level1Out150[26] , 
        \Level1Out150[25] , \Level1Out150[24] , \Level1Out150[23] , 
        \Level1Out150[22] , \Level1Out150[21] , \Level1Out150[20] , 
        \Level1Out150[19] , \Level1Out150[18] , \Level1Out150[17] , 
        \Level1Out150[16] , \Level1Out150[15] , \Level1Out150[14] , 
        \Level1Out150[13] , \Level1Out150[12] , \Level1Out150[11] , 
        \Level1Out150[10] , \Level1Out150[9] , \Level1Out150[8] , 
        \Level1Out150[7] , \Level1Out150[6] , \Level1Out150[5] , 
        \Level1Out150[4] , \Level1Out150[3] , \Level1Out150[2] , 
        \Level1Out150[1] , \Level1Out150[0] }), .In2({\Level1Out151[31] , 
        \Level1Out151[30] , \Level1Out151[29] , \Level1Out151[28] , 
        \Level1Out151[27] , \Level1Out151[26] , \Level1Out151[25] , 
        \Level1Out151[24] , \Level1Out151[23] , \Level1Out151[22] , 
        \Level1Out151[21] , \Level1Out151[20] , \Level1Out151[19] , 
        \Level1Out151[18] , \Level1Out151[17] , \Level1Out151[16] , 
        \Level1Out151[15] , \Level1Out151[14] , \Level1Out151[13] , 
        \Level1Out151[12] , \Level1Out151[11] , \Level1Out151[10] , 
        \Level1Out151[9] , \Level1Out151[8] , \Level1Out151[7] , 
        \Level1Out151[6] , \Level1Out151[5] , \Level1Out151[4] , 
        \Level1Out151[3] , \Level1Out151[2] , \Level1Out151[1] , 
        \Level1Out151[0] }), .Read1(\Level1Load150[0] ), .Read2(
        \Level1Load151[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_252_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load252[0] ), .Out({\Level4Out252[31] , \Level4Out252[30] , 
        \Level4Out252[29] , \Level4Out252[28] , \Level4Out252[27] , 
        \Level4Out252[26] , \Level4Out252[25] , \Level4Out252[24] , 
        \Level4Out252[23] , \Level4Out252[22] , \Level4Out252[21] , 
        \Level4Out252[20] , \Level4Out252[19] , \Level4Out252[18] , 
        \Level4Out252[17] , \Level4Out252[16] , \Level4Out252[15] , 
        \Level4Out252[14] , \Level4Out252[13] , \Level4Out252[12] , 
        \Level4Out252[11] , \Level4Out252[10] , \Level4Out252[9] , 
        \Level4Out252[8] , \Level4Out252[7] , \Level4Out252[6] , 
        \Level4Out252[5] , \Level4Out252[4] , \Level4Out252[3] , 
        \Level4Out252[2] , \Level4Out252[1] , \Level4Out252[0] }), .In1({
        \Level2Out252[31] , \Level2Out252[30] , \Level2Out252[29] , 
        \Level2Out252[28] , \Level2Out252[27] , \Level2Out252[26] , 
        \Level2Out252[25] , \Level2Out252[24] , \Level2Out252[23] , 
        \Level2Out252[22] , \Level2Out252[21] , \Level2Out252[20] , 
        \Level2Out252[19] , \Level2Out252[18] , \Level2Out252[17] , 
        \Level2Out252[16] , \Level2Out252[15] , \Level2Out252[14] , 
        \Level2Out252[13] , \Level2Out252[12] , \Level2Out252[11] , 
        \Level2Out252[10] , \Level2Out252[9] , \Level2Out252[8] , 
        \Level2Out252[7] , \Level2Out252[6] , \Level2Out252[5] , 
        \Level2Out252[4] , \Level2Out252[3] , \Level2Out252[2] , 
        \Level2Out252[1] , \Level2Out252[0] }), .In2({\Level2Out254[31] , 
        \Level2Out254[30] , \Level2Out254[29] , \Level2Out254[28] , 
        \Level2Out254[27] , \Level2Out254[26] , \Level2Out254[25] , 
        \Level2Out254[24] , \Level2Out254[23] , \Level2Out254[22] , 
        \Level2Out254[21] , \Level2Out254[20] , \Level2Out254[19] , 
        \Level2Out254[18] , \Level2Out254[17] , \Level2Out254[16] , 
        \Level2Out254[15] , \Level2Out254[14] , \Level2Out254[13] , 
        \Level2Out254[12] , \Level2Out254[11] , \Level2Out254[10] , 
        \Level2Out254[9] , \Level2Out254[8] , \Level2Out254[7] , 
        \Level2Out254[6] , \Level2Out254[5] , \Level2Out254[4] , 
        \Level2Out254[3] , \Level2Out254[2] , \Level2Out254[1] , 
        \Level2Out254[0] }), .Read1(\Level2Load252[0] ), .Read2(
        \Level2Load254[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_20_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load20[0] ), .Out({\Level4Out20[31] , \Level4Out20[30] , 
        \Level4Out20[29] , \Level4Out20[28] , \Level4Out20[27] , 
        \Level4Out20[26] , \Level4Out20[25] , \Level4Out20[24] , 
        \Level4Out20[23] , \Level4Out20[22] , \Level4Out20[21] , 
        \Level4Out20[20] , \Level4Out20[19] , \Level4Out20[18] , 
        \Level4Out20[17] , \Level4Out20[16] , \Level4Out20[15] , 
        \Level4Out20[14] , \Level4Out20[13] , \Level4Out20[12] , 
        \Level4Out20[11] , \Level4Out20[10] , \Level4Out20[9] , 
        \Level4Out20[8] , \Level4Out20[7] , \Level4Out20[6] , \Level4Out20[5] , 
        \Level4Out20[4] , \Level4Out20[3] , \Level4Out20[2] , \Level4Out20[1] , 
        \Level4Out20[0] }), .In1({\Level2Out20[31] , \Level2Out20[30] , 
        \Level2Out20[29] , \Level2Out20[28] , \Level2Out20[27] , 
        \Level2Out20[26] , \Level2Out20[25] , \Level2Out20[24] , 
        \Level2Out20[23] , \Level2Out20[22] , \Level2Out20[21] , 
        \Level2Out20[20] , \Level2Out20[19] , \Level2Out20[18] , 
        \Level2Out20[17] , \Level2Out20[16] , \Level2Out20[15] , 
        \Level2Out20[14] , \Level2Out20[13] , \Level2Out20[12] , 
        \Level2Out20[11] , \Level2Out20[10] , \Level2Out20[9] , 
        \Level2Out20[8] , \Level2Out20[7] , \Level2Out20[6] , \Level2Out20[5] , 
        \Level2Out20[4] , \Level2Out20[3] , \Level2Out20[2] , \Level2Out20[1] , 
        \Level2Out20[0] }), .In2({\Level2Out22[31] , \Level2Out22[30] , 
        \Level2Out22[29] , \Level2Out22[28] , \Level2Out22[27] , 
        \Level2Out22[26] , \Level2Out22[25] , \Level2Out22[24] , 
        \Level2Out22[23] , \Level2Out22[22] , \Level2Out22[21] , 
        \Level2Out22[20] , \Level2Out22[19] , \Level2Out22[18] , 
        \Level2Out22[17] , \Level2Out22[16] , \Level2Out22[15] , 
        \Level2Out22[14] , \Level2Out22[13] , \Level2Out22[12] , 
        \Level2Out22[11] , \Level2Out22[10] , \Level2Out22[9] , 
        \Level2Out22[8] , \Level2Out22[7] , \Level2Out22[6] , \Level2Out22[5] , 
        \Level2Out22[4] , \Level2Out22[3] , \Level2Out22[2] , \Level2Out22[1] , 
        \Level2Out22[0] }), .Read1(\Level2Load20[0] ), .Read2(
        \Level2Load22[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_219 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink219[31] , \ScanLink219[30] , 
        \ScanLink219[29] , \ScanLink219[28] , \ScanLink219[27] , 
        \ScanLink219[26] , \ScanLink219[25] , \ScanLink219[24] , 
        \ScanLink219[23] , \ScanLink219[22] , \ScanLink219[21] , 
        \ScanLink219[20] , \ScanLink219[19] , \ScanLink219[18] , 
        \ScanLink219[17] , \ScanLink219[16] , \ScanLink219[15] , 
        \ScanLink219[14] , \ScanLink219[13] , \ScanLink219[12] , 
        \ScanLink219[11] , \ScanLink219[10] , \ScanLink219[9] , 
        \ScanLink219[8] , \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , 
        \ScanLink219[4] , \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , 
        \ScanLink219[0] }), .ScanOut({\ScanLink220[31] , \ScanLink220[30] , 
        \ScanLink220[29] , \ScanLink220[28] , \ScanLink220[27] , 
        \ScanLink220[26] , \ScanLink220[25] , \ScanLink220[24] , 
        \ScanLink220[23] , \ScanLink220[22] , \ScanLink220[21] , 
        \ScanLink220[20] , \ScanLink220[19] , \ScanLink220[18] , 
        \ScanLink220[17] , \ScanLink220[16] , \ScanLink220[15] , 
        \ScanLink220[14] , \ScanLink220[13] , \ScanLink220[12] , 
        \ScanLink220[11] , \ScanLink220[10] , \ScanLink220[9] , 
        \ScanLink220[8] , \ScanLink220[7] , \ScanLink220[6] , \ScanLink220[5] , 
        \ScanLink220[4] , \ScanLink220[3] , \ScanLink220[2] , \ScanLink220[1] , 
        \ScanLink220[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load219[0] ), .Out({\Level1Out219[31] , \Level1Out219[30] , 
        \Level1Out219[29] , \Level1Out219[28] , \Level1Out219[27] , 
        \Level1Out219[26] , \Level1Out219[25] , \Level1Out219[24] , 
        \Level1Out219[23] , \Level1Out219[22] , \Level1Out219[21] , 
        \Level1Out219[20] , \Level1Out219[19] , \Level1Out219[18] , 
        \Level1Out219[17] , \Level1Out219[16] , \Level1Out219[15] , 
        \Level1Out219[14] , \Level1Out219[13] , \Level1Out219[12] , 
        \Level1Out219[11] , \Level1Out219[10] , \Level1Out219[9] , 
        \Level1Out219[8] , \Level1Out219[7] , \Level1Out219[6] , 
        \Level1Out219[5] , \Level1Out219[4] , \Level1Out219[3] , 
        \Level1Out219[2] , \Level1Out219[1] , \Level1Out219[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_160_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load160[0] ), .Out({\Level16Out160[31] , \Level16Out160[30] , 
        \Level16Out160[29] , \Level16Out160[28] , \Level16Out160[27] , 
        \Level16Out160[26] , \Level16Out160[25] , \Level16Out160[24] , 
        \Level16Out160[23] , \Level16Out160[22] , \Level16Out160[21] , 
        \Level16Out160[20] , \Level16Out160[19] , \Level16Out160[18] , 
        \Level16Out160[17] , \Level16Out160[16] , \Level16Out160[15] , 
        \Level16Out160[14] , \Level16Out160[13] , \Level16Out160[12] , 
        \Level16Out160[11] , \Level16Out160[10] , \Level16Out160[9] , 
        \Level16Out160[8] , \Level16Out160[7] , \Level16Out160[6] , 
        \Level16Out160[5] , \Level16Out160[4] , \Level16Out160[3] , 
        \Level16Out160[2] , \Level16Out160[1] , \Level16Out160[0] }), .In1({
        \Level8Out160[31] , \Level8Out160[30] , \Level8Out160[29] , 
        \Level8Out160[28] , \Level8Out160[27] , \Level8Out160[26] , 
        \Level8Out160[25] , \Level8Out160[24] , \Level8Out160[23] , 
        \Level8Out160[22] , \Level8Out160[21] , \Level8Out160[20] , 
        \Level8Out160[19] , \Level8Out160[18] , \Level8Out160[17] , 
        \Level8Out160[16] , \Level8Out160[15] , \Level8Out160[14] , 
        \Level8Out160[13] , \Level8Out160[12] , \Level8Out160[11] , 
        \Level8Out160[10] , \Level8Out160[9] , \Level8Out160[8] , 
        \Level8Out160[7] , \Level8Out160[6] , \Level8Out160[5] , 
        \Level8Out160[4] , \Level8Out160[3] , \Level8Out160[2] , 
        \Level8Out160[1] , \Level8Out160[0] }), .In2({\Level8Out168[31] , 
        \Level8Out168[30] , \Level8Out168[29] , \Level8Out168[28] , 
        \Level8Out168[27] , \Level8Out168[26] , \Level8Out168[25] , 
        \Level8Out168[24] , \Level8Out168[23] , \Level8Out168[22] , 
        \Level8Out168[21] , \Level8Out168[20] , \Level8Out168[19] , 
        \Level8Out168[18] , \Level8Out168[17] , \Level8Out168[16] , 
        \Level8Out168[15] , \Level8Out168[14] , \Level8Out168[13] , 
        \Level8Out168[12] , \Level8Out168[11] , \Level8Out168[10] , 
        \Level8Out168[9] , \Level8Out168[8] , \Level8Out168[7] , 
        \Level8Out168[6] , \Level8Out168[5] , \Level8Out168[4] , 
        \Level8Out168[3] , \Level8Out168[2] , \Level8Out168[1] , 
        \Level8Out168[0] }), .Read1(\Level8Load160[0] ), .Read2(
        \Level8Load168[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_92 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink92[31] , \ScanLink92[30] , 
        \ScanLink92[29] , \ScanLink92[28] , \ScanLink92[27] , \ScanLink92[26] , 
        \ScanLink92[25] , \ScanLink92[24] , \ScanLink92[23] , \ScanLink92[22] , 
        \ScanLink92[21] , \ScanLink92[20] , \ScanLink92[19] , \ScanLink92[18] , 
        \ScanLink92[17] , \ScanLink92[16] , \ScanLink92[15] , \ScanLink92[14] , 
        \ScanLink92[13] , \ScanLink92[12] , \ScanLink92[11] , \ScanLink92[10] , 
        \ScanLink92[9] , \ScanLink92[8] , \ScanLink92[7] , \ScanLink92[6] , 
        \ScanLink92[5] , \ScanLink92[4] , \ScanLink92[3] , \ScanLink92[2] , 
        \ScanLink92[1] , \ScanLink92[0] }), .ScanOut({\ScanLink93[31] , 
        \ScanLink93[30] , \ScanLink93[29] , \ScanLink93[28] , \ScanLink93[27] , 
        \ScanLink93[26] , \ScanLink93[25] , \ScanLink93[24] , \ScanLink93[23] , 
        \ScanLink93[22] , \ScanLink93[21] , \ScanLink93[20] , \ScanLink93[19] , 
        \ScanLink93[18] , \ScanLink93[17] , \ScanLink93[16] , \ScanLink93[15] , 
        \ScanLink93[14] , \ScanLink93[13] , \ScanLink93[12] , \ScanLink93[11] , 
        \ScanLink93[10] , \ScanLink93[9] , \ScanLink93[8] , \ScanLink93[7] , 
        \ScanLink93[6] , \ScanLink93[5] , \ScanLink93[4] , \ScanLink93[3] , 
        \ScanLink93[2] , \ScanLink93[1] , \ScanLink93[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load92[0] ), .Out({
        \Level1Out92[31] , \Level1Out92[30] , \Level1Out92[29] , 
        \Level1Out92[28] , \Level1Out92[27] , \Level1Out92[26] , 
        \Level1Out92[25] , \Level1Out92[24] , \Level1Out92[23] , 
        \Level1Out92[22] , \Level1Out92[21] , \Level1Out92[20] , 
        \Level1Out92[19] , \Level1Out92[18] , \Level1Out92[17] , 
        \Level1Out92[16] , \Level1Out92[15] , \Level1Out92[14] , 
        \Level1Out92[13] , \Level1Out92[12] , \Level1Out92[11] , 
        \Level1Out92[10] , \Level1Out92[9] , \Level1Out92[8] , 
        \Level1Out92[7] , \Level1Out92[6] , \Level1Out92[5] , \Level1Out92[4] , 
        \Level1Out92[3] , \Level1Out92[2] , \Level1Out92[1] , \Level1Out92[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_80_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load80[0] ), .Out({\Level2Out80[31] , \Level2Out80[30] , 
        \Level2Out80[29] , \Level2Out80[28] , \Level2Out80[27] , 
        \Level2Out80[26] , \Level2Out80[25] , \Level2Out80[24] , 
        \Level2Out80[23] , \Level2Out80[22] , \Level2Out80[21] , 
        \Level2Out80[20] , \Level2Out80[19] , \Level2Out80[18] , 
        \Level2Out80[17] , \Level2Out80[16] , \Level2Out80[15] , 
        \Level2Out80[14] , \Level2Out80[13] , \Level2Out80[12] , 
        \Level2Out80[11] , \Level2Out80[10] , \Level2Out80[9] , 
        \Level2Out80[8] , \Level2Out80[7] , \Level2Out80[6] , \Level2Out80[5] , 
        \Level2Out80[4] , \Level2Out80[3] , \Level2Out80[2] , \Level2Out80[1] , 
        \Level2Out80[0] }), .In1({\Level1Out80[31] , \Level1Out80[30] , 
        \Level1Out80[29] , \Level1Out80[28] , \Level1Out80[27] , 
        \Level1Out80[26] , \Level1Out80[25] , \Level1Out80[24] , 
        \Level1Out80[23] , \Level1Out80[22] , \Level1Out80[21] , 
        \Level1Out80[20] , \Level1Out80[19] , \Level1Out80[18] , 
        \Level1Out80[17] , \Level1Out80[16] , \Level1Out80[15] , 
        \Level1Out80[14] , \Level1Out80[13] , \Level1Out80[12] , 
        \Level1Out80[11] , \Level1Out80[10] , \Level1Out80[9] , 
        \Level1Out80[8] , \Level1Out80[7] , \Level1Out80[6] , \Level1Out80[5] , 
        \Level1Out80[4] , \Level1Out80[3] , \Level1Out80[2] , \Level1Out80[1] , 
        \Level1Out80[0] }), .In2({\Level1Out81[31] , \Level1Out81[30] , 
        \Level1Out81[29] , \Level1Out81[28] , \Level1Out81[27] , 
        \Level1Out81[26] , \Level1Out81[25] , \Level1Out81[24] , 
        \Level1Out81[23] , \Level1Out81[22] , \Level1Out81[21] , 
        \Level1Out81[20] , \Level1Out81[19] , \Level1Out81[18] , 
        \Level1Out81[17] , \Level1Out81[16] , \Level1Out81[15] , 
        \Level1Out81[14] , \Level1Out81[13] , \Level1Out81[12] , 
        \Level1Out81[11] , \Level1Out81[10] , \Level1Out81[9] , 
        \Level1Out81[8] , \Level1Out81[7] , \Level1Out81[6] , \Level1Out81[5] , 
        \Level1Out81[4] , \Level1Out81[3] , \Level1Out81[2] , \Level1Out81[1] , 
        \Level1Out81[0] }), .Read1(\Level1Load80[0] ), .Read2(
        \Level1Load81[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_208_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load208[0] ), .Out({\Level16Out208[31] , \Level16Out208[30] , 
        \Level16Out208[29] , \Level16Out208[28] , \Level16Out208[27] , 
        \Level16Out208[26] , \Level16Out208[25] , \Level16Out208[24] , 
        \Level16Out208[23] , \Level16Out208[22] , \Level16Out208[21] , 
        \Level16Out208[20] , \Level16Out208[19] , \Level16Out208[18] , 
        \Level16Out208[17] , \Level16Out208[16] , \Level16Out208[15] , 
        \Level16Out208[14] , \Level16Out208[13] , \Level16Out208[12] , 
        \Level16Out208[11] , \Level16Out208[10] , \Level16Out208[9] , 
        \Level16Out208[8] , \Level16Out208[7] , \Level16Out208[6] , 
        \Level16Out208[5] , \Level16Out208[4] , \Level16Out208[3] , 
        \Level16Out208[2] , \Level16Out208[1] , \Level16Out208[0] }), .In1({
        \Level8Out208[31] , \Level8Out208[30] , \Level8Out208[29] , 
        \Level8Out208[28] , \Level8Out208[27] , \Level8Out208[26] , 
        \Level8Out208[25] , \Level8Out208[24] , \Level8Out208[23] , 
        \Level8Out208[22] , \Level8Out208[21] , \Level8Out208[20] , 
        \Level8Out208[19] , \Level8Out208[18] , \Level8Out208[17] , 
        \Level8Out208[16] , \Level8Out208[15] , \Level8Out208[14] , 
        \Level8Out208[13] , \Level8Out208[12] , \Level8Out208[11] , 
        \Level8Out208[10] , \Level8Out208[9] , \Level8Out208[8] , 
        \Level8Out208[7] , \Level8Out208[6] , \Level8Out208[5] , 
        \Level8Out208[4] , \Level8Out208[3] , \Level8Out208[2] , 
        \Level8Out208[1] , \Level8Out208[0] }), .In2({\Level8Out216[31] , 
        \Level8Out216[30] , \Level8Out216[29] , \Level8Out216[28] , 
        \Level8Out216[27] , \Level8Out216[26] , \Level8Out216[25] , 
        \Level8Out216[24] , \Level8Out216[23] , \Level8Out216[22] , 
        \Level8Out216[21] , \Level8Out216[20] , \Level8Out216[19] , 
        \Level8Out216[18] , \Level8Out216[17] , \Level8Out216[16] , 
        \Level8Out216[15] , \Level8Out216[14] , \Level8Out216[13] , 
        \Level8Out216[12] , \Level8Out216[11] , \Level8Out216[10] , 
        \Level8Out216[9] , \Level8Out216[8] , \Level8Out216[7] , 
        \Level8Out216[6] , \Level8Out216[5] , \Level8Out216[4] , 
        \Level8Out216[3] , \Level8Out216[2] , \Level8Out216[1] , 
        \Level8Out216[0] }), .Read1(\Level8Load208[0] ), .Read2(
        \Level8Load216[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_197 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink197[31] , \ScanLink197[30] , 
        \ScanLink197[29] , \ScanLink197[28] , \ScanLink197[27] , 
        \ScanLink197[26] , \ScanLink197[25] , \ScanLink197[24] , 
        \ScanLink197[23] , \ScanLink197[22] , \ScanLink197[21] , 
        \ScanLink197[20] , \ScanLink197[19] , \ScanLink197[18] , 
        \ScanLink197[17] , \ScanLink197[16] , \ScanLink197[15] , 
        \ScanLink197[14] , \ScanLink197[13] , \ScanLink197[12] , 
        \ScanLink197[11] , \ScanLink197[10] , \ScanLink197[9] , 
        \ScanLink197[8] , \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , 
        \ScanLink197[4] , \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , 
        \ScanLink197[0] }), .ScanOut({\ScanLink198[31] , \ScanLink198[30] , 
        \ScanLink198[29] , \ScanLink198[28] , \ScanLink198[27] , 
        \ScanLink198[26] , \ScanLink198[25] , \ScanLink198[24] , 
        \ScanLink198[23] , \ScanLink198[22] , \ScanLink198[21] , 
        \ScanLink198[20] , \ScanLink198[19] , \ScanLink198[18] , 
        \ScanLink198[17] , \ScanLink198[16] , \ScanLink198[15] , 
        \ScanLink198[14] , \ScanLink198[13] , \ScanLink198[12] , 
        \ScanLink198[11] , \ScanLink198[10] , \ScanLink198[9] , 
        \ScanLink198[8] , \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , 
        \ScanLink198[4] , \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , 
        \ScanLink198[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load197[0] ), .Out({\Level1Out197[31] , \Level1Out197[30] , 
        \Level1Out197[29] , \Level1Out197[28] , \Level1Out197[27] , 
        \Level1Out197[26] , \Level1Out197[25] , \Level1Out197[24] , 
        \Level1Out197[23] , \Level1Out197[22] , \Level1Out197[21] , 
        \Level1Out197[20] , \Level1Out197[19] , \Level1Out197[18] , 
        \Level1Out197[17] , \Level1Out197[16] , \Level1Out197[15] , 
        \Level1Out197[14] , \Level1Out197[13] , \Level1Out197[12] , 
        \Level1Out197[11] , \Level1Out197[10] , \Level1Out197[9] , 
        \Level1Out197[8] , \Level1Out197[7] , \Level1Out197[6] , 
        \Level1Out197[5] , \Level1Out197[4] , \Level1Out197[3] , 
        \Level1Out197[2] , \Level1Out197[1] , \Level1Out197[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load0[0] ), .Out({\Level8Out0[31] , \Level8Out0[30] , 
        \Level8Out0[29] , \Level8Out0[28] , \Level8Out0[27] , \Level8Out0[26] , 
        \Level8Out0[25] , \Level8Out0[24] , \Level8Out0[23] , \Level8Out0[22] , 
        \Level8Out0[21] , \Level8Out0[20] , \Level8Out0[19] , \Level8Out0[18] , 
        \Level8Out0[17] , \Level8Out0[16] , \Level8Out0[15] , \Level8Out0[14] , 
        \Level8Out0[13] , \Level8Out0[12] , \Level8Out0[11] , \Level8Out0[10] , 
        \Level8Out0[9] , \Level8Out0[8] , \Level8Out0[7] , \Level8Out0[6] , 
        \Level8Out0[5] , \Level8Out0[4] , \Level8Out0[3] , \Level8Out0[2] , 
        \Level8Out0[1] , \Level8Out0[0] }), .In1({\Level4Out0[31] , 
        \Level4Out0[30] , \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , 
        \Level4Out0[26] , \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , 
        \Level4Out0[22] , \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , 
        \Level4Out0[18] , \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , 
        \Level4Out0[14] , \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , 
        \Level4Out0[10] , \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , 
        \Level4Out0[6] , \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , 
        \Level4Out0[2] , \Level4Out0[1] , \Level4Out0[0] }), .In2({
        \Level4Out4[31] , \Level4Out4[30] , \Level4Out4[29] , \Level4Out4[28] , 
        \Level4Out4[27] , \Level4Out4[26] , \Level4Out4[25] , \Level4Out4[24] , 
        \Level4Out4[23] , \Level4Out4[22] , \Level4Out4[21] , \Level4Out4[20] , 
        \Level4Out4[19] , \Level4Out4[18] , \Level4Out4[17] , \Level4Out4[16] , 
        \Level4Out4[15] , \Level4Out4[14] , \Level4Out4[13] , \Level4Out4[12] , 
        \Level4Out4[11] , \Level4Out4[10] , \Level4Out4[9] , \Level4Out4[8] , 
        \Level4Out4[7] , \Level4Out4[6] , \Level4Out4[5] , \Level4Out4[4] , 
        \Level4Out4[3] , \Level4Out4[2] , \Level4Out4[1] , \Level4Out4[0] }), 
        .Read1(\Level4Load0[0] ), .Read2(\Level4Load4[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_50 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanOut({\ScanLink51[31] , 
        \ScanLink51[30] , \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , 
        \ScanLink51[26] , \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , 
        \ScanLink51[22] , \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , 
        \ScanLink51[18] , \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , 
        \ScanLink51[14] , \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , 
        \ScanLink51[10] , \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , 
        \ScanLink51[6] , \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , 
        \ScanLink51[2] , \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load50[0] ), .Out({
        \Level1Out50[31] , \Level1Out50[30] , \Level1Out50[29] , 
        \Level1Out50[28] , \Level1Out50[27] , \Level1Out50[26] , 
        \Level1Out50[25] , \Level1Out50[24] , \Level1Out50[23] , 
        \Level1Out50[22] , \Level1Out50[21] , \Level1Out50[20] , 
        \Level1Out50[19] , \Level1Out50[18] , \Level1Out50[17] , 
        \Level1Out50[16] , \Level1Out50[15] , \Level1Out50[14] , 
        \Level1Out50[13] , \Level1Out50[12] , \Level1Out50[11] , 
        \Level1Out50[10] , \Level1Out50[9] , \Level1Out50[8] , 
        \Level1Out50[7] , \Level1Out50[6] , \Level1Out50[5] , \Level1Out50[4] , 
        \Level1Out50[3] , \Level1Out50[2] , \Level1Out50[1] , \Level1Out50[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_77 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink77[31] , \ScanLink77[30] , 
        \ScanLink77[29] , \ScanLink77[28] , \ScanLink77[27] , \ScanLink77[26] , 
        \ScanLink77[25] , \ScanLink77[24] , \ScanLink77[23] , \ScanLink77[22] , 
        \ScanLink77[21] , \ScanLink77[20] , \ScanLink77[19] , \ScanLink77[18] , 
        \ScanLink77[17] , \ScanLink77[16] , \ScanLink77[15] , \ScanLink77[14] , 
        \ScanLink77[13] , \ScanLink77[12] , \ScanLink77[11] , \ScanLink77[10] , 
        \ScanLink77[9] , \ScanLink77[8] , \ScanLink77[7] , \ScanLink77[6] , 
        \ScanLink77[5] , \ScanLink77[4] , \ScanLink77[3] , \ScanLink77[2] , 
        \ScanLink77[1] , \ScanLink77[0] }), .ScanOut({\ScanLink78[31] , 
        \ScanLink78[30] , \ScanLink78[29] , \ScanLink78[28] , \ScanLink78[27] , 
        \ScanLink78[26] , \ScanLink78[25] , \ScanLink78[24] , \ScanLink78[23] , 
        \ScanLink78[22] , \ScanLink78[21] , \ScanLink78[20] , \ScanLink78[19] , 
        \ScanLink78[18] , \ScanLink78[17] , \ScanLink78[16] , \ScanLink78[15] , 
        \ScanLink78[14] , \ScanLink78[13] , \ScanLink78[12] , \ScanLink78[11] , 
        \ScanLink78[10] , \ScanLink78[9] , \ScanLink78[8] , \ScanLink78[7] , 
        \ScanLink78[6] , \ScanLink78[5] , \ScanLink78[4] , \ScanLink78[3] , 
        \ScanLink78[2] , \ScanLink78[1] , \ScanLink78[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load77[0] ), .Out({
        \Level1Out77[31] , \Level1Out77[30] , \Level1Out77[29] , 
        \Level1Out77[28] , \Level1Out77[27] , \Level1Out77[26] , 
        \Level1Out77[25] , \Level1Out77[24] , \Level1Out77[23] , 
        \Level1Out77[22] , \Level1Out77[21] , \Level1Out77[20] , 
        \Level1Out77[19] , \Level1Out77[18] , \Level1Out77[17] , 
        \Level1Out77[16] , \Level1Out77[15] , \Level1Out77[14] , 
        \Level1Out77[13] , \Level1Out77[12] , \Level1Out77[11] , 
        \Level1Out77[10] , \Level1Out77[9] , \Level1Out77[8] , 
        \Level1Out77[7] , \Level1Out77[6] , \Level1Out77[5] , \Level1Out77[4] , 
        \Level1Out77[3] , \Level1Out77[2] , \Level1Out77[1] , \Level1Out77[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_72_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load72[0] ), .Out({\Level8Out72[31] , \Level8Out72[30] , 
        \Level8Out72[29] , \Level8Out72[28] , \Level8Out72[27] , 
        \Level8Out72[26] , \Level8Out72[25] , \Level8Out72[24] , 
        \Level8Out72[23] , \Level8Out72[22] , \Level8Out72[21] , 
        \Level8Out72[20] , \Level8Out72[19] , \Level8Out72[18] , 
        \Level8Out72[17] , \Level8Out72[16] , \Level8Out72[15] , 
        \Level8Out72[14] , \Level8Out72[13] , \Level8Out72[12] , 
        \Level8Out72[11] , \Level8Out72[10] , \Level8Out72[9] , 
        \Level8Out72[8] , \Level8Out72[7] , \Level8Out72[6] , \Level8Out72[5] , 
        \Level8Out72[4] , \Level8Out72[3] , \Level8Out72[2] , \Level8Out72[1] , 
        \Level8Out72[0] }), .In1({\Level4Out72[31] , \Level4Out72[30] , 
        \Level4Out72[29] , \Level4Out72[28] , \Level4Out72[27] , 
        \Level4Out72[26] , \Level4Out72[25] , \Level4Out72[24] , 
        \Level4Out72[23] , \Level4Out72[22] , \Level4Out72[21] , 
        \Level4Out72[20] , \Level4Out72[19] , \Level4Out72[18] , 
        \Level4Out72[17] , \Level4Out72[16] , \Level4Out72[15] , 
        \Level4Out72[14] , \Level4Out72[13] , \Level4Out72[12] , 
        \Level4Out72[11] , \Level4Out72[10] , \Level4Out72[9] , 
        \Level4Out72[8] , \Level4Out72[7] , \Level4Out72[6] , \Level4Out72[5] , 
        \Level4Out72[4] , \Level4Out72[3] , \Level4Out72[2] , \Level4Out72[1] , 
        \Level4Out72[0] }), .In2({\Level4Out76[31] , \Level4Out76[30] , 
        \Level4Out76[29] , \Level4Out76[28] , \Level4Out76[27] , 
        \Level4Out76[26] , \Level4Out76[25] , \Level4Out76[24] , 
        \Level4Out76[23] , \Level4Out76[22] , \Level4Out76[21] , 
        \Level4Out76[20] , \Level4Out76[19] , \Level4Out76[18] , 
        \Level4Out76[17] , \Level4Out76[16] , \Level4Out76[15] , 
        \Level4Out76[14] , \Level4Out76[13] , \Level4Out76[12] , 
        \Level4Out76[11] , \Level4Out76[10] , \Level4Out76[9] , 
        \Level4Out76[8] , \Level4Out76[7] , \Level4Out76[6] , \Level4Out76[5] , 
        \Level4Out76[4] , \Level4Out76[3] , \Level4Out76[2] , \Level4Out76[1] , 
        \Level4Out76[0] }), .Read1(\Level4Load72[0] ), .Read2(
        \Level4Load76[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_196_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load196[0] ), .Out({\Level2Out196[31] , \Level2Out196[30] , 
        \Level2Out196[29] , \Level2Out196[28] , \Level2Out196[27] , 
        \Level2Out196[26] , \Level2Out196[25] , \Level2Out196[24] , 
        \Level2Out196[23] , \Level2Out196[22] , \Level2Out196[21] , 
        \Level2Out196[20] , \Level2Out196[19] , \Level2Out196[18] , 
        \Level2Out196[17] , \Level2Out196[16] , \Level2Out196[15] , 
        \Level2Out196[14] , \Level2Out196[13] , \Level2Out196[12] , 
        \Level2Out196[11] , \Level2Out196[10] , \Level2Out196[9] , 
        \Level2Out196[8] , \Level2Out196[7] , \Level2Out196[6] , 
        \Level2Out196[5] , \Level2Out196[4] , \Level2Out196[3] , 
        \Level2Out196[2] , \Level2Out196[1] , \Level2Out196[0] }), .In1({
        \Level1Out196[31] , \Level1Out196[30] , \Level1Out196[29] , 
        \Level1Out196[28] , \Level1Out196[27] , \Level1Out196[26] , 
        \Level1Out196[25] , \Level1Out196[24] , \Level1Out196[23] , 
        \Level1Out196[22] , \Level1Out196[21] , \Level1Out196[20] , 
        \Level1Out196[19] , \Level1Out196[18] , \Level1Out196[17] , 
        \Level1Out196[16] , \Level1Out196[15] , \Level1Out196[14] , 
        \Level1Out196[13] , \Level1Out196[12] , \Level1Out196[11] , 
        \Level1Out196[10] , \Level1Out196[9] , \Level1Out196[8] , 
        \Level1Out196[7] , \Level1Out196[6] , \Level1Out196[5] , 
        \Level1Out196[4] , \Level1Out196[3] , \Level1Out196[2] , 
        \Level1Out196[1] , \Level1Out196[0] }), .In2({\Level1Out197[31] , 
        \Level1Out197[30] , \Level1Out197[29] , \Level1Out197[28] , 
        \Level1Out197[27] , \Level1Out197[26] , \Level1Out197[25] , 
        \Level1Out197[24] , \Level1Out197[23] , \Level1Out197[22] , 
        \Level1Out197[21] , \Level1Out197[20] , \Level1Out197[19] , 
        \Level1Out197[18] , \Level1Out197[17] , \Level1Out197[16] , 
        \Level1Out197[15] , \Level1Out197[14] , \Level1Out197[13] , 
        \Level1Out197[12] , \Level1Out197[11] , \Level1Out197[10] , 
        \Level1Out197[9] , \Level1Out197[8] , \Level1Out197[7] , 
        \Level1Out197[6] , \Level1Out197[5] , \Level1Out197[4] , 
        \Level1Out197[3] , \Level1Out197[2] , \Level1Out197[1] , 
        \Level1Out197[0] }), .Read1(\Level1Load196[0] ), .Read2(
        \Level1Load197[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_200_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load200[0] ), .Out({\Level8Out200[31] , \Level8Out200[30] , 
        \Level8Out200[29] , \Level8Out200[28] , \Level8Out200[27] , 
        \Level8Out200[26] , \Level8Out200[25] , \Level8Out200[24] , 
        \Level8Out200[23] , \Level8Out200[22] , \Level8Out200[21] , 
        \Level8Out200[20] , \Level8Out200[19] , \Level8Out200[18] , 
        \Level8Out200[17] , \Level8Out200[16] , \Level8Out200[15] , 
        \Level8Out200[14] , \Level8Out200[13] , \Level8Out200[12] , 
        \Level8Out200[11] , \Level8Out200[10] , \Level8Out200[9] , 
        \Level8Out200[8] , \Level8Out200[7] , \Level8Out200[6] , 
        \Level8Out200[5] , \Level8Out200[4] , \Level8Out200[3] , 
        \Level8Out200[2] , \Level8Out200[1] , \Level8Out200[0] }), .In1({
        \Level4Out200[31] , \Level4Out200[30] , \Level4Out200[29] , 
        \Level4Out200[28] , \Level4Out200[27] , \Level4Out200[26] , 
        \Level4Out200[25] , \Level4Out200[24] , \Level4Out200[23] , 
        \Level4Out200[22] , \Level4Out200[21] , \Level4Out200[20] , 
        \Level4Out200[19] , \Level4Out200[18] , \Level4Out200[17] , 
        \Level4Out200[16] , \Level4Out200[15] , \Level4Out200[14] , 
        \Level4Out200[13] , \Level4Out200[12] , \Level4Out200[11] , 
        \Level4Out200[10] , \Level4Out200[9] , \Level4Out200[8] , 
        \Level4Out200[7] , \Level4Out200[6] , \Level4Out200[5] , 
        \Level4Out200[4] , \Level4Out200[3] , \Level4Out200[2] , 
        \Level4Out200[1] , \Level4Out200[0] }), .In2({\Level4Out204[31] , 
        \Level4Out204[30] , \Level4Out204[29] , \Level4Out204[28] , 
        \Level4Out204[27] , \Level4Out204[26] , \Level4Out204[25] , 
        \Level4Out204[24] , \Level4Out204[23] , \Level4Out204[22] , 
        \Level4Out204[21] , \Level4Out204[20] , \Level4Out204[19] , 
        \Level4Out204[18] , \Level4Out204[17] , \Level4Out204[16] , 
        \Level4Out204[15] , \Level4Out204[14] , \Level4Out204[13] , 
        \Level4Out204[12] , \Level4Out204[11] , \Level4Out204[10] , 
        \Level4Out204[9] , \Level4Out204[8] , \Level4Out204[7] , 
        \Level4Out204[6] , \Level4Out204[5] , \Level4Out204[4] , 
        \Level4Out204[3] , \Level4Out204[2] , \Level4Out204[1] , 
        \Level4Out204[0] }), .Read1(\Level4Load200[0] ), .Read2(
        \Level4Load204[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_155 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink155[31] , \ScanLink155[30] , 
        \ScanLink155[29] , \ScanLink155[28] , \ScanLink155[27] , 
        \ScanLink155[26] , \ScanLink155[25] , \ScanLink155[24] , 
        \ScanLink155[23] , \ScanLink155[22] , \ScanLink155[21] , 
        \ScanLink155[20] , \ScanLink155[19] , \ScanLink155[18] , 
        \ScanLink155[17] , \ScanLink155[16] , \ScanLink155[15] , 
        \ScanLink155[14] , \ScanLink155[13] , \ScanLink155[12] , 
        \ScanLink155[11] , \ScanLink155[10] , \ScanLink155[9] , 
        \ScanLink155[8] , \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , 
        \ScanLink155[4] , \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , 
        \ScanLink155[0] }), .ScanOut({\ScanLink156[31] , \ScanLink156[30] , 
        \ScanLink156[29] , \ScanLink156[28] , \ScanLink156[27] , 
        \ScanLink156[26] , \ScanLink156[25] , \ScanLink156[24] , 
        \ScanLink156[23] , \ScanLink156[22] , \ScanLink156[21] , 
        \ScanLink156[20] , \ScanLink156[19] , \ScanLink156[18] , 
        \ScanLink156[17] , \ScanLink156[16] , \ScanLink156[15] , 
        \ScanLink156[14] , \ScanLink156[13] , \ScanLink156[12] , 
        \ScanLink156[11] , \ScanLink156[10] , \ScanLink156[9] , 
        \ScanLink156[8] , \ScanLink156[7] , \ScanLink156[6] , \ScanLink156[5] , 
        \ScanLink156[4] , \ScanLink156[3] , \ScanLink156[2] , \ScanLink156[1] , 
        \ScanLink156[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load155[0] ), .Out({\Level1Out155[31] , \Level1Out155[30] , 
        \Level1Out155[29] , \Level1Out155[28] , \Level1Out155[27] , 
        \Level1Out155[26] , \Level1Out155[25] , \Level1Out155[24] , 
        \Level1Out155[23] , \Level1Out155[22] , \Level1Out155[21] , 
        \Level1Out155[20] , \Level1Out155[19] , \Level1Out155[18] , 
        \Level1Out155[17] , \Level1Out155[16] , \Level1Out155[15] , 
        \Level1Out155[14] , \Level1Out155[13] , \Level1Out155[12] , 
        \Level1Out155[11] , \Level1Out155[10] , \Level1Out155[9] , 
        \Level1Out155[8] , \Level1Out155[7] , \Level1Out155[6] , 
        \Level1Out155[5] , \Level1Out155[4] , \Level1Out155[3] , 
        \Level1Out155[2] , \Level1Out155[1] , \Level1Out155[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_172 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink172[31] , \ScanLink172[30] , 
        \ScanLink172[29] , \ScanLink172[28] , \ScanLink172[27] , 
        \ScanLink172[26] , \ScanLink172[25] , \ScanLink172[24] , 
        \ScanLink172[23] , \ScanLink172[22] , \ScanLink172[21] , 
        \ScanLink172[20] , \ScanLink172[19] , \ScanLink172[18] , 
        \ScanLink172[17] , \ScanLink172[16] , \ScanLink172[15] , 
        \ScanLink172[14] , \ScanLink172[13] , \ScanLink172[12] , 
        \ScanLink172[11] , \ScanLink172[10] , \ScanLink172[9] , 
        \ScanLink172[8] , \ScanLink172[7] , \ScanLink172[6] , \ScanLink172[5] , 
        \ScanLink172[4] , \ScanLink172[3] , \ScanLink172[2] , \ScanLink172[1] , 
        \ScanLink172[0] }), .ScanOut({\ScanLink173[31] , \ScanLink173[30] , 
        \ScanLink173[29] , \ScanLink173[28] , \ScanLink173[27] , 
        \ScanLink173[26] , \ScanLink173[25] , \ScanLink173[24] , 
        \ScanLink173[23] , \ScanLink173[22] , \ScanLink173[21] , 
        \ScanLink173[20] , \ScanLink173[19] , \ScanLink173[18] , 
        \ScanLink173[17] , \ScanLink173[16] , \ScanLink173[15] , 
        \ScanLink173[14] , \ScanLink173[13] , \ScanLink173[12] , 
        \ScanLink173[11] , \ScanLink173[10] , \ScanLink173[9] , 
        \ScanLink173[8] , \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , 
        \ScanLink173[4] , \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , 
        \ScanLink173[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load172[0] ), .Out({\Level1Out172[31] , \Level1Out172[30] , 
        \Level1Out172[29] , \Level1Out172[28] , \Level1Out172[27] , 
        \Level1Out172[26] , \Level1Out172[25] , \Level1Out172[24] , 
        \Level1Out172[23] , \Level1Out172[22] , \Level1Out172[21] , 
        \Level1Out172[20] , \Level1Out172[19] , \Level1Out172[18] , 
        \Level1Out172[17] , \Level1Out172[16] , \Level1Out172[15] , 
        \Level1Out172[14] , \Level1Out172[13] , \Level1Out172[12] , 
        \Level1Out172[11] , \Level1Out172[10] , \Level1Out172[9] , 
        \Level1Out172[8] , \Level1Out172[7] , \Level1Out172[6] , 
        \Level1Out172[5] , \Level1Out172[4] , \Level1Out172[3] , 
        \Level1Out172[2] , \Level1Out172[1] , \Level1Out172[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_242 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink242[31] , \ScanLink242[30] , 
        \ScanLink242[29] , \ScanLink242[28] , \ScanLink242[27] , 
        \ScanLink242[26] , \ScanLink242[25] , \ScanLink242[24] , 
        \ScanLink242[23] , \ScanLink242[22] , \ScanLink242[21] , 
        \ScanLink242[20] , \ScanLink242[19] , \ScanLink242[18] , 
        \ScanLink242[17] , \ScanLink242[16] , \ScanLink242[15] , 
        \ScanLink242[14] , \ScanLink242[13] , \ScanLink242[12] , 
        \ScanLink242[11] , \ScanLink242[10] , \ScanLink242[9] , 
        \ScanLink242[8] , \ScanLink242[7] , \ScanLink242[6] , \ScanLink242[5] , 
        \ScanLink242[4] , \ScanLink242[3] , \ScanLink242[2] , \ScanLink242[1] , 
        \ScanLink242[0] }), .ScanOut({\ScanLink243[31] , \ScanLink243[30] , 
        \ScanLink243[29] , \ScanLink243[28] , \ScanLink243[27] , 
        \ScanLink243[26] , \ScanLink243[25] , \ScanLink243[24] , 
        \ScanLink243[23] , \ScanLink243[22] , \ScanLink243[21] , 
        \ScanLink243[20] , \ScanLink243[19] , \ScanLink243[18] , 
        \ScanLink243[17] , \ScanLink243[16] , \ScanLink243[15] , 
        \ScanLink243[14] , \ScanLink243[13] , \ScanLink243[12] , 
        \ScanLink243[11] , \ScanLink243[10] , \ScanLink243[9] , 
        \ScanLink243[8] , \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , 
        \ScanLink243[4] , \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , 
        \ScanLink243[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load242[0] ), .Out({\Level1Out242[31] , \Level1Out242[30] , 
        \Level1Out242[29] , \Level1Out242[28] , \Level1Out242[27] , 
        \Level1Out242[26] , \Level1Out242[25] , \Level1Out242[24] , 
        \Level1Out242[23] , \Level1Out242[22] , \Level1Out242[21] , 
        \Level1Out242[20] , \Level1Out242[19] , \Level1Out242[18] , 
        \Level1Out242[17] , \Level1Out242[16] , \Level1Out242[15] , 
        \Level1Out242[14] , \Level1Out242[13] , \Level1Out242[12] , 
        \Level1Out242[11] , \Level1Out242[10] , \Level1Out242[9] , 
        \Level1Out242[8] , \Level1Out242[7] , \Level1Out242[6] , 
        \Level1Out242[5] , \Level1Out242[4] , \Level1Out242[3] , 
        \Level1Out242[2] , \Level1Out242[1] , \Level1Out242[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_46_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load46[0] ), .Out({\Level2Out46[31] , \Level2Out46[30] , 
        \Level2Out46[29] , \Level2Out46[28] , \Level2Out46[27] , 
        \Level2Out46[26] , \Level2Out46[25] , \Level2Out46[24] , 
        \Level2Out46[23] , \Level2Out46[22] , \Level2Out46[21] , 
        \Level2Out46[20] , \Level2Out46[19] , \Level2Out46[18] , 
        \Level2Out46[17] , \Level2Out46[16] , \Level2Out46[15] , 
        \Level2Out46[14] , \Level2Out46[13] , \Level2Out46[12] , 
        \Level2Out46[11] , \Level2Out46[10] , \Level2Out46[9] , 
        \Level2Out46[8] , \Level2Out46[7] , \Level2Out46[6] , \Level2Out46[5] , 
        \Level2Out46[4] , \Level2Out46[3] , \Level2Out46[2] , \Level2Out46[1] , 
        \Level2Out46[0] }), .In1({\Level1Out46[31] , \Level1Out46[30] , 
        \Level1Out46[29] , \Level1Out46[28] , \Level1Out46[27] , 
        \Level1Out46[26] , \Level1Out46[25] , \Level1Out46[24] , 
        \Level1Out46[23] , \Level1Out46[22] , \Level1Out46[21] , 
        \Level1Out46[20] , \Level1Out46[19] , \Level1Out46[18] , 
        \Level1Out46[17] , \Level1Out46[16] , \Level1Out46[15] , 
        \Level1Out46[14] , \Level1Out46[13] , \Level1Out46[12] , 
        \Level1Out46[11] , \Level1Out46[10] , \Level1Out46[9] , 
        \Level1Out46[8] , \Level1Out46[7] , \Level1Out46[6] , \Level1Out46[5] , 
        \Level1Out46[4] , \Level1Out46[3] , \Level1Out46[2] , \Level1Out46[1] , 
        \Level1Out46[0] }), .In2({\Level1Out47[31] , \Level1Out47[30] , 
        \Level1Out47[29] , \Level1Out47[28] , \Level1Out47[27] , 
        \Level1Out47[26] , \Level1Out47[25] , \Level1Out47[24] , 
        \Level1Out47[23] , \Level1Out47[22] , \Level1Out47[21] , 
        \Level1Out47[20] , \Level1Out47[19] , \Level1Out47[18] , 
        \Level1Out47[17] , \Level1Out47[16] , \Level1Out47[15] , 
        \Level1Out47[14] , \Level1Out47[13] , \Level1Out47[12] , 
        \Level1Out47[11] , \Level1Out47[10] , \Level1Out47[9] , 
        \Level1Out47[8] , \Level1Out47[7] , \Level1Out47[6] , \Level1Out47[5] , 
        \Level1Out47[4] , \Level1Out47[3] , \Level1Out47[2] , \Level1Out47[1] , 
        \Level1Out47[0] }), .Read1(\Level1Load46[0] ), .Read2(
        \Level1Load47[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_234_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load234[0] ), .Out({\Level2Out234[31] , \Level2Out234[30] , 
        \Level2Out234[29] , \Level2Out234[28] , \Level2Out234[27] , 
        \Level2Out234[26] , \Level2Out234[25] , \Level2Out234[24] , 
        \Level2Out234[23] , \Level2Out234[22] , \Level2Out234[21] , 
        \Level2Out234[20] , \Level2Out234[19] , \Level2Out234[18] , 
        \Level2Out234[17] , \Level2Out234[16] , \Level2Out234[15] , 
        \Level2Out234[14] , \Level2Out234[13] , \Level2Out234[12] , 
        \Level2Out234[11] , \Level2Out234[10] , \Level2Out234[9] , 
        \Level2Out234[8] , \Level2Out234[7] , \Level2Out234[6] , 
        \Level2Out234[5] , \Level2Out234[4] , \Level2Out234[3] , 
        \Level2Out234[2] , \Level2Out234[1] , \Level2Out234[0] }), .In1({
        \Level1Out234[31] , \Level1Out234[30] , \Level1Out234[29] , 
        \Level1Out234[28] , \Level1Out234[27] , \Level1Out234[26] , 
        \Level1Out234[25] , \Level1Out234[24] , \Level1Out234[23] , 
        \Level1Out234[22] , \Level1Out234[21] , \Level1Out234[20] , 
        \Level1Out234[19] , \Level1Out234[18] , \Level1Out234[17] , 
        \Level1Out234[16] , \Level1Out234[15] , \Level1Out234[14] , 
        \Level1Out234[13] , \Level1Out234[12] , \Level1Out234[11] , 
        \Level1Out234[10] , \Level1Out234[9] , \Level1Out234[8] , 
        \Level1Out234[7] , \Level1Out234[6] , \Level1Out234[5] , 
        \Level1Out234[4] , \Level1Out234[3] , \Level1Out234[2] , 
        \Level1Out234[1] , \Level1Out234[0] }), .In2({\Level1Out235[31] , 
        \Level1Out235[30] , \Level1Out235[29] , \Level1Out235[28] , 
        \Level1Out235[27] , \Level1Out235[26] , \Level1Out235[25] , 
        \Level1Out235[24] , \Level1Out235[23] , \Level1Out235[22] , 
        \Level1Out235[21] , \Level1Out235[20] , \Level1Out235[19] , 
        \Level1Out235[18] , \Level1Out235[17] , \Level1Out235[16] , 
        \Level1Out235[15] , \Level1Out235[14] , \Level1Out235[13] , 
        \Level1Out235[12] , \Level1Out235[11] , \Level1Out235[10] , 
        \Level1Out235[9] , \Level1Out235[8] , \Level1Out235[7] , 
        \Level1Out235[6] , \Level1Out235[5] , \Level1Out235[4] , 
        \Level1Out235[3] , \Level1Out235[2] , \Level1Out235[1] , 
        \Level1Out235[0] }), .Read1(\Level1Load234[0] ), .Read2(
        \Level1Load235[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_136_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load136[0] ), .Out({\Level4Out136[31] , \Level4Out136[30] , 
        \Level4Out136[29] , \Level4Out136[28] , \Level4Out136[27] , 
        \Level4Out136[26] , \Level4Out136[25] , \Level4Out136[24] , 
        \Level4Out136[23] , \Level4Out136[22] , \Level4Out136[21] , 
        \Level4Out136[20] , \Level4Out136[19] , \Level4Out136[18] , 
        \Level4Out136[17] , \Level4Out136[16] , \Level4Out136[15] , 
        \Level4Out136[14] , \Level4Out136[13] , \Level4Out136[12] , 
        \Level4Out136[11] , \Level4Out136[10] , \Level4Out136[9] , 
        \Level4Out136[8] , \Level4Out136[7] , \Level4Out136[6] , 
        \Level4Out136[5] , \Level4Out136[4] , \Level4Out136[3] , 
        \Level4Out136[2] , \Level4Out136[1] , \Level4Out136[0] }), .In1({
        \Level2Out136[31] , \Level2Out136[30] , \Level2Out136[29] , 
        \Level2Out136[28] , \Level2Out136[27] , \Level2Out136[26] , 
        \Level2Out136[25] , \Level2Out136[24] , \Level2Out136[23] , 
        \Level2Out136[22] , \Level2Out136[21] , \Level2Out136[20] , 
        \Level2Out136[19] , \Level2Out136[18] , \Level2Out136[17] , 
        \Level2Out136[16] , \Level2Out136[15] , \Level2Out136[14] , 
        \Level2Out136[13] , \Level2Out136[12] , \Level2Out136[11] , 
        \Level2Out136[10] , \Level2Out136[9] , \Level2Out136[8] , 
        \Level2Out136[7] , \Level2Out136[6] , \Level2Out136[5] , 
        \Level2Out136[4] , \Level2Out136[3] , \Level2Out136[2] , 
        \Level2Out136[1] , \Level2Out136[0] }), .In2({\Level2Out138[31] , 
        \Level2Out138[30] , \Level2Out138[29] , \Level2Out138[28] , 
        \Level2Out138[27] , \Level2Out138[26] , \Level2Out138[25] , 
        \Level2Out138[24] , \Level2Out138[23] , \Level2Out138[22] , 
        \Level2Out138[21] , \Level2Out138[20] , \Level2Out138[19] , 
        \Level2Out138[18] , \Level2Out138[17] , \Level2Out138[16] , 
        \Level2Out138[15] , \Level2Out138[14] , \Level2Out138[13] , 
        \Level2Out138[12] , \Level2Out138[11] , \Level2Out138[10] , 
        \Level2Out138[9] , \Level2Out138[8] , \Level2Out138[7] , 
        \Level2Out138[6] , \Level2Out138[5] , \Level2Out138[4] , 
        \Level2Out138[3] , \Level2Out138[2] , \Level2Out138[1] , 
        \Level2Out138[0] }), .Read1(\Level2Load136[0] ), .Read2(
        \Level2Load138[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_228_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load228[0] ), .Out({\Level4Out228[31] , \Level4Out228[30] , 
        \Level4Out228[29] , \Level4Out228[28] , \Level4Out228[27] , 
        \Level4Out228[26] , \Level4Out228[25] , \Level4Out228[24] , 
        \Level4Out228[23] , \Level4Out228[22] , \Level4Out228[21] , 
        \Level4Out228[20] , \Level4Out228[19] , \Level4Out228[18] , 
        \Level4Out228[17] , \Level4Out228[16] , \Level4Out228[15] , 
        \Level4Out228[14] , \Level4Out228[13] , \Level4Out228[12] , 
        \Level4Out228[11] , \Level4Out228[10] , \Level4Out228[9] , 
        \Level4Out228[8] , \Level4Out228[7] , \Level4Out228[6] , 
        \Level4Out228[5] , \Level4Out228[4] , \Level4Out228[3] , 
        \Level4Out228[2] , \Level4Out228[1] , \Level4Out228[0] }), .In1({
        \Level2Out228[31] , \Level2Out228[30] , \Level2Out228[29] , 
        \Level2Out228[28] , \Level2Out228[27] , \Level2Out228[26] , 
        \Level2Out228[25] , \Level2Out228[24] , \Level2Out228[23] , 
        \Level2Out228[22] , \Level2Out228[21] , \Level2Out228[20] , 
        \Level2Out228[19] , \Level2Out228[18] , \Level2Out228[17] , 
        \Level2Out228[16] , \Level2Out228[15] , \Level2Out228[14] , 
        \Level2Out228[13] , \Level2Out228[12] , \Level2Out228[11] , 
        \Level2Out228[10] , \Level2Out228[9] , \Level2Out228[8] , 
        \Level2Out228[7] , \Level2Out228[6] , \Level2Out228[5] , 
        \Level2Out228[4] , \Level2Out228[3] , \Level2Out228[2] , 
        \Level2Out228[1] , \Level2Out228[0] }), .In2({\Level2Out230[31] , 
        \Level2Out230[30] , \Level2Out230[29] , \Level2Out230[28] , 
        \Level2Out230[27] , \Level2Out230[26] , \Level2Out230[25] , 
        \Level2Out230[24] , \Level2Out230[23] , \Level2Out230[22] , 
        \Level2Out230[21] , \Level2Out230[20] , \Level2Out230[19] , 
        \Level2Out230[18] , \Level2Out230[17] , \Level2Out230[16] , 
        \Level2Out230[15] , \Level2Out230[14] , \Level2Out230[13] , 
        \Level2Out230[12] , \Level2Out230[11] , \Level2Out230[10] , 
        \Level2Out230[9] , \Level2Out230[8] , \Level2Out230[7] , 
        \Level2Out230[6] , \Level2Out230[5] , \Level2Out230[4] , 
        \Level2Out230[3] , \Level2Out230[2] , \Level2Out230[1] , 
        \Level2Out230[0] }), .Read1(\Level2Load228[0] ), .Read2(
        \Level2Load230[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_100_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load100[0] ), .Out({\Level2Out100[31] , \Level2Out100[30] , 
        \Level2Out100[29] , \Level2Out100[28] , \Level2Out100[27] , 
        \Level2Out100[26] , \Level2Out100[25] , \Level2Out100[24] , 
        \Level2Out100[23] , \Level2Out100[22] , \Level2Out100[21] , 
        \Level2Out100[20] , \Level2Out100[19] , \Level2Out100[18] , 
        \Level2Out100[17] , \Level2Out100[16] , \Level2Out100[15] , 
        \Level2Out100[14] , \Level2Out100[13] , \Level2Out100[12] , 
        \Level2Out100[11] , \Level2Out100[10] , \Level2Out100[9] , 
        \Level2Out100[8] , \Level2Out100[7] , \Level2Out100[6] , 
        \Level2Out100[5] , \Level2Out100[4] , \Level2Out100[3] , 
        \Level2Out100[2] , \Level2Out100[1] , \Level2Out100[0] }), .In1({
        \Level1Out100[31] , \Level1Out100[30] , \Level1Out100[29] , 
        \Level1Out100[28] , \Level1Out100[27] , \Level1Out100[26] , 
        \Level1Out100[25] , \Level1Out100[24] , \Level1Out100[23] , 
        \Level1Out100[22] , \Level1Out100[21] , \Level1Out100[20] , 
        \Level1Out100[19] , \Level1Out100[18] , \Level1Out100[17] , 
        \Level1Out100[16] , \Level1Out100[15] , \Level1Out100[14] , 
        \Level1Out100[13] , \Level1Out100[12] , \Level1Out100[11] , 
        \Level1Out100[10] , \Level1Out100[9] , \Level1Out100[8] , 
        \Level1Out100[7] , \Level1Out100[6] , \Level1Out100[5] , 
        \Level1Out100[4] , \Level1Out100[3] , \Level1Out100[2] , 
        \Level1Out100[1] , \Level1Out100[0] }), .In2({\Level1Out101[31] , 
        \Level1Out101[30] , \Level1Out101[29] , \Level1Out101[28] , 
        \Level1Out101[27] , \Level1Out101[26] , \Level1Out101[25] , 
        \Level1Out101[24] , \Level1Out101[23] , \Level1Out101[22] , 
        \Level1Out101[21] , \Level1Out101[20] , \Level1Out101[19] , 
        \Level1Out101[18] , \Level1Out101[17] , \Level1Out101[16] , 
        \Level1Out101[15] , \Level1Out101[14] , \Level1Out101[13] , 
        \Level1Out101[12] , \Level1Out101[11] , \Level1Out101[10] , 
        \Level1Out101[9] , \Level1Out101[8] , \Level1Out101[7] , 
        \Level1Out101[6] , \Level1Out101[5] , \Level1Out101[4] , 
        \Level1Out101[3] , \Level1Out101[2] , \Level1Out101[1] , 
        \Level1Out101[0] }), .Read1(\Level1Load100[0] ), .Read2(
        \Level1Load101[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load192[0] ), .Out({\Level4Out192[31] , \Level4Out192[30] , 
        \Level4Out192[29] , \Level4Out192[28] , \Level4Out192[27] , 
        \Level4Out192[26] , \Level4Out192[25] , \Level4Out192[24] , 
        \Level4Out192[23] , \Level4Out192[22] , \Level4Out192[21] , 
        \Level4Out192[20] , \Level4Out192[19] , \Level4Out192[18] , 
        \Level4Out192[17] , \Level4Out192[16] , \Level4Out192[15] , 
        \Level4Out192[14] , \Level4Out192[13] , \Level4Out192[12] , 
        \Level4Out192[11] , \Level4Out192[10] , \Level4Out192[9] , 
        \Level4Out192[8] , \Level4Out192[7] , \Level4Out192[6] , 
        \Level4Out192[5] , \Level4Out192[4] , \Level4Out192[3] , 
        \Level4Out192[2] , \Level4Out192[1] , \Level4Out192[0] }), .In1({
        \Level2Out192[31] , \Level2Out192[30] , \Level2Out192[29] , 
        \Level2Out192[28] , \Level2Out192[27] , \Level2Out192[26] , 
        \Level2Out192[25] , \Level2Out192[24] , \Level2Out192[23] , 
        \Level2Out192[22] , \Level2Out192[21] , \Level2Out192[20] , 
        \Level2Out192[19] , \Level2Out192[18] , \Level2Out192[17] , 
        \Level2Out192[16] , \Level2Out192[15] , \Level2Out192[14] , 
        \Level2Out192[13] , \Level2Out192[12] , \Level2Out192[11] , 
        \Level2Out192[10] , \Level2Out192[9] , \Level2Out192[8] , 
        \Level2Out192[7] , \Level2Out192[6] , \Level2Out192[5] , 
        \Level2Out192[4] , \Level2Out192[3] , \Level2Out192[2] , 
        \Level2Out192[1] , \Level2Out192[0] }), .In2({\Level2Out194[31] , 
        \Level2Out194[30] , \Level2Out194[29] , \Level2Out194[28] , 
        \Level2Out194[27] , \Level2Out194[26] , \Level2Out194[25] , 
        \Level2Out194[24] , \Level2Out194[23] , \Level2Out194[22] , 
        \Level2Out194[21] , \Level2Out194[20] , \Level2Out194[19] , 
        \Level2Out194[18] , \Level2Out194[17] , \Level2Out194[16] , 
        \Level2Out194[15] , \Level2Out194[14] , \Level2Out194[13] , 
        \Level2Out194[12] , \Level2Out194[11] , \Level2Out194[10] , 
        \Level2Out194[9] , \Level2Out194[8] , \Level2Out194[7] , 
        \Level2Out194[6] , \Level2Out194[5] , \Level2Out194[4] , 
        \Level2Out194[3] , \Level2Out194[2] , \Level2Out194[1] , 
        \Level2Out194[0] }), .Read1(\Level2Load192[0] ), .Read2(
        \Level2Load194[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load40[0] ), .Out({\Level8Out40[31] , \Level8Out40[30] , 
        \Level8Out40[29] , \Level8Out40[28] , \Level8Out40[27] , 
        \Level8Out40[26] , \Level8Out40[25] , \Level8Out40[24] , 
        \Level8Out40[23] , \Level8Out40[22] , \Level8Out40[21] , 
        \Level8Out40[20] , \Level8Out40[19] , \Level8Out40[18] , 
        \Level8Out40[17] , \Level8Out40[16] , \Level8Out40[15] , 
        \Level8Out40[14] , \Level8Out40[13] , \Level8Out40[12] , 
        \Level8Out40[11] , \Level8Out40[10] , \Level8Out40[9] , 
        \Level8Out40[8] , \Level8Out40[7] , \Level8Out40[6] , \Level8Out40[5] , 
        \Level8Out40[4] , \Level8Out40[3] , \Level8Out40[2] , \Level8Out40[1] , 
        \Level8Out40[0] }), .In1({\Level4Out40[31] , \Level4Out40[30] , 
        \Level4Out40[29] , \Level4Out40[28] , \Level4Out40[27] , 
        \Level4Out40[26] , \Level4Out40[25] , \Level4Out40[24] , 
        \Level4Out40[23] , \Level4Out40[22] , \Level4Out40[21] , 
        \Level4Out40[20] , \Level4Out40[19] , \Level4Out40[18] , 
        \Level4Out40[17] , \Level4Out40[16] , \Level4Out40[15] , 
        \Level4Out40[14] , \Level4Out40[13] , \Level4Out40[12] , 
        \Level4Out40[11] , \Level4Out40[10] , \Level4Out40[9] , 
        \Level4Out40[8] , \Level4Out40[7] , \Level4Out40[6] , \Level4Out40[5] , 
        \Level4Out40[4] , \Level4Out40[3] , \Level4Out40[2] , \Level4Out40[1] , 
        \Level4Out40[0] }), .In2({\Level4Out44[31] , \Level4Out44[30] , 
        \Level4Out44[29] , \Level4Out44[28] , \Level4Out44[27] , 
        \Level4Out44[26] , \Level4Out44[25] , \Level4Out44[24] , 
        \Level4Out44[23] , \Level4Out44[22] , \Level4Out44[21] , 
        \Level4Out44[20] , \Level4Out44[19] , \Level4Out44[18] , 
        \Level4Out44[17] , \Level4Out44[16] , \Level4Out44[15] , 
        \Level4Out44[14] , \Level4Out44[13] , \Level4Out44[12] , 
        \Level4Out44[11] , \Level4Out44[10] , \Level4Out44[9] , 
        \Level4Out44[8] , \Level4Out44[7] , \Level4Out44[6] , \Level4Out44[5] , 
        \Level4Out44[4] , \Level4Out44[3] , \Level4Out44[2] , \Level4Out44[1] , 
        \Level4Out44[0] }), .Read1(\Level4Load40[0] ), .Read2(
        \Level4Load44[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_232_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load232[0] ), .Out({\Level8Out232[31] , \Level8Out232[30] , 
        \Level8Out232[29] , \Level8Out232[28] , \Level8Out232[27] , 
        \Level8Out232[26] , \Level8Out232[25] , \Level8Out232[24] , 
        \Level8Out232[23] , \Level8Out232[22] , \Level8Out232[21] , 
        \Level8Out232[20] , \Level8Out232[19] , \Level8Out232[18] , 
        \Level8Out232[17] , \Level8Out232[16] , \Level8Out232[15] , 
        \Level8Out232[14] , \Level8Out232[13] , \Level8Out232[12] , 
        \Level8Out232[11] , \Level8Out232[10] , \Level8Out232[9] , 
        \Level8Out232[8] , \Level8Out232[7] , \Level8Out232[6] , 
        \Level8Out232[5] , \Level8Out232[4] , \Level8Out232[3] , 
        \Level8Out232[2] , \Level8Out232[1] , \Level8Out232[0] }), .In1({
        \Level4Out232[31] , \Level4Out232[30] , \Level4Out232[29] , 
        \Level4Out232[28] , \Level4Out232[27] , \Level4Out232[26] , 
        \Level4Out232[25] , \Level4Out232[24] , \Level4Out232[23] , 
        \Level4Out232[22] , \Level4Out232[21] , \Level4Out232[20] , 
        \Level4Out232[19] , \Level4Out232[18] , \Level4Out232[17] , 
        \Level4Out232[16] , \Level4Out232[15] , \Level4Out232[14] , 
        \Level4Out232[13] , \Level4Out232[12] , \Level4Out232[11] , 
        \Level4Out232[10] , \Level4Out232[9] , \Level4Out232[8] , 
        \Level4Out232[7] , \Level4Out232[6] , \Level4Out232[5] , 
        \Level4Out232[4] , \Level4Out232[3] , \Level4Out232[2] , 
        \Level4Out232[1] , \Level4Out232[0] }), .In2({\Level4Out236[31] , 
        \Level4Out236[30] , \Level4Out236[29] , \Level4Out236[28] , 
        \Level4Out236[27] , \Level4Out236[26] , \Level4Out236[25] , 
        \Level4Out236[24] , \Level4Out236[23] , \Level4Out236[22] , 
        \Level4Out236[21] , \Level4Out236[20] , \Level4Out236[19] , 
        \Level4Out236[18] , \Level4Out236[17] , \Level4Out236[16] , 
        \Level4Out236[15] , \Level4Out236[14] , \Level4Out236[13] , 
        \Level4Out236[12] , \Level4Out236[11] , \Level4Out236[10] , 
        \Level4Out236[9] , \Level4Out236[8] , \Level4Out236[7] , 
        \Level4Out236[6] , \Level4Out236[5] , \Level4Out236[4] , 
        \Level4Out236[3] , \Level4Out236[2] , \Level4Out236[1] , 
        \Level4Out236[0] }), .Read1(\Level4Load232[0] ), .Read2(
        \Level4Load236[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanOut({\ScanLink12[31] , 
        \ScanLink12[30] , \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , 
        \ScanLink12[26] , \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , 
        \ScanLink12[22] , \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , 
        \ScanLink12[18] , \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , 
        \ScanLink12[14] , \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , 
        \ScanLink12[10] , \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , 
        \ScanLink12[6] , \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , 
        \ScanLink12[2] , \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load11[0] ), .Out({
        \Level1Out11[31] , \Level1Out11[30] , \Level1Out11[29] , 
        \Level1Out11[28] , \Level1Out11[27] , \Level1Out11[26] , 
        \Level1Out11[25] , \Level1Out11[24] , \Level1Out11[23] , 
        \Level1Out11[22] , \Level1Out11[21] , \Level1Out11[20] , 
        \Level1Out11[19] , \Level1Out11[18] , \Level1Out11[17] , 
        \Level1Out11[16] , \Level1Out11[15] , \Level1Out11[14] , 
        \Level1Out11[13] , \Level1Out11[12] , \Level1Out11[11] , 
        \Level1Out11[10] , \Level1Out11[9] , \Level1Out11[8] , 
        \Level1Out11[7] , \Level1Out11[6] , \Level1Out11[5] , \Level1Out11[4] , 
        \Level1Out11[3] , \Level1Out11[2] , \Level1Out11[1] , \Level1Out11[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_25 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanOut({\ScanLink26[31] , 
        \ScanLink26[30] , \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , 
        \ScanLink26[26] , \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , 
        \ScanLink26[22] , \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , 
        \ScanLink26[18] , \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , 
        \ScanLink26[14] , \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , 
        \ScanLink26[10] , \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , 
        \ScanLink26[6] , \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , 
        \ScanLink26[2] , \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load25[0] ), .Out({
        \Level1Out25[31] , \Level1Out25[30] , \Level1Out25[29] , 
        \Level1Out25[28] , \Level1Out25[27] , \Level1Out25[26] , 
        \Level1Out25[25] , \Level1Out25[24] , \Level1Out25[23] , 
        \Level1Out25[22] , \Level1Out25[21] , \Level1Out25[20] , 
        \Level1Out25[19] , \Level1Out25[18] , \Level1Out25[17] , 
        \Level1Out25[16] , \Level1Out25[15] , \Level1Out25[14] , 
        \Level1Out25[13] , \Level1Out25[12] , \Level1Out25[11] , 
        \Level1Out25[10] , \Level1Out25[9] , \Level1Out25[8] , 
        \Level1Out25[7] , \Level1Out25[6] , \Level1Out25[5] , \Level1Out25[4] , 
        \Level1Out25[3] , \Level1Out25[2] , \Level1Out25[1] , \Level1Out25[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_169 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink169[31] , \ScanLink169[30] , 
        \ScanLink169[29] , \ScanLink169[28] , \ScanLink169[27] , 
        \ScanLink169[26] , \ScanLink169[25] , \ScanLink169[24] , 
        \ScanLink169[23] , \ScanLink169[22] , \ScanLink169[21] , 
        \ScanLink169[20] , \ScanLink169[19] , \ScanLink169[18] , 
        \ScanLink169[17] , \ScanLink169[16] , \ScanLink169[15] , 
        \ScanLink169[14] , \ScanLink169[13] , \ScanLink169[12] , 
        \ScanLink169[11] , \ScanLink169[10] , \ScanLink169[9] , 
        \ScanLink169[8] , \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , 
        \ScanLink169[4] , \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , 
        \ScanLink169[0] }), .ScanOut({\ScanLink170[31] , \ScanLink170[30] , 
        \ScanLink170[29] , \ScanLink170[28] , \ScanLink170[27] , 
        \ScanLink170[26] , \ScanLink170[25] , \ScanLink170[24] , 
        \ScanLink170[23] , \ScanLink170[22] , \ScanLink170[21] , 
        \ScanLink170[20] , \ScanLink170[19] , \ScanLink170[18] , 
        \ScanLink170[17] , \ScanLink170[16] , \ScanLink170[15] , 
        \ScanLink170[14] , \ScanLink170[13] , \ScanLink170[12] , 
        \ScanLink170[11] , \ScanLink170[10] , \ScanLink170[9] , 
        \ScanLink170[8] , \ScanLink170[7] , \ScanLink170[6] , \ScanLink170[5] , 
        \ScanLink170[4] , \ScanLink170[3] , \ScanLink170[2] , \ScanLink170[1] , 
        \ScanLink170[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load169[0] ), .Out({\Level1Out169[31] , \Level1Out169[30] , 
        \Level1Out169[29] , \Level1Out169[28] , \Level1Out169[27] , 
        \Level1Out169[26] , \Level1Out169[25] , \Level1Out169[24] , 
        \Level1Out169[23] , \Level1Out169[22] , \Level1Out169[21] , 
        \Level1Out169[20] , \Level1Out169[19] , \Level1Out169[18] , 
        \Level1Out169[17] , \Level1Out169[16] , \Level1Out169[15] , 
        \Level1Out169[14] , \Level1Out169[13] , \Level1Out169[12] , 
        \Level1Out169[11] , \Level1Out169[10] , \Level1Out169[9] , 
        \Level1Out169[8] , \Level1Out169[7] , \Level1Out169[6] , 
        \Level1Out169[5] , \Level1Out169[4] , \Level1Out169[3] , 
        \Level1Out169[2] , \Level1Out169[1] , \Level1Out169[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_74_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load74[0] ), .Out({\Level2Out74[31] , \Level2Out74[30] , 
        \Level2Out74[29] , \Level2Out74[28] , \Level2Out74[27] , 
        \Level2Out74[26] , \Level2Out74[25] , \Level2Out74[24] , 
        \Level2Out74[23] , \Level2Out74[22] , \Level2Out74[21] , 
        \Level2Out74[20] , \Level2Out74[19] , \Level2Out74[18] , 
        \Level2Out74[17] , \Level2Out74[16] , \Level2Out74[15] , 
        \Level2Out74[14] , \Level2Out74[13] , \Level2Out74[12] , 
        \Level2Out74[11] , \Level2Out74[10] , \Level2Out74[9] , 
        \Level2Out74[8] , \Level2Out74[7] , \Level2Out74[6] , \Level2Out74[5] , 
        \Level2Out74[4] , \Level2Out74[3] , \Level2Out74[2] , \Level2Out74[1] , 
        \Level2Out74[0] }), .In1({\Level1Out74[31] , \Level1Out74[30] , 
        \Level1Out74[29] , \Level1Out74[28] , \Level1Out74[27] , 
        \Level1Out74[26] , \Level1Out74[25] , \Level1Out74[24] , 
        \Level1Out74[23] , \Level1Out74[22] , \Level1Out74[21] , 
        \Level1Out74[20] , \Level1Out74[19] , \Level1Out74[18] , 
        \Level1Out74[17] , \Level1Out74[16] , \Level1Out74[15] , 
        \Level1Out74[14] , \Level1Out74[13] , \Level1Out74[12] , 
        \Level1Out74[11] , \Level1Out74[10] , \Level1Out74[9] , 
        \Level1Out74[8] , \Level1Out74[7] , \Level1Out74[6] , \Level1Out74[5] , 
        \Level1Out74[4] , \Level1Out74[3] , \Level1Out74[2] , \Level1Out74[1] , 
        \Level1Out74[0] }), .In2({\Level1Out75[31] , \Level1Out75[30] , 
        \Level1Out75[29] , \Level1Out75[28] , \Level1Out75[27] , 
        \Level1Out75[26] , \Level1Out75[25] , \Level1Out75[24] , 
        \Level1Out75[23] , \Level1Out75[22] , \Level1Out75[21] , 
        \Level1Out75[20] , \Level1Out75[19] , \Level1Out75[18] , 
        \Level1Out75[17] , \Level1Out75[16] , \Level1Out75[15] , 
        \Level1Out75[14] , \Level1Out75[13] , \Level1Out75[12] , 
        \Level1Out75[11] , \Level1Out75[10] , \Level1Out75[9] , 
        \Level1Out75[8] , \Level1Out75[7] , \Level1Out75[6] , \Level1Out75[5] , 
        \Level1Out75[4] , \Level1Out75[3] , \Level1Out75[2] , \Level1Out75[1] , 
        \Level1Out75[0] }), .Read1(\Level1Load74[0] ), .Read2(
        \Level1Load75[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_118_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load118[0] ), .Out({\Level2Out118[31] , \Level2Out118[30] , 
        \Level2Out118[29] , \Level2Out118[28] , \Level2Out118[27] , 
        \Level2Out118[26] , \Level2Out118[25] , \Level2Out118[24] , 
        \Level2Out118[23] , \Level2Out118[22] , \Level2Out118[21] , 
        \Level2Out118[20] , \Level2Out118[19] , \Level2Out118[18] , 
        \Level2Out118[17] , \Level2Out118[16] , \Level2Out118[15] , 
        \Level2Out118[14] , \Level2Out118[13] , \Level2Out118[12] , 
        \Level2Out118[11] , \Level2Out118[10] , \Level2Out118[9] , 
        \Level2Out118[8] , \Level2Out118[7] , \Level2Out118[6] , 
        \Level2Out118[5] , \Level2Out118[4] , \Level2Out118[3] , 
        \Level2Out118[2] , \Level2Out118[1] , \Level2Out118[0] }), .In1({
        \Level1Out118[31] , \Level1Out118[30] , \Level1Out118[29] , 
        \Level1Out118[28] , \Level1Out118[27] , \Level1Out118[26] , 
        \Level1Out118[25] , \Level1Out118[24] , \Level1Out118[23] , 
        \Level1Out118[22] , \Level1Out118[21] , \Level1Out118[20] , 
        \Level1Out118[19] , \Level1Out118[18] , \Level1Out118[17] , 
        \Level1Out118[16] , \Level1Out118[15] , \Level1Out118[14] , 
        \Level1Out118[13] , \Level1Out118[12] , \Level1Out118[11] , 
        \Level1Out118[10] , \Level1Out118[9] , \Level1Out118[8] , 
        \Level1Out118[7] , \Level1Out118[6] , \Level1Out118[5] , 
        \Level1Out118[4] , \Level1Out118[3] , \Level1Out118[2] , 
        \Level1Out118[1] , \Level1Out118[0] }), .In2({\Level1Out119[31] , 
        \Level1Out119[30] , \Level1Out119[29] , \Level1Out119[28] , 
        \Level1Out119[27] , \Level1Out119[26] , \Level1Out119[25] , 
        \Level1Out119[24] , \Level1Out119[23] , \Level1Out119[22] , 
        \Level1Out119[21] , \Level1Out119[20] , \Level1Out119[19] , 
        \Level1Out119[18] , \Level1Out119[17] , \Level1Out119[16] , 
        \Level1Out119[15] , \Level1Out119[14] , \Level1Out119[13] , 
        \Level1Out119[12] , \Level1Out119[11] , \Level1Out119[10] , 
        \Level1Out119[9] , \Level1Out119[8] , \Level1Out119[7] , 
        \Level1Out119[6] , \Level1Out119[5] , \Level1Out119[4] , 
        \Level1Out119[3] , \Level1Out119[2] , \Level1Out119[1] , 
        \Level1Out119[0] }), .Read1(\Level1Load118[0] ), .Read2(
        \Level1Load119[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_132_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load132[0] ), .Out({\Level2Out132[31] , \Level2Out132[30] , 
        \Level2Out132[29] , \Level2Out132[28] , \Level2Out132[27] , 
        \Level2Out132[26] , \Level2Out132[25] , \Level2Out132[24] , 
        \Level2Out132[23] , \Level2Out132[22] , \Level2Out132[21] , 
        \Level2Out132[20] , \Level2Out132[19] , \Level2Out132[18] , 
        \Level2Out132[17] , \Level2Out132[16] , \Level2Out132[15] , 
        \Level2Out132[14] , \Level2Out132[13] , \Level2Out132[12] , 
        \Level2Out132[11] , \Level2Out132[10] , \Level2Out132[9] , 
        \Level2Out132[8] , \Level2Out132[7] , \Level2Out132[6] , 
        \Level2Out132[5] , \Level2Out132[4] , \Level2Out132[3] , 
        \Level2Out132[2] , \Level2Out132[1] , \Level2Out132[0] }), .In1({
        \Level1Out132[31] , \Level1Out132[30] , \Level1Out132[29] , 
        \Level1Out132[28] , \Level1Out132[27] , \Level1Out132[26] , 
        \Level1Out132[25] , \Level1Out132[24] , \Level1Out132[23] , 
        \Level1Out132[22] , \Level1Out132[21] , \Level1Out132[20] , 
        \Level1Out132[19] , \Level1Out132[18] , \Level1Out132[17] , 
        \Level1Out132[16] , \Level1Out132[15] , \Level1Out132[14] , 
        \Level1Out132[13] , \Level1Out132[12] , \Level1Out132[11] , 
        \Level1Out132[10] , \Level1Out132[9] , \Level1Out132[8] , 
        \Level1Out132[7] , \Level1Out132[6] , \Level1Out132[5] , 
        \Level1Out132[4] , \Level1Out132[3] , \Level1Out132[2] , 
        \Level1Out132[1] , \Level1Out132[0] }), .In2({\Level1Out133[31] , 
        \Level1Out133[30] , \Level1Out133[29] , \Level1Out133[28] , 
        \Level1Out133[27] , \Level1Out133[26] , \Level1Out133[25] , 
        \Level1Out133[24] , \Level1Out133[23] , \Level1Out133[22] , 
        \Level1Out133[21] , \Level1Out133[20] , \Level1Out133[19] , 
        \Level1Out133[18] , \Level1Out133[17] , \Level1Out133[16] , 
        \Level1Out133[15] , \Level1Out133[14] , \Level1Out133[13] , 
        \Level1Out133[12] , \Level1Out133[11] , \Level1Out133[10] , 
        \Level1Out133[9] , \Level1Out133[8] , \Level1Out133[7] , 
        \Level1Out133[6] , \Level1Out133[5] , \Level1Out133[4] , 
        \Level1Out133[3] , \Level1Out133[2] , \Level1Out133[1] , 
        \Level1Out133[0] }), .Read1(\Level1Load132[0] ), .Read2(
        \Level1Load133[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_206_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load206[0] ), .Out({\Level2Out206[31] , \Level2Out206[30] , 
        \Level2Out206[29] , \Level2Out206[28] , \Level2Out206[27] , 
        \Level2Out206[26] , \Level2Out206[25] , \Level2Out206[24] , 
        \Level2Out206[23] , \Level2Out206[22] , \Level2Out206[21] , 
        \Level2Out206[20] , \Level2Out206[19] , \Level2Out206[18] , 
        \Level2Out206[17] , \Level2Out206[16] , \Level2Out206[15] , 
        \Level2Out206[14] , \Level2Out206[13] , \Level2Out206[12] , 
        \Level2Out206[11] , \Level2Out206[10] , \Level2Out206[9] , 
        \Level2Out206[8] , \Level2Out206[7] , \Level2Out206[6] , 
        \Level2Out206[5] , \Level2Out206[4] , \Level2Out206[3] , 
        \Level2Out206[2] , \Level2Out206[1] , \Level2Out206[0] }), .In1({
        \Level1Out206[31] , \Level1Out206[30] , \Level1Out206[29] , 
        \Level1Out206[28] , \Level1Out206[27] , \Level1Out206[26] , 
        \Level1Out206[25] , \Level1Out206[24] , \Level1Out206[23] , 
        \Level1Out206[22] , \Level1Out206[21] , \Level1Out206[20] , 
        \Level1Out206[19] , \Level1Out206[18] , \Level1Out206[17] , 
        \Level1Out206[16] , \Level1Out206[15] , \Level1Out206[14] , 
        \Level1Out206[13] , \Level1Out206[12] , \Level1Out206[11] , 
        \Level1Out206[10] , \Level1Out206[9] , \Level1Out206[8] , 
        \Level1Out206[7] , \Level1Out206[6] , \Level1Out206[5] , 
        \Level1Out206[4] , \Level1Out206[3] , \Level1Out206[2] , 
        \Level1Out206[1] , \Level1Out206[0] }), .In2({\Level1Out207[31] , 
        \Level1Out207[30] , \Level1Out207[29] , \Level1Out207[28] , 
        \Level1Out207[27] , \Level1Out207[26] , \Level1Out207[25] , 
        \Level1Out207[24] , \Level1Out207[23] , \Level1Out207[22] , 
        \Level1Out207[21] , \Level1Out207[20] , \Level1Out207[19] , 
        \Level1Out207[18] , \Level1Out207[17] , \Level1Out207[16] , 
        \Level1Out207[15] , \Level1Out207[14] , \Level1Out207[13] , 
        \Level1Out207[12] , \Level1Out207[11] , \Level1Out207[10] , 
        \Level1Out207[9] , \Level1Out207[8] , \Level1Out207[7] , 
        \Level1Out207[6] , \Level1Out207[5] , \Level1Out207[4] , 
        \Level1Out207[3] , \Level1Out207[2] , \Level1Out207[1] , 
        \Level1Out207[0] }), .Read1(\Level1Load206[0] ), .Read2(
        \Level1Load207[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_68_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load68[0] ), .Out({\Level4Out68[31] , \Level4Out68[30] , 
        \Level4Out68[29] , \Level4Out68[28] , \Level4Out68[27] , 
        \Level4Out68[26] , \Level4Out68[25] , \Level4Out68[24] , 
        \Level4Out68[23] , \Level4Out68[22] , \Level4Out68[21] , 
        \Level4Out68[20] , \Level4Out68[19] , \Level4Out68[18] , 
        \Level4Out68[17] , \Level4Out68[16] , \Level4Out68[15] , 
        \Level4Out68[14] , \Level4Out68[13] , \Level4Out68[12] , 
        \Level4Out68[11] , \Level4Out68[10] , \Level4Out68[9] , 
        \Level4Out68[8] , \Level4Out68[7] , \Level4Out68[6] , \Level4Out68[5] , 
        \Level4Out68[4] , \Level4Out68[3] , \Level4Out68[2] , \Level4Out68[1] , 
        \Level4Out68[0] }), .In1({\Level2Out68[31] , \Level2Out68[30] , 
        \Level2Out68[29] , \Level2Out68[28] , \Level2Out68[27] , 
        \Level2Out68[26] , \Level2Out68[25] , \Level2Out68[24] , 
        \Level2Out68[23] , \Level2Out68[22] , \Level2Out68[21] , 
        \Level2Out68[20] , \Level2Out68[19] , \Level2Out68[18] , 
        \Level2Out68[17] , \Level2Out68[16] , \Level2Out68[15] , 
        \Level2Out68[14] , \Level2Out68[13] , \Level2Out68[12] , 
        \Level2Out68[11] , \Level2Out68[10] , \Level2Out68[9] , 
        \Level2Out68[8] , \Level2Out68[7] , \Level2Out68[6] , \Level2Out68[5] , 
        \Level2Out68[4] , \Level2Out68[3] , \Level2Out68[2] , \Level2Out68[1] , 
        \Level2Out68[0] }), .In2({\Level2Out70[31] , \Level2Out70[30] , 
        \Level2Out70[29] , \Level2Out70[28] , \Level2Out70[27] , 
        \Level2Out70[26] , \Level2Out70[25] , \Level2Out70[24] , 
        \Level2Out70[23] , \Level2Out70[22] , \Level2Out70[21] , 
        \Level2Out70[20] , \Level2Out70[19] , \Level2Out70[18] , 
        \Level2Out70[17] , \Level2Out70[16] , \Level2Out70[15] , 
        \Level2Out70[14] , \Level2Out70[13] , \Level2Out70[12] , 
        \Level2Out70[11] , \Level2Out70[10] , \Level2Out70[9] , 
        \Level2Out70[8] , \Level2Out70[7] , \Level2Out70[6] , \Level2Out70[5] , 
        \Level2Out70[4] , \Level2Out70[3] , \Level2Out70[2] , \Level2Out70[1] , 
        \Level2Out70[0] }), .Read1(\Level2Load68[0] ), .Read2(
        \Level2Load70[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_104_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load104[0] ), .Out({\Level4Out104[31] , \Level4Out104[30] , 
        \Level4Out104[29] , \Level4Out104[28] , \Level4Out104[27] , 
        \Level4Out104[26] , \Level4Out104[25] , \Level4Out104[24] , 
        \Level4Out104[23] , \Level4Out104[22] , \Level4Out104[21] , 
        \Level4Out104[20] , \Level4Out104[19] , \Level4Out104[18] , 
        \Level4Out104[17] , \Level4Out104[16] , \Level4Out104[15] , 
        \Level4Out104[14] , \Level4Out104[13] , \Level4Out104[12] , 
        \Level4Out104[11] , \Level4Out104[10] , \Level4Out104[9] , 
        \Level4Out104[8] , \Level4Out104[7] , \Level4Out104[6] , 
        \Level4Out104[5] , \Level4Out104[4] , \Level4Out104[3] , 
        \Level4Out104[2] , \Level4Out104[1] , \Level4Out104[0] }), .In1({
        \Level2Out104[31] , \Level2Out104[30] , \Level2Out104[29] , 
        \Level2Out104[28] , \Level2Out104[27] , \Level2Out104[26] , 
        \Level2Out104[25] , \Level2Out104[24] , \Level2Out104[23] , 
        \Level2Out104[22] , \Level2Out104[21] , \Level2Out104[20] , 
        \Level2Out104[19] , \Level2Out104[18] , \Level2Out104[17] , 
        \Level2Out104[16] , \Level2Out104[15] , \Level2Out104[14] , 
        \Level2Out104[13] , \Level2Out104[12] , \Level2Out104[11] , 
        \Level2Out104[10] , \Level2Out104[9] , \Level2Out104[8] , 
        \Level2Out104[7] , \Level2Out104[6] , \Level2Out104[5] , 
        \Level2Out104[4] , \Level2Out104[3] , \Level2Out104[2] , 
        \Level2Out104[1] , \Level2Out104[0] }), .In2({\Level2Out106[31] , 
        \Level2Out106[30] , \Level2Out106[29] , \Level2Out106[28] , 
        \Level2Out106[27] , \Level2Out106[26] , \Level2Out106[25] , 
        \Level2Out106[24] , \Level2Out106[23] , \Level2Out106[22] , 
        \Level2Out106[21] , \Level2Out106[20] , \Level2Out106[19] , 
        \Level2Out106[18] , \Level2Out106[17] , \Level2Out106[16] , 
        \Level2Out106[15] , \Level2Out106[14] , \Level2Out106[13] , 
        \Level2Out106[12] , \Level2Out106[11] , \Level2Out106[10] , 
        \Level2Out106[9] , \Level2Out106[8] , \Level2Out106[7] , 
        \Level2Out106[6] , \Level2Out106[5] , \Level2Out106[4] , 
        \Level2Out106[3] , \Level2Out106[2] , \Level2Out106[1] , 
        \Level2Out106[0] }), .Read1(\Level2Load104[0] ), .Read2(
        \Level2Load106[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_43 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanOut({\ScanLink44[31] , 
        \ScanLink44[30] , \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , 
        \ScanLink44[26] , \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , 
        \ScanLink44[22] , \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , 
        \ScanLink44[18] , \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , 
        \ScanLink44[14] , \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , 
        \ScanLink44[10] , \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , 
        \ScanLink44[6] , \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , 
        \ScanLink44[2] , \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load43[0] ), .Out({
        \Level1Out43[31] , \Level1Out43[30] , \Level1Out43[29] , 
        \Level1Out43[28] , \Level1Out43[27] , \Level1Out43[26] , 
        \Level1Out43[25] , \Level1Out43[24] , \Level1Out43[23] , 
        \Level1Out43[22] , \Level1Out43[21] , \Level1Out43[20] , 
        \Level1Out43[19] , \Level1Out43[18] , \Level1Out43[17] , 
        \Level1Out43[16] , \Level1Out43[15] , \Level1Out43[14] , 
        \Level1Out43[13] , \Level1Out43[12] , \Level1Out43[11] , 
        \Level1Out43[10] , \Level1Out43[9] , \Level1Out43[8] , 
        \Level1Out43[7] , \Level1Out43[6] , \Level1Out43[5] , \Level1Out43[4] , 
        \Level1Out43[3] , \Level1Out43[2] , \Level1Out43[1] , \Level1Out43[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_64 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink64[31] , \ScanLink64[30] , 
        \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , 
        \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , 
        \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , 
        \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , 
        \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , 
        \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , 
        \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , 
        \ScanLink64[1] , \ScanLink64[0] }), .ScanOut({\ScanLink65[31] , 
        \ScanLink65[30] , \ScanLink65[29] , \ScanLink65[28] , \ScanLink65[27] , 
        \ScanLink65[26] , \ScanLink65[25] , \ScanLink65[24] , \ScanLink65[23] , 
        \ScanLink65[22] , \ScanLink65[21] , \ScanLink65[20] , \ScanLink65[19] , 
        \ScanLink65[18] , \ScanLink65[17] , \ScanLink65[16] , \ScanLink65[15] , 
        \ScanLink65[14] , \ScanLink65[13] , \ScanLink65[12] , \ScanLink65[11] , 
        \ScanLink65[10] , \ScanLink65[9] , \ScanLink65[8] , \ScanLink65[7] , 
        \ScanLink65[6] , \ScanLink65[5] , \ScanLink65[4] , \ScanLink65[3] , 
        \ScanLink65[2] , \ScanLink65[1] , \ScanLink65[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load64[0] ), .Out({
        \Level1Out64[31] , \Level1Out64[30] , \Level1Out64[29] , 
        \Level1Out64[28] , \Level1Out64[27] , \Level1Out64[26] , 
        \Level1Out64[25] , \Level1Out64[24] , \Level1Out64[23] , 
        \Level1Out64[22] , \Level1Out64[21] , \Level1Out64[20] , 
        \Level1Out64[19] , \Level1Out64[18] , \Level1Out64[17] , 
        \Level1Out64[16] , \Level1Out64[15] , \Level1Out64[14] , 
        \Level1Out64[13] , \Level1Out64[12] , \Level1Out64[11] , 
        \Level1Out64[10] , \Level1Out64[9] , \Level1Out64[8] , 
        \Level1Out64[7] , \Level1Out64[6] , \Level1Out64[5] , \Level1Out64[4] , 
        \Level1Out64[3] , \Level1Out64[2] , \Level1Out64[1] , \Level1Out64[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_81 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink81[31] , \ScanLink81[30] , 
        \ScanLink81[29] , \ScanLink81[28] , \ScanLink81[27] , \ScanLink81[26] , 
        \ScanLink81[25] , \ScanLink81[24] , \ScanLink81[23] , \ScanLink81[22] , 
        \ScanLink81[21] , \ScanLink81[20] , \ScanLink81[19] , \ScanLink81[18] , 
        \ScanLink81[17] , \ScanLink81[16] , \ScanLink81[15] , \ScanLink81[14] , 
        \ScanLink81[13] , \ScanLink81[12] , \ScanLink81[11] , \ScanLink81[10] , 
        \ScanLink81[9] , \ScanLink81[8] , \ScanLink81[7] , \ScanLink81[6] , 
        \ScanLink81[5] , \ScanLink81[4] , \ScanLink81[3] , \ScanLink81[2] , 
        \ScanLink81[1] , \ScanLink81[0] }), .ScanOut({\ScanLink82[31] , 
        \ScanLink82[30] , \ScanLink82[29] , \ScanLink82[28] , \ScanLink82[27] , 
        \ScanLink82[26] , \ScanLink82[25] , \ScanLink82[24] , \ScanLink82[23] , 
        \ScanLink82[22] , \ScanLink82[21] , \ScanLink82[20] , \ScanLink82[19] , 
        \ScanLink82[18] , \ScanLink82[17] , \ScanLink82[16] , \ScanLink82[15] , 
        \ScanLink82[14] , \ScanLink82[13] , \ScanLink82[12] , \ScanLink82[11] , 
        \ScanLink82[10] , \ScanLink82[9] , \ScanLink82[8] , \ScanLink82[7] , 
        \ScanLink82[6] , \ScanLink82[5] , \ScanLink82[4] , \ScanLink82[3] , 
        \ScanLink82[2] , \ScanLink82[1] , \ScanLink82[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load81[0] ), .Out({
        \Level1Out81[31] , \Level1Out81[30] , \Level1Out81[29] , 
        \Level1Out81[28] , \Level1Out81[27] , \Level1Out81[26] , 
        \Level1Out81[25] , \Level1Out81[24] , \Level1Out81[23] , 
        \Level1Out81[22] , \Level1Out81[21] , \Level1Out81[20] , 
        \Level1Out81[19] , \Level1Out81[18] , \Level1Out81[17] , 
        \Level1Out81[16] , \Level1Out81[15] , \Level1Out81[14] , 
        \Level1Out81[13] , \Level1Out81[12] , \Level1Out81[11] , 
        \Level1Out81[10] , \Level1Out81[9] , \Level1Out81[8] , 
        \Level1Out81[7] , \Level1Out81[6] , \Level1Out81[5] , \Level1Out81[4] , 
        \Level1Out81[3] , \Level1Out81[2] , \Level1Out81[1] , \Level1Out81[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_89 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink89[31] , \ScanLink89[30] , 
        \ScanLink89[29] , \ScanLink89[28] , \ScanLink89[27] , \ScanLink89[26] , 
        \ScanLink89[25] , \ScanLink89[24] , \ScanLink89[23] , \ScanLink89[22] , 
        \ScanLink89[21] , \ScanLink89[20] , \ScanLink89[19] , \ScanLink89[18] , 
        \ScanLink89[17] , \ScanLink89[16] , \ScanLink89[15] , \ScanLink89[14] , 
        \ScanLink89[13] , \ScanLink89[12] , \ScanLink89[11] , \ScanLink89[10] , 
        \ScanLink89[9] , \ScanLink89[8] , \ScanLink89[7] , \ScanLink89[6] , 
        \ScanLink89[5] , \ScanLink89[4] , \ScanLink89[3] , \ScanLink89[2] , 
        \ScanLink89[1] , \ScanLink89[0] }), .ScanOut({\ScanLink90[31] , 
        \ScanLink90[30] , \ScanLink90[29] , \ScanLink90[28] , \ScanLink90[27] , 
        \ScanLink90[26] , \ScanLink90[25] , \ScanLink90[24] , \ScanLink90[23] , 
        \ScanLink90[22] , \ScanLink90[21] , \ScanLink90[20] , \ScanLink90[19] , 
        \ScanLink90[18] , \ScanLink90[17] , \ScanLink90[16] , \ScanLink90[15] , 
        \ScanLink90[14] , \ScanLink90[13] , \ScanLink90[12] , \ScanLink90[11] , 
        \ScanLink90[10] , \ScanLink90[9] , \ScanLink90[8] , \ScanLink90[7] , 
        \ScanLink90[6] , \ScanLink90[5] , \ScanLink90[4] , \ScanLink90[3] , 
        \ScanLink90[2] , \ScanLink90[1] , \ScanLink90[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load89[0] ), .Out({
        \Level1Out89[31] , \Level1Out89[30] , \Level1Out89[29] , 
        \Level1Out89[28] , \Level1Out89[27] , \Level1Out89[26] , 
        \Level1Out89[25] , \Level1Out89[24] , \Level1Out89[23] , 
        \Level1Out89[22] , \Level1Out89[21] , \Level1Out89[20] , 
        \Level1Out89[19] , \Level1Out89[18] , \Level1Out89[17] , 
        \Level1Out89[16] , \Level1Out89[15] , \Level1Out89[14] , 
        \Level1Out89[13] , \Level1Out89[12] , \Level1Out89[11] , 
        \Level1Out89[10] , \Level1Out89[9] , \Level1Out89[8] , 
        \Level1Out89[7] , \Level1Out89[6] , \Level1Out89[5] , \Level1Out89[4] , 
        \Level1Out89[3] , \Level1Out89[2] , \Level1Out89[1] , \Level1Out89[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_107 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink107[31] , \ScanLink107[30] , 
        \ScanLink107[29] , \ScanLink107[28] , \ScanLink107[27] , 
        \ScanLink107[26] , \ScanLink107[25] , \ScanLink107[24] , 
        \ScanLink107[23] , \ScanLink107[22] , \ScanLink107[21] , 
        \ScanLink107[20] , \ScanLink107[19] , \ScanLink107[18] , 
        \ScanLink107[17] , \ScanLink107[16] , \ScanLink107[15] , 
        \ScanLink107[14] , \ScanLink107[13] , \ScanLink107[12] , 
        \ScanLink107[11] , \ScanLink107[10] , \ScanLink107[9] , 
        \ScanLink107[8] , \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , 
        \ScanLink107[4] , \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , 
        \ScanLink107[0] }), .ScanOut({\ScanLink108[31] , \ScanLink108[30] , 
        \ScanLink108[29] , \ScanLink108[28] , \ScanLink108[27] , 
        \ScanLink108[26] , \ScanLink108[25] , \ScanLink108[24] , 
        \ScanLink108[23] , \ScanLink108[22] , \ScanLink108[21] , 
        \ScanLink108[20] , \ScanLink108[19] , \ScanLink108[18] , 
        \ScanLink108[17] , \ScanLink108[16] , \ScanLink108[15] , 
        \ScanLink108[14] , \ScanLink108[13] , \ScanLink108[12] , 
        \ScanLink108[11] , \ScanLink108[10] , \ScanLink108[9] , 
        \ScanLink108[8] , \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , 
        \ScanLink108[4] , \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , 
        \ScanLink108[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load107[0] ), .Out({\Level1Out107[31] , \Level1Out107[30] , 
        \Level1Out107[29] , \Level1Out107[28] , \Level1Out107[27] , 
        \Level1Out107[26] , \Level1Out107[25] , \Level1Out107[24] , 
        \Level1Out107[23] , \Level1Out107[22] , \Level1Out107[21] , 
        \Level1Out107[20] , \Level1Out107[19] , \Level1Out107[18] , 
        \Level1Out107[17] , \Level1Out107[16] , \Level1Out107[15] , 
        \Level1Out107[14] , \Level1Out107[13] , \Level1Out107[12] , 
        \Level1Out107[11] , \Level1Out107[10] , \Level1Out107[9] , 
        \Level1Out107[8] , \Level1Out107[7] , \Level1Out107[6] , 
        \Level1Out107[5] , \Level1Out107[4] , \Level1Out107[3] , 
        \Level1Out107[2] , \Level1Out107[1] , \Level1Out107[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_237 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink237[31] , \ScanLink237[30] , 
        \ScanLink237[29] , \ScanLink237[28] , \ScanLink237[27] , 
        \ScanLink237[26] , \ScanLink237[25] , \ScanLink237[24] , 
        \ScanLink237[23] , \ScanLink237[22] , \ScanLink237[21] , 
        \ScanLink237[20] , \ScanLink237[19] , \ScanLink237[18] , 
        \ScanLink237[17] , \ScanLink237[16] , \ScanLink237[15] , 
        \ScanLink237[14] , \ScanLink237[13] , \ScanLink237[12] , 
        \ScanLink237[11] , \ScanLink237[10] , \ScanLink237[9] , 
        \ScanLink237[8] , \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , 
        \ScanLink237[4] , \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , 
        \ScanLink237[0] }), .ScanOut({\ScanLink238[31] , \ScanLink238[30] , 
        \ScanLink238[29] , \ScanLink238[28] , \ScanLink238[27] , 
        \ScanLink238[26] , \ScanLink238[25] , \ScanLink238[24] , 
        \ScanLink238[23] , \ScanLink238[22] , \ScanLink238[21] , 
        \ScanLink238[20] , \ScanLink238[19] , \ScanLink238[18] , 
        \ScanLink238[17] , \ScanLink238[16] , \ScanLink238[15] , 
        \ScanLink238[14] , \ScanLink238[13] , \ScanLink238[12] , 
        \ScanLink238[11] , \ScanLink238[10] , \ScanLink238[9] , 
        \ScanLink238[8] , \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , 
        \ScanLink238[4] , \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , 
        \ScanLink238[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load237[0] ), .Out({\Level1Out237[31] , \Level1Out237[30] , 
        \Level1Out237[29] , \Level1Out237[28] , \Level1Out237[27] , 
        \Level1Out237[26] , \Level1Out237[25] , \Level1Out237[24] , 
        \Level1Out237[23] , \Level1Out237[22] , \Level1Out237[21] , 
        \Level1Out237[20] , \Level1Out237[19] , \Level1Out237[18] , 
        \Level1Out237[17] , \Level1Out237[16] , \Level1Out237[15] , 
        \Level1Out237[14] , \Level1Out237[13] , \Level1Out237[12] , 
        \Level1Out237[11] , \Level1Out237[10] , \Level1Out237[9] , 
        \Level1Out237[8] , \Level1Out237[7] , \Level1Out237[6] , 
        \Level1Out237[5] , \Level1Out237[4] , \Level1Out237[3] , 
        \Level1Out237[2] , \Level1Out237[1] , \Level1Out237[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_176_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load176[0] ), .Out({\Level16Out176[31] , \Level16Out176[30] , 
        \Level16Out176[29] , \Level16Out176[28] , \Level16Out176[27] , 
        \Level16Out176[26] , \Level16Out176[25] , \Level16Out176[24] , 
        \Level16Out176[23] , \Level16Out176[22] , \Level16Out176[21] , 
        \Level16Out176[20] , \Level16Out176[19] , \Level16Out176[18] , 
        \Level16Out176[17] , \Level16Out176[16] , \Level16Out176[15] , 
        \Level16Out176[14] , \Level16Out176[13] , \Level16Out176[12] , 
        \Level16Out176[11] , \Level16Out176[10] , \Level16Out176[9] , 
        \Level16Out176[8] , \Level16Out176[7] , \Level16Out176[6] , 
        \Level16Out176[5] , \Level16Out176[4] , \Level16Out176[3] , 
        \Level16Out176[2] , \Level16Out176[1] , \Level16Out176[0] }), .In1({
        \Level8Out176[31] , \Level8Out176[30] , \Level8Out176[29] , 
        \Level8Out176[28] , \Level8Out176[27] , \Level8Out176[26] , 
        \Level8Out176[25] , \Level8Out176[24] , \Level8Out176[23] , 
        \Level8Out176[22] , \Level8Out176[21] , \Level8Out176[20] , 
        \Level8Out176[19] , \Level8Out176[18] , \Level8Out176[17] , 
        \Level8Out176[16] , \Level8Out176[15] , \Level8Out176[14] , 
        \Level8Out176[13] , \Level8Out176[12] , \Level8Out176[11] , 
        \Level8Out176[10] , \Level8Out176[9] , \Level8Out176[8] , 
        \Level8Out176[7] , \Level8Out176[6] , \Level8Out176[5] , 
        \Level8Out176[4] , \Level8Out176[3] , \Level8Out176[2] , 
        \Level8Out176[1] , \Level8Out176[0] }), .In2({\Level8Out184[31] , 
        \Level8Out184[30] , \Level8Out184[29] , \Level8Out184[28] , 
        \Level8Out184[27] , \Level8Out184[26] , \Level8Out184[25] , 
        \Level8Out184[24] , \Level8Out184[23] , \Level8Out184[22] , 
        \Level8Out184[21] , \Level8Out184[20] , \Level8Out184[19] , 
        \Level8Out184[18] , \Level8Out184[17] , \Level8Out184[16] , 
        \Level8Out184[15] , \Level8Out184[14] , \Level8Out184[13] , 
        \Level8Out184[12] , \Level8Out184[11] , \Level8Out184[10] , 
        \Level8Out184[9] , \Level8Out184[8] , \Level8Out184[7] , 
        \Level8Out184[6] , \Level8Out184[5] , \Level8Out184[4] , 
        \Level8Out184[3] , \Level8Out184[2] , \Level8Out184[1] , 
        \Level8Out184[0] }), .Read1(\Level8Load176[0] ), .Read2(
        \Level8Load184[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load6[0] ), .Out({\Level2Out6[31] , \Level2Out6[30] , 
        \Level2Out6[29] , \Level2Out6[28] , \Level2Out6[27] , \Level2Out6[26] , 
        \Level2Out6[25] , \Level2Out6[24] , \Level2Out6[23] , \Level2Out6[22] , 
        \Level2Out6[21] , \Level2Out6[20] , \Level2Out6[19] , \Level2Out6[18] , 
        \Level2Out6[17] , \Level2Out6[16] , \Level2Out6[15] , \Level2Out6[14] , 
        \Level2Out6[13] , \Level2Out6[12] , \Level2Out6[11] , \Level2Out6[10] , 
        \Level2Out6[9] , \Level2Out6[8] , \Level2Out6[7] , \Level2Out6[6] , 
        \Level2Out6[5] , \Level2Out6[4] , \Level2Out6[3] , \Level2Out6[2] , 
        \Level2Out6[1] , \Level2Out6[0] }), .In1({\Level1Out6[31] , 
        \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , \Level1Out6[27] , 
        \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , \Level1Out6[23] , 
        \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , \Level1Out6[19] , 
        \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , \Level1Out6[15] , 
        \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , \Level1Out6[11] , 
        \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , \Level1Out6[7] , 
        \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , \Level1Out6[3] , 
        \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] }), .In2({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] }), 
        .Read1(\Level1Load6[0] ), .Read2(\Level1Load7[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load32[0] ), .Out({\Level16Out32[31] , \Level16Out32[30] , 
        \Level16Out32[29] , \Level16Out32[28] , \Level16Out32[27] , 
        \Level16Out32[26] , \Level16Out32[25] , \Level16Out32[24] , 
        \Level16Out32[23] , \Level16Out32[22] , \Level16Out32[21] , 
        \Level16Out32[20] , \Level16Out32[19] , \Level16Out32[18] , 
        \Level16Out32[17] , \Level16Out32[16] , \Level16Out32[15] , 
        \Level16Out32[14] , \Level16Out32[13] , \Level16Out32[12] , 
        \Level16Out32[11] , \Level16Out32[10] , \Level16Out32[9] , 
        \Level16Out32[8] , \Level16Out32[7] , \Level16Out32[6] , 
        \Level16Out32[5] , \Level16Out32[4] , \Level16Out32[3] , 
        \Level16Out32[2] , \Level16Out32[1] , \Level16Out32[0] }), .In1({
        \Level8Out32[31] , \Level8Out32[30] , \Level8Out32[29] , 
        \Level8Out32[28] , \Level8Out32[27] , \Level8Out32[26] , 
        \Level8Out32[25] , \Level8Out32[24] , \Level8Out32[23] , 
        \Level8Out32[22] , \Level8Out32[21] , \Level8Out32[20] , 
        \Level8Out32[19] , \Level8Out32[18] , \Level8Out32[17] , 
        \Level8Out32[16] , \Level8Out32[15] , \Level8Out32[14] , 
        \Level8Out32[13] , \Level8Out32[12] , \Level8Out32[11] , 
        \Level8Out32[10] , \Level8Out32[9] , \Level8Out32[8] , 
        \Level8Out32[7] , \Level8Out32[6] , \Level8Out32[5] , \Level8Out32[4] , 
        \Level8Out32[3] , \Level8Out32[2] , \Level8Out32[1] , \Level8Out32[0] 
        }), .In2({\Level8Out40[31] , \Level8Out40[30] , \Level8Out40[29] , 
        \Level8Out40[28] , \Level8Out40[27] , \Level8Out40[26] , 
        \Level8Out40[25] , \Level8Out40[24] , \Level8Out40[23] , 
        \Level8Out40[22] , \Level8Out40[21] , \Level8Out40[20] , 
        \Level8Out40[19] , \Level8Out40[18] , \Level8Out40[17] , 
        \Level8Out40[16] , \Level8Out40[15] , \Level8Out40[14] , 
        \Level8Out40[13] , \Level8Out40[12] , \Level8Out40[11] , 
        \Level8Out40[10] , \Level8Out40[9] , \Level8Out40[8] , 
        \Level8Out40[7] , \Level8Out40[6] , \Level8Out40[5] , \Level8Out40[4] , 
        \Level8Out40[3] , \Level8Out40[2] , \Level8Out40[1] , \Level8Out40[0] 
        }), .Read1(\Level8Load32[0] ), .Read2(\Level8Load40[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_120 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink120[31] , \ScanLink120[30] , 
        \ScanLink120[29] , \ScanLink120[28] , \ScanLink120[27] , 
        \ScanLink120[26] , \ScanLink120[25] , \ScanLink120[24] , 
        \ScanLink120[23] , \ScanLink120[22] , \ScanLink120[21] , 
        \ScanLink120[20] , \ScanLink120[19] , \ScanLink120[18] , 
        \ScanLink120[17] , \ScanLink120[16] , \ScanLink120[15] , 
        \ScanLink120[14] , \ScanLink120[13] , \ScanLink120[12] , 
        \ScanLink120[11] , \ScanLink120[10] , \ScanLink120[9] , 
        \ScanLink120[8] , \ScanLink120[7] , \ScanLink120[6] , \ScanLink120[5] , 
        \ScanLink120[4] , \ScanLink120[3] , \ScanLink120[2] , \ScanLink120[1] , 
        \ScanLink120[0] }), .ScanOut({\ScanLink121[31] , \ScanLink121[30] , 
        \ScanLink121[29] , \ScanLink121[28] , \ScanLink121[27] , 
        \ScanLink121[26] , \ScanLink121[25] , \ScanLink121[24] , 
        \ScanLink121[23] , \ScanLink121[22] , \ScanLink121[21] , 
        \ScanLink121[20] , \ScanLink121[19] , \ScanLink121[18] , 
        \ScanLink121[17] , \ScanLink121[16] , \ScanLink121[15] , 
        \ScanLink121[14] , \ScanLink121[13] , \ScanLink121[12] , 
        \ScanLink121[11] , \ScanLink121[10] , \ScanLink121[9] , 
        \ScanLink121[8] , \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , 
        \ScanLink121[4] , \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , 
        \ScanLink121[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load120[0] ), .Out({\Level1Out120[31] , \Level1Out120[30] , 
        \Level1Out120[29] , \Level1Out120[28] , \Level1Out120[27] , 
        \Level1Out120[26] , \Level1Out120[25] , \Level1Out120[24] , 
        \Level1Out120[23] , \Level1Out120[22] , \Level1Out120[21] , 
        \Level1Out120[20] , \Level1Out120[19] , \Level1Out120[18] , 
        \Level1Out120[17] , \Level1Out120[16] , \Level1Out120[15] , 
        \Level1Out120[14] , \Level1Out120[13] , \Level1Out120[12] , 
        \Level1Out120[11] , \Level1Out120[10] , \Level1Out120[9] , 
        \Level1Out120[8] , \Level1Out120[7] , \Level1Out120[6] , 
        \Level1Out120[5] , \Level1Out120[4] , \Level1Out120[3] , 
        \Level1Out120[2] , \Level1Out120[1] , \Level1Out120[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_128 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink128[31] , \ScanLink128[30] , 
        \ScanLink128[29] , \ScanLink128[28] , \ScanLink128[27] , 
        \ScanLink128[26] , \ScanLink128[25] , \ScanLink128[24] , 
        \ScanLink128[23] , \ScanLink128[22] , \ScanLink128[21] , 
        \ScanLink128[20] , \ScanLink128[19] , \ScanLink128[18] , 
        \ScanLink128[17] , \ScanLink128[16] , \ScanLink128[15] , 
        \ScanLink128[14] , \ScanLink128[13] , \ScanLink128[12] , 
        \ScanLink128[11] , \ScanLink128[10] , \ScanLink128[9] , 
        \ScanLink128[8] , \ScanLink128[7] , \ScanLink128[6] , \ScanLink128[5] , 
        \ScanLink128[4] , \ScanLink128[3] , \ScanLink128[2] , \ScanLink128[1] , 
        \ScanLink128[0] }), .ScanOut({\ScanLink129[31] , \ScanLink129[30] , 
        \ScanLink129[29] , \ScanLink129[28] , \ScanLink129[27] , 
        \ScanLink129[26] , \ScanLink129[25] , \ScanLink129[24] , 
        \ScanLink129[23] , \ScanLink129[22] , \ScanLink129[21] , 
        \ScanLink129[20] , \ScanLink129[19] , \ScanLink129[18] , 
        \ScanLink129[17] , \ScanLink129[16] , \ScanLink129[15] , 
        \ScanLink129[14] , \ScanLink129[13] , \ScanLink129[12] , 
        \ScanLink129[11] , \ScanLink129[10] , \ScanLink129[9] , 
        \ScanLink129[8] , \ScanLink129[7] , \ScanLink129[6] , \ScanLink129[5] , 
        \ScanLink129[4] , \ScanLink129[3] , \ScanLink129[2] , \ScanLink129[1] , 
        \ScanLink129[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load128[0] ), .Out({\Level1Out128[31] , \Level1Out128[30] , 
        \Level1Out128[29] , \Level1Out128[28] , \Level1Out128[27] , 
        \Level1Out128[26] , \Level1Out128[25] , \Level1Out128[24] , 
        \Level1Out128[23] , \Level1Out128[22] , \Level1Out128[21] , 
        \Level1Out128[20] , \Level1Out128[19] , \Level1Out128[18] , 
        \Level1Out128[17] , \Level1Out128[16] , \Level1Out128[15] , 
        \Level1Out128[14] , \Level1Out128[13] , \Level1Out128[12] , 
        \Level1Out128[11] , \Level1Out128[10] , \Level1Out128[9] , 
        \Level1Out128[8] , \Level1Out128[7] , \Level1Out128[6] , 
        \Level1Out128[5] , \Level1Out128[4] , \Level1Out128[3] , 
        \Level1Out128[2] , \Level1Out128[1] , \Level1Out128[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_184 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink184[31] , \ScanLink184[30] , 
        \ScanLink184[29] , \ScanLink184[28] , \ScanLink184[27] , 
        \ScanLink184[26] , \ScanLink184[25] , \ScanLink184[24] , 
        \ScanLink184[23] , \ScanLink184[22] , \ScanLink184[21] , 
        \ScanLink184[20] , \ScanLink184[19] , \ScanLink184[18] , 
        \ScanLink184[17] , \ScanLink184[16] , \ScanLink184[15] , 
        \ScanLink184[14] , \ScanLink184[13] , \ScanLink184[12] , 
        \ScanLink184[11] , \ScanLink184[10] , \ScanLink184[9] , 
        \ScanLink184[8] , \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , 
        \ScanLink184[4] , \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , 
        \ScanLink184[0] }), .ScanOut({\ScanLink185[31] , \ScanLink185[30] , 
        \ScanLink185[29] , \ScanLink185[28] , \ScanLink185[27] , 
        \ScanLink185[26] , \ScanLink185[25] , \ScanLink185[24] , 
        \ScanLink185[23] , \ScanLink185[22] , \ScanLink185[21] , 
        \ScanLink185[20] , \ScanLink185[19] , \ScanLink185[18] , 
        \ScanLink185[17] , \ScanLink185[16] , \ScanLink185[15] , 
        \ScanLink185[14] , \ScanLink185[13] , \ScanLink185[12] , 
        \ScanLink185[11] , \ScanLink185[10] , \ScanLink185[9] , 
        \ScanLink185[8] , \ScanLink185[7] , \ScanLink185[6] , \ScanLink185[5] , 
        \ScanLink185[4] , \ScanLink185[3] , \ScanLink185[2] , \ScanLink185[1] , 
        \ScanLink185[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load184[0] ), .Out({\Level1Out184[31] , \Level1Out184[30] , 
        \Level1Out184[29] , \Level1Out184[28] , \Level1Out184[27] , 
        \Level1Out184[26] , \Level1Out184[25] , \Level1Out184[24] , 
        \Level1Out184[23] , \Level1Out184[22] , \Level1Out184[21] , 
        \Level1Out184[20] , \Level1Out184[19] , \Level1Out184[18] , 
        \Level1Out184[17] , \Level1Out184[16] , \Level1Out184[15] , 
        \Level1Out184[14] , \Level1Out184[13] , \Level1Out184[12] , 
        \Level1Out184[11] , \Level1Out184[10] , \Level1Out184[9] , 
        \Level1Out184[8] , \Level1Out184[7] , \Level1Out184[6] , 
        \Level1Out184[5] , \Level1Out184[4] , \Level1Out184[3] , 
        \Level1Out184[2] , \Level1Out184[1] , \Level1Out184[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_210 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink210[31] , \ScanLink210[30] , 
        \ScanLink210[29] , \ScanLink210[28] , \ScanLink210[27] , 
        \ScanLink210[26] , \ScanLink210[25] , \ScanLink210[24] , 
        \ScanLink210[23] , \ScanLink210[22] , \ScanLink210[21] , 
        \ScanLink210[20] , \ScanLink210[19] , \ScanLink210[18] , 
        \ScanLink210[17] , \ScanLink210[16] , \ScanLink210[15] , 
        \ScanLink210[14] , \ScanLink210[13] , \ScanLink210[12] , 
        \ScanLink210[11] , \ScanLink210[10] , \ScanLink210[9] , 
        \ScanLink210[8] , \ScanLink210[7] , \ScanLink210[6] , \ScanLink210[5] , 
        \ScanLink210[4] , \ScanLink210[3] , \ScanLink210[2] , \ScanLink210[1] , 
        \ScanLink210[0] }), .ScanOut({\ScanLink211[31] , \ScanLink211[30] , 
        \ScanLink211[29] , \ScanLink211[28] , \ScanLink211[27] , 
        \ScanLink211[26] , \ScanLink211[25] , \ScanLink211[24] , 
        \ScanLink211[23] , \ScanLink211[22] , \ScanLink211[21] , 
        \ScanLink211[20] , \ScanLink211[19] , \ScanLink211[18] , 
        \ScanLink211[17] , \ScanLink211[16] , \ScanLink211[15] , 
        \ScanLink211[14] , \ScanLink211[13] , \ScanLink211[12] , 
        \ScanLink211[11] , \ScanLink211[10] , \ScanLink211[9] , 
        \ScanLink211[8] , \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , 
        \ScanLink211[4] , \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , 
        \ScanLink211[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load210[0] ), .Out({\Level1Out210[31] , \Level1Out210[30] , 
        \Level1Out210[29] , \Level1Out210[28] , \Level1Out210[27] , 
        \Level1Out210[26] , \Level1Out210[25] , \Level1Out210[24] , 
        \Level1Out210[23] , \Level1Out210[22] , \Level1Out210[21] , 
        \Level1Out210[20] , \Level1Out210[19] , \Level1Out210[18] , 
        \Level1Out210[17] , \Level1Out210[16] , \Level1Out210[15] , 
        \Level1Out210[14] , \Level1Out210[13] , \Level1Out210[12] , 
        \Level1Out210[11] , \Level1Out210[10] , \Level1Out210[9] , 
        \Level1Out210[8] , \Level1Out210[7] , \Level1Out210[6] , 
        \Level1Out210[5] , \Level1Out210[4] , \Level1Out210[3] , 
        \Level1Out210[2] , \Level1Out210[1] , \Level1Out210[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_218 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink218[31] , \ScanLink218[30] , 
        \ScanLink218[29] , \ScanLink218[28] , \ScanLink218[27] , 
        \ScanLink218[26] , \ScanLink218[25] , \ScanLink218[24] , 
        \ScanLink218[23] , \ScanLink218[22] , \ScanLink218[21] , 
        \ScanLink218[20] , \ScanLink218[19] , \ScanLink218[18] , 
        \ScanLink218[17] , \ScanLink218[16] , \ScanLink218[15] , 
        \ScanLink218[14] , \ScanLink218[13] , \ScanLink218[12] , 
        \ScanLink218[11] , \ScanLink218[10] , \ScanLink218[9] , 
        \ScanLink218[8] , \ScanLink218[7] , \ScanLink218[6] , \ScanLink218[5] , 
        \ScanLink218[4] , \ScanLink218[3] , \ScanLink218[2] , \ScanLink218[1] , 
        \ScanLink218[0] }), .ScanOut({\ScanLink219[31] , \ScanLink219[30] , 
        \ScanLink219[29] , \ScanLink219[28] , \ScanLink219[27] , 
        \ScanLink219[26] , \ScanLink219[25] , \ScanLink219[24] , 
        \ScanLink219[23] , \ScanLink219[22] , \ScanLink219[21] , 
        \ScanLink219[20] , \ScanLink219[19] , \ScanLink219[18] , 
        \ScanLink219[17] , \ScanLink219[16] , \ScanLink219[15] , 
        \ScanLink219[14] , \ScanLink219[13] , \ScanLink219[12] , 
        \ScanLink219[11] , \ScanLink219[10] , \ScanLink219[9] , 
        \ScanLink219[8] , \ScanLink219[7] , \ScanLink219[6] , \ScanLink219[5] , 
        \ScanLink219[4] , \ScanLink219[3] , \ScanLink219[2] , \ScanLink219[1] , 
        \ScanLink219[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load218[0] ), .Out({\Level1Out218[31] , \Level1Out218[30] , 
        \Level1Out218[29] , \Level1Out218[28] , \Level1Out218[27] , 
        \Level1Out218[26] , \Level1Out218[25] , \Level1Out218[24] , 
        \Level1Out218[23] , \Level1Out218[22] , \Level1Out218[21] , 
        \Level1Out218[20] , \Level1Out218[19] , \Level1Out218[18] , 
        \Level1Out218[17] , \Level1Out218[16] , \Level1Out218[15] , 
        \Level1Out218[14] , \Level1Out218[13] , \Level1Out218[12] , 
        \Level1Out218[11] , \Level1Out218[10] , \Level1Out218[9] , 
        \Level1Out218[8] , \Level1Out218[7] , \Level1Out218[6] , 
        \Level1Out218[5] , \Level1Out218[4] , \Level1Out218[3] , 
        \Level1Out218[2] , \Level1Out218[1] , \Level1Out218[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_146 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink146[31] , \ScanLink146[30] , 
        \ScanLink146[29] , \ScanLink146[28] , \ScanLink146[27] , 
        \ScanLink146[26] , \ScanLink146[25] , \ScanLink146[24] , 
        \ScanLink146[23] , \ScanLink146[22] , \ScanLink146[21] , 
        \ScanLink146[20] , \ScanLink146[19] , \ScanLink146[18] , 
        \ScanLink146[17] , \ScanLink146[16] , \ScanLink146[15] , 
        \ScanLink146[14] , \ScanLink146[13] , \ScanLink146[12] , 
        \ScanLink146[11] , \ScanLink146[10] , \ScanLink146[9] , 
        \ScanLink146[8] , \ScanLink146[7] , \ScanLink146[6] , \ScanLink146[5] , 
        \ScanLink146[4] , \ScanLink146[3] , \ScanLink146[2] , \ScanLink146[1] , 
        \ScanLink146[0] }), .ScanOut({\ScanLink147[31] , \ScanLink147[30] , 
        \ScanLink147[29] , \ScanLink147[28] , \ScanLink147[27] , 
        \ScanLink147[26] , \ScanLink147[25] , \ScanLink147[24] , 
        \ScanLink147[23] , \ScanLink147[22] , \ScanLink147[21] , 
        \ScanLink147[20] , \ScanLink147[19] , \ScanLink147[18] , 
        \ScanLink147[17] , \ScanLink147[16] , \ScanLink147[15] , 
        \ScanLink147[14] , \ScanLink147[13] , \ScanLink147[12] , 
        \ScanLink147[11] , \ScanLink147[10] , \ScanLink147[9] , 
        \ScanLink147[8] , \ScanLink147[7] , \ScanLink147[6] , \ScanLink147[5] , 
        \ScanLink147[4] , \ScanLink147[3] , \ScanLink147[2] , \ScanLink147[1] , 
        \ScanLink147[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load146[0] ), .Out({\Level1Out146[31] , \Level1Out146[30] , 
        \Level1Out146[29] , \Level1Out146[28] , \Level1Out146[27] , 
        \Level1Out146[26] , \Level1Out146[25] , \Level1Out146[24] , 
        \Level1Out146[23] , \Level1Out146[22] , \Level1Out146[21] , 
        \Level1Out146[20] , \Level1Out146[19] , \Level1Out146[18] , 
        \Level1Out146[17] , \Level1Out146[16] , \Level1Out146[15] , 
        \Level1Out146[14] , \Level1Out146[13] , \Level1Out146[12] , 
        \Level1Out146[11] , \Level1Out146[10] , \Level1Out146[9] , 
        \Level1Out146[8] , \Level1Out146[7] , \Level1Out146[6] , 
        \Level1Out146[5] , \Level1Out146[4] , \Level1Out146[3] , 
        \Level1Out146[2] , \Level1Out146[1] , \Level1Out146[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_161 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink161[31] , \ScanLink161[30] , 
        \ScanLink161[29] , \ScanLink161[28] , \ScanLink161[27] , 
        \ScanLink161[26] , \ScanLink161[25] , \ScanLink161[24] , 
        \ScanLink161[23] , \ScanLink161[22] , \ScanLink161[21] , 
        \ScanLink161[20] , \ScanLink161[19] , \ScanLink161[18] , 
        \ScanLink161[17] , \ScanLink161[16] , \ScanLink161[15] , 
        \ScanLink161[14] , \ScanLink161[13] , \ScanLink161[12] , 
        \ScanLink161[11] , \ScanLink161[10] , \ScanLink161[9] , 
        \ScanLink161[8] , \ScanLink161[7] , \ScanLink161[6] , \ScanLink161[5] , 
        \ScanLink161[4] , \ScanLink161[3] , \ScanLink161[2] , \ScanLink161[1] , 
        \ScanLink161[0] }), .ScanOut({\ScanLink162[31] , \ScanLink162[30] , 
        \ScanLink162[29] , \ScanLink162[28] , \ScanLink162[27] , 
        \ScanLink162[26] , \ScanLink162[25] , \ScanLink162[24] , 
        \ScanLink162[23] , \ScanLink162[22] , \ScanLink162[21] , 
        \ScanLink162[20] , \ScanLink162[19] , \ScanLink162[18] , 
        \ScanLink162[17] , \ScanLink162[16] , \ScanLink162[15] , 
        \ScanLink162[14] , \ScanLink162[13] , \ScanLink162[12] , 
        \ScanLink162[11] , \ScanLink162[10] , \ScanLink162[9] , 
        \ScanLink162[8] , \ScanLink162[7] , \ScanLink162[6] , \ScanLink162[5] , 
        \ScanLink162[4] , \ScanLink162[3] , \ScanLink162[2] , \ScanLink162[1] , 
        \ScanLink162[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load161[0] ), .Out({\Level1Out161[31] , \Level1Out161[30] , 
        \Level1Out161[29] , \Level1Out161[28] , \Level1Out161[27] , 
        \Level1Out161[26] , \Level1Out161[25] , \Level1Out161[24] , 
        \Level1Out161[23] , \Level1Out161[22] , \Level1Out161[21] , 
        \Level1Out161[20] , \Level1Out161[19] , \Level1Out161[18] , 
        \Level1Out161[17] , \Level1Out161[16] , \Level1Out161[15] , 
        \Level1Out161[14] , \Level1Out161[13] , \Level1Out161[12] , 
        \Level1Out161[11] , \Level1Out161[10] , \Level1Out161[9] , 
        \Level1Out161[8] , \Level1Out161[7] , \Level1Out161[6] , 
        \Level1Out161[5] , \Level1Out161[4] , \Level1Out161[3] , 
        \Level1Out161[2] , \Level1Out161[1] , \Level1Out161[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_158_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load158[0] ), .Out({\Level2Out158[31] , \Level2Out158[30] , 
        \Level2Out158[29] , \Level2Out158[28] , \Level2Out158[27] , 
        \Level2Out158[26] , \Level2Out158[25] , \Level2Out158[24] , 
        \Level2Out158[23] , \Level2Out158[22] , \Level2Out158[21] , 
        \Level2Out158[20] , \Level2Out158[19] , \Level2Out158[18] , 
        \Level2Out158[17] , \Level2Out158[16] , \Level2Out158[15] , 
        \Level2Out158[14] , \Level2Out158[13] , \Level2Out158[12] , 
        \Level2Out158[11] , \Level2Out158[10] , \Level2Out158[9] , 
        \Level2Out158[8] , \Level2Out158[7] , \Level2Out158[6] , 
        \Level2Out158[5] , \Level2Out158[4] , \Level2Out158[3] , 
        \Level2Out158[2] , \Level2Out158[1] , \Level2Out158[0] }), .In1({
        \Level1Out158[31] , \Level1Out158[30] , \Level1Out158[29] , 
        \Level1Out158[28] , \Level1Out158[27] , \Level1Out158[26] , 
        \Level1Out158[25] , \Level1Out158[24] , \Level1Out158[23] , 
        \Level1Out158[22] , \Level1Out158[21] , \Level1Out158[20] , 
        \Level1Out158[19] , \Level1Out158[18] , \Level1Out158[17] , 
        \Level1Out158[16] , \Level1Out158[15] , \Level1Out158[14] , 
        \Level1Out158[13] , \Level1Out158[12] , \Level1Out158[11] , 
        \Level1Out158[10] , \Level1Out158[9] , \Level1Out158[8] , 
        \Level1Out158[7] , \Level1Out158[6] , \Level1Out158[5] , 
        \Level1Out158[4] , \Level1Out158[3] , \Level1Out158[2] , 
        \Level1Out158[1] , \Level1Out158[0] }), .In2({\Level1Out159[31] , 
        \Level1Out159[30] , \Level1Out159[29] , \Level1Out159[28] , 
        \Level1Out159[27] , \Level1Out159[26] , \Level1Out159[25] , 
        \Level1Out159[24] , \Level1Out159[23] , \Level1Out159[22] , 
        \Level1Out159[21] , \Level1Out159[20] , \Level1Out159[19] , 
        \Level1Out159[18] , \Level1Out159[17] , \Level1Out159[16] , 
        \Level1Out159[15] , \Level1Out159[14] , \Level1Out159[13] , 
        \Level1Out159[12] , \Level1Out159[11] , \Level1Out159[10] , 
        \Level1Out159[9] , \Level1Out159[8] , \Level1Out159[7] , 
        \Level1Out159[6] , \Level1Out159[5] , \Level1Out159[4] , 
        \Level1Out159[3] , \Level1Out159[2] , \Level1Out159[1] , 
        \Level1Out159[0] }), .Read1(\Level1Load158[0] ), .Read2(
        \Level1Load159[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_144_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load144[0] ), .Out({\Level4Out144[31] , \Level4Out144[30] , 
        \Level4Out144[29] , \Level4Out144[28] , \Level4Out144[27] , 
        \Level4Out144[26] , \Level4Out144[25] , \Level4Out144[24] , 
        \Level4Out144[23] , \Level4Out144[22] , \Level4Out144[21] , 
        \Level4Out144[20] , \Level4Out144[19] , \Level4Out144[18] , 
        \Level4Out144[17] , \Level4Out144[16] , \Level4Out144[15] , 
        \Level4Out144[14] , \Level4Out144[13] , \Level4Out144[12] , 
        \Level4Out144[11] , \Level4Out144[10] , \Level4Out144[9] , 
        \Level4Out144[8] , \Level4Out144[7] , \Level4Out144[6] , 
        \Level4Out144[5] , \Level4Out144[4] , \Level4Out144[3] , 
        \Level4Out144[2] , \Level4Out144[1] , \Level4Out144[0] }), .In1({
        \Level2Out144[31] , \Level2Out144[30] , \Level2Out144[29] , 
        \Level2Out144[28] , \Level2Out144[27] , \Level2Out144[26] , 
        \Level2Out144[25] , \Level2Out144[24] , \Level2Out144[23] , 
        \Level2Out144[22] , \Level2Out144[21] , \Level2Out144[20] , 
        \Level2Out144[19] , \Level2Out144[18] , \Level2Out144[17] , 
        \Level2Out144[16] , \Level2Out144[15] , \Level2Out144[14] , 
        \Level2Out144[13] , \Level2Out144[12] , \Level2Out144[11] , 
        \Level2Out144[10] , \Level2Out144[9] , \Level2Out144[8] , 
        \Level2Out144[7] , \Level2Out144[6] , \Level2Out144[5] , 
        \Level2Out144[4] , \Level2Out144[3] , \Level2Out144[2] , 
        \Level2Out144[1] , \Level2Out144[0] }), .In2({\Level2Out146[31] , 
        \Level2Out146[30] , \Level2Out146[29] , \Level2Out146[28] , 
        \Level2Out146[27] , \Level2Out146[26] , \Level2Out146[25] , 
        \Level2Out146[24] , \Level2Out146[23] , \Level2Out146[22] , 
        \Level2Out146[21] , \Level2Out146[20] , \Level2Out146[19] , 
        \Level2Out146[18] , \Level2Out146[17] , \Level2Out146[16] , 
        \Level2Out146[15] , \Level2Out146[14] , \Level2Out146[13] , 
        \Level2Out146[12] , \Level2Out146[11] , \Level2Out146[10] , 
        \Level2Out146[9] , \Level2Out146[8] , \Level2Out146[7] , 
        \Level2Out146[6] , \Level2Out146[5] , \Level2Out146[4] , 
        \Level2Out146[3] , \Level2Out146[2] , \Level2Out146[1] , 
        \Level2Out146[0] }), .Read1(\Level2Load144[0] ), .Read2(
        \Level2Load146[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_246_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load246[0] ), .Out({\Level2Out246[31] , \Level2Out246[30] , 
        \Level2Out246[29] , \Level2Out246[28] , \Level2Out246[27] , 
        \Level2Out246[26] , \Level2Out246[25] , \Level2Out246[24] , 
        \Level2Out246[23] , \Level2Out246[22] , \Level2Out246[21] , 
        \Level2Out246[20] , \Level2Out246[19] , \Level2Out246[18] , 
        \Level2Out246[17] , \Level2Out246[16] , \Level2Out246[15] , 
        \Level2Out246[14] , \Level2Out246[13] , \Level2Out246[12] , 
        \Level2Out246[11] , \Level2Out246[10] , \Level2Out246[9] , 
        \Level2Out246[8] , \Level2Out246[7] , \Level2Out246[6] , 
        \Level2Out246[5] , \Level2Out246[4] , \Level2Out246[3] , 
        \Level2Out246[2] , \Level2Out246[1] , \Level2Out246[0] }), .In1({
        \Level1Out246[31] , \Level1Out246[30] , \Level1Out246[29] , 
        \Level1Out246[28] , \Level1Out246[27] , \Level1Out246[26] , 
        \Level1Out246[25] , \Level1Out246[24] , \Level1Out246[23] , 
        \Level1Out246[22] , \Level1Out246[21] , \Level1Out246[20] , 
        \Level1Out246[19] , \Level1Out246[18] , \Level1Out246[17] , 
        \Level1Out246[16] , \Level1Out246[15] , \Level1Out246[14] , 
        \Level1Out246[13] , \Level1Out246[12] , \Level1Out246[11] , 
        \Level1Out246[10] , \Level1Out246[9] , \Level1Out246[8] , 
        \Level1Out246[7] , \Level1Out246[6] , \Level1Out246[5] , 
        \Level1Out246[4] , \Level1Out246[3] , \Level1Out246[2] , 
        \Level1Out246[1] , \Level1Out246[0] }), .In2({\Level1Out247[31] , 
        \Level1Out247[30] , \Level1Out247[29] , \Level1Out247[28] , 
        \Level1Out247[27] , \Level1Out247[26] , \Level1Out247[25] , 
        \Level1Out247[24] , \Level1Out247[23] , \Level1Out247[22] , 
        \Level1Out247[21] , \Level1Out247[20] , \Level1Out247[19] , 
        \Level1Out247[18] , \Level1Out247[17] , \Level1Out247[16] , 
        \Level1Out247[15] , \Level1Out247[14] , \Level1Out247[13] , 
        \Level1Out247[12] , \Level1Out247[11] , \Level1Out247[10] , 
        \Level1Out247[9] , \Level1Out247[8] , \Level1Out247[7] , 
        \Level1Out247[6] , \Level1Out247[5] , \Level1Out247[4] , 
        \Level1Out247[3] , \Level1Out247[2] , \Level1Out247[1] , 
        \Level1Out247[0] }), .Read1(\Level1Load246[0] ), .Read2(
        \Level1Load247[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_251 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink251[31] , \ScanLink251[30] , 
        \ScanLink251[29] , \ScanLink251[28] , \ScanLink251[27] , 
        \ScanLink251[26] , \ScanLink251[25] , \ScanLink251[24] , 
        \ScanLink251[23] , \ScanLink251[22] , \ScanLink251[21] , 
        \ScanLink251[20] , \ScanLink251[19] , \ScanLink251[18] , 
        \ScanLink251[17] , \ScanLink251[16] , \ScanLink251[15] , 
        \ScanLink251[14] , \ScanLink251[13] , \ScanLink251[12] , 
        \ScanLink251[11] , \ScanLink251[10] , \ScanLink251[9] , 
        \ScanLink251[8] , \ScanLink251[7] , \ScanLink251[6] , \ScanLink251[5] , 
        \ScanLink251[4] , \ScanLink251[3] , \ScanLink251[2] , \ScanLink251[1] , 
        \ScanLink251[0] }), .ScanOut({\ScanLink252[31] , \ScanLink252[30] , 
        \ScanLink252[29] , \ScanLink252[28] , \ScanLink252[27] , 
        \ScanLink252[26] , \ScanLink252[25] , \ScanLink252[24] , 
        \ScanLink252[23] , \ScanLink252[22] , \ScanLink252[21] , 
        \ScanLink252[20] , \ScanLink252[19] , \ScanLink252[18] , 
        \ScanLink252[17] , \ScanLink252[16] , \ScanLink252[15] , 
        \ScanLink252[14] , \ScanLink252[13] , \ScanLink252[12] , 
        \ScanLink252[11] , \ScanLink252[10] , \ScanLink252[9] , 
        \ScanLink252[8] , \ScanLink252[7] , \ScanLink252[6] , \ScanLink252[5] , 
        \ScanLink252[4] , \ScanLink252[3] , \ScanLink252[2] , \ScanLink252[1] , 
        \ScanLink252[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load251[0] ), .Out({\Level1Out251[31] , \Level1Out251[30] , 
        \Level1Out251[29] , \Level1Out251[28] , \Level1Out251[27] , 
        \Level1Out251[26] , \Level1Out251[25] , \Level1Out251[24] , 
        \Level1Out251[23] , \Level1Out251[22] , \Level1Out251[21] , 
        \Level1Out251[20] , \Level1Out251[19] , \Level1Out251[18] , 
        \Level1Out251[17] , \Level1Out251[16] , \Level1Out251[15] , 
        \Level1Out251[14] , \Level1Out251[13] , \Level1Out251[12] , 
        \Level1Out251[11] , \Level1Out251[10] , \Level1Out251[9] , 
        \Level1Out251[8] , \Level1Out251[7] , \Level1Out251[6] , 
        \Level1Out251[5] , \Level1Out251[4] , \Level1Out251[3] , 
        \Level1Out251[2] , \Level1Out251[1] , \Level1Out251[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_34_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load34[0] ), .Out({\Level2Out34[31] , \Level2Out34[30] , 
        \Level2Out34[29] , \Level2Out34[28] , \Level2Out34[27] , 
        \Level2Out34[26] , \Level2Out34[25] , \Level2Out34[24] , 
        \Level2Out34[23] , \Level2Out34[22] , \Level2Out34[21] , 
        \Level2Out34[20] , \Level2Out34[19] , \Level2Out34[18] , 
        \Level2Out34[17] , \Level2Out34[16] , \Level2Out34[15] , 
        \Level2Out34[14] , \Level2Out34[13] , \Level2Out34[12] , 
        \Level2Out34[11] , \Level2Out34[10] , \Level2Out34[9] , 
        \Level2Out34[8] , \Level2Out34[7] , \Level2Out34[6] , \Level2Out34[5] , 
        \Level2Out34[4] , \Level2Out34[3] , \Level2Out34[2] , \Level2Out34[1] , 
        \Level2Out34[0] }), .In1({\Level1Out34[31] , \Level1Out34[30] , 
        \Level1Out34[29] , \Level1Out34[28] , \Level1Out34[27] , 
        \Level1Out34[26] , \Level1Out34[25] , \Level1Out34[24] , 
        \Level1Out34[23] , \Level1Out34[22] , \Level1Out34[21] , 
        \Level1Out34[20] , \Level1Out34[19] , \Level1Out34[18] , 
        \Level1Out34[17] , \Level1Out34[16] , \Level1Out34[15] , 
        \Level1Out34[14] , \Level1Out34[13] , \Level1Out34[12] , 
        \Level1Out34[11] , \Level1Out34[10] , \Level1Out34[9] , 
        \Level1Out34[8] , \Level1Out34[7] , \Level1Out34[6] , \Level1Out34[5] , 
        \Level1Out34[4] , \Level1Out34[3] , \Level1Out34[2] , \Level1Out34[1] , 
        \Level1Out34[0] }), .In2({\Level1Out35[31] , \Level1Out35[30] , 
        \Level1Out35[29] , \Level1Out35[28] , \Level1Out35[27] , 
        \Level1Out35[26] , \Level1Out35[25] , \Level1Out35[24] , 
        \Level1Out35[23] , \Level1Out35[22] , \Level1Out35[21] , 
        \Level1Out35[20] , \Level1Out35[19] , \Level1Out35[18] , 
        \Level1Out35[17] , \Level1Out35[16] , \Level1Out35[15] , 
        \Level1Out35[14] , \Level1Out35[13] , \Level1Out35[12] , 
        \Level1Out35[11] , \Level1Out35[10] , \Level1Out35[9] , 
        \Level1Out35[8] , \Level1Out35[7] , \Level1Out35[6] , \Level1Out35[5] , 
        \Level1Out35[4] , \Level1Out35[3] , \Level1Out35[2] , \Level1Out35[1] , 
        \Level1Out35[0] }), .Read1(\Level1Load34[0] ), .Read2(
        \Level1Load35[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_96_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load96[0] ), .Out({\Level8Out96[31] , \Level8Out96[30] , 
        \Level8Out96[29] , \Level8Out96[28] , \Level8Out96[27] , 
        \Level8Out96[26] , \Level8Out96[25] , \Level8Out96[24] , 
        \Level8Out96[23] , \Level8Out96[22] , \Level8Out96[21] , 
        \Level8Out96[20] , \Level8Out96[19] , \Level8Out96[18] , 
        \Level8Out96[17] , \Level8Out96[16] , \Level8Out96[15] , 
        \Level8Out96[14] , \Level8Out96[13] , \Level8Out96[12] , 
        \Level8Out96[11] , \Level8Out96[10] , \Level8Out96[9] , 
        \Level8Out96[8] , \Level8Out96[7] , \Level8Out96[6] , \Level8Out96[5] , 
        \Level8Out96[4] , \Level8Out96[3] , \Level8Out96[2] , \Level8Out96[1] , 
        \Level8Out96[0] }), .In1({\Level4Out96[31] , \Level4Out96[30] , 
        \Level4Out96[29] , \Level4Out96[28] , \Level4Out96[27] , 
        \Level4Out96[26] , \Level4Out96[25] , \Level4Out96[24] , 
        \Level4Out96[23] , \Level4Out96[22] , \Level4Out96[21] , 
        \Level4Out96[20] , \Level4Out96[19] , \Level4Out96[18] , 
        \Level4Out96[17] , \Level4Out96[16] , \Level4Out96[15] , 
        \Level4Out96[14] , \Level4Out96[13] , \Level4Out96[12] , 
        \Level4Out96[11] , \Level4Out96[10] , \Level4Out96[9] , 
        \Level4Out96[8] , \Level4Out96[7] , \Level4Out96[6] , \Level4Out96[5] , 
        \Level4Out96[4] , \Level4Out96[3] , \Level4Out96[2] , \Level4Out96[1] , 
        \Level4Out96[0] }), .In2({\Level4Out100[31] , \Level4Out100[30] , 
        \Level4Out100[29] , \Level4Out100[28] , \Level4Out100[27] , 
        \Level4Out100[26] , \Level4Out100[25] , \Level4Out100[24] , 
        \Level4Out100[23] , \Level4Out100[22] , \Level4Out100[21] , 
        \Level4Out100[20] , \Level4Out100[19] , \Level4Out100[18] , 
        \Level4Out100[17] , \Level4Out100[16] , \Level4Out100[15] , 
        \Level4Out100[14] , \Level4Out100[13] , \Level4Out100[12] , 
        \Level4Out100[11] , \Level4Out100[10] , \Level4Out100[9] , 
        \Level4Out100[8] , \Level4Out100[7] , \Level4Out100[6] , 
        \Level4Out100[5] , \Level4Out100[4] , \Level4Out100[3] , 
        \Level4Out100[2] , \Level4Out100[1] , \Level4Out100[0] }), .Read1(
        \Level4Load96[0] ), .Read2(\Level4Load100[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_28_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load28[0] ), .Out({\Level4Out28[31] , \Level4Out28[30] , 
        \Level4Out28[29] , \Level4Out28[28] , \Level4Out28[27] , 
        \Level4Out28[26] , \Level4Out28[25] , \Level4Out28[24] , 
        \Level4Out28[23] , \Level4Out28[22] , \Level4Out28[21] , 
        \Level4Out28[20] , \Level4Out28[19] , \Level4Out28[18] , 
        \Level4Out28[17] , \Level4Out28[16] , \Level4Out28[15] , 
        \Level4Out28[14] , \Level4Out28[13] , \Level4Out28[12] , 
        \Level4Out28[11] , \Level4Out28[10] , \Level4Out28[9] , 
        \Level4Out28[8] , \Level4Out28[7] , \Level4Out28[6] , \Level4Out28[5] , 
        \Level4Out28[4] , \Level4Out28[3] , \Level4Out28[2] , \Level4Out28[1] , 
        \Level4Out28[0] }), .In1({\Level2Out28[31] , \Level2Out28[30] , 
        \Level2Out28[29] , \Level2Out28[28] , \Level2Out28[27] , 
        \Level2Out28[26] , \Level2Out28[25] , \Level2Out28[24] , 
        \Level2Out28[23] , \Level2Out28[22] , \Level2Out28[21] , 
        \Level2Out28[20] , \Level2Out28[19] , \Level2Out28[18] , 
        \Level2Out28[17] , \Level2Out28[16] , \Level2Out28[15] , 
        \Level2Out28[14] , \Level2Out28[13] , \Level2Out28[12] , 
        \Level2Out28[11] , \Level2Out28[10] , \Level2Out28[9] , 
        \Level2Out28[8] , \Level2Out28[7] , \Level2Out28[6] , \Level2Out28[5] , 
        \Level2Out28[4] , \Level2Out28[3] , \Level2Out28[2] , \Level2Out28[1] , 
        \Level2Out28[0] }), .In2({\Level2Out30[31] , \Level2Out30[30] , 
        \Level2Out30[29] , \Level2Out30[28] , \Level2Out30[27] , 
        \Level2Out30[26] , \Level2Out30[25] , \Level2Out30[24] , 
        \Level2Out30[23] , \Level2Out30[22] , \Level2Out30[21] , 
        \Level2Out30[20] , \Level2Out30[19] , \Level2Out30[18] , 
        \Level2Out30[17] , \Level2Out30[16] , \Level2Out30[15] , 
        \Level2Out30[14] , \Level2Out30[13] , \Level2Out30[12] , 
        \Level2Out30[11] , \Level2Out30[10] , \Level2Out30[9] , 
        \Level2Out30[8] , \Level2Out30[7] , \Level2Out30[6] , \Level2Out30[5] , 
        \Level2Out30[4] , \Level2Out30[3] , \Level2Out30[2] , \Level2Out30[1] , 
        \Level2Out30[0] }), .Read1(\Level2Load28[0] ), .Read2(
        \Level2Load30[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_172_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load172[0] ), .Out({\Level2Out172[31] , \Level2Out172[30] , 
        \Level2Out172[29] , \Level2Out172[28] , \Level2Out172[27] , 
        \Level2Out172[26] , \Level2Out172[25] , \Level2Out172[24] , 
        \Level2Out172[23] , \Level2Out172[22] , \Level2Out172[21] , 
        \Level2Out172[20] , \Level2Out172[19] , \Level2Out172[18] , 
        \Level2Out172[17] , \Level2Out172[16] , \Level2Out172[15] , 
        \Level2Out172[14] , \Level2Out172[13] , \Level2Out172[12] , 
        \Level2Out172[11] , \Level2Out172[10] , \Level2Out172[9] , 
        \Level2Out172[8] , \Level2Out172[7] , \Level2Out172[6] , 
        \Level2Out172[5] , \Level2Out172[4] , \Level2Out172[3] , 
        \Level2Out172[2] , \Level2Out172[1] , \Level2Out172[0] }), .In1({
        \Level1Out172[31] , \Level1Out172[30] , \Level1Out172[29] , 
        \Level1Out172[28] , \Level1Out172[27] , \Level1Out172[26] , 
        \Level1Out172[25] , \Level1Out172[24] , \Level1Out172[23] , 
        \Level1Out172[22] , \Level1Out172[21] , \Level1Out172[20] , 
        \Level1Out172[19] , \Level1Out172[18] , \Level1Out172[17] , 
        \Level1Out172[16] , \Level1Out172[15] , \Level1Out172[14] , 
        \Level1Out172[13] , \Level1Out172[12] , \Level1Out172[11] , 
        \Level1Out172[10] , \Level1Out172[9] , \Level1Out172[8] , 
        \Level1Out172[7] , \Level1Out172[6] , \Level1Out172[5] , 
        \Level1Out172[4] , \Level1Out172[3] , \Level1Out172[2] , 
        \Level1Out172[1] , \Level1Out172[0] }), .In2({\Level1Out173[31] , 
        \Level1Out173[30] , \Level1Out173[29] , \Level1Out173[28] , 
        \Level1Out173[27] , \Level1Out173[26] , \Level1Out173[25] , 
        \Level1Out173[24] , \Level1Out173[23] , \Level1Out173[22] , 
        \Level1Out173[21] , \Level1Out173[20] , \Level1Out173[19] , 
        \Level1Out173[18] , \Level1Out173[17] , \Level1Out173[16] , 
        \Level1Out173[15] , \Level1Out173[14] , \Level1Out173[13] , 
        \Level1Out173[12] , \Level1Out173[11] , \Level1Out173[10] , 
        \Level1Out173[9] , \Level1Out173[8] , \Level1Out173[7] , 
        \Level1Out173[6] , \Level1Out173[5] , \Level1Out173[4] , 
        \Level1Out173[3] , \Level1Out173[2] , \Level1Out173[1] , 
        \Level1Out173[0] }), .Read1(\Level1Load172[0] ), .Read2(
        \Level1Load173[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_88_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load88[0] ), .Out({\Level2Out88[31] , \Level2Out88[30] , 
        \Level2Out88[29] , \Level2Out88[28] , \Level2Out88[27] , 
        \Level2Out88[26] , \Level2Out88[25] , \Level2Out88[24] , 
        \Level2Out88[23] , \Level2Out88[22] , \Level2Out88[21] , 
        \Level2Out88[20] , \Level2Out88[19] , \Level2Out88[18] , 
        \Level2Out88[17] , \Level2Out88[16] , \Level2Out88[15] , 
        \Level2Out88[14] , \Level2Out88[13] , \Level2Out88[12] , 
        \Level2Out88[11] , \Level2Out88[10] , \Level2Out88[9] , 
        \Level2Out88[8] , \Level2Out88[7] , \Level2Out88[6] , \Level2Out88[5] , 
        \Level2Out88[4] , \Level2Out88[3] , \Level2Out88[2] , \Level2Out88[1] , 
        \Level2Out88[0] }), .In1({\Level1Out88[31] , \Level1Out88[30] , 
        \Level1Out88[29] , \Level1Out88[28] , \Level1Out88[27] , 
        \Level1Out88[26] , \Level1Out88[25] , \Level1Out88[24] , 
        \Level1Out88[23] , \Level1Out88[22] , \Level1Out88[21] , 
        \Level1Out88[20] , \Level1Out88[19] , \Level1Out88[18] , 
        \Level1Out88[17] , \Level1Out88[16] , \Level1Out88[15] , 
        \Level1Out88[14] , \Level1Out88[13] , \Level1Out88[12] , 
        \Level1Out88[11] , \Level1Out88[10] , \Level1Out88[9] , 
        \Level1Out88[8] , \Level1Out88[7] , \Level1Out88[6] , \Level1Out88[5] , 
        \Level1Out88[4] , \Level1Out88[3] , \Level1Out88[2] , \Level1Out88[1] , 
        \Level1Out88[0] }), .In2({\Level1Out89[31] , \Level1Out89[30] , 
        \Level1Out89[29] , \Level1Out89[28] , \Level1Out89[27] , 
        \Level1Out89[26] , \Level1Out89[25] , \Level1Out89[24] , 
        \Level1Out89[23] , \Level1Out89[22] , \Level1Out89[21] , 
        \Level1Out89[20] , \Level1Out89[19] , \Level1Out89[18] , 
        \Level1Out89[17] , \Level1Out89[16] , \Level1Out89[15] , 
        \Level1Out89[14] , \Level1Out89[13] , \Level1Out89[12] , 
        \Level1Out89[11] , \Level1Out89[10] , \Level1Out89[9] , 
        \Level1Out89[8] , \Level1Out89[7] , \Level1Out89[6] , \Level1Out89[5] , 
        \Level1Out89[4] , \Level1Out89[3] , \Level1Out89[2] , \Level1Out89[1] , 
        \Level1Out89[0] }), .Read1(\Level1Load88[0] ), .Read2(
        \Level1Load89[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_58 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanOut({\ScanLink59[31] , 
        \ScanLink59[30] , \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , 
        \ScanLink59[26] , \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , 
        \ScanLink59[22] , \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , 
        \ScanLink59[18] , \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , 
        \ScanLink59[14] , \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , 
        \ScanLink59[10] , \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , 
        \ScanLink59[6] , \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , 
        \ScanLink59[2] , \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load58[0] ), .Out({
        \Level1Out58[31] , \Level1Out58[30] , \Level1Out58[29] , 
        \Level1Out58[28] , \Level1Out58[27] , \Level1Out58[26] , 
        \Level1Out58[25] , \Level1Out58[24] , \Level1Out58[23] , 
        \Level1Out58[22] , \Level1Out58[21] , \Level1Out58[20] , 
        \Level1Out58[19] , \Level1Out58[18] , \Level1Out58[17] , 
        \Level1Out58[16] , \Level1Out58[15] , \Level1Out58[14] , 
        \Level1Out58[13] , \Level1Out58[12] , \Level1Out58[11] , 
        \Level1Out58[10] , \Level1Out58[9] , \Level1Out58[8] , 
        \Level1Out58[7] , \Level1Out58[6] , \Level1Out58[5] , \Level1Out58[4] , 
        \Level1Out58[3] , \Level1Out58[2] , \Level1Out58[1] , \Level1Out58[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_114 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink114[31] , \ScanLink114[30] , 
        \ScanLink114[29] , \ScanLink114[28] , \ScanLink114[27] , 
        \ScanLink114[26] , \ScanLink114[25] , \ScanLink114[24] , 
        \ScanLink114[23] , \ScanLink114[22] , \ScanLink114[21] , 
        \ScanLink114[20] , \ScanLink114[19] , \ScanLink114[18] , 
        \ScanLink114[17] , \ScanLink114[16] , \ScanLink114[15] , 
        \ScanLink114[14] , \ScanLink114[13] , \ScanLink114[12] , 
        \ScanLink114[11] , \ScanLink114[10] , \ScanLink114[9] , 
        \ScanLink114[8] , \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , 
        \ScanLink114[4] , \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , 
        \ScanLink114[0] }), .ScanOut({\ScanLink115[31] , \ScanLink115[30] , 
        \ScanLink115[29] , \ScanLink115[28] , \ScanLink115[27] , 
        \ScanLink115[26] , \ScanLink115[25] , \ScanLink115[24] , 
        \ScanLink115[23] , \ScanLink115[22] , \ScanLink115[21] , 
        \ScanLink115[20] , \ScanLink115[19] , \ScanLink115[18] , 
        \ScanLink115[17] , \ScanLink115[16] , \ScanLink115[15] , 
        \ScanLink115[14] , \ScanLink115[13] , \ScanLink115[12] , 
        \ScanLink115[11] , \ScanLink115[10] , \ScanLink115[9] , 
        \ScanLink115[8] , \ScanLink115[7] , \ScanLink115[6] , \ScanLink115[5] , 
        \ScanLink115[4] , \ScanLink115[3] , \ScanLink115[2] , \ScanLink115[1] , 
        \ScanLink115[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load114[0] ), .Out({\Level1Out114[31] , \Level1Out114[30] , 
        \Level1Out114[29] , \Level1Out114[28] , \Level1Out114[27] , 
        \Level1Out114[26] , \Level1Out114[25] , \Level1Out114[24] , 
        \Level1Out114[23] , \Level1Out114[22] , \Level1Out114[21] , 
        \Level1Out114[20] , \Level1Out114[19] , \Level1Out114[18] , 
        \Level1Out114[17] , \Level1Out114[16] , \Level1Out114[15] , 
        \Level1Out114[14] , \Level1Out114[13] , \Level1Out114[12] , 
        \Level1Out114[11] , \Level1Out114[10] , \Level1Out114[9] , 
        \Level1Out114[8] , \Level1Out114[7] , \Level1Out114[6] , 
        \Level1Out114[5] , \Level1Out114[4] , \Level1Out114[3] , 
        \Level1Out114[2] , \Level1Out114[1] , \Level1Out114[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_224 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink224[31] , \ScanLink224[30] , 
        \ScanLink224[29] , \ScanLink224[28] , \ScanLink224[27] , 
        \ScanLink224[26] , \ScanLink224[25] , \ScanLink224[24] , 
        \ScanLink224[23] , \ScanLink224[22] , \ScanLink224[21] , 
        \ScanLink224[20] , \ScanLink224[19] , \ScanLink224[18] , 
        \ScanLink224[17] , \ScanLink224[16] , \ScanLink224[15] , 
        \ScanLink224[14] , \ScanLink224[13] , \ScanLink224[12] , 
        \ScanLink224[11] , \ScanLink224[10] , \ScanLink224[9] , 
        \ScanLink224[8] , \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , 
        \ScanLink224[4] , \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , 
        \ScanLink224[0] }), .ScanOut({\ScanLink225[31] , \ScanLink225[30] , 
        \ScanLink225[29] , \ScanLink225[28] , \ScanLink225[27] , 
        \ScanLink225[26] , \ScanLink225[25] , \ScanLink225[24] , 
        \ScanLink225[23] , \ScanLink225[22] , \ScanLink225[21] , 
        \ScanLink225[20] , \ScanLink225[19] , \ScanLink225[18] , 
        \ScanLink225[17] , \ScanLink225[16] , \ScanLink225[15] , 
        \ScanLink225[14] , \ScanLink225[13] , \ScanLink225[12] , 
        \ScanLink225[11] , \ScanLink225[10] , \ScanLink225[9] , 
        \ScanLink225[8] , \ScanLink225[7] , \ScanLink225[6] , \ScanLink225[5] , 
        \ScanLink225[4] , \ScanLink225[3] , \ScanLink225[2] , \ScanLink225[1] , 
        \ScanLink225[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load224[0] ), .Out({\Level1Out224[31] , \Level1Out224[30] , 
        \Level1Out224[29] , \Level1Out224[28] , \Level1Out224[27] , 
        \Level1Out224[26] , \Level1Out224[25] , \Level1Out224[24] , 
        \Level1Out224[23] , \Level1Out224[22] , \Level1Out224[21] , 
        \Level1Out224[20] , \Level1Out224[19] , \Level1Out224[18] , 
        \Level1Out224[17] , \Level1Out224[16] , \Level1Out224[15] , 
        \Level1Out224[14] , \Level1Out224[13] , \Level1Out224[12] , 
        \Level1Out224[11] , \Level1Out224[10] , \Level1Out224[9] , 
        \Level1Out224[8] , \Level1Out224[7] , \Level1Out224[6] , 
        \Level1Out224[5] , \Level1Out224[4] , \Level1Out224[3] , 
        \Level1Out224[2] , \Level1Out224[1] , \Level1Out224[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_90_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load90[0] ), .Out({\Level2Out90[31] , \Level2Out90[30] , 
        \Level2Out90[29] , \Level2Out90[28] , \Level2Out90[27] , 
        \Level2Out90[26] , \Level2Out90[25] , \Level2Out90[24] , 
        \Level2Out90[23] , \Level2Out90[22] , \Level2Out90[21] , 
        \Level2Out90[20] , \Level2Out90[19] , \Level2Out90[18] , 
        \Level2Out90[17] , \Level2Out90[16] , \Level2Out90[15] , 
        \Level2Out90[14] , \Level2Out90[13] , \Level2Out90[12] , 
        \Level2Out90[11] , \Level2Out90[10] , \Level2Out90[9] , 
        \Level2Out90[8] , \Level2Out90[7] , \Level2Out90[6] , \Level2Out90[5] , 
        \Level2Out90[4] , \Level2Out90[3] , \Level2Out90[2] , \Level2Out90[1] , 
        \Level2Out90[0] }), .In1({\Level1Out90[31] , \Level1Out90[30] , 
        \Level1Out90[29] , \Level1Out90[28] , \Level1Out90[27] , 
        \Level1Out90[26] , \Level1Out90[25] , \Level1Out90[24] , 
        \Level1Out90[23] , \Level1Out90[22] , \Level1Out90[21] , 
        \Level1Out90[20] , \Level1Out90[19] , \Level1Out90[18] , 
        \Level1Out90[17] , \Level1Out90[16] , \Level1Out90[15] , 
        \Level1Out90[14] , \Level1Out90[13] , \Level1Out90[12] , 
        \Level1Out90[11] , \Level1Out90[10] , \Level1Out90[9] , 
        \Level1Out90[8] , \Level1Out90[7] , \Level1Out90[6] , \Level1Out90[5] , 
        \Level1Out90[4] , \Level1Out90[3] , \Level1Out90[2] , \Level1Out90[1] , 
        \Level1Out90[0] }), .In2({\Level1Out91[31] , \Level1Out91[30] , 
        \Level1Out91[29] , \Level1Out91[28] , \Level1Out91[27] , 
        \Level1Out91[26] , \Level1Out91[25] , \Level1Out91[24] , 
        \Level1Out91[23] , \Level1Out91[22] , \Level1Out91[21] , 
        \Level1Out91[20] , \Level1Out91[19] , \Level1Out91[18] , 
        \Level1Out91[17] , \Level1Out91[16] , \Level1Out91[15] , 
        \Level1Out91[14] , \Level1Out91[13] , \Level1Out91[12] , 
        \Level1Out91[11] , \Level1Out91[10] , \Level1Out91[9] , 
        \Level1Out91[8] , \Level1Out91[7] , \Level1Out91[6] , \Level1Out91[5] , 
        \Level1Out91[4] , \Level1Out91[3] , \Level1Out91[2] , \Level1Out91[1] , 
        \Level1Out91[0] }), .Read1(\Level1Load90[0] ), .Read2(
        \Level1Load91[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_140_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load140[0] ), .Out({\Level2Out140[31] , \Level2Out140[30] , 
        \Level2Out140[29] , \Level2Out140[28] , \Level2Out140[27] , 
        \Level2Out140[26] , \Level2Out140[25] , \Level2Out140[24] , 
        \Level2Out140[23] , \Level2Out140[22] , \Level2Out140[21] , 
        \Level2Out140[20] , \Level2Out140[19] , \Level2Out140[18] , 
        \Level2Out140[17] , \Level2Out140[16] , \Level2Out140[15] , 
        \Level2Out140[14] , \Level2Out140[13] , \Level2Out140[12] , 
        \Level2Out140[11] , \Level2Out140[10] , \Level2Out140[9] , 
        \Level2Out140[8] , \Level2Out140[7] , \Level2Out140[6] , 
        \Level2Out140[5] , \Level2Out140[4] , \Level2Out140[3] , 
        \Level2Out140[2] , \Level2Out140[1] , \Level2Out140[0] }), .In1({
        \Level1Out140[31] , \Level1Out140[30] , \Level1Out140[29] , 
        \Level1Out140[28] , \Level1Out140[27] , \Level1Out140[26] , 
        \Level1Out140[25] , \Level1Out140[24] , \Level1Out140[23] , 
        \Level1Out140[22] , \Level1Out140[21] , \Level1Out140[20] , 
        \Level1Out140[19] , \Level1Out140[18] , \Level1Out140[17] , 
        \Level1Out140[16] , \Level1Out140[15] , \Level1Out140[14] , 
        \Level1Out140[13] , \Level1Out140[12] , \Level1Out140[11] , 
        \Level1Out140[10] , \Level1Out140[9] , \Level1Out140[8] , 
        \Level1Out140[7] , \Level1Out140[6] , \Level1Out140[5] , 
        \Level1Out140[4] , \Level1Out140[3] , \Level1Out140[2] , 
        \Level1Out140[1] , \Level1Out140[0] }), .In2({\Level1Out141[31] , 
        \Level1Out141[30] , \Level1Out141[29] , \Level1Out141[28] , 
        \Level1Out141[27] , \Level1Out141[26] , \Level1Out141[25] , 
        \Level1Out141[24] , \Level1Out141[23] , \Level1Out141[22] , 
        \Level1Out141[21] , \Level1Out141[20] , \Level1Out141[19] , 
        \Level1Out141[18] , \Level1Out141[17] , \Level1Out141[16] , 
        \Level1Out141[15] , \Level1Out141[14] , \Level1Out141[13] , 
        \Level1Out141[12] , \Level1Out141[11] , \Level1Out141[10] , 
        \Level1Out141[9] , \Level1Out141[8] , \Level1Out141[7] , 
        \Level1Out141[6] , \Level1Out141[5] , \Level1Out141[4] , 
        \Level1Out141[3] , \Level1Out141[2] , \Level1Out141[1] , 
        \Level1Out141[0] }), .Read1(\Level1Load140[0] ), .Read2(
        \Level1Load141[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_176_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load176[0] ), .Out({\Level4Out176[31] , \Level4Out176[30] , 
        \Level4Out176[29] , \Level4Out176[28] , \Level4Out176[27] , 
        \Level4Out176[26] , \Level4Out176[25] , \Level4Out176[24] , 
        \Level4Out176[23] , \Level4Out176[22] , \Level4Out176[21] , 
        \Level4Out176[20] , \Level4Out176[19] , \Level4Out176[18] , 
        \Level4Out176[17] , \Level4Out176[16] , \Level4Out176[15] , 
        \Level4Out176[14] , \Level4Out176[13] , \Level4Out176[12] , 
        \Level4Out176[11] , \Level4Out176[10] , \Level4Out176[9] , 
        \Level4Out176[8] , \Level4Out176[7] , \Level4Out176[6] , 
        \Level4Out176[5] , \Level4Out176[4] , \Level4Out176[3] , 
        \Level4Out176[2] , \Level4Out176[1] , \Level4Out176[0] }), .In1({
        \Level2Out176[31] , \Level2Out176[30] , \Level2Out176[29] , 
        \Level2Out176[28] , \Level2Out176[27] , \Level2Out176[26] , 
        \Level2Out176[25] , \Level2Out176[24] , \Level2Out176[23] , 
        \Level2Out176[22] , \Level2Out176[21] , \Level2Out176[20] , 
        \Level2Out176[19] , \Level2Out176[18] , \Level2Out176[17] , 
        \Level2Out176[16] , \Level2Out176[15] , \Level2Out176[14] , 
        \Level2Out176[13] , \Level2Out176[12] , \Level2Out176[11] , 
        \Level2Out176[10] , \Level2Out176[9] , \Level2Out176[8] , 
        \Level2Out176[7] , \Level2Out176[6] , \Level2Out176[5] , 
        \Level2Out176[4] , \Level2Out176[3] , \Level2Out176[2] , 
        \Level2Out176[1] , \Level2Out176[0] }), .In2({\Level2Out178[31] , 
        \Level2Out178[30] , \Level2Out178[29] , \Level2Out178[28] , 
        \Level2Out178[27] , \Level2Out178[26] , \Level2Out178[25] , 
        \Level2Out178[24] , \Level2Out178[23] , \Level2Out178[22] , 
        \Level2Out178[21] , \Level2Out178[20] , \Level2Out178[19] , 
        \Level2Out178[18] , \Level2Out178[17] , \Level2Out178[16] , 
        \Level2Out178[15] , \Level2Out178[14] , \Level2Out178[13] , 
        \Level2Out178[12] , \Level2Out178[11] , \Level2Out178[10] , 
        \Level2Out178[9] , \Level2Out178[8] , \Level2Out178[7] , 
        \Level2Out178[6] , \Level2Out178[5] , \Level2Out178[4] , 
        \Level2Out178[3] , \Level2Out178[2] , \Level2Out178[1] , 
        \Level2Out178[0] }), .Read1(\Level2Load176[0] ), .Read2(
        \Level2Load178[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load32[0] ), .Out({\Level8Out32[31] , \Level8Out32[30] , 
        \Level8Out32[29] , \Level8Out32[28] , \Level8Out32[27] , 
        \Level8Out32[26] , \Level8Out32[25] , \Level8Out32[24] , 
        \Level8Out32[23] , \Level8Out32[22] , \Level8Out32[21] , 
        \Level8Out32[20] , \Level8Out32[19] , \Level8Out32[18] , 
        \Level8Out32[17] , \Level8Out32[16] , \Level8Out32[15] , 
        \Level8Out32[14] , \Level8Out32[13] , \Level8Out32[12] , 
        \Level8Out32[11] , \Level8Out32[10] , \Level8Out32[9] , 
        \Level8Out32[8] , \Level8Out32[7] , \Level8Out32[6] , \Level8Out32[5] , 
        \Level8Out32[4] , \Level8Out32[3] , \Level8Out32[2] , \Level8Out32[1] , 
        \Level8Out32[0] }), .In1({\Level4Out32[31] , \Level4Out32[30] , 
        \Level4Out32[29] , \Level4Out32[28] , \Level4Out32[27] , 
        \Level4Out32[26] , \Level4Out32[25] , \Level4Out32[24] , 
        \Level4Out32[23] , \Level4Out32[22] , \Level4Out32[21] , 
        \Level4Out32[20] , \Level4Out32[19] , \Level4Out32[18] , 
        \Level4Out32[17] , \Level4Out32[16] , \Level4Out32[15] , 
        \Level4Out32[14] , \Level4Out32[13] , \Level4Out32[12] , 
        \Level4Out32[11] , \Level4Out32[10] , \Level4Out32[9] , 
        \Level4Out32[8] , \Level4Out32[7] , \Level4Out32[6] , \Level4Out32[5] , 
        \Level4Out32[4] , \Level4Out32[3] , \Level4Out32[2] , \Level4Out32[1] , 
        \Level4Out32[0] }), .In2({\Level4Out36[31] , \Level4Out36[30] , 
        \Level4Out36[29] , \Level4Out36[28] , \Level4Out36[27] , 
        \Level4Out36[26] , \Level4Out36[25] , \Level4Out36[24] , 
        \Level4Out36[23] , \Level4Out36[22] , \Level4Out36[21] , 
        \Level4Out36[20] , \Level4Out36[19] , \Level4Out36[18] , 
        \Level4Out36[17] , \Level4Out36[16] , \Level4Out36[15] , 
        \Level4Out36[14] , \Level4Out36[13] , \Level4Out36[12] , 
        \Level4Out36[11] , \Level4Out36[10] , \Level4Out36[9] , 
        \Level4Out36[8] , \Level4Out36[7] , \Level4Out36[6] , \Level4Out36[5] , 
        \Level4Out36[4] , \Level4Out36[3] , \Level4Out36[2] , \Level4Out36[1] , 
        \Level4Out36[0] }), .Read1(\Level4Load32[0] ), .Read2(
        \Level4Load36[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_240_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load240[0] ), .Out({\Level8Out240[31] , \Level8Out240[30] , 
        \Level8Out240[29] , \Level8Out240[28] , \Level8Out240[27] , 
        \Level8Out240[26] , \Level8Out240[25] , \Level8Out240[24] , 
        \Level8Out240[23] , \Level8Out240[22] , \Level8Out240[21] , 
        \Level8Out240[20] , \Level8Out240[19] , \Level8Out240[18] , 
        \Level8Out240[17] , \Level8Out240[16] , \Level8Out240[15] , 
        \Level8Out240[14] , \Level8Out240[13] , \Level8Out240[12] , 
        \Level8Out240[11] , \Level8Out240[10] , \Level8Out240[9] , 
        \Level8Out240[8] , \Level8Out240[7] , \Level8Out240[6] , 
        \Level8Out240[5] , \Level8Out240[4] , \Level8Out240[3] , 
        \Level8Out240[2] , \Level8Out240[1] , \Level8Out240[0] }), .In1({
        \Level4Out240[31] , \Level4Out240[30] , \Level4Out240[29] , 
        \Level4Out240[28] , \Level4Out240[27] , \Level4Out240[26] , 
        \Level4Out240[25] , \Level4Out240[24] , \Level4Out240[23] , 
        \Level4Out240[22] , \Level4Out240[21] , \Level4Out240[20] , 
        \Level4Out240[19] , \Level4Out240[18] , \Level4Out240[17] , 
        \Level4Out240[16] , \Level4Out240[15] , \Level4Out240[14] , 
        \Level4Out240[13] , \Level4Out240[12] , \Level4Out240[11] , 
        \Level4Out240[10] , \Level4Out240[9] , \Level4Out240[8] , 
        \Level4Out240[7] , \Level4Out240[6] , \Level4Out240[5] , 
        \Level4Out240[4] , \Level4Out240[3] , \Level4Out240[2] , 
        \Level4Out240[1] , \Level4Out240[0] }), .In2({\Level4Out244[31] , 
        \Level4Out244[30] , \Level4Out244[29] , \Level4Out244[28] , 
        \Level4Out244[27] , \Level4Out244[26] , \Level4Out244[25] , 
        \Level4Out244[24] , \Level4Out244[23] , \Level4Out244[22] , 
        \Level4Out244[21] , \Level4Out244[20] , \Level4Out244[19] , 
        \Level4Out244[18] , \Level4Out244[17] , \Level4Out244[16] , 
        \Level4Out244[15] , \Level4Out244[14] , \Level4Out244[13] , 
        \Level4Out244[12] , \Level4Out244[11] , \Level4Out244[10] , 
        \Level4Out244[9] , \Level4Out244[8] , \Level4Out244[7] , 
        \Level4Out244[6] , \Level4Out244[5] , \Level4Out244[4] , 
        \Level4Out244[3] , \Level4Out244[2] , \Level4Out244[1] , 
        \Level4Out244[0] }), .Read1(\Level4Load240[0] ), .Read2(
        \Level4Load244[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_133 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink133[31] , \ScanLink133[30] , 
        \ScanLink133[29] , \ScanLink133[28] , \ScanLink133[27] , 
        \ScanLink133[26] , \ScanLink133[25] , \ScanLink133[24] , 
        \ScanLink133[23] , \ScanLink133[22] , \ScanLink133[21] , 
        \ScanLink133[20] , \ScanLink133[19] , \ScanLink133[18] , 
        \ScanLink133[17] , \ScanLink133[16] , \ScanLink133[15] , 
        \ScanLink133[14] , \ScanLink133[13] , \ScanLink133[12] , 
        \ScanLink133[11] , \ScanLink133[10] , \ScanLink133[9] , 
        \ScanLink133[8] , \ScanLink133[7] , \ScanLink133[6] , \ScanLink133[5] , 
        \ScanLink133[4] , \ScanLink133[3] , \ScanLink133[2] , \ScanLink133[1] , 
        \ScanLink133[0] }), .ScanOut({\ScanLink134[31] , \ScanLink134[30] , 
        \ScanLink134[29] , \ScanLink134[28] , \ScanLink134[27] , 
        \ScanLink134[26] , \ScanLink134[25] , \ScanLink134[24] , 
        \ScanLink134[23] , \ScanLink134[22] , \ScanLink134[21] , 
        \ScanLink134[20] , \ScanLink134[19] , \ScanLink134[18] , 
        \ScanLink134[17] , \ScanLink134[16] , \ScanLink134[15] , 
        \ScanLink134[14] , \ScanLink134[13] , \ScanLink134[12] , 
        \ScanLink134[11] , \ScanLink134[10] , \ScanLink134[9] , 
        \ScanLink134[8] , \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , 
        \ScanLink134[4] , \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , 
        \ScanLink134[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load133[0] ), .Out({\Level1Out133[31] , \Level1Out133[30] , 
        \Level1Out133[29] , \Level1Out133[28] , \Level1Out133[27] , 
        \Level1Out133[26] , \Level1Out133[25] , \Level1Out133[24] , 
        \Level1Out133[23] , \Level1Out133[22] , \Level1Out133[21] , 
        \Level1Out133[20] , \Level1Out133[19] , \Level1Out133[18] , 
        \Level1Out133[17] , \Level1Out133[16] , \Level1Out133[15] , 
        \Level1Out133[14] , \Level1Out133[13] , \Level1Out133[12] , 
        \Level1Out133[11] , \Level1Out133[10] , \Level1Out133[9] , 
        \Level1Out133[8] , \Level1Out133[7] , \Level1Out133[6] , 
        \Level1Out133[5] , \Level1Out133[4] , \Level1Out133[3] , 
        \Level1Out133[2] , \Level1Out133[1] , \Level1Out133[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_203 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink203[31] , \ScanLink203[30] , 
        \ScanLink203[29] , \ScanLink203[28] , \ScanLink203[27] , 
        \ScanLink203[26] , \ScanLink203[25] , \ScanLink203[24] , 
        \ScanLink203[23] , \ScanLink203[22] , \ScanLink203[21] , 
        \ScanLink203[20] , \ScanLink203[19] , \ScanLink203[18] , 
        \ScanLink203[17] , \ScanLink203[16] , \ScanLink203[15] , 
        \ScanLink203[14] , \ScanLink203[13] , \ScanLink203[12] , 
        \ScanLink203[11] , \ScanLink203[10] , \ScanLink203[9] , 
        \ScanLink203[8] , \ScanLink203[7] , \ScanLink203[6] , \ScanLink203[5] , 
        \ScanLink203[4] , \ScanLink203[3] , \ScanLink203[2] , \ScanLink203[1] , 
        \ScanLink203[0] }), .ScanOut({\ScanLink204[31] , \ScanLink204[30] , 
        \ScanLink204[29] , \ScanLink204[28] , \ScanLink204[27] , 
        \ScanLink204[26] , \ScanLink204[25] , \ScanLink204[24] , 
        \ScanLink204[23] , \ScanLink204[22] , \ScanLink204[21] , 
        \ScanLink204[20] , \ScanLink204[19] , \ScanLink204[18] , 
        \ScanLink204[17] , \ScanLink204[16] , \ScanLink204[15] , 
        \ScanLink204[14] , \ScanLink204[13] , \ScanLink204[12] , 
        \ScanLink204[11] , \ScanLink204[10] , \ScanLink204[9] , 
        \ScanLink204[8] , \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , 
        \ScanLink204[4] , \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , 
        \ScanLink204[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load203[0] ), .Out({\Level1Out203[31] , \Level1Out203[30] , 
        \Level1Out203[29] , \Level1Out203[28] , \Level1Out203[27] , 
        \Level1Out203[26] , \Level1Out203[25] , \Level1Out203[24] , 
        \Level1Out203[23] , \Level1Out203[22] , \Level1Out203[21] , 
        \Level1Out203[20] , \Level1Out203[19] , \Level1Out203[18] , 
        \Level1Out203[17] , \Level1Out203[16] , \Level1Out203[15] , 
        \Level1Out203[14] , \Level1Out203[13] , \Level1Out203[12] , 
        \Level1Out203[11] , \Level1Out203[10] , \Level1Out203[9] , 
        \Level1Out203[8] , \Level1Out203[7] , \Level1Out203[6] , 
        \Level1Out203[5] , \Level1Out203[4] , \Level1Out203[3] , 
        \Level1Out203[2] , \Level1Out203[1] , \Level1Out203[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_24 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanOut({\ScanLink25[31] , 
        \ScanLink25[30] , \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , 
        \ScanLink25[26] , \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , 
        \ScanLink25[22] , \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , 
        \ScanLink25[18] , \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , 
        \ScanLink25[14] , \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , 
        \ScanLink25[10] , \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , 
        \ScanLink25[6] , \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , 
        \ScanLink25[2] , \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load24[0] ), .Out({
        \Level1Out24[31] , \Level1Out24[30] , \Level1Out24[29] , 
        \Level1Out24[28] , \Level1Out24[27] , \Level1Out24[26] , 
        \Level1Out24[25] , \Level1Out24[24] , \Level1Out24[23] , 
        \Level1Out24[22] , \Level1Out24[21] , \Level1Out24[20] , 
        \Level1Out24[19] , \Level1Out24[18] , \Level1Out24[17] , 
        \Level1Out24[16] , \Level1Out24[15] , \Level1Out24[14] , 
        \Level1Out24[13] , \Level1Out24[12] , \Level1Out24[11] , 
        \Level1Out24[10] , \Level1Out24[9] , \Level1Out24[8] , 
        \Level1Out24[7] , \Level1Out24[6] , \Level1Out24[5] , \Level1Out24[4] , 
        \Level1Out24[3] , \Level1Out24[2] , \Level1Out24[1] , \Level1Out24[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_36 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanOut({\ScanLink37[31] , 
        \ScanLink37[30] , \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , 
        \ScanLink37[26] , \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , 
        \ScanLink37[22] , \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , 
        \ScanLink37[18] , \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , 
        \ScanLink37[14] , \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , 
        \ScanLink37[10] , \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , 
        \ScanLink37[6] , \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , 
        \ScanLink37[2] , \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load36[0] ), .Out({
        \Level1Out36[31] , \Level1Out36[30] , \Level1Out36[29] , 
        \Level1Out36[28] , \Level1Out36[27] , \Level1Out36[26] , 
        \Level1Out36[25] , \Level1Out36[24] , \Level1Out36[23] , 
        \Level1Out36[22] , \Level1Out36[21] , \Level1Out36[20] , 
        \Level1Out36[19] , \Level1Out36[18] , \Level1Out36[17] , 
        \Level1Out36[16] , \Level1Out36[15] , \Level1Out36[14] , 
        \Level1Out36[13] , \Level1Out36[12] , \Level1Out36[11] , 
        \Level1Out36[10] , \Level1Out36[9] , \Level1Out36[8] , 
        \Level1Out36[7] , \Level1Out36[6] , \Level1Out36[5] , \Level1Out36[4] , 
        \Level1Out36[3] , \Level1Out36[2] , \Level1Out36[1] , \Level1Out36[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load48[0] ), .Out({\Level8Out48[31] , \Level8Out48[30] , 
        \Level8Out48[29] , \Level8Out48[28] , \Level8Out48[27] , 
        \Level8Out48[26] , \Level8Out48[25] , \Level8Out48[24] , 
        \Level8Out48[23] , \Level8Out48[22] , \Level8Out48[21] , 
        \Level8Out48[20] , \Level8Out48[19] , \Level8Out48[18] , 
        \Level8Out48[17] , \Level8Out48[16] , \Level8Out48[15] , 
        \Level8Out48[14] , \Level8Out48[13] , \Level8Out48[12] , 
        \Level8Out48[11] , \Level8Out48[10] , \Level8Out48[9] , 
        \Level8Out48[8] , \Level8Out48[7] , \Level8Out48[6] , \Level8Out48[5] , 
        \Level8Out48[4] , \Level8Out48[3] , \Level8Out48[2] , \Level8Out48[1] , 
        \Level8Out48[0] }), .In1({\Level4Out48[31] , \Level4Out48[30] , 
        \Level4Out48[29] , \Level4Out48[28] , \Level4Out48[27] , 
        \Level4Out48[26] , \Level4Out48[25] , \Level4Out48[24] , 
        \Level4Out48[23] , \Level4Out48[22] , \Level4Out48[21] , 
        \Level4Out48[20] , \Level4Out48[19] , \Level4Out48[18] , 
        \Level4Out48[17] , \Level4Out48[16] , \Level4Out48[15] , 
        \Level4Out48[14] , \Level4Out48[13] , \Level4Out48[12] , 
        \Level4Out48[11] , \Level4Out48[10] , \Level4Out48[9] , 
        \Level4Out48[8] , \Level4Out48[7] , \Level4Out48[6] , \Level4Out48[5] , 
        \Level4Out48[4] , \Level4Out48[3] , \Level4Out48[2] , \Level4Out48[1] , 
        \Level4Out48[0] }), .In2({\Level4Out52[31] , \Level4Out52[30] , 
        \Level4Out52[29] , \Level4Out52[28] , \Level4Out52[27] , 
        \Level4Out52[26] , \Level4Out52[25] , \Level4Out52[24] , 
        \Level4Out52[23] , \Level4Out52[22] , \Level4Out52[21] , 
        \Level4Out52[20] , \Level4Out52[19] , \Level4Out52[18] , 
        \Level4Out52[17] , \Level4Out52[16] , \Level4Out52[15] , 
        \Level4Out52[14] , \Level4Out52[13] , \Level4Out52[12] , 
        \Level4Out52[11] , \Level4Out52[10] , \Level4Out52[9] , 
        \Level4Out52[8] , \Level4Out52[7] , \Level4Out52[6] , \Level4Out52[5] , 
        \Level4Out52[4] , \Level4Out52[3] , \Level4Out52[2] , \Level4Out52[1] , 
        \Level4Out52[0] }), .Read1(\Level4Load48[0] ), .Read2(
        \Level4Load52[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_88 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink88[31] , \ScanLink88[30] , 
        \ScanLink88[29] , \ScanLink88[28] , \ScanLink88[27] , \ScanLink88[26] , 
        \ScanLink88[25] , \ScanLink88[24] , \ScanLink88[23] , \ScanLink88[22] , 
        \ScanLink88[21] , \ScanLink88[20] , \ScanLink88[19] , \ScanLink88[18] , 
        \ScanLink88[17] , \ScanLink88[16] , \ScanLink88[15] , \ScanLink88[14] , 
        \ScanLink88[13] , \ScanLink88[12] , \ScanLink88[11] , \ScanLink88[10] , 
        \ScanLink88[9] , \ScanLink88[8] , \ScanLink88[7] , \ScanLink88[6] , 
        \ScanLink88[5] , \ScanLink88[4] , \ScanLink88[3] , \ScanLink88[2] , 
        \ScanLink88[1] , \ScanLink88[0] }), .ScanOut({\ScanLink89[31] , 
        \ScanLink89[30] , \ScanLink89[29] , \ScanLink89[28] , \ScanLink89[27] , 
        \ScanLink89[26] , \ScanLink89[25] , \ScanLink89[24] , \ScanLink89[23] , 
        \ScanLink89[22] , \ScanLink89[21] , \ScanLink89[20] , \ScanLink89[19] , 
        \ScanLink89[18] , \ScanLink89[17] , \ScanLink89[16] , \ScanLink89[15] , 
        \ScanLink89[14] , \ScanLink89[13] , \ScanLink89[12] , \ScanLink89[11] , 
        \ScanLink89[10] , \ScanLink89[9] , \ScanLink89[8] , \ScanLink89[7] , 
        \ScanLink89[6] , \ScanLink89[5] , \ScanLink89[4] , \ScanLink89[3] , 
        \ScanLink89[2] , \ScanLink89[1] , \ScanLink89[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load88[0] ), .Out({
        \Level1Out88[31] , \Level1Out88[30] , \Level1Out88[29] , 
        \Level1Out88[28] , \Level1Out88[27] , \Level1Out88[26] , 
        \Level1Out88[25] , \Level1Out88[24] , \Level1Out88[23] , 
        \Level1Out88[22] , \Level1Out88[21] , \Level1Out88[20] , 
        \Level1Out88[19] , \Level1Out88[18] , \Level1Out88[17] , 
        \Level1Out88[16] , \Level1Out88[15] , \Level1Out88[14] , 
        \Level1Out88[13] , \Level1Out88[12] , \Level1Out88[11] , 
        \Level1Out88[10] , \Level1Out88[9] , \Level1Out88[8] , 
        \Level1Out88[7] , \Level1Out88[6] , \Level1Out88[5] , \Level1Out88[4] , 
        \Level1Out88[3] , \Level1Out88[2] , \Level1Out88[1] , \Level1Out88[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_236 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink236[31] , \ScanLink236[30] , 
        \ScanLink236[29] , \ScanLink236[28] , \ScanLink236[27] , 
        \ScanLink236[26] , \ScanLink236[25] , \ScanLink236[24] , 
        \ScanLink236[23] , \ScanLink236[22] , \ScanLink236[21] , 
        \ScanLink236[20] , \ScanLink236[19] , \ScanLink236[18] , 
        \ScanLink236[17] , \ScanLink236[16] , \ScanLink236[15] , 
        \ScanLink236[14] , \ScanLink236[13] , \ScanLink236[12] , 
        \ScanLink236[11] , \ScanLink236[10] , \ScanLink236[9] , 
        \ScanLink236[8] , \ScanLink236[7] , \ScanLink236[6] , \ScanLink236[5] , 
        \ScanLink236[4] , \ScanLink236[3] , \ScanLink236[2] , \ScanLink236[1] , 
        \ScanLink236[0] }), .ScanOut({\ScanLink237[31] , \ScanLink237[30] , 
        \ScanLink237[29] , \ScanLink237[28] , \ScanLink237[27] , 
        \ScanLink237[26] , \ScanLink237[25] , \ScanLink237[24] , 
        \ScanLink237[23] , \ScanLink237[22] , \ScanLink237[21] , 
        \ScanLink237[20] , \ScanLink237[19] , \ScanLink237[18] , 
        \ScanLink237[17] , \ScanLink237[16] , \ScanLink237[15] , 
        \ScanLink237[14] , \ScanLink237[13] , \ScanLink237[12] , 
        \ScanLink237[11] , \ScanLink237[10] , \ScanLink237[9] , 
        \ScanLink237[8] , \ScanLink237[7] , \ScanLink237[6] , \ScanLink237[5] , 
        \ScanLink237[4] , \ScanLink237[3] , \ScanLink237[2] , \ScanLink237[1] , 
        \ScanLink237[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load236[0] ), .Out({\Level1Out236[31] , \Level1Out236[30] , 
        \Level1Out236[29] , \Level1Out236[28] , \Level1Out236[27] , 
        \Level1Out236[26] , \Level1Out236[25] , \Level1Out236[24] , 
        \Level1Out236[23] , \Level1Out236[22] , \Level1Out236[21] , 
        \Level1Out236[20] , \Level1Out236[19] , \Level1Out236[18] , 
        \Level1Out236[17] , \Level1Out236[16] , \Level1Out236[15] , 
        \Level1Out236[14] , \Level1Out236[13] , \Level1Out236[12] , 
        \Level1Out236[11] , \Level1Out236[10] , \Level1Out236[9] , 
        \Level1Out236[8] , \Level1Out236[7] , \Level1Out236[6] , 
        \Level1Out236[5] , \Level1Out236[4] , \Level1Out236[3] , 
        \Level1Out236[2] , \Level1Out236[1] , \Level1Out236[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_186_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load186[0] ), .Out({\Level2Out186[31] , \Level2Out186[30] , 
        \Level2Out186[29] , \Level2Out186[28] , \Level2Out186[27] , 
        \Level2Out186[26] , \Level2Out186[25] , \Level2Out186[24] , 
        \Level2Out186[23] , \Level2Out186[22] , \Level2Out186[21] , 
        \Level2Out186[20] , \Level2Out186[19] , \Level2Out186[18] , 
        \Level2Out186[17] , \Level2Out186[16] , \Level2Out186[15] , 
        \Level2Out186[14] , \Level2Out186[13] , \Level2Out186[12] , 
        \Level2Out186[11] , \Level2Out186[10] , \Level2Out186[9] , 
        \Level2Out186[8] , \Level2Out186[7] , \Level2Out186[6] , 
        \Level2Out186[5] , \Level2Out186[4] , \Level2Out186[3] , 
        \Level2Out186[2] , \Level2Out186[1] , \Level2Out186[0] }), .In1({
        \Level1Out186[31] , \Level1Out186[30] , \Level1Out186[29] , 
        \Level1Out186[28] , \Level1Out186[27] , \Level1Out186[26] , 
        \Level1Out186[25] , \Level1Out186[24] , \Level1Out186[23] , 
        \Level1Out186[22] , \Level1Out186[21] , \Level1Out186[20] , 
        \Level1Out186[19] , \Level1Out186[18] , \Level1Out186[17] , 
        \Level1Out186[16] , \Level1Out186[15] , \Level1Out186[14] , 
        \Level1Out186[13] , \Level1Out186[12] , \Level1Out186[11] , 
        \Level1Out186[10] , \Level1Out186[9] , \Level1Out186[8] , 
        \Level1Out186[7] , \Level1Out186[6] , \Level1Out186[5] , 
        \Level1Out186[4] , \Level1Out186[3] , \Level1Out186[2] , 
        \Level1Out186[1] , \Level1Out186[0] }), .In2({\Level1Out187[31] , 
        \Level1Out187[30] , \Level1Out187[29] , \Level1Out187[28] , 
        \Level1Out187[27] , \Level1Out187[26] , \Level1Out187[25] , 
        \Level1Out187[24] , \Level1Out187[23] , \Level1Out187[22] , 
        \Level1Out187[21] , \Level1Out187[20] , \Level1Out187[19] , 
        \Level1Out187[18] , \Level1Out187[17] , \Level1Out187[16] , 
        \Level1Out187[15] , \Level1Out187[14] , \Level1Out187[13] , 
        \Level1Out187[12] , \Level1Out187[11] , \Level1Out187[10] , 
        \Level1Out187[9] , \Level1Out187[8] , \Level1Out187[7] , 
        \Level1Out187[6] , \Level1Out187[5] , \Level1Out187[4] , 
        \Level1Out187[3] , \Level1Out187[2] , \Level1Out187[1] , 
        \Level1Out187[0] }), .Read1(\Level1Load186[0] ), .Read2(
        \Level1Load187[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_16 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load192[0] ), .Out({\Level16Out192[31] , \Level16Out192[30] , 
        \Level16Out192[29] , \Level16Out192[28] , \Level16Out192[27] , 
        \Level16Out192[26] , \Level16Out192[25] , \Level16Out192[24] , 
        \Level16Out192[23] , \Level16Out192[22] , \Level16Out192[21] , 
        \Level16Out192[20] , \Level16Out192[19] , \Level16Out192[18] , 
        \Level16Out192[17] , \Level16Out192[16] , \Level16Out192[15] , 
        \Level16Out192[14] , \Level16Out192[13] , \Level16Out192[12] , 
        \Level16Out192[11] , \Level16Out192[10] , \Level16Out192[9] , 
        \Level16Out192[8] , \Level16Out192[7] , \Level16Out192[6] , 
        \Level16Out192[5] , \Level16Out192[4] , \Level16Out192[3] , 
        \Level16Out192[2] , \Level16Out192[1] , \Level16Out192[0] }), .In1({
        \Level8Out192[31] , \Level8Out192[30] , \Level8Out192[29] , 
        \Level8Out192[28] , \Level8Out192[27] , \Level8Out192[26] , 
        \Level8Out192[25] , \Level8Out192[24] , \Level8Out192[23] , 
        \Level8Out192[22] , \Level8Out192[21] , \Level8Out192[20] , 
        \Level8Out192[19] , \Level8Out192[18] , \Level8Out192[17] , 
        \Level8Out192[16] , \Level8Out192[15] , \Level8Out192[14] , 
        \Level8Out192[13] , \Level8Out192[12] , \Level8Out192[11] , 
        \Level8Out192[10] , \Level8Out192[9] , \Level8Out192[8] , 
        \Level8Out192[7] , \Level8Out192[6] , \Level8Out192[5] , 
        \Level8Out192[4] , \Level8Out192[3] , \Level8Out192[2] , 
        \Level8Out192[1] , \Level8Out192[0] }), .In2({\Level8Out200[31] , 
        \Level8Out200[30] , \Level8Out200[29] , \Level8Out200[28] , 
        \Level8Out200[27] , \Level8Out200[26] , \Level8Out200[25] , 
        \Level8Out200[24] , \Level8Out200[23] , \Level8Out200[22] , 
        \Level8Out200[21] , \Level8Out200[20] , \Level8Out200[19] , 
        \Level8Out200[18] , \Level8Out200[17] , \Level8Out200[16] , 
        \Level8Out200[15] , \Level8Out200[14] , \Level8Out200[13] , 
        \Level8Out200[12] , \Level8Out200[11] , \Level8Out200[10] , 
        \Level8Out200[9] , \Level8Out200[8] , \Level8Out200[7] , 
        \Level8Out200[6] , \Level8Out200[5] , \Level8Out200[4] , 
        \Level8Out200[3] , \Level8Out200[2] , \Level8Out200[1] , 
        \Level8Out200[0] }), .Read1(\Level8Load192[0] ), .Read2(
        \Level8Load200[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load56[0] ), .Out({\Level2Out56[31] , \Level2Out56[30] , 
        \Level2Out56[29] , \Level2Out56[28] , \Level2Out56[27] , 
        \Level2Out56[26] , \Level2Out56[25] , \Level2Out56[24] , 
        \Level2Out56[23] , \Level2Out56[22] , \Level2Out56[21] , 
        \Level2Out56[20] , \Level2Out56[19] , \Level2Out56[18] , 
        \Level2Out56[17] , \Level2Out56[16] , \Level2Out56[15] , 
        \Level2Out56[14] , \Level2Out56[13] , \Level2Out56[12] , 
        \Level2Out56[11] , \Level2Out56[10] , \Level2Out56[9] , 
        \Level2Out56[8] , \Level2Out56[7] , \Level2Out56[6] , \Level2Out56[5] , 
        \Level2Out56[4] , \Level2Out56[3] , \Level2Out56[2] , \Level2Out56[1] , 
        \Level2Out56[0] }), .In1({\Level1Out56[31] , \Level1Out56[30] , 
        \Level1Out56[29] , \Level1Out56[28] , \Level1Out56[27] , 
        \Level1Out56[26] , \Level1Out56[25] , \Level1Out56[24] , 
        \Level1Out56[23] , \Level1Out56[22] , \Level1Out56[21] , 
        \Level1Out56[20] , \Level1Out56[19] , \Level1Out56[18] , 
        \Level1Out56[17] , \Level1Out56[16] , \Level1Out56[15] , 
        \Level1Out56[14] , \Level1Out56[13] , \Level1Out56[12] , 
        \Level1Out56[11] , \Level1Out56[10] , \Level1Out56[9] , 
        \Level1Out56[8] , \Level1Out56[7] , \Level1Out56[6] , \Level1Out56[5] , 
        \Level1Out56[4] , \Level1Out56[3] , \Level1Out56[2] , \Level1Out56[1] , 
        \Level1Out56[0] }), .In2({\Level1Out57[31] , \Level1Out57[30] , 
        \Level1Out57[29] , \Level1Out57[28] , \Level1Out57[27] , 
        \Level1Out57[26] , \Level1Out57[25] , \Level1Out57[24] , 
        \Level1Out57[23] , \Level1Out57[22] , \Level1Out57[21] , 
        \Level1Out57[20] , \Level1Out57[19] , \Level1Out57[18] , 
        \Level1Out57[17] , \Level1Out57[16] , \Level1Out57[15] , 
        \Level1Out57[14] , \Level1Out57[13] , \Level1Out57[12] , 
        \Level1Out57[11] , \Level1Out57[10] , \Level1Out57[9] , 
        \Level1Out57[8] , \Level1Out57[7] , \Level1Out57[6] , \Level1Out57[5] , 
        \Level1Out57[4] , \Level1Out57[3] , \Level1Out57[2] , \Level1Out57[1] , 
        \Level1Out57[0] }), .Read1(\Level1Load56[0] ), .Read2(
        \Level1Load57[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_106 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink106[31] , \ScanLink106[30] , 
        \ScanLink106[29] , \ScanLink106[28] , \ScanLink106[27] , 
        \ScanLink106[26] , \ScanLink106[25] , \ScanLink106[24] , 
        \ScanLink106[23] , \ScanLink106[22] , \ScanLink106[21] , 
        \ScanLink106[20] , \ScanLink106[19] , \ScanLink106[18] , 
        \ScanLink106[17] , \ScanLink106[16] , \ScanLink106[15] , 
        \ScanLink106[14] , \ScanLink106[13] , \ScanLink106[12] , 
        \ScanLink106[11] , \ScanLink106[10] , \ScanLink106[9] , 
        \ScanLink106[8] , \ScanLink106[7] , \ScanLink106[6] , \ScanLink106[5] , 
        \ScanLink106[4] , \ScanLink106[3] , \ScanLink106[2] , \ScanLink106[1] , 
        \ScanLink106[0] }), .ScanOut({\ScanLink107[31] , \ScanLink107[30] , 
        \ScanLink107[29] , \ScanLink107[28] , \ScanLink107[27] , 
        \ScanLink107[26] , \ScanLink107[25] , \ScanLink107[24] , 
        \ScanLink107[23] , \ScanLink107[22] , \ScanLink107[21] , 
        \ScanLink107[20] , \ScanLink107[19] , \ScanLink107[18] , 
        \ScanLink107[17] , \ScanLink107[16] , \ScanLink107[15] , 
        \ScanLink107[14] , \ScanLink107[13] , \ScanLink107[12] , 
        \ScanLink107[11] , \ScanLink107[10] , \ScanLink107[9] , 
        \ScanLink107[8] , \ScanLink107[7] , \ScanLink107[6] , \ScanLink107[5] , 
        \ScanLink107[4] , \ScanLink107[3] , \ScanLink107[2] , \ScanLink107[1] , 
        \ScanLink107[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load106[0] ), .Out({\Level1Out106[31] , \Level1Out106[30] , 
        \Level1Out106[29] , \Level1Out106[28] , \Level1Out106[27] , 
        \Level1Out106[26] , \Level1Out106[25] , \Level1Out106[24] , 
        \Level1Out106[23] , \Level1Out106[22] , \Level1Out106[21] , 
        \Level1Out106[20] , \Level1Out106[19] , \Level1Out106[18] , 
        \Level1Out106[17] , \Level1Out106[16] , \Level1Out106[15] , 
        \Level1Out106[14] , \Level1Out106[13] , \Level1Out106[12] , 
        \Level1Out106[11] , \Level1Out106[10] , \Level1Out106[9] , 
        \Level1Out106[8] , \Level1Out106[7] , \Level1Out106[6] , 
        \Level1Out106[5] , \Level1Out106[4] , \Level1Out106[3] , 
        \Level1Out106[2] , \Level1Out106[1] , \Level1Out106[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_121 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink121[31] , \ScanLink121[30] , 
        \ScanLink121[29] , \ScanLink121[28] , \ScanLink121[27] , 
        \ScanLink121[26] , \ScanLink121[25] , \ScanLink121[24] , 
        \ScanLink121[23] , \ScanLink121[22] , \ScanLink121[21] , 
        \ScanLink121[20] , \ScanLink121[19] , \ScanLink121[18] , 
        \ScanLink121[17] , \ScanLink121[16] , \ScanLink121[15] , 
        \ScanLink121[14] , \ScanLink121[13] , \ScanLink121[12] , 
        \ScanLink121[11] , \ScanLink121[10] , \ScanLink121[9] , 
        \ScanLink121[8] , \ScanLink121[7] , \ScanLink121[6] , \ScanLink121[5] , 
        \ScanLink121[4] , \ScanLink121[3] , \ScanLink121[2] , \ScanLink121[1] , 
        \ScanLink121[0] }), .ScanOut({\ScanLink122[31] , \ScanLink122[30] , 
        \ScanLink122[29] , \ScanLink122[28] , \ScanLink122[27] , 
        \ScanLink122[26] , \ScanLink122[25] , \ScanLink122[24] , 
        \ScanLink122[23] , \ScanLink122[22] , \ScanLink122[21] , 
        \ScanLink122[20] , \ScanLink122[19] , \ScanLink122[18] , 
        \ScanLink122[17] , \ScanLink122[16] , \ScanLink122[15] , 
        \ScanLink122[14] , \ScanLink122[13] , \ScanLink122[12] , 
        \ScanLink122[11] , \ScanLink122[10] , \ScanLink122[9] , 
        \ScanLink122[8] , \ScanLink122[7] , \ScanLink122[6] , \ScanLink122[5] , 
        \ScanLink122[4] , \ScanLink122[3] , \ScanLink122[2] , \ScanLink122[1] , 
        \ScanLink122[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load121[0] ), .Out({\Level1Out121[31] , \Level1Out121[30] , 
        \Level1Out121[29] , \Level1Out121[28] , \Level1Out121[27] , 
        \Level1Out121[26] , \Level1Out121[25] , \Level1Out121[24] , 
        \Level1Out121[23] , \Level1Out121[22] , \Level1Out121[21] , 
        \Level1Out121[20] , \Level1Out121[19] , \Level1Out121[18] , 
        \Level1Out121[17] , \Level1Out121[16] , \Level1Out121[15] , 
        \Level1Out121[14] , \Level1Out121[13] , \Level1Out121[12] , 
        \Level1Out121[11] , \Level1Out121[10] , \Level1Out121[9] , 
        \Level1Out121[8] , \Level1Out121[7] , \Level1Out121[6] , 
        \Level1Out121[5] , \Level1Out121[4] , \Level1Out121[3] , 
        \Level1Out121[2] , \Level1Out121[1] , \Level1Out121[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_110_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load110[0] ), .Out({\Level2Out110[31] , \Level2Out110[30] , 
        \Level2Out110[29] , \Level2Out110[28] , \Level2Out110[27] , 
        \Level2Out110[26] , \Level2Out110[25] , \Level2Out110[24] , 
        \Level2Out110[23] , \Level2Out110[22] , \Level2Out110[21] , 
        \Level2Out110[20] , \Level2Out110[19] , \Level2Out110[18] , 
        \Level2Out110[17] , \Level2Out110[16] , \Level2Out110[15] , 
        \Level2Out110[14] , \Level2Out110[13] , \Level2Out110[12] , 
        \Level2Out110[11] , \Level2Out110[10] , \Level2Out110[9] , 
        \Level2Out110[8] , \Level2Out110[7] , \Level2Out110[6] , 
        \Level2Out110[5] , \Level2Out110[4] , \Level2Out110[3] , 
        \Level2Out110[2] , \Level2Out110[1] , \Level2Out110[0] }), .In1({
        \Level1Out110[31] , \Level1Out110[30] , \Level1Out110[29] , 
        \Level1Out110[28] , \Level1Out110[27] , \Level1Out110[26] , 
        \Level1Out110[25] , \Level1Out110[24] , \Level1Out110[23] , 
        \Level1Out110[22] , \Level1Out110[21] , \Level1Out110[20] , 
        \Level1Out110[19] , \Level1Out110[18] , \Level1Out110[17] , 
        \Level1Out110[16] , \Level1Out110[15] , \Level1Out110[14] , 
        \Level1Out110[13] , \Level1Out110[12] , \Level1Out110[11] , 
        \Level1Out110[10] , \Level1Out110[9] , \Level1Out110[8] , 
        \Level1Out110[7] , \Level1Out110[6] , \Level1Out110[5] , 
        \Level1Out110[4] , \Level1Out110[3] , \Level1Out110[2] , 
        \Level1Out110[1] , \Level1Out110[0] }), .In2({\Level1Out111[31] , 
        \Level1Out111[30] , \Level1Out111[29] , \Level1Out111[28] , 
        \Level1Out111[27] , \Level1Out111[26] , \Level1Out111[25] , 
        \Level1Out111[24] , \Level1Out111[23] , \Level1Out111[22] , 
        \Level1Out111[21] , \Level1Out111[20] , \Level1Out111[19] , 
        \Level1Out111[18] , \Level1Out111[17] , \Level1Out111[16] , 
        \Level1Out111[15] , \Level1Out111[14] , \Level1Out111[13] , 
        \Level1Out111[12] , \Level1Out111[11] , \Level1Out111[10] , 
        \Level1Out111[9] , \Level1Out111[8] , \Level1Out111[7] , 
        \Level1Out111[6] , \Level1Out111[5] , \Level1Out111[4] , 
        \Level1Out111[3] , \Level1Out111[2] , \Level1Out111[1] , 
        \Level1Out111[0] }), .Read1(\Level1Load110[0] ), .Read2(
        \Level1Load111[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_224_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load224[0] ), .Out({\Level2Out224[31] , \Level2Out224[30] , 
        \Level2Out224[29] , \Level2Out224[28] , \Level2Out224[27] , 
        \Level2Out224[26] , \Level2Out224[25] , \Level2Out224[24] , 
        \Level2Out224[23] , \Level2Out224[22] , \Level2Out224[21] , 
        \Level2Out224[20] , \Level2Out224[19] , \Level2Out224[18] , 
        \Level2Out224[17] , \Level2Out224[16] , \Level2Out224[15] , 
        \Level2Out224[14] , \Level2Out224[13] , \Level2Out224[12] , 
        \Level2Out224[11] , \Level2Out224[10] , \Level2Out224[9] , 
        \Level2Out224[8] , \Level2Out224[7] , \Level2Out224[6] , 
        \Level2Out224[5] , \Level2Out224[4] , \Level2Out224[3] , 
        \Level2Out224[2] , \Level2Out224[1] , \Level2Out224[0] }), .In1({
        \Level1Out224[31] , \Level1Out224[30] , \Level1Out224[29] , 
        \Level1Out224[28] , \Level1Out224[27] , \Level1Out224[26] , 
        \Level1Out224[25] , \Level1Out224[24] , \Level1Out224[23] , 
        \Level1Out224[22] , \Level1Out224[21] , \Level1Out224[20] , 
        \Level1Out224[19] , \Level1Out224[18] , \Level1Out224[17] , 
        \Level1Out224[16] , \Level1Out224[15] , \Level1Out224[14] , 
        \Level1Out224[13] , \Level1Out224[12] , \Level1Out224[11] , 
        \Level1Out224[10] , \Level1Out224[9] , \Level1Out224[8] , 
        \Level1Out224[7] , \Level1Out224[6] , \Level1Out224[5] , 
        \Level1Out224[4] , \Level1Out224[3] , \Level1Out224[2] , 
        \Level1Out224[1] , \Level1Out224[0] }), .In2({\Level1Out225[31] , 
        \Level1Out225[30] , \Level1Out225[29] , \Level1Out225[28] , 
        \Level1Out225[27] , \Level1Out225[26] , \Level1Out225[25] , 
        \Level1Out225[24] , \Level1Out225[23] , \Level1Out225[22] , 
        \Level1Out225[21] , \Level1Out225[20] , \Level1Out225[19] , 
        \Level1Out225[18] , \Level1Out225[17] , \Level1Out225[16] , 
        \Level1Out225[15] , \Level1Out225[14] , \Level1Out225[13] , 
        \Level1Out225[12] , \Level1Out225[11] , \Level1Out225[10] , 
        \Level1Out225[9] , \Level1Out225[8] , \Level1Out225[7] , 
        \Level1Out225[6] , \Level1Out225[5] , \Level1Out225[4] , 
        \Level1Out225[3] , \Level1Out225[2] , \Level1Out225[1] , 
        \Level1Out225[0] }), .Read1(\Level1Load224[0] ), .Read2(
        \Level1Load225[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_211 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink211[31] , \ScanLink211[30] , 
        \ScanLink211[29] , \ScanLink211[28] , \ScanLink211[27] , 
        \ScanLink211[26] , \ScanLink211[25] , \ScanLink211[24] , 
        \ScanLink211[23] , \ScanLink211[22] , \ScanLink211[21] , 
        \ScanLink211[20] , \ScanLink211[19] , \ScanLink211[18] , 
        \ScanLink211[17] , \ScanLink211[16] , \ScanLink211[15] , 
        \ScanLink211[14] , \ScanLink211[13] , \ScanLink211[12] , 
        \ScanLink211[11] , \ScanLink211[10] , \ScanLink211[9] , 
        \ScanLink211[8] , \ScanLink211[7] , \ScanLink211[6] , \ScanLink211[5] , 
        \ScanLink211[4] , \ScanLink211[3] , \ScanLink211[2] , \ScanLink211[1] , 
        \ScanLink211[0] }), .ScanOut({\ScanLink212[31] , \ScanLink212[30] , 
        \ScanLink212[29] , \ScanLink212[28] , \ScanLink212[27] , 
        \ScanLink212[26] , \ScanLink212[25] , \ScanLink212[24] , 
        \ScanLink212[23] , \ScanLink212[22] , \ScanLink212[21] , 
        \ScanLink212[20] , \ScanLink212[19] , \ScanLink212[18] , 
        \ScanLink212[17] , \ScanLink212[16] , \ScanLink212[15] , 
        \ScanLink212[14] , \ScanLink212[13] , \ScanLink212[12] , 
        \ScanLink212[11] , \ScanLink212[10] , \ScanLink212[9] , 
        \ScanLink212[8] , \ScanLink212[7] , \ScanLink212[6] , \ScanLink212[5] , 
        \ScanLink212[4] , \ScanLink212[3] , \ScanLink212[2] , \ScanLink212[1] , 
        \ScanLink212[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load211[0] ), .Out({\Level1Out211[31] , \Level1Out211[30] , 
        \Level1Out211[29] , \Level1Out211[28] , \Level1Out211[27] , 
        \Level1Out211[26] , \Level1Out211[25] , \Level1Out211[24] , 
        \Level1Out211[23] , \Level1Out211[22] , \Level1Out211[21] , 
        \Level1Out211[20] , \Level1Out211[19] , \Level1Out211[18] , 
        \Level1Out211[17] , \Level1Out211[16] , \Level1Out211[15] , 
        \Level1Out211[14] , \Level1Out211[13] , \Level1Out211[12] , 
        \Level1Out211[11] , \Level1Out211[10] , \Level1Out211[9] , 
        \Level1Out211[8] , \Level1Out211[7] , \Level1Out211[6] , 
        \Level1Out211[5] , \Level1Out211[4] , \Level1Out211[3] , 
        \Level1Out211[2] , \Level1Out211[1] , \Level1Out211[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_60_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load60[0] ), .Out({\Level4Out60[31] , \Level4Out60[30] , 
        \Level4Out60[29] , \Level4Out60[28] , \Level4Out60[27] , 
        \Level4Out60[26] , \Level4Out60[25] , \Level4Out60[24] , 
        \Level4Out60[23] , \Level4Out60[22] , \Level4Out60[21] , 
        \Level4Out60[20] , \Level4Out60[19] , \Level4Out60[18] , 
        \Level4Out60[17] , \Level4Out60[16] , \Level4Out60[15] , 
        \Level4Out60[14] , \Level4Out60[13] , \Level4Out60[12] , 
        \Level4Out60[11] , \Level4Out60[10] , \Level4Out60[9] , 
        \Level4Out60[8] , \Level4Out60[7] , \Level4Out60[6] , \Level4Out60[5] , 
        \Level4Out60[4] , \Level4Out60[3] , \Level4Out60[2] , \Level4Out60[1] , 
        \Level4Out60[0] }), .In1({\Level2Out60[31] , \Level2Out60[30] , 
        \Level2Out60[29] , \Level2Out60[28] , \Level2Out60[27] , 
        \Level2Out60[26] , \Level2Out60[25] , \Level2Out60[24] , 
        \Level2Out60[23] , \Level2Out60[22] , \Level2Out60[21] , 
        \Level2Out60[20] , \Level2Out60[19] , \Level2Out60[18] , 
        \Level2Out60[17] , \Level2Out60[16] , \Level2Out60[15] , 
        \Level2Out60[14] , \Level2Out60[13] , \Level2Out60[12] , 
        \Level2Out60[11] , \Level2Out60[10] , \Level2Out60[9] , 
        \Level2Out60[8] , \Level2Out60[7] , \Level2Out60[6] , \Level2Out60[5] , 
        \Level2Out60[4] , \Level2Out60[3] , \Level2Out60[2] , \Level2Out60[1] , 
        \Level2Out60[0] }), .In2({\Level2Out62[31] , \Level2Out62[30] , 
        \Level2Out62[29] , \Level2Out62[28] , \Level2Out62[27] , 
        \Level2Out62[26] , \Level2Out62[25] , \Level2Out62[24] , 
        \Level2Out62[23] , \Level2Out62[22] , \Level2Out62[21] , 
        \Level2Out62[20] , \Level2Out62[19] , \Level2Out62[18] , 
        \Level2Out62[17] , \Level2Out62[16] , \Level2Out62[15] , 
        \Level2Out62[14] , \Level2Out62[13] , \Level2Out62[12] , 
        \Level2Out62[11] , \Level2Out62[10] , \Level2Out62[9] , 
        \Level2Out62[8] , \Level2Out62[7] , \Level2Out62[6] , \Level2Out62[5] , 
        \Level2Out62[4] , \Level2Out62[3] , \Level2Out62[2] , \Level2Out62[1] , 
        \Level2Out62[0] }), .Read1(\Level2Load60[0] ), .Read2(
        \Level2Load62[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_212_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load212[0] ), .Out({\Level4Out212[31] , \Level4Out212[30] , 
        \Level4Out212[29] , \Level4Out212[28] , \Level4Out212[27] , 
        \Level4Out212[26] , \Level4Out212[25] , \Level4Out212[24] , 
        \Level4Out212[23] , \Level4Out212[22] , \Level4Out212[21] , 
        \Level4Out212[20] , \Level4Out212[19] , \Level4Out212[18] , 
        \Level4Out212[17] , \Level4Out212[16] , \Level4Out212[15] , 
        \Level4Out212[14] , \Level4Out212[13] , \Level4Out212[12] , 
        \Level4Out212[11] , \Level4Out212[10] , \Level4Out212[9] , 
        \Level4Out212[8] , \Level4Out212[7] , \Level4Out212[6] , 
        \Level4Out212[5] , \Level4Out212[4] , \Level4Out212[3] , 
        \Level4Out212[2] , \Level4Out212[1] , \Level4Out212[0] }), .In1({
        \Level2Out212[31] , \Level2Out212[30] , \Level2Out212[29] , 
        \Level2Out212[28] , \Level2Out212[27] , \Level2Out212[26] , 
        \Level2Out212[25] , \Level2Out212[24] , \Level2Out212[23] , 
        \Level2Out212[22] , \Level2Out212[21] , \Level2Out212[20] , 
        \Level2Out212[19] , \Level2Out212[18] , \Level2Out212[17] , 
        \Level2Out212[16] , \Level2Out212[15] , \Level2Out212[14] , 
        \Level2Out212[13] , \Level2Out212[12] , \Level2Out212[11] , 
        \Level2Out212[10] , \Level2Out212[9] , \Level2Out212[8] , 
        \Level2Out212[7] , \Level2Out212[6] , \Level2Out212[5] , 
        \Level2Out212[4] , \Level2Out212[3] , \Level2Out212[2] , 
        \Level2Out212[1] , \Level2Out212[0] }), .In2({\Level2Out214[31] , 
        \Level2Out214[30] , \Level2Out214[29] , \Level2Out214[28] , 
        \Level2Out214[27] , \Level2Out214[26] , \Level2Out214[25] , 
        \Level2Out214[24] , \Level2Out214[23] , \Level2Out214[22] , 
        \Level2Out214[21] , \Level2Out214[20] , \Level2Out214[19] , 
        \Level2Out214[18] , \Level2Out214[17] , \Level2Out214[16] , 
        \Level2Out214[15] , \Level2Out214[14] , \Level2Out214[13] , 
        \Level2Out214[12] , \Level2Out214[11] , \Level2Out214[10] , 
        \Level2Out214[9] , \Level2Out214[8] , \Level2Out214[7] , 
        \Level2Out214[6] , \Level2Out214[5] , \Level2Out214[4] , 
        \Level2Out214[3] , \Level2Out214[2] , \Level2Out214[1] , 
        \Level2Out214[0] }), .Read1(\Level2Load212[0] ), .Read2(
        \Level2Load214[0] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Top_Node ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink256[31] , \ScanLink256[30] , 
        \ScanLink256[29] , \ScanLink256[28] , \ScanLink256[27] , 
        \ScanLink256[26] , \ScanLink256[25] , \ScanLink256[24] , 
        \ScanLink256[23] , \ScanLink256[22] , \ScanLink256[21] , 
        \ScanLink256[20] , \ScanLink256[19] , \ScanLink256[18] , 
        \ScanLink256[17] , \ScanLink256[16] , \ScanLink256[15] , 
        \ScanLink256[14] , \ScanLink256[13] , \ScanLink256[12] , 
        \ScanLink256[11] , \ScanLink256[10] , \ScanLink256[9] , 
        \ScanLink256[8] , \ScanLink256[7] , \ScanLink256[6] , \ScanLink256[5] , 
        \ScanLink256[4] , \ScanLink256[3] , \ScanLink256[2] , \ScanLink256[1] , 
        \ScanLink256[0] }), .ScanOut({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b0), .Id(1'b1), .In1({\Level128Out0[31] , \Level128Out0[30] , 
        \Level128Out0[29] , \Level128Out0[28] , \Level128Out0[27] , 
        \Level128Out0[26] , \Level128Out0[25] , \Level128Out0[24] , 
        \Level128Out0[23] , \Level128Out0[22] , \Level128Out0[21] , 
        \Level128Out0[20] , \Level128Out0[19] , \Level128Out0[18] , 
        \Level128Out0[17] , \Level128Out0[16] , \Level128Out0[15] , 
        \Level128Out0[14] , \Level128Out0[13] , \Level128Out0[12] , 
        \Level128Out0[11] , \Level128Out0[10] , \Level128Out0[9] , 
        \Level128Out0[8] , \Level128Out0[7] , \Level128Out0[6] , 
        \Level128Out0[5] , \Level128Out0[4] , \Level128Out0[3] , 
        \Level128Out0[2] , \Level128Out0[1] , \Level128Out0[0] }), .In2({
        \Level128Out128[31] , \Level128Out128[30] , \Level128Out128[29] , 
        \Level128Out128[28] , \Level128Out128[27] , \Level128Out128[26] , 
        \Level128Out128[25] , \Level128Out128[24] , \Level128Out128[23] , 
        \Level128Out128[22] , \Level128Out128[21] , \Level128Out128[20] , 
        \Level128Out128[19] , \Level128Out128[18] , \Level128Out128[17] , 
        \Level128Out128[16] , \Level128Out128[15] , \Level128Out128[14] , 
        \Level128Out128[13] , \Level128Out128[12] , \Level128Out128[11] , 
        \Level128Out128[10] , \Level128Out128[9] , \Level128Out128[8] , 
        \Level128Out128[7] , \Level128Out128[6] , \Level128Out128[5] , 
        \Level128Out128[4] , \Level128Out128[3] , \Level128Out128[2] , 
        \Level128Out128[1] , \Level128Out128[0] }), .Read1(\Level128Load0[0] ), 
        .Read2(\Level128Load128[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_18 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanOut({\ScanLink19[31] , 
        \ScanLink19[30] , \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , 
        \ScanLink19[26] , \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , 
        \ScanLink19[22] , \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , 
        \ScanLink19[18] , \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , 
        \ScanLink19[14] , \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , 
        \ScanLink19[10] , \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , 
        \ScanLink19[6] , \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , 
        \ScanLink19[2] , \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load18[0] ), .Out({
        \Level1Out18[31] , \Level1Out18[30] , \Level1Out18[29] , 
        \Level1Out18[28] , \Level1Out18[27] , \Level1Out18[26] , 
        \Level1Out18[25] , \Level1Out18[24] , \Level1Out18[23] , 
        \Level1Out18[22] , \Level1Out18[21] , \Level1Out18[20] , 
        \Level1Out18[19] , \Level1Out18[18] , \Level1Out18[17] , 
        \Level1Out18[16] , \Level1Out18[15] , \Level1Out18[14] , 
        \Level1Out18[13] , \Level1Out18[12] , \Level1Out18[11] , 
        \Level1Out18[10] , \Level1Out18[9] , \Level1Out18[8] , 
        \Level1Out18[7] , \Level1Out18[6] , \Level1Out18[5] , \Level1Out18[4] , 
        \Level1Out18[3] , \Level1Out18[2] , \Level1Out18[1] , \Level1Out18[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_51 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanOut({\ScanLink52[31] , 
        \ScanLink52[30] , \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , 
        \ScanLink52[26] , \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , 
        \ScanLink52[22] , \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , 
        \ScanLink52[18] , \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , 
        \ScanLink52[14] , \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , 
        \ScanLink52[10] , \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , 
        \ScanLink52[6] , \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , 
        \ScanLink52[2] , \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load51[0] ), .Out({
        \Level1Out51[31] , \Level1Out51[30] , \Level1Out51[29] , 
        \Level1Out51[28] , \Level1Out51[27] , \Level1Out51[26] , 
        \Level1Out51[25] , \Level1Out51[24] , \Level1Out51[23] , 
        \Level1Out51[22] , \Level1Out51[21] , \Level1Out51[20] , 
        \Level1Out51[19] , \Level1Out51[18] , \Level1Out51[17] , 
        \Level1Out51[16] , \Level1Out51[15] , \Level1Out51[14] , 
        \Level1Out51[13] , \Level1Out51[12] , \Level1Out51[11] , 
        \Level1Out51[10] , \Level1Out51[9] , \Level1Out51[8] , 
        \Level1Out51[7] , \Level1Out51[6] , \Level1Out51[5] , \Level1Out51[4] , 
        \Level1Out51[3] , \Level1Out51[2] , \Level1Out51[1] , \Level1Out51[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_76 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink76[31] , \ScanLink76[30] , 
        \ScanLink76[29] , \ScanLink76[28] , \ScanLink76[27] , \ScanLink76[26] , 
        \ScanLink76[25] , \ScanLink76[24] , \ScanLink76[23] , \ScanLink76[22] , 
        \ScanLink76[21] , \ScanLink76[20] , \ScanLink76[19] , \ScanLink76[18] , 
        \ScanLink76[17] , \ScanLink76[16] , \ScanLink76[15] , \ScanLink76[14] , 
        \ScanLink76[13] , \ScanLink76[12] , \ScanLink76[11] , \ScanLink76[10] , 
        \ScanLink76[9] , \ScanLink76[8] , \ScanLink76[7] , \ScanLink76[6] , 
        \ScanLink76[5] , \ScanLink76[4] , \ScanLink76[3] , \ScanLink76[2] , 
        \ScanLink76[1] , \ScanLink76[0] }), .ScanOut({\ScanLink77[31] , 
        \ScanLink77[30] , \ScanLink77[29] , \ScanLink77[28] , \ScanLink77[27] , 
        \ScanLink77[26] , \ScanLink77[25] , \ScanLink77[24] , \ScanLink77[23] , 
        \ScanLink77[22] , \ScanLink77[21] , \ScanLink77[20] , \ScanLink77[19] , 
        \ScanLink77[18] , \ScanLink77[17] , \ScanLink77[16] , \ScanLink77[15] , 
        \ScanLink77[14] , \ScanLink77[13] , \ScanLink77[12] , \ScanLink77[11] , 
        \ScanLink77[10] , \ScanLink77[9] , \ScanLink77[8] , \ScanLink77[7] , 
        \ScanLink77[6] , \ScanLink77[5] , \ScanLink77[4] , \ScanLink77[3] , 
        \ScanLink77[2] , \ScanLink77[1] , \ScanLink77[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load76[0] ), .Out({
        \Level1Out76[31] , \Level1Out76[30] , \Level1Out76[29] , 
        \Level1Out76[28] , \Level1Out76[27] , \Level1Out76[26] , 
        \Level1Out76[25] , \Level1Out76[24] , \Level1Out76[23] , 
        \Level1Out76[22] , \Level1Out76[21] , \Level1Out76[20] , 
        \Level1Out76[19] , \Level1Out76[18] , \Level1Out76[17] , 
        \Level1Out76[16] , \Level1Out76[15] , \Level1Out76[14] , 
        \Level1Out76[13] , \Level1Out76[12] , \Level1Out76[11] , 
        \Level1Out76[10] , \Level1Out76[9] , \Level1Out76[8] , 
        \Level1Out76[7] , \Level1Out76[6] , \Level1Out76[5] , \Level1Out76[4] , 
        \Level1Out76[3] , \Level1Out76[2] , \Level1Out76[1] , \Level1Out76[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_168 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink168[31] , \ScanLink168[30] , 
        \ScanLink168[29] , \ScanLink168[28] , \ScanLink168[27] , 
        \ScanLink168[26] , \ScanLink168[25] , \ScanLink168[24] , 
        \ScanLink168[23] , \ScanLink168[22] , \ScanLink168[21] , 
        \ScanLink168[20] , \ScanLink168[19] , \ScanLink168[18] , 
        \ScanLink168[17] , \ScanLink168[16] , \ScanLink168[15] , 
        \ScanLink168[14] , \ScanLink168[13] , \ScanLink168[12] , 
        \ScanLink168[11] , \ScanLink168[10] , \ScanLink168[9] , 
        \ScanLink168[8] , \ScanLink168[7] , \ScanLink168[6] , \ScanLink168[5] , 
        \ScanLink168[4] , \ScanLink168[3] , \ScanLink168[2] , \ScanLink168[1] , 
        \ScanLink168[0] }), .ScanOut({\ScanLink169[31] , \ScanLink169[30] , 
        \ScanLink169[29] , \ScanLink169[28] , \ScanLink169[27] , 
        \ScanLink169[26] , \ScanLink169[25] , \ScanLink169[24] , 
        \ScanLink169[23] , \ScanLink169[22] , \ScanLink169[21] , 
        \ScanLink169[20] , \ScanLink169[19] , \ScanLink169[18] , 
        \ScanLink169[17] , \ScanLink169[16] , \ScanLink169[15] , 
        \ScanLink169[14] , \ScanLink169[13] , \ScanLink169[12] , 
        \ScanLink169[11] , \ScanLink169[10] , \ScanLink169[9] , 
        \ScanLink169[8] , \ScanLink169[7] , \ScanLink169[6] , \ScanLink169[5] , 
        \ScanLink169[4] , \ScanLink169[3] , \ScanLink169[2] , \ScanLink169[1] , 
        \ScanLink169[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load168[0] ), .Out({\Level1Out168[31] , \Level1Out168[30] , 
        \Level1Out168[29] , \Level1Out168[28] , \Level1Out168[27] , 
        \Level1Out168[26] , \Level1Out168[25] , \Level1Out168[24] , 
        \Level1Out168[23] , \Level1Out168[22] , \Level1Out168[21] , 
        \Level1Out168[20] , \Level1Out168[19] , \Level1Out168[18] , 
        \Level1Out168[17] , \Level1Out168[16] , \Level1Out168[15] , 
        \Level1Out168[14] , \Level1Out168[13] , \Level1Out168[12] , 
        \Level1Out168[11] , \Level1Out168[10] , \Level1Out168[9] , 
        \Level1Out168[8] , \Level1Out168[7] , \Level1Out168[6] , 
        \Level1Out168[5] , \Level1Out168[4] , \Level1Out168[3] , 
        \Level1Out168[2] , \Level1Out168[1] , \Level1Out168[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load8[0] ), .Out({\Level8Out8[31] , \Level8Out8[30] , 
        \Level8Out8[29] , \Level8Out8[28] , \Level8Out8[27] , \Level8Out8[26] , 
        \Level8Out8[25] , \Level8Out8[24] , \Level8Out8[23] , \Level8Out8[22] , 
        \Level8Out8[21] , \Level8Out8[20] , \Level8Out8[19] , \Level8Out8[18] , 
        \Level8Out8[17] , \Level8Out8[16] , \Level8Out8[15] , \Level8Out8[14] , 
        \Level8Out8[13] , \Level8Out8[12] , \Level8Out8[11] , \Level8Out8[10] , 
        \Level8Out8[9] , \Level8Out8[8] , \Level8Out8[7] , \Level8Out8[6] , 
        \Level8Out8[5] , \Level8Out8[4] , \Level8Out8[3] , \Level8Out8[2] , 
        \Level8Out8[1] , \Level8Out8[0] }), .In1({\Level4Out8[31] , 
        \Level4Out8[30] , \Level4Out8[29] , \Level4Out8[28] , \Level4Out8[27] , 
        \Level4Out8[26] , \Level4Out8[25] , \Level4Out8[24] , \Level4Out8[23] , 
        \Level4Out8[22] , \Level4Out8[21] , \Level4Out8[20] , \Level4Out8[19] , 
        \Level4Out8[18] , \Level4Out8[17] , \Level4Out8[16] , \Level4Out8[15] , 
        \Level4Out8[14] , \Level4Out8[13] , \Level4Out8[12] , \Level4Out8[11] , 
        \Level4Out8[10] , \Level4Out8[9] , \Level4Out8[8] , \Level4Out8[7] , 
        \Level4Out8[6] , \Level4Out8[5] , \Level4Out8[4] , \Level4Out8[3] , 
        \Level4Out8[2] , \Level4Out8[1] , \Level4Out8[0] }), .In2({
        \Level4Out12[31] , \Level4Out12[30] , \Level4Out12[29] , 
        \Level4Out12[28] , \Level4Out12[27] , \Level4Out12[26] , 
        \Level4Out12[25] , \Level4Out12[24] , \Level4Out12[23] , 
        \Level4Out12[22] , \Level4Out12[21] , \Level4Out12[20] , 
        \Level4Out12[19] , \Level4Out12[18] , \Level4Out12[17] , 
        \Level4Out12[16] , \Level4Out12[15] , \Level4Out12[14] , 
        \Level4Out12[13] , \Level4Out12[12] , \Level4Out12[11] , 
        \Level4Out12[10] , \Level4Out12[9] , \Level4Out12[8] , 
        \Level4Out12[7] , \Level4Out12[6] , \Level4Out12[5] , \Level4Out12[4] , 
        \Level4Out12[3] , \Level4Out12[2] , \Level4Out12[1] , \Level4Out12[0] 
        }), .Read1(\Level4Load8[0] ), .Read2(\Level4Load12[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_93 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink93[31] , \ScanLink93[30] , 
        \ScanLink93[29] , \ScanLink93[28] , \ScanLink93[27] , \ScanLink93[26] , 
        \ScanLink93[25] , \ScanLink93[24] , \ScanLink93[23] , \ScanLink93[22] , 
        \ScanLink93[21] , \ScanLink93[20] , \ScanLink93[19] , \ScanLink93[18] , 
        \ScanLink93[17] , \ScanLink93[16] , \ScanLink93[15] , \ScanLink93[14] , 
        \ScanLink93[13] , \ScanLink93[12] , \ScanLink93[11] , \ScanLink93[10] , 
        \ScanLink93[9] , \ScanLink93[8] , \ScanLink93[7] , \ScanLink93[6] , 
        \ScanLink93[5] , \ScanLink93[4] , \ScanLink93[3] , \ScanLink93[2] , 
        \ScanLink93[1] , \ScanLink93[0] }), .ScanOut({\ScanLink94[31] , 
        \ScanLink94[30] , \ScanLink94[29] , \ScanLink94[28] , \ScanLink94[27] , 
        \ScanLink94[26] , \ScanLink94[25] , \ScanLink94[24] , \ScanLink94[23] , 
        \ScanLink94[22] , \ScanLink94[21] , \ScanLink94[20] , \ScanLink94[19] , 
        \ScanLink94[18] , \ScanLink94[17] , \ScanLink94[16] , \ScanLink94[15] , 
        \ScanLink94[14] , \ScanLink94[13] , \ScanLink94[12] , \ScanLink94[11] , 
        \ScanLink94[10] , \ScanLink94[9] , \ScanLink94[8] , \ScanLink94[7] , 
        \ScanLink94[6] , \ScanLink94[5] , \ScanLink94[4] , \ScanLink94[3] , 
        \ScanLink94[2] , \ScanLink94[1] , \ScanLink94[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load93[0] ), .Out({
        \Level1Out93[31] , \Level1Out93[30] , \Level1Out93[29] , 
        \Level1Out93[28] , \Level1Out93[27] , \Level1Out93[26] , 
        \Level1Out93[25] , \Level1Out93[24] , \Level1Out93[23] , 
        \Level1Out93[22] , \Level1Out93[21] , \Level1Out93[20] , 
        \Level1Out93[19] , \Level1Out93[18] , \Level1Out93[17] , 
        \Level1Out93[16] , \Level1Out93[15] , \Level1Out93[14] , 
        \Level1Out93[13] , \Level1Out93[12] , \Level1Out93[11] , 
        \Level1Out93[10] , \Level1Out93[9] , \Level1Out93[8] , 
        \Level1Out93[7] , \Level1Out93[6] , \Level1Out93[5] , \Level1Out93[4] , 
        \Level1Out93[3] , \Level1Out93[2] , \Level1Out93[1] , \Level1Out93[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_154 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink154[31] , \ScanLink154[30] , 
        \ScanLink154[29] , \ScanLink154[28] , \ScanLink154[27] , 
        \ScanLink154[26] , \ScanLink154[25] , \ScanLink154[24] , 
        \ScanLink154[23] , \ScanLink154[22] , \ScanLink154[21] , 
        \ScanLink154[20] , \ScanLink154[19] , \ScanLink154[18] , 
        \ScanLink154[17] , \ScanLink154[16] , \ScanLink154[15] , 
        \ScanLink154[14] , \ScanLink154[13] , \ScanLink154[12] , 
        \ScanLink154[11] , \ScanLink154[10] , \ScanLink154[9] , 
        \ScanLink154[8] , \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , 
        \ScanLink154[4] , \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , 
        \ScanLink154[0] }), .ScanOut({\ScanLink155[31] , \ScanLink155[30] , 
        \ScanLink155[29] , \ScanLink155[28] , \ScanLink155[27] , 
        \ScanLink155[26] , \ScanLink155[25] , \ScanLink155[24] , 
        \ScanLink155[23] , \ScanLink155[22] , \ScanLink155[21] , 
        \ScanLink155[20] , \ScanLink155[19] , \ScanLink155[18] , 
        \ScanLink155[17] , \ScanLink155[16] , \ScanLink155[15] , 
        \ScanLink155[14] , \ScanLink155[13] , \ScanLink155[12] , 
        \ScanLink155[11] , \ScanLink155[10] , \ScanLink155[9] , 
        \ScanLink155[8] , \ScanLink155[7] , \ScanLink155[6] , \ScanLink155[5] , 
        \ScanLink155[4] , \ScanLink155[3] , \ScanLink155[2] , \ScanLink155[1] , 
        \ScanLink155[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load154[0] ), .Out({\Level1Out154[31] , \Level1Out154[30] , 
        \Level1Out154[29] , \Level1Out154[28] , \Level1Out154[27] , 
        \Level1Out154[26] , \Level1Out154[25] , \Level1Out154[24] , 
        \Level1Out154[23] , \Level1Out154[22] , \Level1Out154[21] , 
        \Level1Out154[20] , \Level1Out154[19] , \Level1Out154[18] , 
        \Level1Out154[17] , \Level1Out154[16] , \Level1Out154[15] , 
        \Level1Out154[14] , \Level1Out154[13] , \Level1Out154[12] , 
        \Level1Out154[11] , \Level1Out154[10] , \Level1Out154[9] , 
        \Level1Out154[8] , \Level1Out154[7] , \Level1Out154[6] , 
        \Level1Out154[5] , \Level1Out154[4] , \Level1Out154[3] , 
        \Level1Out154[2] , \Level1Out154[1] , \Level1Out154[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_173 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink173[31] , \ScanLink173[30] , 
        \ScanLink173[29] , \ScanLink173[28] , \ScanLink173[27] , 
        \ScanLink173[26] , \ScanLink173[25] , \ScanLink173[24] , 
        \ScanLink173[23] , \ScanLink173[22] , \ScanLink173[21] , 
        \ScanLink173[20] , \ScanLink173[19] , \ScanLink173[18] , 
        \ScanLink173[17] , \ScanLink173[16] , \ScanLink173[15] , 
        \ScanLink173[14] , \ScanLink173[13] , \ScanLink173[12] , 
        \ScanLink173[11] , \ScanLink173[10] , \ScanLink173[9] , 
        \ScanLink173[8] , \ScanLink173[7] , \ScanLink173[6] , \ScanLink173[5] , 
        \ScanLink173[4] , \ScanLink173[3] , \ScanLink173[2] , \ScanLink173[1] , 
        \ScanLink173[0] }), .ScanOut({\ScanLink174[31] , \ScanLink174[30] , 
        \ScanLink174[29] , \ScanLink174[28] , \ScanLink174[27] , 
        \ScanLink174[26] , \ScanLink174[25] , \ScanLink174[24] , 
        \ScanLink174[23] , \ScanLink174[22] , \ScanLink174[21] , 
        \ScanLink174[20] , \ScanLink174[19] , \ScanLink174[18] , 
        \ScanLink174[17] , \ScanLink174[16] , \ScanLink174[15] , 
        \ScanLink174[14] , \ScanLink174[13] , \ScanLink174[12] , 
        \ScanLink174[11] , \ScanLink174[10] , \ScanLink174[9] , 
        \ScanLink174[8] , \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , 
        \ScanLink174[4] , \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , 
        \ScanLink174[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load173[0] ), .Out({\Level1Out173[31] , \Level1Out173[30] , 
        \Level1Out173[29] , \Level1Out173[28] , \Level1Out173[27] , 
        \Level1Out173[26] , \Level1Out173[25] , \Level1Out173[24] , 
        \Level1Out173[23] , \Level1Out173[22] , \Level1Out173[21] , 
        \Level1Out173[20] , \Level1Out173[19] , \Level1Out173[18] , 
        \Level1Out173[17] , \Level1Out173[16] , \Level1Out173[15] , 
        \Level1Out173[14] , \Level1Out173[13] , \Level1Out173[12] , 
        \Level1Out173[11] , \Level1Out173[10] , \Level1Out173[9] , 
        \Level1Out173[8] , \Level1Out173[7] , \Level1Out173[6] , 
        \Level1Out173[5] , \Level1Out173[4] , \Level1Out173[3] , 
        \Level1Out173[2] , \Level1Out173[1] , \Level1Out173[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_243 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink243[31] , \ScanLink243[30] , 
        \ScanLink243[29] , \ScanLink243[28] , \ScanLink243[27] , 
        \ScanLink243[26] , \ScanLink243[25] , \ScanLink243[24] , 
        \ScanLink243[23] , \ScanLink243[22] , \ScanLink243[21] , 
        \ScanLink243[20] , \ScanLink243[19] , \ScanLink243[18] , 
        \ScanLink243[17] , \ScanLink243[16] , \ScanLink243[15] , 
        \ScanLink243[14] , \ScanLink243[13] , \ScanLink243[12] , 
        \ScanLink243[11] , \ScanLink243[10] , \ScanLink243[9] , 
        \ScanLink243[8] , \ScanLink243[7] , \ScanLink243[6] , \ScanLink243[5] , 
        \ScanLink243[4] , \ScanLink243[3] , \ScanLink243[2] , \ScanLink243[1] , 
        \ScanLink243[0] }), .ScanOut({\ScanLink244[31] , \ScanLink244[30] , 
        \ScanLink244[29] , \ScanLink244[28] , \ScanLink244[27] , 
        \ScanLink244[26] , \ScanLink244[25] , \ScanLink244[24] , 
        \ScanLink244[23] , \ScanLink244[22] , \ScanLink244[21] , 
        \ScanLink244[20] , \ScanLink244[19] , \ScanLink244[18] , 
        \ScanLink244[17] , \ScanLink244[16] , \ScanLink244[15] , 
        \ScanLink244[14] , \ScanLink244[13] , \ScanLink244[12] , 
        \ScanLink244[11] , \ScanLink244[10] , \ScanLink244[9] , 
        \ScanLink244[8] , \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , 
        \ScanLink244[4] , \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , 
        \ScanLink244[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load243[0] ), .Out({\Level1Out243[31] , \Level1Out243[30] , 
        \Level1Out243[29] , \Level1Out243[28] , \Level1Out243[27] , 
        \Level1Out243[26] , \Level1Out243[25] , \Level1Out243[24] , 
        \Level1Out243[23] , \Level1Out243[22] , \Level1Out243[21] , 
        \Level1Out243[20] , \Level1Out243[19] , \Level1Out243[18] , 
        \Level1Out243[17] , \Level1Out243[16] , \Level1Out243[15] , 
        \Level1Out243[14] , \Level1Out243[13] , \Level1Out243[12] , 
        \Level1Out243[11] , \Level1Out243[10] , \Level1Out243[9] , 
        \Level1Out243[8] , \Level1Out243[7] , \Level1Out243[6] , 
        \Level1Out243[5] , \Level1Out243[4] , \Level1Out243[3] , 
        \Level1Out243[2] , \Level1Out243[1] , \Level1Out243[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_208_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load208[0] ), .Out({\Level8Out208[31] , \Level8Out208[30] , 
        \Level8Out208[29] , \Level8Out208[28] , \Level8Out208[27] , 
        \Level8Out208[26] , \Level8Out208[25] , \Level8Out208[24] , 
        \Level8Out208[23] , \Level8Out208[22] , \Level8Out208[21] , 
        \Level8Out208[20] , \Level8Out208[19] , \Level8Out208[18] , 
        \Level8Out208[17] , \Level8Out208[16] , \Level8Out208[15] , 
        \Level8Out208[14] , \Level8Out208[13] , \Level8Out208[12] , 
        \Level8Out208[11] , \Level8Out208[10] , \Level8Out208[9] , 
        \Level8Out208[8] , \Level8Out208[7] , \Level8Out208[6] , 
        \Level8Out208[5] , \Level8Out208[4] , \Level8Out208[3] , 
        \Level8Out208[2] , \Level8Out208[1] , \Level8Out208[0] }), .In1({
        \Level4Out208[31] , \Level4Out208[30] , \Level4Out208[29] , 
        \Level4Out208[28] , \Level4Out208[27] , \Level4Out208[26] , 
        \Level4Out208[25] , \Level4Out208[24] , \Level4Out208[23] , 
        \Level4Out208[22] , \Level4Out208[21] , \Level4Out208[20] , 
        \Level4Out208[19] , \Level4Out208[18] , \Level4Out208[17] , 
        \Level4Out208[16] , \Level4Out208[15] , \Level4Out208[14] , 
        \Level4Out208[13] , \Level4Out208[12] , \Level4Out208[11] , 
        \Level4Out208[10] , \Level4Out208[9] , \Level4Out208[8] , 
        \Level4Out208[7] , \Level4Out208[6] , \Level4Out208[5] , 
        \Level4Out208[4] , \Level4Out208[3] , \Level4Out208[2] , 
        \Level4Out208[1] , \Level4Out208[0] }), .In2({\Level4Out212[31] , 
        \Level4Out212[30] , \Level4Out212[29] , \Level4Out212[28] , 
        \Level4Out212[27] , \Level4Out212[26] , \Level4Out212[25] , 
        \Level4Out212[24] , \Level4Out212[23] , \Level4Out212[22] , 
        \Level4Out212[21] , \Level4Out212[20] , \Level4Out212[19] , 
        \Level4Out212[18] , \Level4Out212[17] , \Level4Out212[16] , 
        \Level4Out212[15] , \Level4Out212[14] , \Level4Out212[13] , 
        \Level4Out212[12] , \Level4Out212[11] , \Level4Out212[10] , 
        \Level4Out212[9] , \Level4Out212[8] , \Level4Out212[7] , 
        \Level4Out212[6] , \Level4Out212[5] , \Level4Out212[4] , 
        \Level4Out212[3] , \Level4Out212[2] , \Level4Out212[1] , 
        \Level4Out212[0] }), .Read1(\Level4Load208[0] ), .Read2(
        \Level4Load212[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_122_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load122[0] ), .Out({\Level2Out122[31] , \Level2Out122[30] , 
        \Level2Out122[29] , \Level2Out122[28] , \Level2Out122[27] , 
        \Level2Out122[26] , \Level2Out122[25] , \Level2Out122[24] , 
        \Level2Out122[23] , \Level2Out122[22] , \Level2Out122[21] , 
        \Level2Out122[20] , \Level2Out122[19] , \Level2Out122[18] , 
        \Level2Out122[17] , \Level2Out122[16] , \Level2Out122[15] , 
        \Level2Out122[14] , \Level2Out122[13] , \Level2Out122[12] , 
        \Level2Out122[11] , \Level2Out122[10] , \Level2Out122[9] , 
        \Level2Out122[8] , \Level2Out122[7] , \Level2Out122[6] , 
        \Level2Out122[5] , \Level2Out122[4] , \Level2Out122[3] , 
        \Level2Out122[2] , \Level2Out122[1] , \Level2Out122[0] }), .In1({
        \Level1Out122[31] , \Level1Out122[30] , \Level1Out122[29] , 
        \Level1Out122[28] , \Level1Out122[27] , \Level1Out122[26] , 
        \Level1Out122[25] , \Level1Out122[24] , \Level1Out122[23] , 
        \Level1Out122[22] , \Level1Out122[21] , \Level1Out122[20] , 
        \Level1Out122[19] , \Level1Out122[18] , \Level1Out122[17] , 
        \Level1Out122[16] , \Level1Out122[15] , \Level1Out122[14] , 
        \Level1Out122[13] , \Level1Out122[12] , \Level1Out122[11] , 
        \Level1Out122[10] , \Level1Out122[9] , \Level1Out122[8] , 
        \Level1Out122[7] , \Level1Out122[6] , \Level1Out122[5] , 
        \Level1Out122[4] , \Level1Out122[3] , \Level1Out122[2] , 
        \Level1Out122[1] , \Level1Out122[0] }), .In2({\Level1Out123[31] , 
        \Level1Out123[30] , \Level1Out123[29] , \Level1Out123[28] , 
        \Level1Out123[27] , \Level1Out123[26] , \Level1Out123[25] , 
        \Level1Out123[24] , \Level1Out123[23] , \Level1Out123[22] , 
        \Level1Out123[21] , \Level1Out123[20] , \Level1Out123[19] , 
        \Level1Out123[18] , \Level1Out123[17] , \Level1Out123[16] , 
        \Level1Out123[15] , \Level1Out123[14] , \Level1Out123[13] , 
        \Level1Out123[12] , \Level1Out123[11] , \Level1Out123[10] , 
        \Level1Out123[9] , \Level1Out123[8] , \Level1Out123[7] , 
        \Level1Out123[6] , \Level1Out123[5] , \Level1Out123[4] , 
        \Level1Out123[3] , \Level1Out123[2] , \Level1Out123[1] , 
        \Level1Out123[0] }), .Read1(\Level1Load122[0] ), .Read2(
        \Level1Load123[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_220_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load220[0] ), .Out({\Level4Out220[31] , \Level4Out220[30] , 
        \Level4Out220[29] , \Level4Out220[28] , \Level4Out220[27] , 
        \Level4Out220[26] , \Level4Out220[25] , \Level4Out220[24] , 
        \Level4Out220[23] , \Level4Out220[22] , \Level4Out220[21] , 
        \Level4Out220[20] , \Level4Out220[19] , \Level4Out220[18] , 
        \Level4Out220[17] , \Level4Out220[16] , \Level4Out220[15] , 
        \Level4Out220[14] , \Level4Out220[13] , \Level4Out220[12] , 
        \Level4Out220[11] , \Level4Out220[10] , \Level4Out220[9] , 
        \Level4Out220[8] , \Level4Out220[7] , \Level4Out220[6] , 
        \Level4Out220[5] , \Level4Out220[4] , \Level4Out220[3] , 
        \Level4Out220[2] , \Level4Out220[1] , \Level4Out220[0] }), .In1({
        \Level2Out220[31] , \Level2Out220[30] , \Level2Out220[29] , 
        \Level2Out220[28] , \Level2Out220[27] , \Level2Out220[26] , 
        \Level2Out220[25] , \Level2Out220[24] , \Level2Out220[23] , 
        \Level2Out220[22] , \Level2Out220[21] , \Level2Out220[20] , 
        \Level2Out220[19] , \Level2Out220[18] , \Level2Out220[17] , 
        \Level2Out220[16] , \Level2Out220[15] , \Level2Out220[14] , 
        \Level2Out220[13] , \Level2Out220[12] , \Level2Out220[11] , 
        \Level2Out220[10] , \Level2Out220[9] , \Level2Out220[8] , 
        \Level2Out220[7] , \Level2Out220[6] , \Level2Out220[5] , 
        \Level2Out220[4] , \Level2Out220[3] , \Level2Out220[2] , 
        \Level2Out220[1] , \Level2Out220[0] }), .In2({\Level2Out222[31] , 
        \Level2Out222[30] , \Level2Out222[29] , \Level2Out222[28] , 
        \Level2Out222[27] , \Level2Out222[26] , \Level2Out222[25] , 
        \Level2Out222[24] , \Level2Out222[23] , \Level2Out222[22] , 
        \Level2Out222[21] , \Level2Out222[20] , \Level2Out222[19] , 
        \Level2Out222[18] , \Level2Out222[17] , \Level2Out222[16] , 
        \Level2Out222[15] , \Level2Out222[14] , \Level2Out222[13] , 
        \Level2Out222[12] , \Level2Out222[11] , \Level2Out222[10] , 
        \Level2Out222[9] , \Level2Out222[8] , \Level2Out222[7] , 
        \Level2Out222[6] , \Level2Out222[5] , \Level2Out222[4] , 
        \Level2Out222[3] , \Level2Out222[2] , \Level2Out222[1] , 
        \Level2Out222[0] }), .Read1(\Level2Load220[0] ), .Read2(
        \Level2Load222[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_52_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load52[0] ), .Out({\Level4Out52[31] , \Level4Out52[30] , 
        \Level4Out52[29] , \Level4Out52[28] , \Level4Out52[27] , 
        \Level4Out52[26] , \Level4Out52[25] , \Level4Out52[24] , 
        \Level4Out52[23] , \Level4Out52[22] , \Level4Out52[21] , 
        \Level4Out52[20] , \Level4Out52[19] , \Level4Out52[18] , 
        \Level4Out52[17] , \Level4Out52[16] , \Level4Out52[15] , 
        \Level4Out52[14] , \Level4Out52[13] , \Level4Out52[12] , 
        \Level4Out52[11] , \Level4Out52[10] , \Level4Out52[9] , 
        \Level4Out52[8] , \Level4Out52[7] , \Level4Out52[6] , \Level4Out52[5] , 
        \Level4Out52[4] , \Level4Out52[3] , \Level4Out52[2] , \Level4Out52[1] , 
        \Level4Out52[0] }), .In1({\Level2Out52[31] , \Level2Out52[30] , 
        \Level2Out52[29] , \Level2Out52[28] , \Level2Out52[27] , 
        \Level2Out52[26] , \Level2Out52[25] , \Level2Out52[24] , 
        \Level2Out52[23] , \Level2Out52[22] , \Level2Out52[21] , 
        \Level2Out52[20] , \Level2Out52[19] , \Level2Out52[18] , 
        \Level2Out52[17] , \Level2Out52[16] , \Level2Out52[15] , 
        \Level2Out52[14] , \Level2Out52[13] , \Level2Out52[12] , 
        \Level2Out52[11] , \Level2Out52[10] , \Level2Out52[9] , 
        \Level2Out52[8] , \Level2Out52[7] , \Level2Out52[6] , \Level2Out52[5] , 
        \Level2Out52[4] , \Level2Out52[3] , \Level2Out52[2] , \Level2Out52[1] , 
        \Level2Out52[0] }), .In2({\Level2Out54[31] , \Level2Out54[30] , 
        \Level2Out54[29] , \Level2Out54[28] , \Level2Out54[27] , 
        \Level2Out54[26] , \Level2Out54[25] , \Level2Out54[24] , 
        \Level2Out54[23] , \Level2Out54[22] , \Level2Out54[21] , 
        \Level2Out54[20] , \Level2Out54[19] , \Level2Out54[18] , 
        \Level2Out54[17] , \Level2Out54[16] , \Level2Out54[15] , 
        \Level2Out54[14] , \Level2Out54[13] , \Level2Out54[12] , 
        \Level2Out54[11] , \Level2Out54[10] , \Level2Out54[9] , 
        \Level2Out54[8] , \Level2Out54[7] , \Level2Out54[6] , \Level2Out54[5] , 
        \Level2Out54[4] , \Level2Out54[3] , \Level2Out54[2] , \Level2Out54[1] , 
        \Level2Out54[0] }), .Read1(\Level2Load52[0] ), .Read2(
        \Level2Load54[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_38 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanOut({\ScanLink39[31] , 
        \ScanLink39[30] , \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , 
        \ScanLink39[26] , \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , 
        \ScanLink39[22] , \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , 
        \ScanLink39[18] , \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , 
        \ScanLink39[14] , \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , 
        \ScanLink39[10] , \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , 
        \ScanLink39[6] , \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , 
        \ScanLink39[2] , \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load38[0] ), .Out({
        \Level1Out38[31] , \Level1Out38[30] , \Level1Out38[29] , 
        \Level1Out38[28] , \Level1Out38[27] , \Level1Out38[26] , 
        \Level1Out38[25] , \Level1Out38[24] , \Level1Out38[23] , 
        \Level1Out38[22] , \Level1Out38[21] , \Level1Out38[20] , 
        \Level1Out38[19] , \Level1Out38[18] , \Level1Out38[17] , 
        \Level1Out38[16] , \Level1Out38[15] , \Level1Out38[14] , 
        \Level1Out38[13] , \Level1Out38[12] , \Level1Out38[11] , 
        \Level1Out38[10] , \Level1Out38[9] , \Level1Out38[8] , 
        \Level1Out38[7] , \Level1Out38[6] , \Level1Out38[5] , \Level1Out38[4] , 
        \Level1Out38[3] , \Level1Out38[2] , \Level1Out38[1] , \Level1Out38[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_94 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink94[31] , \ScanLink94[30] , 
        \ScanLink94[29] , \ScanLink94[28] , \ScanLink94[27] , \ScanLink94[26] , 
        \ScanLink94[25] , \ScanLink94[24] , \ScanLink94[23] , \ScanLink94[22] , 
        \ScanLink94[21] , \ScanLink94[20] , \ScanLink94[19] , \ScanLink94[18] , 
        \ScanLink94[17] , \ScanLink94[16] , \ScanLink94[15] , \ScanLink94[14] , 
        \ScanLink94[13] , \ScanLink94[12] , \ScanLink94[11] , \ScanLink94[10] , 
        \ScanLink94[9] , \ScanLink94[8] , \ScanLink94[7] , \ScanLink94[6] , 
        \ScanLink94[5] , \ScanLink94[4] , \ScanLink94[3] , \ScanLink94[2] , 
        \ScanLink94[1] , \ScanLink94[0] }), .ScanOut({\ScanLink95[31] , 
        \ScanLink95[30] , \ScanLink95[29] , \ScanLink95[28] , \ScanLink95[27] , 
        \ScanLink95[26] , \ScanLink95[25] , \ScanLink95[24] , \ScanLink95[23] , 
        \ScanLink95[22] , \ScanLink95[21] , \ScanLink95[20] , \ScanLink95[19] , 
        \ScanLink95[18] , \ScanLink95[17] , \ScanLink95[16] , \ScanLink95[15] , 
        \ScanLink95[14] , \ScanLink95[13] , \ScanLink95[12] , \ScanLink95[11] , 
        \ScanLink95[10] , \ScanLink95[9] , \ScanLink95[8] , \ScanLink95[7] , 
        \ScanLink95[6] , \ScanLink95[5] , \ScanLink95[4] , \ScanLink95[3] , 
        \ScanLink95[2] , \ScanLink95[1] , \ScanLink95[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load94[0] ), .Out({
        \Level1Out94[31] , \Level1Out94[30] , \Level1Out94[29] , 
        \Level1Out94[28] , \Level1Out94[27] , \Level1Out94[26] , 
        \Level1Out94[25] , \Level1Out94[24] , \Level1Out94[23] , 
        \Level1Out94[22] , \Level1Out94[21] , \Level1Out94[20] , 
        \Level1Out94[19] , \Level1Out94[18] , \Level1Out94[17] , 
        \Level1Out94[16] , \Level1Out94[15] , \Level1Out94[14] , 
        \Level1Out94[13] , \Level1Out94[12] , \Level1Out94[11] , 
        \Level1Out94[10] , \Level1Out94[9] , \Level1Out94[8] , 
        \Level1Out94[7] , \Level1Out94[6] , \Level1Out94[5] , \Level1Out94[4] , 
        \Level1Out94[3] , \Level1Out94[2] , \Level1Out94[1] , \Level1Out94[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_196 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink196[31] , \ScanLink196[30] , 
        \ScanLink196[29] , \ScanLink196[28] , \ScanLink196[27] , 
        \ScanLink196[26] , \ScanLink196[25] , \ScanLink196[24] , 
        \ScanLink196[23] , \ScanLink196[22] , \ScanLink196[21] , 
        \ScanLink196[20] , \ScanLink196[19] , \ScanLink196[18] , 
        \ScanLink196[17] , \ScanLink196[16] , \ScanLink196[15] , 
        \ScanLink196[14] , \ScanLink196[13] , \ScanLink196[12] , 
        \ScanLink196[11] , \ScanLink196[10] , \ScanLink196[9] , 
        \ScanLink196[8] , \ScanLink196[7] , \ScanLink196[6] , \ScanLink196[5] , 
        \ScanLink196[4] , \ScanLink196[3] , \ScanLink196[2] , \ScanLink196[1] , 
        \ScanLink196[0] }), .ScanOut({\ScanLink197[31] , \ScanLink197[30] , 
        \ScanLink197[29] , \ScanLink197[28] , \ScanLink197[27] , 
        \ScanLink197[26] , \ScanLink197[25] , \ScanLink197[24] , 
        \ScanLink197[23] , \ScanLink197[22] , \ScanLink197[21] , 
        \ScanLink197[20] , \ScanLink197[19] , \ScanLink197[18] , 
        \ScanLink197[17] , \ScanLink197[16] , \ScanLink197[15] , 
        \ScanLink197[14] , \ScanLink197[13] , \ScanLink197[12] , 
        \ScanLink197[11] , \ScanLink197[10] , \ScanLink197[9] , 
        \ScanLink197[8] , \ScanLink197[7] , \ScanLink197[6] , \ScanLink197[5] , 
        \ScanLink197[4] , \ScanLink197[3] , \ScanLink197[2] , \ScanLink197[1] , 
        \ScanLink197[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load196[0] ), .Out({\Level1Out196[31] , \Level1Out196[30] , 
        \Level1Out196[29] , \Level1Out196[28] , \Level1Out196[27] , 
        \Level1Out196[26] , \Level1Out196[25] , \Level1Out196[24] , 
        \Level1Out196[23] , \Level1Out196[22] , \Level1Out196[21] , 
        \Level1Out196[20] , \Level1Out196[19] , \Level1Out196[18] , 
        \Level1Out196[17] , \Level1Out196[16] , \Level1Out196[15] , 
        \Level1Out196[14] , \Level1Out196[13] , \Level1Out196[12] , 
        \Level1Out196[11] , \Level1Out196[10] , \Level1Out196[9] , 
        \Level1Out196[8] , \Level1Out196[7] , \Level1Out196[6] , 
        \Level1Out196[5] , \Level1Out196[4] , \Level1Out196[3] , 
        \Level1Out196[2] , \Level1Out196[1] , \Level1Out196[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_64_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load64[0] ), .Out({\Level2Out64[31] , \Level2Out64[30] , 
        \Level2Out64[29] , \Level2Out64[28] , \Level2Out64[27] , 
        \Level2Out64[26] , \Level2Out64[25] , \Level2Out64[24] , 
        \Level2Out64[23] , \Level2Out64[22] , \Level2Out64[21] , 
        \Level2Out64[20] , \Level2Out64[19] , \Level2Out64[18] , 
        \Level2Out64[17] , \Level2Out64[16] , \Level2Out64[15] , 
        \Level2Out64[14] , \Level2Out64[13] , \Level2Out64[12] , 
        \Level2Out64[11] , \Level2Out64[10] , \Level2Out64[9] , 
        \Level2Out64[8] , \Level2Out64[7] , \Level2Out64[6] , \Level2Out64[5] , 
        \Level2Out64[4] , \Level2Out64[3] , \Level2Out64[2] , \Level2Out64[1] , 
        \Level2Out64[0] }), .In1({\Level1Out64[31] , \Level1Out64[30] , 
        \Level1Out64[29] , \Level1Out64[28] , \Level1Out64[27] , 
        \Level1Out64[26] , \Level1Out64[25] , \Level1Out64[24] , 
        \Level1Out64[23] , \Level1Out64[22] , \Level1Out64[21] , 
        \Level1Out64[20] , \Level1Out64[19] , \Level1Out64[18] , 
        \Level1Out64[17] , \Level1Out64[16] , \Level1Out64[15] , 
        \Level1Out64[14] , \Level1Out64[13] , \Level1Out64[12] , 
        \Level1Out64[11] , \Level1Out64[10] , \Level1Out64[9] , 
        \Level1Out64[8] , \Level1Out64[7] , \Level1Out64[6] , \Level1Out64[5] , 
        \Level1Out64[4] , \Level1Out64[3] , \Level1Out64[2] , \Level1Out64[1] , 
        \Level1Out64[0] }), .In2({\Level1Out65[31] , \Level1Out65[30] , 
        \Level1Out65[29] , \Level1Out65[28] , \Level1Out65[27] , 
        \Level1Out65[26] , \Level1Out65[25] , \Level1Out65[24] , 
        \Level1Out65[23] , \Level1Out65[22] , \Level1Out65[21] , 
        \Level1Out65[20] , \Level1Out65[19] , \Level1Out65[18] , 
        \Level1Out65[17] , \Level1Out65[16] , \Level1Out65[15] , 
        \Level1Out65[14] , \Level1Out65[13] , \Level1Out65[12] , 
        \Level1Out65[11] , \Level1Out65[10] , \Level1Out65[9] , 
        \Level1Out65[8] , \Level1Out65[7] , \Level1Out65[6] , \Level1Out65[5] , 
        \Level1Out65[4] , \Level1Out65[3] , \Level1Out65[2] , \Level1Out65[1] , 
        \Level1Out65[0] }), .Read1(\Level1Load64[0] ), .Read2(
        \Level1Load65[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_108_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load108[0] ), .Out({\Level2Out108[31] , \Level2Out108[30] , 
        \Level2Out108[29] , \Level2Out108[28] , \Level2Out108[27] , 
        \Level2Out108[26] , \Level2Out108[25] , \Level2Out108[24] , 
        \Level2Out108[23] , \Level2Out108[22] , \Level2Out108[21] , 
        \Level2Out108[20] , \Level2Out108[19] , \Level2Out108[18] , 
        \Level2Out108[17] , \Level2Out108[16] , \Level2Out108[15] , 
        \Level2Out108[14] , \Level2Out108[13] , \Level2Out108[12] , 
        \Level2Out108[11] , \Level2Out108[10] , \Level2Out108[9] , 
        \Level2Out108[8] , \Level2Out108[7] , \Level2Out108[6] , 
        \Level2Out108[5] , \Level2Out108[4] , \Level2Out108[3] , 
        \Level2Out108[2] , \Level2Out108[1] , \Level2Out108[0] }), .In1({
        \Level1Out108[31] , \Level1Out108[30] , \Level1Out108[29] , 
        \Level1Out108[28] , \Level1Out108[27] , \Level1Out108[26] , 
        \Level1Out108[25] , \Level1Out108[24] , \Level1Out108[23] , 
        \Level1Out108[22] , \Level1Out108[21] , \Level1Out108[20] , 
        \Level1Out108[19] , \Level1Out108[18] , \Level1Out108[17] , 
        \Level1Out108[16] , \Level1Out108[15] , \Level1Out108[14] , 
        \Level1Out108[13] , \Level1Out108[12] , \Level1Out108[11] , 
        \Level1Out108[10] , \Level1Out108[9] , \Level1Out108[8] , 
        \Level1Out108[7] , \Level1Out108[6] , \Level1Out108[5] , 
        \Level1Out108[4] , \Level1Out108[3] , \Level1Out108[2] , 
        \Level1Out108[1] , \Level1Out108[0] }), .In2({\Level1Out109[31] , 
        \Level1Out109[30] , \Level1Out109[29] , \Level1Out109[28] , 
        \Level1Out109[27] , \Level1Out109[26] , \Level1Out109[25] , 
        \Level1Out109[24] , \Level1Out109[23] , \Level1Out109[22] , 
        \Level1Out109[21] , \Level1Out109[20] , \Level1Out109[19] , 
        \Level1Out109[18] , \Level1Out109[17] , \Level1Out109[16] , 
        \Level1Out109[15] , \Level1Out109[14] , \Level1Out109[13] , 
        \Level1Out109[12] , \Level1Out109[11] , \Level1Out109[10] , 
        \Level1Out109[9] , \Level1Out109[8] , \Level1Out109[7] , 
        \Level1Out109[6] , \Level1Out109[5] , \Level1Out109[4] , 
        \Level1Out109[3] , \Level1Out109[2] , \Level1Out109[1] , 
        \Level1Out109[0] }), .Read1(\Level1Load108[0] ), .Read2(
        \Level1Load109[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_216_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load216[0] ), .Out({\Level2Out216[31] , \Level2Out216[30] , 
        \Level2Out216[29] , \Level2Out216[28] , \Level2Out216[27] , 
        \Level2Out216[26] , \Level2Out216[25] , \Level2Out216[24] , 
        \Level2Out216[23] , \Level2Out216[22] , \Level2Out216[21] , 
        \Level2Out216[20] , \Level2Out216[19] , \Level2Out216[18] , 
        \Level2Out216[17] , \Level2Out216[16] , \Level2Out216[15] , 
        \Level2Out216[14] , \Level2Out216[13] , \Level2Out216[12] , 
        \Level2Out216[11] , \Level2Out216[10] , \Level2Out216[9] , 
        \Level2Out216[8] , \Level2Out216[7] , \Level2Out216[6] , 
        \Level2Out216[5] , \Level2Out216[4] , \Level2Out216[3] , 
        \Level2Out216[2] , \Level2Out216[1] , \Level2Out216[0] }), .In1({
        \Level1Out216[31] , \Level1Out216[30] , \Level1Out216[29] , 
        \Level1Out216[28] , \Level1Out216[27] , \Level1Out216[26] , 
        \Level1Out216[25] , \Level1Out216[24] , \Level1Out216[23] , 
        \Level1Out216[22] , \Level1Out216[21] , \Level1Out216[20] , 
        \Level1Out216[19] , \Level1Out216[18] , \Level1Out216[17] , 
        \Level1Out216[16] , \Level1Out216[15] , \Level1Out216[14] , 
        \Level1Out216[13] , \Level1Out216[12] , \Level1Out216[11] , 
        \Level1Out216[10] , \Level1Out216[9] , \Level1Out216[8] , 
        \Level1Out216[7] , \Level1Out216[6] , \Level1Out216[5] , 
        \Level1Out216[4] , \Level1Out216[3] , \Level1Out216[2] , 
        \Level1Out216[1] , \Level1Out216[0] }), .In2({\Level1Out217[31] , 
        \Level1Out217[30] , \Level1Out217[29] , \Level1Out217[28] , 
        \Level1Out217[27] , \Level1Out217[26] , \Level1Out217[25] , 
        \Level1Out217[24] , \Level1Out217[23] , \Level1Out217[22] , 
        \Level1Out217[21] , \Level1Out217[20] , \Level1Out217[19] , 
        \Level1Out217[18] , \Level1Out217[17] , \Level1Out217[16] , 
        \Level1Out217[15] , \Level1Out217[14] , \Level1Out217[13] , 
        \Level1Out217[12] , \Level1Out217[11] , \Level1Out217[10] , 
        \Level1Out217[9] , \Level1Out217[8] , \Level1Out217[7] , 
        \Level1Out217[6] , \Level1Out217[5] , \Level1Out217[4] , 
        \Level1Out217[3] , \Level1Out217[2] , \Level1Out217[1] , 
        \Level1Out217[0] }), .Read1(\Level1Load216[0] ), .Read2(
        \Level1Load217[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_191 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink191[31] , \ScanLink191[30] , 
        \ScanLink191[29] , \ScanLink191[28] , \ScanLink191[27] , 
        \ScanLink191[26] , \ScanLink191[25] , \ScanLink191[24] , 
        \ScanLink191[23] , \ScanLink191[22] , \ScanLink191[21] , 
        \ScanLink191[20] , \ScanLink191[19] , \ScanLink191[18] , 
        \ScanLink191[17] , \ScanLink191[16] , \ScanLink191[15] , 
        \ScanLink191[14] , \ScanLink191[13] , \ScanLink191[12] , 
        \ScanLink191[11] , \ScanLink191[10] , \ScanLink191[9] , 
        \ScanLink191[8] , \ScanLink191[7] , \ScanLink191[6] , \ScanLink191[5] , 
        \ScanLink191[4] , \ScanLink191[3] , \ScanLink191[2] , \ScanLink191[1] , 
        \ScanLink191[0] }), .ScanOut({\ScanLink192[31] , \ScanLink192[30] , 
        \ScanLink192[29] , \ScanLink192[28] , \ScanLink192[27] , 
        \ScanLink192[26] , \ScanLink192[25] , \ScanLink192[24] , 
        \ScanLink192[23] , \ScanLink192[22] , \ScanLink192[21] , 
        \ScanLink192[20] , \ScanLink192[19] , \ScanLink192[18] , 
        \ScanLink192[17] , \ScanLink192[16] , \ScanLink192[15] , 
        \ScanLink192[14] , \ScanLink192[13] , \ScanLink192[12] , 
        \ScanLink192[11] , \ScanLink192[10] , \ScanLink192[9] , 
        \ScanLink192[8] , \ScanLink192[7] , \ScanLink192[6] , \ScanLink192[5] , 
        \ScanLink192[4] , \ScanLink192[3] , \ScanLink192[2] , \ScanLink192[1] , 
        \ScanLink192[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load191[0] ), .Out({\Level1Out191[31] , \Level1Out191[30] , 
        \Level1Out191[29] , \Level1Out191[28] , \Level1Out191[27] , 
        \Level1Out191[26] , \Level1Out191[25] , \Level1Out191[24] , 
        \Level1Out191[23] , \Level1Out191[22] , \Level1Out191[21] , 
        \Level1Out191[20] , \Level1Out191[19] , \Level1Out191[18] , 
        \Level1Out191[17] , \Level1Out191[16] , \Level1Out191[15] , 
        \Level1Out191[14] , \Level1Out191[13] , \Level1Out191[12] , 
        \Level1Out191[11] , \Level1Out191[10] , \Level1Out191[9] , 
        \Level1Out191[8] , \Level1Out191[7] , \Level1Out191[6] , 
        \Level1Out191[5] , \Level1Out191[4] , \Level1Out191[3] , 
        \Level1Out191[2] , \Level1Out191[1] , \Level1Out191[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_224_32 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load224[0] ), .Out({\Level32Out224[31] , \Level32Out224[30] , 
        \Level32Out224[29] , \Level32Out224[28] , \Level32Out224[27] , 
        \Level32Out224[26] , \Level32Out224[25] , \Level32Out224[24] , 
        \Level32Out224[23] , \Level32Out224[22] , \Level32Out224[21] , 
        \Level32Out224[20] , \Level32Out224[19] , \Level32Out224[18] , 
        \Level32Out224[17] , \Level32Out224[16] , \Level32Out224[15] , 
        \Level32Out224[14] , \Level32Out224[13] , \Level32Out224[12] , 
        \Level32Out224[11] , \Level32Out224[10] , \Level32Out224[9] , 
        \Level32Out224[8] , \Level32Out224[7] , \Level32Out224[6] , 
        \Level32Out224[5] , \Level32Out224[4] , \Level32Out224[3] , 
        \Level32Out224[2] , \Level32Out224[1] , \Level32Out224[0] }), .In1({
        \Level16Out224[31] , \Level16Out224[30] , \Level16Out224[29] , 
        \Level16Out224[28] , \Level16Out224[27] , \Level16Out224[26] , 
        \Level16Out224[25] , \Level16Out224[24] , \Level16Out224[23] , 
        \Level16Out224[22] , \Level16Out224[21] , \Level16Out224[20] , 
        \Level16Out224[19] , \Level16Out224[18] , \Level16Out224[17] , 
        \Level16Out224[16] , \Level16Out224[15] , \Level16Out224[14] , 
        \Level16Out224[13] , \Level16Out224[12] , \Level16Out224[11] , 
        \Level16Out224[10] , \Level16Out224[9] , \Level16Out224[8] , 
        \Level16Out224[7] , \Level16Out224[6] , \Level16Out224[5] , 
        \Level16Out224[4] , \Level16Out224[3] , \Level16Out224[2] , 
        \Level16Out224[1] , \Level16Out224[0] }), .In2({\Level16Out240[31] , 
        \Level16Out240[30] , \Level16Out240[29] , \Level16Out240[28] , 
        \Level16Out240[27] , \Level16Out240[26] , \Level16Out240[25] , 
        \Level16Out240[24] , \Level16Out240[23] , \Level16Out240[22] , 
        \Level16Out240[21] , \Level16Out240[20] , \Level16Out240[19] , 
        \Level16Out240[18] , \Level16Out240[17] , \Level16Out240[16] , 
        \Level16Out240[15] , \Level16Out240[14] , \Level16Out240[13] , 
        \Level16Out240[12] , \Level16Out240[11] , \Level16Out240[10] , 
        \Level16Out240[9] , \Level16Out240[8] , \Level16Out240[7] , 
        \Level16Out240[6] , \Level16Out240[5] , \Level16Out240[4] , 
        \Level16Out240[3] , \Level16Out240[2] , \Level16Out240[1] , 
        \Level16Out240[0] }), .Read1(\Level16Load224[0] ), .Read2(
        \Level16Load240[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_56 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanOut({\ScanLink57[31] , 
        \ScanLink57[30] , \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , 
        \ScanLink57[26] , \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , 
        \ScanLink57[22] , \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , 
        \ScanLink57[18] , \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , 
        \ScanLink57[14] , \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , 
        \ScanLink57[10] , \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , 
        \ScanLink57[6] , \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , 
        \ScanLink57[2] , \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load56[0] ), .Out({
        \Level1Out56[31] , \Level1Out56[30] , \Level1Out56[29] , 
        \Level1Out56[28] , \Level1Out56[27] , \Level1Out56[26] , 
        \Level1Out56[25] , \Level1Out56[24] , \Level1Out56[23] , 
        \Level1Out56[22] , \Level1Out56[21] , \Level1Out56[20] , 
        \Level1Out56[19] , \Level1Out56[18] , \Level1Out56[17] , 
        \Level1Out56[16] , \Level1Out56[15] , \Level1Out56[14] , 
        \Level1Out56[13] , \Level1Out56[12] , \Level1Out56[11] , 
        \Level1Out56[10] , \Level1Out56[9] , \Level1Out56[8] , 
        \Level1Out56[7] , \Level1Out56[6] , \Level1Out56[5] , \Level1Out56[4] , 
        \Level1Out56[3] , \Level1Out56[2] , \Level1Out56[1] , \Level1Out56[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load2[0] ), .Out({\Level2Out2[31] , \Level2Out2[30] , 
        \Level2Out2[29] , \Level2Out2[28] , \Level2Out2[27] , \Level2Out2[26] , 
        \Level2Out2[25] , \Level2Out2[24] , \Level2Out2[23] , \Level2Out2[22] , 
        \Level2Out2[21] , \Level2Out2[20] , \Level2Out2[19] , \Level2Out2[18] , 
        \Level2Out2[17] , \Level2Out2[16] , \Level2Out2[15] , \Level2Out2[14] , 
        \Level2Out2[13] , \Level2Out2[12] , \Level2Out2[11] , \Level2Out2[10] , 
        \Level2Out2[9] , \Level2Out2[8] , \Level2Out2[7] , \Level2Out2[6] , 
        \Level2Out2[5] , \Level2Out2[4] , \Level2Out2[3] , \Level2Out2[2] , 
        \Level2Out2[1] , \Level2Out2[0] }), .In1({\Level1Out2[31] , 
        \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , \Level1Out2[27] , 
        \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , \Level1Out2[23] , 
        \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , \Level1Out2[19] , 
        \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , \Level1Out2[15] , 
        \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , \Level1Out2[11] , 
        \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , \Level1Out2[7] , 
        \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , \Level1Out2[3] , 
        \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] }), .In2({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] }), 
        .Read1(\Level1Load2[0] ), .Read2(\Level1Load3[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_71 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink71[31] , \ScanLink71[30] , 
        \ScanLink71[29] , \ScanLink71[28] , \ScanLink71[27] , \ScanLink71[26] , 
        \ScanLink71[25] , \ScanLink71[24] , \ScanLink71[23] , \ScanLink71[22] , 
        \ScanLink71[21] , \ScanLink71[20] , \ScanLink71[19] , \ScanLink71[18] , 
        \ScanLink71[17] , \ScanLink71[16] , \ScanLink71[15] , \ScanLink71[14] , 
        \ScanLink71[13] , \ScanLink71[12] , \ScanLink71[11] , \ScanLink71[10] , 
        \ScanLink71[9] , \ScanLink71[8] , \ScanLink71[7] , \ScanLink71[6] , 
        \ScanLink71[5] , \ScanLink71[4] , \ScanLink71[3] , \ScanLink71[2] , 
        \ScanLink71[1] , \ScanLink71[0] }), .ScanOut({\ScanLink72[31] , 
        \ScanLink72[30] , \ScanLink72[29] , \ScanLink72[28] , \ScanLink72[27] , 
        \ScanLink72[26] , \ScanLink72[25] , \ScanLink72[24] , \ScanLink72[23] , 
        \ScanLink72[22] , \ScanLink72[21] , \ScanLink72[20] , \ScanLink72[19] , 
        \ScanLink72[18] , \ScanLink72[17] , \ScanLink72[16] , \ScanLink72[15] , 
        \ScanLink72[14] , \ScanLink72[13] , \ScanLink72[12] , \ScanLink72[11] , 
        \ScanLink72[10] , \ScanLink72[9] , \ScanLink72[8] , \ScanLink72[7] , 
        \ScanLink72[6] , \ScanLink72[5] , \ScanLink72[4] , \ScanLink72[3] , 
        \ScanLink72[2] , \ScanLink72[1] , \ScanLink72[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load71[0] ), .Out({
        \Level1Out71[31] , \Level1Out71[30] , \Level1Out71[29] , 
        \Level1Out71[28] , \Level1Out71[27] , \Level1Out71[26] , 
        \Level1Out71[25] , \Level1Out71[24] , \Level1Out71[23] , 
        \Level1Out71[22] , \Level1Out71[21] , \Level1Out71[20] , 
        \Level1Out71[19] , \Level1Out71[18] , \Level1Out71[17] , 
        \Level1Out71[16] , \Level1Out71[15] , \Level1Out71[14] , 
        \Level1Out71[13] , \Level1Out71[12] , \Level1Out71[11] , 
        \Level1Out71[10] , \Level1Out71[9] , \Level1Out71[8] , 
        \Level1Out71[7] , \Level1Out71[6] , \Level1Out71[5] , \Level1Out71[4] , 
        \Level1Out71[3] , \Level1Out71[2] , \Level1Out71[1] , \Level1Out71[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_196_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load196[0] ), .Out({\Level4Out196[31] , \Level4Out196[30] , 
        \Level4Out196[29] , \Level4Out196[28] , \Level4Out196[27] , 
        \Level4Out196[26] , \Level4Out196[25] , \Level4Out196[24] , 
        \Level4Out196[23] , \Level4Out196[22] , \Level4Out196[21] , 
        \Level4Out196[20] , \Level4Out196[19] , \Level4Out196[18] , 
        \Level4Out196[17] , \Level4Out196[16] , \Level4Out196[15] , 
        \Level4Out196[14] , \Level4Out196[13] , \Level4Out196[12] , 
        \Level4Out196[11] , \Level4Out196[10] , \Level4Out196[9] , 
        \Level4Out196[8] , \Level4Out196[7] , \Level4Out196[6] , 
        \Level4Out196[5] , \Level4Out196[4] , \Level4Out196[3] , 
        \Level4Out196[2] , \Level4Out196[1] , \Level4Out196[0] }), .In1({
        \Level2Out196[31] , \Level2Out196[30] , \Level2Out196[29] , 
        \Level2Out196[28] , \Level2Out196[27] , \Level2Out196[26] , 
        \Level2Out196[25] , \Level2Out196[24] , \Level2Out196[23] , 
        \Level2Out196[22] , \Level2Out196[21] , \Level2Out196[20] , 
        \Level2Out196[19] , \Level2Out196[18] , \Level2Out196[17] , 
        \Level2Out196[16] , \Level2Out196[15] , \Level2Out196[14] , 
        \Level2Out196[13] , \Level2Out196[12] , \Level2Out196[11] , 
        \Level2Out196[10] , \Level2Out196[9] , \Level2Out196[8] , 
        \Level2Out196[7] , \Level2Out196[6] , \Level2Out196[5] , 
        \Level2Out196[4] , \Level2Out196[3] , \Level2Out196[2] , 
        \Level2Out196[1] , \Level2Out196[0] }), .In2({\Level2Out198[31] , 
        \Level2Out198[30] , \Level2Out198[29] , \Level2Out198[28] , 
        \Level2Out198[27] , \Level2Out198[26] , \Level2Out198[25] , 
        \Level2Out198[24] , \Level2Out198[23] , \Level2Out198[22] , 
        \Level2Out198[21] , \Level2Out198[20] , \Level2Out198[19] , 
        \Level2Out198[18] , \Level2Out198[17] , \Level2Out198[16] , 
        \Level2Out198[15] , \Level2Out198[14] , \Level2Out198[13] , 
        \Level2Out198[12] , \Level2Out198[11] , \Level2Out198[10] , 
        \Level2Out198[9] , \Level2Out198[8] , \Level2Out198[7] , 
        \Level2Out198[6] , \Level2Out198[5] , \Level2Out198[4] , 
        \Level2Out198[3] , \Level2Out198[2] , \Level2Out198[1] , 
        \Level2Out198[0] }), .Read1(\Level2Load196[0] ), .Read2(
        \Level2Load198[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load128[0] ), .Out({\Level8Out128[31] , \Level8Out128[30] , 
        \Level8Out128[29] , \Level8Out128[28] , \Level8Out128[27] , 
        \Level8Out128[26] , \Level8Out128[25] , \Level8Out128[24] , 
        \Level8Out128[23] , \Level8Out128[22] , \Level8Out128[21] , 
        \Level8Out128[20] , \Level8Out128[19] , \Level8Out128[18] , 
        \Level8Out128[17] , \Level8Out128[16] , \Level8Out128[15] , 
        \Level8Out128[14] , \Level8Out128[13] , \Level8Out128[12] , 
        \Level8Out128[11] , \Level8Out128[10] , \Level8Out128[9] , 
        \Level8Out128[8] , \Level8Out128[7] , \Level8Out128[6] , 
        \Level8Out128[5] , \Level8Out128[4] , \Level8Out128[3] , 
        \Level8Out128[2] , \Level8Out128[1] , \Level8Out128[0] }), .In1({
        \Level4Out128[31] , \Level4Out128[30] , \Level4Out128[29] , 
        \Level4Out128[28] , \Level4Out128[27] , \Level4Out128[26] , 
        \Level4Out128[25] , \Level4Out128[24] , \Level4Out128[23] , 
        \Level4Out128[22] , \Level4Out128[21] , \Level4Out128[20] , 
        \Level4Out128[19] , \Level4Out128[18] , \Level4Out128[17] , 
        \Level4Out128[16] , \Level4Out128[15] , \Level4Out128[14] , 
        \Level4Out128[13] , \Level4Out128[12] , \Level4Out128[11] , 
        \Level4Out128[10] , \Level4Out128[9] , \Level4Out128[8] , 
        \Level4Out128[7] , \Level4Out128[6] , \Level4Out128[5] , 
        \Level4Out128[4] , \Level4Out128[3] , \Level4Out128[2] , 
        \Level4Out128[1] , \Level4Out128[0] }), .In2({\Level4Out132[31] , 
        \Level4Out132[30] , \Level4Out132[29] , \Level4Out132[28] , 
        \Level4Out132[27] , \Level4Out132[26] , \Level4Out132[25] , 
        \Level4Out132[24] , \Level4Out132[23] , \Level4Out132[22] , 
        \Level4Out132[21] , \Level4Out132[20] , \Level4Out132[19] , 
        \Level4Out132[18] , \Level4Out132[17] , \Level4Out132[16] , 
        \Level4Out132[15] , \Level4Out132[14] , \Level4Out132[13] , 
        \Level4Out132[12] , \Level4Out132[11] , \Level4Out132[10] , 
        \Level4Out132[9] , \Level4Out132[8] , \Level4Out132[7] , 
        \Level4Out132[6] , \Level4Out132[5] , \Level4Out132[4] , 
        \Level4Out132[3] , \Level4Out132[2] , \Level4Out132[1] , 
        \Level4Out132[0] }), .Read1(\Level4Load128[0] ), .Read2(
        \Level4Load132[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_64 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level64Load192[0] ), .Out({\Level64Out192[31] , \Level64Out192[30] , 
        \Level64Out192[29] , \Level64Out192[28] , \Level64Out192[27] , 
        \Level64Out192[26] , \Level64Out192[25] , \Level64Out192[24] , 
        \Level64Out192[23] , \Level64Out192[22] , \Level64Out192[21] , 
        \Level64Out192[20] , \Level64Out192[19] , \Level64Out192[18] , 
        \Level64Out192[17] , \Level64Out192[16] , \Level64Out192[15] , 
        \Level64Out192[14] , \Level64Out192[13] , \Level64Out192[12] , 
        \Level64Out192[11] , \Level64Out192[10] , \Level64Out192[9] , 
        \Level64Out192[8] , \Level64Out192[7] , \Level64Out192[6] , 
        \Level64Out192[5] , \Level64Out192[4] , \Level64Out192[3] , 
        \Level64Out192[2] , \Level64Out192[1] , \Level64Out192[0] }), .In1({
        \Level32Out192[31] , \Level32Out192[30] , \Level32Out192[29] , 
        \Level32Out192[28] , \Level32Out192[27] , \Level32Out192[26] , 
        \Level32Out192[25] , \Level32Out192[24] , \Level32Out192[23] , 
        \Level32Out192[22] , \Level32Out192[21] , \Level32Out192[20] , 
        \Level32Out192[19] , \Level32Out192[18] , \Level32Out192[17] , 
        \Level32Out192[16] , \Level32Out192[15] , \Level32Out192[14] , 
        \Level32Out192[13] , \Level32Out192[12] , \Level32Out192[11] , 
        \Level32Out192[10] , \Level32Out192[9] , \Level32Out192[8] , 
        \Level32Out192[7] , \Level32Out192[6] , \Level32Out192[5] , 
        \Level32Out192[4] , \Level32Out192[3] , \Level32Out192[2] , 
        \Level32Out192[1] , \Level32Out192[0] }), .In2({\Level32Out224[31] , 
        \Level32Out224[30] , \Level32Out224[29] , \Level32Out224[28] , 
        \Level32Out224[27] , \Level32Out224[26] , \Level32Out224[25] , 
        \Level32Out224[24] , \Level32Out224[23] , \Level32Out224[22] , 
        \Level32Out224[21] , \Level32Out224[20] , \Level32Out224[19] , 
        \Level32Out224[18] , \Level32Out224[17] , \Level32Out224[16] , 
        \Level32Out224[15] , \Level32Out224[14] , \Level32Out224[13] , 
        \Level32Out224[12] , \Level32Out224[11] , \Level32Out224[10] , 
        \Level32Out224[9] , \Level32Out224[8] , \Level32Out224[7] , 
        \Level32Out224[6] , \Level32Out224[5] , \Level32Out224[4] , 
        \Level32Out224[3] , \Level32Out224[2] , \Level32Out224[1] , 
        \Level32Out224[0] }), .Read1(\Level32Load192[0] ), .Read2(
        \Level32Load224[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_153 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink153[31] , \ScanLink153[30] , 
        \ScanLink153[29] , \ScanLink153[28] , \ScanLink153[27] , 
        \ScanLink153[26] , \ScanLink153[25] , \ScanLink153[24] , 
        \ScanLink153[23] , \ScanLink153[22] , \ScanLink153[21] , 
        \ScanLink153[20] , \ScanLink153[19] , \ScanLink153[18] , 
        \ScanLink153[17] , \ScanLink153[16] , \ScanLink153[15] , 
        \ScanLink153[14] , \ScanLink153[13] , \ScanLink153[12] , 
        \ScanLink153[11] , \ScanLink153[10] , \ScanLink153[9] , 
        \ScanLink153[8] , \ScanLink153[7] , \ScanLink153[6] , \ScanLink153[5] , 
        \ScanLink153[4] , \ScanLink153[3] , \ScanLink153[2] , \ScanLink153[1] , 
        \ScanLink153[0] }), .ScanOut({\ScanLink154[31] , \ScanLink154[30] , 
        \ScanLink154[29] , \ScanLink154[28] , \ScanLink154[27] , 
        \ScanLink154[26] , \ScanLink154[25] , \ScanLink154[24] , 
        \ScanLink154[23] , \ScanLink154[22] , \ScanLink154[21] , 
        \ScanLink154[20] , \ScanLink154[19] , \ScanLink154[18] , 
        \ScanLink154[17] , \ScanLink154[16] , \ScanLink154[15] , 
        \ScanLink154[14] , \ScanLink154[13] , \ScanLink154[12] , 
        \ScanLink154[11] , \ScanLink154[10] , \ScanLink154[9] , 
        \ScanLink154[8] , \ScanLink154[7] , \ScanLink154[6] , \ScanLink154[5] , 
        \ScanLink154[4] , \ScanLink154[3] , \ScanLink154[2] , \ScanLink154[1] , 
        \ScanLink154[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load153[0] ), .Out({\Level1Out153[31] , \Level1Out153[30] , 
        \Level1Out153[29] , \Level1Out153[28] , \Level1Out153[27] , 
        \Level1Out153[26] , \Level1Out153[25] , \Level1Out153[24] , 
        \Level1Out153[23] , \Level1Out153[22] , \Level1Out153[21] , 
        \Level1Out153[20] , \Level1Out153[19] , \Level1Out153[18] , 
        \Level1Out153[17] , \Level1Out153[16] , \Level1Out153[15] , 
        \Level1Out153[14] , \Level1Out153[13] , \Level1Out153[12] , 
        \Level1Out153[11] , \Level1Out153[10] , \Level1Out153[9] , 
        \Level1Out153[8] , \Level1Out153[7] , \Level1Out153[6] , 
        \Level1Out153[5] , \Level1Out153[4] , \Level1Out153[3] , 
        \Level1Out153[2] , \Level1Out153[1] , \Level1Out153[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_202_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load202[0] ), .Out({\Level2Out202[31] , \Level2Out202[30] , 
        \Level2Out202[29] , \Level2Out202[28] , \Level2Out202[27] , 
        \Level2Out202[26] , \Level2Out202[25] , \Level2Out202[24] , 
        \Level2Out202[23] , \Level2Out202[22] , \Level2Out202[21] , 
        \Level2Out202[20] , \Level2Out202[19] , \Level2Out202[18] , 
        \Level2Out202[17] , \Level2Out202[16] , \Level2Out202[15] , 
        \Level2Out202[14] , \Level2Out202[13] , \Level2Out202[12] , 
        \Level2Out202[11] , \Level2Out202[10] , \Level2Out202[9] , 
        \Level2Out202[8] , \Level2Out202[7] , \Level2Out202[6] , 
        \Level2Out202[5] , \Level2Out202[4] , \Level2Out202[3] , 
        \Level2Out202[2] , \Level2Out202[1] , \Level2Out202[0] }), .In1({
        \Level1Out202[31] , \Level1Out202[30] , \Level1Out202[29] , 
        \Level1Out202[28] , \Level1Out202[27] , \Level1Out202[26] , 
        \Level1Out202[25] , \Level1Out202[24] , \Level1Out202[23] , 
        \Level1Out202[22] , \Level1Out202[21] , \Level1Out202[20] , 
        \Level1Out202[19] , \Level1Out202[18] , \Level1Out202[17] , 
        \Level1Out202[16] , \Level1Out202[15] , \Level1Out202[14] , 
        \Level1Out202[13] , \Level1Out202[12] , \Level1Out202[11] , 
        \Level1Out202[10] , \Level1Out202[9] , \Level1Out202[8] , 
        \Level1Out202[7] , \Level1Out202[6] , \Level1Out202[5] , 
        \Level1Out202[4] , \Level1Out202[3] , \Level1Out202[2] , 
        \Level1Out202[1] , \Level1Out202[0] }), .In2({\Level1Out203[31] , 
        \Level1Out203[30] , \Level1Out203[29] , \Level1Out203[28] , 
        \Level1Out203[27] , \Level1Out203[26] , \Level1Out203[25] , 
        \Level1Out203[24] , \Level1Out203[23] , \Level1Out203[22] , 
        \Level1Out203[21] , \Level1Out203[20] , \Level1Out203[19] , 
        \Level1Out203[18] , \Level1Out203[17] , \Level1Out203[16] , 
        \Level1Out203[15] , \Level1Out203[14] , \Level1Out203[13] , 
        \Level1Out203[12] , \Level1Out203[11] , \Level1Out203[10] , 
        \Level1Out203[9] , \Level1Out203[8] , \Level1Out203[7] , 
        \Level1Out203[6] , \Level1Out203[5] , \Level1Out203[4] , 
        \Level1Out203[3] , \Level1Out203[2] , \Level1Out203[1] , 
        \Level1Out203[0] }), .Read1(\Level1Load202[0] ), .Read2(
        \Level1Load203[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_174 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink174[31] , \ScanLink174[30] , 
        \ScanLink174[29] , \ScanLink174[28] , \ScanLink174[27] , 
        \ScanLink174[26] , \ScanLink174[25] , \ScanLink174[24] , 
        \ScanLink174[23] , \ScanLink174[22] , \ScanLink174[21] , 
        \ScanLink174[20] , \ScanLink174[19] , \ScanLink174[18] , 
        \ScanLink174[17] , \ScanLink174[16] , \ScanLink174[15] , 
        \ScanLink174[14] , \ScanLink174[13] , \ScanLink174[12] , 
        \ScanLink174[11] , \ScanLink174[10] , \ScanLink174[9] , 
        \ScanLink174[8] , \ScanLink174[7] , \ScanLink174[6] , \ScanLink174[5] , 
        \ScanLink174[4] , \ScanLink174[3] , \ScanLink174[2] , \ScanLink174[1] , 
        \ScanLink174[0] }), .ScanOut({\ScanLink175[31] , \ScanLink175[30] , 
        \ScanLink175[29] , \ScanLink175[28] , \ScanLink175[27] , 
        \ScanLink175[26] , \ScanLink175[25] , \ScanLink175[24] , 
        \ScanLink175[23] , \ScanLink175[22] , \ScanLink175[21] , 
        \ScanLink175[20] , \ScanLink175[19] , \ScanLink175[18] , 
        \ScanLink175[17] , \ScanLink175[16] , \ScanLink175[15] , 
        \ScanLink175[14] , \ScanLink175[13] , \ScanLink175[12] , 
        \ScanLink175[11] , \ScanLink175[10] , \ScanLink175[9] , 
        \ScanLink175[8] , \ScanLink175[7] , \ScanLink175[6] , \ScanLink175[5] , 
        \ScanLink175[4] , \ScanLink175[3] , \ScanLink175[2] , \ScanLink175[1] , 
        \ScanLink175[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load174[0] ), .Out({\Level1Out174[31] , \Level1Out174[30] , 
        \Level1Out174[29] , \Level1Out174[28] , \Level1Out174[27] , 
        \Level1Out174[26] , \Level1Out174[25] , \Level1Out174[24] , 
        \Level1Out174[23] , \Level1Out174[22] , \Level1Out174[21] , 
        \Level1Out174[20] , \Level1Out174[19] , \Level1Out174[18] , 
        \Level1Out174[17] , \Level1Out174[16] , \Level1Out174[15] , 
        \Level1Out174[14] , \Level1Out174[13] , \Level1Out174[12] , 
        \Level1Out174[11] , \Level1Out174[10] , \Level1Out174[9] , 
        \Level1Out174[8] , \Level1Out174[7] , \Level1Out174[6] , 
        \Level1Out174[5] , \Level1Out174[4] , \Level1Out174[3] , 
        \Level1Out174[2] , \Level1Out174[1] , \Level1Out174[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_244 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink244[31] , \ScanLink244[30] , 
        \ScanLink244[29] , \ScanLink244[28] , \ScanLink244[27] , 
        \ScanLink244[26] , \ScanLink244[25] , \ScanLink244[24] , 
        \ScanLink244[23] , \ScanLink244[22] , \ScanLink244[21] , 
        \ScanLink244[20] , \ScanLink244[19] , \ScanLink244[18] , 
        \ScanLink244[17] , \ScanLink244[16] , \ScanLink244[15] , 
        \ScanLink244[14] , \ScanLink244[13] , \ScanLink244[12] , 
        \ScanLink244[11] , \ScanLink244[10] , \ScanLink244[9] , 
        \ScanLink244[8] , \ScanLink244[7] , \ScanLink244[6] , \ScanLink244[5] , 
        \ScanLink244[4] , \ScanLink244[3] , \ScanLink244[2] , \ScanLink244[1] , 
        \ScanLink244[0] }), .ScanOut({\ScanLink245[31] , \ScanLink245[30] , 
        \ScanLink245[29] , \ScanLink245[28] , \ScanLink245[27] , 
        \ScanLink245[26] , \ScanLink245[25] , \ScanLink245[24] , 
        \ScanLink245[23] , \ScanLink245[22] , \ScanLink245[21] , 
        \ScanLink245[20] , \ScanLink245[19] , \ScanLink245[18] , 
        \ScanLink245[17] , \ScanLink245[16] , \ScanLink245[15] , 
        \ScanLink245[14] , \ScanLink245[13] , \ScanLink245[12] , 
        \ScanLink245[11] , \ScanLink245[10] , \ScanLink245[9] , 
        \ScanLink245[8] , \ScanLink245[7] , \ScanLink245[6] , \ScanLink245[5] , 
        \ScanLink245[4] , \ScanLink245[3] , \ScanLink245[2] , \ScanLink245[1] , 
        \ScanLink245[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load244[0] ), .Out({\Level1Out244[31] , \Level1Out244[30] , 
        \Level1Out244[29] , \Level1Out244[28] , \Level1Out244[27] , 
        \Level1Out244[26] , \Level1Out244[25] , \Level1Out244[24] , 
        \Level1Out244[23] , \Level1Out244[22] , \Level1Out244[21] , 
        \Level1Out244[20] , \Level1Out244[19] , \Level1Out244[18] , 
        \Level1Out244[17] , \Level1Out244[16] , \Level1Out244[15] , 
        \Level1Out244[14] , \Level1Out244[13] , \Level1Out244[12] , 
        \Level1Out244[11] , \Level1Out244[10] , \Level1Out244[9] , 
        \Level1Out244[8] , \Level1Out244[7] , \Level1Out244[6] , 
        \Level1Out244[5] , \Level1Out244[4] , \Level1Out244[3] , 
        \Level1Out244[2] , \Level1Out244[1] , \Level1Out244[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_70_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load70[0] ), .Out({\Level2Out70[31] , \Level2Out70[30] , 
        \Level2Out70[29] , \Level2Out70[28] , \Level2Out70[27] , 
        \Level2Out70[26] , \Level2Out70[25] , \Level2Out70[24] , 
        \Level2Out70[23] , \Level2Out70[22] , \Level2Out70[21] , 
        \Level2Out70[20] , \Level2Out70[19] , \Level2Out70[18] , 
        \Level2Out70[17] , \Level2Out70[16] , \Level2Out70[15] , 
        \Level2Out70[14] , \Level2Out70[13] , \Level2Out70[12] , 
        \Level2Out70[11] , \Level2Out70[10] , \Level2Out70[9] , 
        \Level2Out70[8] , \Level2Out70[7] , \Level2Out70[6] , \Level2Out70[5] , 
        \Level2Out70[4] , \Level2Out70[3] , \Level2Out70[2] , \Level2Out70[1] , 
        \Level2Out70[0] }), .In1({\Level1Out70[31] , \Level1Out70[30] , 
        \Level1Out70[29] , \Level1Out70[28] , \Level1Out70[27] , 
        \Level1Out70[26] , \Level1Out70[25] , \Level1Out70[24] , 
        \Level1Out70[23] , \Level1Out70[22] , \Level1Out70[21] , 
        \Level1Out70[20] , \Level1Out70[19] , \Level1Out70[18] , 
        \Level1Out70[17] , \Level1Out70[16] , \Level1Out70[15] , 
        \Level1Out70[14] , \Level1Out70[13] , \Level1Out70[12] , 
        \Level1Out70[11] , \Level1Out70[10] , \Level1Out70[9] , 
        \Level1Out70[8] , \Level1Out70[7] , \Level1Out70[6] , \Level1Out70[5] , 
        \Level1Out70[4] , \Level1Out70[3] , \Level1Out70[2] , \Level1Out70[1] , 
        \Level1Out70[0] }), .In2({\Level1Out71[31] , \Level1Out71[30] , 
        \Level1Out71[29] , \Level1Out71[28] , \Level1Out71[27] , 
        \Level1Out71[26] , \Level1Out71[25] , \Level1Out71[24] , 
        \Level1Out71[23] , \Level1Out71[22] , \Level1Out71[21] , 
        \Level1Out71[20] , \Level1Out71[19] , \Level1Out71[18] , 
        \Level1Out71[17] , \Level1Out71[16] , \Level1Out71[15] , 
        \Level1Out71[14] , \Level1Out71[13] , \Level1Out71[12] , 
        \Level1Out71[11] , \Level1Out71[10] , \Level1Out71[9] , 
        \Level1Out71[8] , \Level1Out71[7] , \Level1Out71[6] , \Level1Out71[5] , 
        \Level1Out71[4] , \Level1Out71[3] , \Level1Out71[2] , \Level1Out71[1] , 
        \Level1Out71[0] }), .Read1(\Level1Load70[0] ), .Read2(
        \Level1Load71[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_100_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load100[0] ), .Out({\Level4Out100[31] , \Level4Out100[30] , 
        \Level4Out100[29] , \Level4Out100[28] , \Level4Out100[27] , 
        \Level4Out100[26] , \Level4Out100[25] , \Level4Out100[24] , 
        \Level4Out100[23] , \Level4Out100[22] , \Level4Out100[21] , 
        \Level4Out100[20] , \Level4Out100[19] , \Level4Out100[18] , 
        \Level4Out100[17] , \Level4Out100[16] , \Level4Out100[15] , 
        \Level4Out100[14] , \Level4Out100[13] , \Level4Out100[12] , 
        \Level4Out100[11] , \Level4Out100[10] , \Level4Out100[9] , 
        \Level4Out100[8] , \Level4Out100[7] , \Level4Out100[6] , 
        \Level4Out100[5] , \Level4Out100[4] , \Level4Out100[3] , 
        \Level4Out100[2] , \Level4Out100[1] , \Level4Out100[0] }), .In1({
        \Level2Out100[31] , \Level2Out100[30] , \Level2Out100[29] , 
        \Level2Out100[28] , \Level2Out100[27] , \Level2Out100[26] , 
        \Level2Out100[25] , \Level2Out100[24] , \Level2Out100[23] , 
        \Level2Out100[22] , \Level2Out100[21] , \Level2Out100[20] , 
        \Level2Out100[19] , \Level2Out100[18] , \Level2Out100[17] , 
        \Level2Out100[16] , \Level2Out100[15] , \Level2Out100[14] , 
        \Level2Out100[13] , \Level2Out100[12] , \Level2Out100[11] , 
        \Level2Out100[10] , \Level2Out100[9] , \Level2Out100[8] , 
        \Level2Out100[7] , \Level2Out100[6] , \Level2Out100[5] , 
        \Level2Out100[4] , \Level2Out100[3] , \Level2Out100[2] , 
        \Level2Out100[1] , \Level2Out100[0] }), .In2({\Level2Out102[31] , 
        \Level2Out102[30] , \Level2Out102[29] , \Level2Out102[28] , 
        \Level2Out102[27] , \Level2Out102[26] , \Level2Out102[25] , 
        \Level2Out102[24] , \Level2Out102[23] , \Level2Out102[22] , 
        \Level2Out102[21] , \Level2Out102[20] , \Level2Out102[19] , 
        \Level2Out102[18] , \Level2Out102[17] , \Level2Out102[16] , 
        \Level2Out102[15] , \Level2Out102[14] , \Level2Out102[13] , 
        \Level2Out102[12] , \Level2Out102[11] , \Level2Out102[10] , 
        \Level2Out102[9] , \Level2Out102[8] , \Level2Out102[7] , 
        \Level2Out102[6] , \Level2Out102[5] , \Level2Out102[4] , 
        \Level2Out102[3] , \Level2Out102[2] , \Level2Out102[1] , 
        \Level2Out102[0] }), .Read1(\Level2Load100[0] ), .Read2(
        \Level2Load102[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_136_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load136[0] ), .Out({\Level2Out136[31] , \Level2Out136[30] , 
        \Level2Out136[29] , \Level2Out136[28] , \Level2Out136[27] , 
        \Level2Out136[26] , \Level2Out136[25] , \Level2Out136[24] , 
        \Level2Out136[23] , \Level2Out136[22] , \Level2Out136[21] , 
        \Level2Out136[20] , \Level2Out136[19] , \Level2Out136[18] , 
        \Level2Out136[17] , \Level2Out136[16] , \Level2Out136[15] , 
        \Level2Out136[14] , \Level2Out136[13] , \Level2Out136[12] , 
        \Level2Out136[11] , \Level2Out136[10] , \Level2Out136[9] , 
        \Level2Out136[8] , \Level2Out136[7] , \Level2Out136[6] , 
        \Level2Out136[5] , \Level2Out136[4] , \Level2Out136[3] , 
        \Level2Out136[2] , \Level2Out136[1] , \Level2Out136[0] }), .In1({
        \Level1Out136[31] , \Level1Out136[30] , \Level1Out136[29] , 
        \Level1Out136[28] , \Level1Out136[27] , \Level1Out136[26] , 
        \Level1Out136[25] , \Level1Out136[24] , \Level1Out136[23] , 
        \Level1Out136[22] , \Level1Out136[21] , \Level1Out136[20] , 
        \Level1Out136[19] , \Level1Out136[18] , \Level1Out136[17] , 
        \Level1Out136[16] , \Level1Out136[15] , \Level1Out136[14] , 
        \Level1Out136[13] , \Level1Out136[12] , \Level1Out136[11] , 
        \Level1Out136[10] , \Level1Out136[9] , \Level1Out136[8] , 
        \Level1Out136[7] , \Level1Out136[6] , \Level1Out136[5] , 
        \Level1Out136[4] , \Level1Out136[3] , \Level1Out136[2] , 
        \Level1Out136[1] , \Level1Out136[0] }), .In2({\Level1Out137[31] , 
        \Level1Out137[30] , \Level1Out137[29] , \Level1Out137[28] , 
        \Level1Out137[27] , \Level1Out137[26] , \Level1Out137[25] , 
        \Level1Out137[24] , \Level1Out137[23] , \Level1Out137[22] , 
        \Level1Out137[21] , \Level1Out137[20] , \Level1Out137[19] , 
        \Level1Out137[18] , \Level1Out137[17] , \Level1Out137[16] , 
        \Level1Out137[15] , \Level1Out137[14] , \Level1Out137[13] , 
        \Level1Out137[12] , \Level1Out137[11] , \Level1Out137[10] , 
        \Level1Out137[9] , \Level1Out137[8] , \Level1Out137[7] , 
        \Level1Out137[6] , \Level1Out137[5] , \Level1Out137[4] , 
        \Level1Out137[3] , \Level1Out137[2] , \Level1Out137[1] , 
        \Level1Out137[0] }), .Read1(\Level1Load136[0] ), .Read2(
        \Level1Load137[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_228_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load228[0] ), .Out({\Level2Out228[31] , \Level2Out228[30] , 
        \Level2Out228[29] , \Level2Out228[28] , \Level2Out228[27] , 
        \Level2Out228[26] , \Level2Out228[25] , \Level2Out228[24] , 
        \Level2Out228[23] , \Level2Out228[22] , \Level2Out228[21] , 
        \Level2Out228[20] , \Level2Out228[19] , \Level2Out228[18] , 
        \Level2Out228[17] , \Level2Out228[16] , \Level2Out228[15] , 
        \Level2Out228[14] , \Level2Out228[13] , \Level2Out228[12] , 
        \Level2Out228[11] , \Level2Out228[10] , \Level2Out228[9] , 
        \Level2Out228[8] , \Level2Out228[7] , \Level2Out228[6] , 
        \Level2Out228[5] , \Level2Out228[4] , \Level2Out228[3] , 
        \Level2Out228[2] , \Level2Out228[1] , \Level2Out228[0] }), .In1({
        \Level1Out228[31] , \Level1Out228[30] , \Level1Out228[29] , 
        \Level1Out228[28] , \Level1Out228[27] , \Level1Out228[26] , 
        \Level1Out228[25] , \Level1Out228[24] , \Level1Out228[23] , 
        \Level1Out228[22] , \Level1Out228[21] , \Level1Out228[20] , 
        \Level1Out228[19] , \Level1Out228[18] , \Level1Out228[17] , 
        \Level1Out228[16] , \Level1Out228[15] , \Level1Out228[14] , 
        \Level1Out228[13] , \Level1Out228[12] , \Level1Out228[11] , 
        \Level1Out228[10] , \Level1Out228[9] , \Level1Out228[8] , 
        \Level1Out228[7] , \Level1Out228[6] , \Level1Out228[5] , 
        \Level1Out228[4] , \Level1Out228[3] , \Level1Out228[2] , 
        \Level1Out228[1] , \Level1Out228[0] }), .In2({\Level1Out229[31] , 
        \Level1Out229[30] , \Level1Out229[29] , \Level1Out229[28] , 
        \Level1Out229[27] , \Level1Out229[26] , \Level1Out229[25] , 
        \Level1Out229[24] , \Level1Out229[23] , \Level1Out229[22] , 
        \Level1Out229[21] , \Level1Out229[20] , \Level1Out229[19] , 
        \Level1Out229[18] , \Level1Out229[17] , \Level1Out229[16] , 
        \Level1Out229[15] , \Level1Out229[14] , \Level1Out229[13] , 
        \Level1Out229[12] , \Level1Out229[11] , \Level1Out229[10] , 
        \Level1Out229[9] , \Level1Out229[8] , \Level1Out229[7] , 
        \Level1Out229[6] , \Level1Out229[5] , \Level1Out229[4] , 
        \Level1Out229[3] , \Level1Out229[2] , \Level1Out229[1] , 
        \Level1Out229[0] }), .Read1(\Level1Load228[0] ), .Read2(
        \Level1Load229[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_192_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load192[0] ), .Out({\Level2Out192[31] , \Level2Out192[30] , 
        \Level2Out192[29] , \Level2Out192[28] , \Level2Out192[27] , 
        \Level2Out192[26] , \Level2Out192[25] , \Level2Out192[24] , 
        \Level2Out192[23] , \Level2Out192[22] , \Level2Out192[21] , 
        \Level2Out192[20] , \Level2Out192[19] , \Level2Out192[18] , 
        \Level2Out192[17] , \Level2Out192[16] , \Level2Out192[15] , 
        \Level2Out192[14] , \Level2Out192[13] , \Level2Out192[12] , 
        \Level2Out192[11] , \Level2Out192[10] , \Level2Out192[9] , 
        \Level2Out192[8] , \Level2Out192[7] , \Level2Out192[6] , 
        \Level2Out192[5] , \Level2Out192[4] , \Level2Out192[3] , 
        \Level2Out192[2] , \Level2Out192[1] , \Level2Out192[0] }), .In1({
        \Level1Out192[31] , \Level1Out192[30] , \Level1Out192[29] , 
        \Level1Out192[28] , \Level1Out192[27] , \Level1Out192[26] , 
        \Level1Out192[25] , \Level1Out192[24] , \Level1Out192[23] , 
        \Level1Out192[22] , \Level1Out192[21] , \Level1Out192[20] , 
        \Level1Out192[19] , \Level1Out192[18] , \Level1Out192[17] , 
        \Level1Out192[16] , \Level1Out192[15] , \Level1Out192[14] , 
        \Level1Out192[13] , \Level1Out192[12] , \Level1Out192[11] , 
        \Level1Out192[10] , \Level1Out192[9] , \Level1Out192[8] , 
        \Level1Out192[7] , \Level1Out192[6] , \Level1Out192[5] , 
        \Level1Out192[4] , \Level1Out192[3] , \Level1Out192[2] , 
        \Level1Out192[1] , \Level1Out192[0] }), .In2({\Level1Out193[31] , 
        \Level1Out193[30] , \Level1Out193[29] , \Level1Out193[28] , 
        \Level1Out193[27] , \Level1Out193[26] , \Level1Out193[25] , 
        \Level1Out193[24] , \Level1Out193[23] , \Level1Out193[22] , 
        \Level1Out193[21] , \Level1Out193[20] , \Level1Out193[19] , 
        \Level1Out193[18] , \Level1Out193[17] , \Level1Out193[16] , 
        \Level1Out193[15] , \Level1Out193[14] , \Level1Out193[13] , 
        \Level1Out193[12] , \Level1Out193[11] , \Level1Out193[10] , 
        \Level1Out193[9] , \Level1Out193[8] , \Level1Out193[7] , 
        \Level1Out193[6] , \Level1Out193[5] , \Level1Out193[4] , 
        \Level1Out193[3] , \Level1Out193[2] , \Level1Out193[1] , 
        \Level1Out193[0] }), .Read1(\Level1Load192[0] ), .Read2(
        \Level1Load193[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_16 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanOut({\ScanLink17[31] , 
        \ScanLink17[30] , \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , 
        \ScanLink17[26] , \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , 
        \ScanLink17[22] , \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , 
        \ScanLink17[18] , \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , 
        \ScanLink17[14] , \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , 
        \ScanLink17[10] , \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , 
        \ScanLink17[6] , \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , 
        \ScanLink17[2] , \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load16[0] ), .Out({
        \Level1Out16[31] , \Level1Out16[30] , \Level1Out16[29] , 
        \Level1Out16[28] , \Level1Out16[27] , \Level1Out16[26] , 
        \Level1Out16[25] , \Level1Out16[24] , \Level1Out16[23] , 
        \Level1Out16[22] , \Level1Out16[21] , \Level1Out16[20] , 
        \Level1Out16[19] , \Level1Out16[18] , \Level1Out16[17] , 
        \Level1Out16[16] , \Level1Out16[15] , \Level1Out16[14] , 
        \Level1Out16[13] , \Level1Out16[12] , \Level1Out16[11] , 
        \Level1Out16[10] , \Level1Out16[9] , \Level1Out16[8] , 
        \Level1Out16[7] , \Level1Out16[6] , \Level1Out16[5] , \Level1Out16[4] , 
        \Level1Out16[3] , \Level1Out16[2] , \Level1Out16[1] , \Level1Out16[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_23 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanOut({\ScanLink24[31] , 
        \ScanLink24[30] , \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , 
        \ScanLink24[26] , \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , 
        \ScanLink24[22] , \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , 
        \ScanLink24[18] , \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , 
        \ScanLink24[14] , \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , 
        \ScanLink24[10] , \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , 
        \ScanLink24[6] , \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , 
        \ScanLink24[2] , \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load23[0] ), .Out({
        \Level1Out23[31] , \Level1Out23[30] , \Level1Out23[29] , 
        \Level1Out23[28] , \Level1Out23[27] , \Level1Out23[26] , 
        \Level1Out23[25] , \Level1Out23[24] , \Level1Out23[23] , 
        \Level1Out23[22] , \Level1Out23[21] , \Level1Out23[20] , 
        \Level1Out23[19] , \Level1Out23[18] , \Level1Out23[17] , 
        \Level1Out23[16] , \Level1Out23[15] , \Level1Out23[14] , 
        \Level1Out23[13] , \Level1Out23[12] , \Level1Out23[11] , 
        \Level1Out23[10] , \Level1Out23[9] , \Level1Out23[8] , 
        \Level1Out23[7] , \Level1Out23[6] , \Level1Out23[5] , \Level1Out23[4] , 
        \Level1Out23[3] , \Level1Out23[2] , \Level1Out23[1] , \Level1Out23[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_148 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink148[31] , \ScanLink148[30] , 
        \ScanLink148[29] , \ScanLink148[28] , \ScanLink148[27] , 
        \ScanLink148[26] , \ScanLink148[25] , \ScanLink148[24] , 
        \ScanLink148[23] , \ScanLink148[22] , \ScanLink148[21] , 
        \ScanLink148[20] , \ScanLink148[19] , \ScanLink148[18] , 
        \ScanLink148[17] , \ScanLink148[16] , \ScanLink148[15] , 
        \ScanLink148[14] , \ScanLink148[13] , \ScanLink148[12] , 
        \ScanLink148[11] , \ScanLink148[10] , \ScanLink148[9] , 
        \ScanLink148[8] , \ScanLink148[7] , \ScanLink148[6] , \ScanLink148[5] , 
        \ScanLink148[4] , \ScanLink148[3] , \ScanLink148[2] , \ScanLink148[1] , 
        \ScanLink148[0] }), .ScanOut({\ScanLink149[31] , \ScanLink149[30] , 
        \ScanLink149[29] , \ScanLink149[28] , \ScanLink149[27] , 
        \ScanLink149[26] , \ScanLink149[25] , \ScanLink149[24] , 
        \ScanLink149[23] , \ScanLink149[22] , \ScanLink149[21] , 
        \ScanLink149[20] , \ScanLink149[19] , \ScanLink149[18] , 
        \ScanLink149[17] , \ScanLink149[16] , \ScanLink149[15] , 
        \ScanLink149[14] , \ScanLink149[13] , \ScanLink149[12] , 
        \ScanLink149[11] , \ScanLink149[10] , \ScanLink149[9] , 
        \ScanLink149[8] , \ScanLink149[7] , \ScanLink149[6] , \ScanLink149[5] , 
        \ScanLink149[4] , \ScanLink149[3] , \ScanLink149[2] , \ScanLink149[1] , 
        \ScanLink149[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load148[0] ), .Out({\Level1Out148[31] , \Level1Out148[30] , 
        \Level1Out148[29] , \Level1Out148[28] , \Level1Out148[27] , 
        \Level1Out148[26] , \Level1Out148[25] , \Level1Out148[24] , 
        \Level1Out148[23] , \Level1Out148[22] , \Level1Out148[21] , 
        \Level1Out148[20] , \Level1Out148[19] , \Level1Out148[18] , 
        \Level1Out148[17] , \Level1Out148[16] , \Level1Out148[15] , 
        \Level1Out148[14] , \Level1Out148[13] , \Level1Out148[12] , 
        \Level1Out148[11] , \Level1Out148[10] , \Level1Out148[9] , 
        \Level1Out148[8] , \Level1Out148[7] , \Level1Out148[6] , 
        \Level1Out148[5] , \Level1Out148[4] , \Level1Out148[3] , 
        \Level1Out148[2] , \Level1Out148[1] , \Level1Out148[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_42_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load42[0] ), .Out({\Level2Out42[31] , \Level2Out42[30] , 
        \Level2Out42[29] , \Level2Out42[28] , \Level2Out42[27] , 
        \Level2Out42[26] , \Level2Out42[25] , \Level2Out42[24] , 
        \Level2Out42[23] , \Level2Out42[22] , \Level2Out42[21] , 
        \Level2Out42[20] , \Level2Out42[19] , \Level2Out42[18] , 
        \Level2Out42[17] , \Level2Out42[16] , \Level2Out42[15] , 
        \Level2Out42[14] , \Level2Out42[13] , \Level2Out42[12] , 
        \Level2Out42[11] , \Level2Out42[10] , \Level2Out42[9] , 
        \Level2Out42[8] , \Level2Out42[7] , \Level2Out42[6] , \Level2Out42[5] , 
        \Level2Out42[4] , \Level2Out42[3] , \Level2Out42[2] , \Level2Out42[1] , 
        \Level2Out42[0] }), .In1({\Level1Out42[31] , \Level1Out42[30] , 
        \Level1Out42[29] , \Level1Out42[28] , \Level1Out42[27] , 
        \Level1Out42[26] , \Level1Out42[25] , \Level1Out42[24] , 
        \Level1Out42[23] , \Level1Out42[22] , \Level1Out42[21] , 
        \Level1Out42[20] , \Level1Out42[19] , \Level1Out42[18] , 
        \Level1Out42[17] , \Level1Out42[16] , \Level1Out42[15] , 
        \Level1Out42[14] , \Level1Out42[13] , \Level1Out42[12] , 
        \Level1Out42[11] , \Level1Out42[10] , \Level1Out42[9] , 
        \Level1Out42[8] , \Level1Out42[7] , \Level1Out42[6] , \Level1Out42[5] , 
        \Level1Out42[4] , \Level1Out42[3] , \Level1Out42[2] , \Level1Out42[1] , 
        \Level1Out42[0] }), .In2({\Level1Out43[31] , \Level1Out43[30] , 
        \Level1Out43[29] , \Level1Out43[28] , \Level1Out43[27] , 
        \Level1Out43[26] , \Level1Out43[25] , \Level1Out43[24] , 
        \Level1Out43[23] , \Level1Out43[22] , \Level1Out43[21] , 
        \Level1Out43[20] , \Level1Out43[19] , \Level1Out43[18] , 
        \Level1Out43[17] , \Level1Out43[16] , \Level1Out43[15] , 
        \Level1Out43[14] , \Level1Out43[13] , \Level1Out43[12] , 
        \Level1Out43[11] , \Level1Out43[10] , \Level1Out43[9] , 
        \Level1Out43[8] , \Level1Out43[7] , \Level1Out43[6] , \Level1Out43[5] , 
        \Level1Out43[4] , \Level1Out43[3] , \Level1Out43[2] , \Level1Out43[1] , 
        \Level1Out43[0] }), .Read1(\Level1Load42[0] ), .Read2(
        \Level1Load43[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_68_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load68[0] ), .Out({\Level2Out68[31] , \Level2Out68[30] , 
        \Level2Out68[29] , \Level2Out68[28] , \Level2Out68[27] , 
        \Level2Out68[26] , \Level2Out68[25] , \Level2Out68[24] , 
        \Level2Out68[23] , \Level2Out68[22] , \Level2Out68[21] , 
        \Level2Out68[20] , \Level2Out68[19] , \Level2Out68[18] , 
        \Level2Out68[17] , \Level2Out68[16] , \Level2Out68[15] , 
        \Level2Out68[14] , \Level2Out68[13] , \Level2Out68[12] , 
        \Level2Out68[11] , \Level2Out68[10] , \Level2Out68[9] , 
        \Level2Out68[8] , \Level2Out68[7] , \Level2Out68[6] , \Level2Out68[5] , 
        \Level2Out68[4] , \Level2Out68[3] , \Level2Out68[2] , \Level2Out68[1] , 
        \Level2Out68[0] }), .In1({\Level1Out68[31] , \Level1Out68[30] , 
        \Level1Out68[29] , \Level1Out68[28] , \Level1Out68[27] , 
        \Level1Out68[26] , \Level1Out68[25] , \Level1Out68[24] , 
        \Level1Out68[23] , \Level1Out68[22] , \Level1Out68[21] , 
        \Level1Out68[20] , \Level1Out68[19] , \Level1Out68[18] , 
        \Level1Out68[17] , \Level1Out68[16] , \Level1Out68[15] , 
        \Level1Out68[14] , \Level1Out68[13] , \Level1Out68[12] , 
        \Level1Out68[11] , \Level1Out68[10] , \Level1Out68[9] , 
        \Level1Out68[8] , \Level1Out68[7] , \Level1Out68[6] , \Level1Out68[5] , 
        \Level1Out68[4] , \Level1Out68[3] , \Level1Out68[2] , \Level1Out68[1] , 
        \Level1Out68[0] }), .In2({\Level1Out69[31] , \Level1Out69[30] , 
        \Level1Out69[29] , \Level1Out69[28] , \Level1Out69[27] , 
        \Level1Out69[26] , \Level1Out69[25] , \Level1Out69[24] , 
        \Level1Out69[23] , \Level1Out69[22] , \Level1Out69[21] , 
        \Level1Out69[20] , \Level1Out69[19] , \Level1Out69[18] , 
        \Level1Out69[17] , \Level1Out69[16] , \Level1Out69[15] , 
        \Level1Out69[14] , \Level1Out69[13] , \Level1Out69[12] , 
        \Level1Out69[11] , \Level1Out69[10] , \Level1Out69[9] , 
        \Level1Out69[8] , \Level1Out69[7] , \Level1Out69[6] , \Level1Out69[5] , 
        \Level1Out69[4] , \Level1Out69[3] , \Level1Out69[2] , \Level1Out69[1] , 
        \Level1Out69[0] }), .Read1(\Level1Load68[0] ), .Read2(
        \Level1Load69[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_104_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load104[0] ), .Out({\Level2Out104[31] , \Level2Out104[30] , 
        \Level2Out104[29] , \Level2Out104[28] , \Level2Out104[27] , 
        \Level2Out104[26] , \Level2Out104[25] , \Level2Out104[24] , 
        \Level2Out104[23] , \Level2Out104[22] , \Level2Out104[21] , 
        \Level2Out104[20] , \Level2Out104[19] , \Level2Out104[18] , 
        \Level2Out104[17] , \Level2Out104[16] , \Level2Out104[15] , 
        \Level2Out104[14] , \Level2Out104[13] , \Level2Out104[12] , 
        \Level2Out104[11] , \Level2Out104[10] , \Level2Out104[9] , 
        \Level2Out104[8] , \Level2Out104[7] , \Level2Out104[6] , 
        \Level2Out104[5] , \Level2Out104[4] , \Level2Out104[3] , 
        \Level2Out104[2] , \Level2Out104[1] , \Level2Out104[0] }), .In1({
        \Level1Out104[31] , \Level1Out104[30] , \Level1Out104[29] , 
        \Level1Out104[28] , \Level1Out104[27] , \Level1Out104[26] , 
        \Level1Out104[25] , \Level1Out104[24] , \Level1Out104[23] , 
        \Level1Out104[22] , \Level1Out104[21] , \Level1Out104[20] , 
        \Level1Out104[19] , \Level1Out104[18] , \Level1Out104[17] , 
        \Level1Out104[16] , \Level1Out104[15] , \Level1Out104[14] , 
        \Level1Out104[13] , \Level1Out104[12] , \Level1Out104[11] , 
        \Level1Out104[10] , \Level1Out104[9] , \Level1Out104[8] , 
        \Level1Out104[7] , \Level1Out104[6] , \Level1Out104[5] , 
        \Level1Out104[4] , \Level1Out104[3] , \Level1Out104[2] , 
        \Level1Out104[1] , \Level1Out104[0] }), .In2({\Level1Out105[31] , 
        \Level1Out105[30] , \Level1Out105[29] , \Level1Out105[28] , 
        \Level1Out105[27] , \Level1Out105[26] , \Level1Out105[25] , 
        \Level1Out105[24] , \Level1Out105[23] , \Level1Out105[22] , 
        \Level1Out105[21] , \Level1Out105[20] , \Level1Out105[19] , 
        \Level1Out105[18] , \Level1Out105[17] , \Level1Out105[16] , 
        \Level1Out105[15] , \Level1Out105[14] , \Level1Out105[13] , 
        \Level1Out105[12] , \Level1Out105[11] , \Level1Out105[10] , 
        \Level1Out105[9] , \Level1Out105[8] , \Level1Out105[7] , 
        \Level1Out105[6] , \Level1Out105[5] , \Level1Out105[4] , 
        \Level1Out105[3] , \Level1Out105[2] , \Level1Out105[1] , 
        \Level1Out105[0] }), .Read1(\Level1Load104[0] ), .Read2(
        \Level1Load105[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_230_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load230[0] ), .Out({\Level2Out230[31] , \Level2Out230[30] , 
        \Level2Out230[29] , \Level2Out230[28] , \Level2Out230[27] , 
        \Level2Out230[26] , \Level2Out230[25] , \Level2Out230[24] , 
        \Level2Out230[23] , \Level2Out230[22] , \Level2Out230[21] , 
        \Level2Out230[20] , \Level2Out230[19] , \Level2Out230[18] , 
        \Level2Out230[17] , \Level2Out230[16] , \Level2Out230[15] , 
        \Level2Out230[14] , \Level2Out230[13] , \Level2Out230[12] , 
        \Level2Out230[11] , \Level2Out230[10] , \Level2Out230[9] , 
        \Level2Out230[8] , \Level2Out230[7] , \Level2Out230[6] , 
        \Level2Out230[5] , \Level2Out230[4] , \Level2Out230[3] , 
        \Level2Out230[2] , \Level2Out230[1] , \Level2Out230[0] }), .In1({
        \Level1Out230[31] , \Level1Out230[30] , \Level1Out230[29] , 
        \Level1Out230[28] , \Level1Out230[27] , \Level1Out230[26] , 
        \Level1Out230[25] , \Level1Out230[24] , \Level1Out230[23] , 
        \Level1Out230[22] , \Level1Out230[21] , \Level1Out230[20] , 
        \Level1Out230[19] , \Level1Out230[18] , \Level1Out230[17] , 
        \Level1Out230[16] , \Level1Out230[15] , \Level1Out230[14] , 
        \Level1Out230[13] , \Level1Out230[12] , \Level1Out230[11] , 
        \Level1Out230[10] , \Level1Out230[9] , \Level1Out230[8] , 
        \Level1Out230[7] , \Level1Out230[6] , \Level1Out230[5] , 
        \Level1Out230[4] , \Level1Out230[3] , \Level1Out230[2] , 
        \Level1Out230[1] , \Level1Out230[0] }), .In2({\Level1Out231[31] , 
        \Level1Out231[30] , \Level1Out231[29] , \Level1Out231[28] , 
        \Level1Out231[27] , \Level1Out231[26] , \Level1Out231[25] , 
        \Level1Out231[24] , \Level1Out231[23] , \Level1Out231[22] , 
        \Level1Out231[21] , \Level1Out231[20] , \Level1Out231[19] , 
        \Level1Out231[18] , \Level1Out231[17] , \Level1Out231[16] , 
        \Level1Out231[15] , \Level1Out231[14] , \Level1Out231[13] , 
        \Level1Out231[12] , \Level1Out231[11] , \Level1Out231[10] , 
        \Level1Out231[9] , \Level1Out231[8] , \Level1Out231[7] , 
        \Level1Out231[6] , \Level1Out231[5] , \Level1Out231[4] , 
        \Level1Out231[3] , \Level1Out231[2] , \Level1Out231[1] , 
        \Level1Out231[0] }), .Read1(\Level1Load230[0] ), .Read2(
        \Level1Load231[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_132_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load132[0] ), .Out({\Level4Out132[31] , \Level4Out132[30] , 
        \Level4Out132[29] , \Level4Out132[28] , \Level4Out132[27] , 
        \Level4Out132[26] , \Level4Out132[25] , \Level4Out132[24] , 
        \Level4Out132[23] , \Level4Out132[22] , \Level4Out132[21] , 
        \Level4Out132[20] , \Level4Out132[19] , \Level4Out132[18] , 
        \Level4Out132[17] , \Level4Out132[16] , \Level4Out132[15] , 
        \Level4Out132[14] , \Level4Out132[13] , \Level4Out132[12] , 
        \Level4Out132[11] , \Level4Out132[10] , \Level4Out132[9] , 
        \Level4Out132[8] , \Level4Out132[7] , \Level4Out132[6] , 
        \Level4Out132[5] , \Level4Out132[4] , \Level4Out132[3] , 
        \Level4Out132[2] , \Level4Out132[1] , \Level4Out132[0] }), .In1({
        \Level2Out132[31] , \Level2Out132[30] , \Level2Out132[29] , 
        \Level2Out132[28] , \Level2Out132[27] , \Level2Out132[26] , 
        \Level2Out132[25] , \Level2Out132[24] , \Level2Out132[23] , 
        \Level2Out132[22] , \Level2Out132[21] , \Level2Out132[20] , 
        \Level2Out132[19] , \Level2Out132[18] , \Level2Out132[17] , 
        \Level2Out132[16] , \Level2Out132[15] , \Level2Out132[14] , 
        \Level2Out132[13] , \Level2Out132[12] , \Level2Out132[11] , 
        \Level2Out132[10] , \Level2Out132[9] , \Level2Out132[8] , 
        \Level2Out132[7] , \Level2Out132[6] , \Level2Out132[5] , 
        \Level2Out132[4] , \Level2Out132[3] , \Level2Out132[2] , 
        \Level2Out132[1] , \Level2Out132[0] }), .In2({\Level2Out134[31] , 
        \Level2Out134[30] , \Level2Out134[29] , \Level2Out134[28] , 
        \Level2Out134[27] , \Level2Out134[26] , \Level2Out134[25] , 
        \Level2Out134[24] , \Level2Out134[23] , \Level2Out134[22] , 
        \Level2Out134[21] , \Level2Out134[20] , \Level2Out134[19] , 
        \Level2Out134[18] , \Level2Out134[17] , \Level2Out134[16] , 
        \Level2Out134[15] , \Level2Out134[14] , \Level2Out134[13] , 
        \Level2Out134[12] , \Level2Out134[11] , \Level2Out134[10] , 
        \Level2Out134[9] , \Level2Out134[8] , \Level2Out134[7] , 
        \Level2Out134[6] , \Level2Out134[5] , \Level2Out134[4] , 
        \Level2Out134[3] , \Level2Out134[2] , \Level2Out134[1] , 
        \Level2Out134[0] }), .Read1(\Level2Load132[0] ), .Read2(
        \Level2Load134[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_128_32 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load128[0] ), .Out({\Level32Out128[31] , \Level32Out128[30] , 
        \Level32Out128[29] , \Level32Out128[28] , \Level32Out128[27] , 
        \Level32Out128[26] , \Level32Out128[25] , \Level32Out128[24] , 
        \Level32Out128[23] , \Level32Out128[22] , \Level32Out128[21] , 
        \Level32Out128[20] , \Level32Out128[19] , \Level32Out128[18] , 
        \Level32Out128[17] , \Level32Out128[16] , \Level32Out128[15] , 
        \Level32Out128[14] , \Level32Out128[13] , \Level32Out128[12] , 
        \Level32Out128[11] , \Level32Out128[10] , \Level32Out128[9] , 
        \Level32Out128[8] , \Level32Out128[7] , \Level32Out128[6] , 
        \Level32Out128[5] , \Level32Out128[4] , \Level32Out128[3] , 
        \Level32Out128[2] , \Level32Out128[1] , \Level32Out128[0] }), .In1({
        \Level16Out128[31] , \Level16Out128[30] , \Level16Out128[29] , 
        \Level16Out128[28] , \Level16Out128[27] , \Level16Out128[26] , 
        \Level16Out128[25] , \Level16Out128[24] , \Level16Out128[23] , 
        \Level16Out128[22] , \Level16Out128[21] , \Level16Out128[20] , 
        \Level16Out128[19] , \Level16Out128[18] , \Level16Out128[17] , 
        \Level16Out128[16] , \Level16Out128[15] , \Level16Out128[14] , 
        \Level16Out128[13] , \Level16Out128[12] , \Level16Out128[11] , 
        \Level16Out128[10] , \Level16Out128[9] , \Level16Out128[8] , 
        \Level16Out128[7] , \Level16Out128[6] , \Level16Out128[5] , 
        \Level16Out128[4] , \Level16Out128[3] , \Level16Out128[2] , 
        \Level16Out128[1] , \Level16Out128[0] }), .In2({\Level16Out144[31] , 
        \Level16Out144[30] , \Level16Out144[29] , \Level16Out144[28] , 
        \Level16Out144[27] , \Level16Out144[26] , \Level16Out144[25] , 
        \Level16Out144[24] , \Level16Out144[23] , \Level16Out144[22] , 
        \Level16Out144[21] , \Level16Out144[20] , \Level16Out144[19] , 
        \Level16Out144[18] , \Level16Out144[17] , \Level16Out144[16] , 
        \Level16Out144[15] , \Level16Out144[14] , \Level16Out144[13] , 
        \Level16Out144[12] , \Level16Out144[11] , \Level16Out144[10] , 
        \Level16Out144[9] , \Level16Out144[8] , \Level16Out144[7] , 
        \Level16Out144[6] , \Level16Out144[5] , \Level16Out144[4] , 
        \Level16Out144[3] , \Level16Out144[2] , \Level16Out144[1] , 
        \Level16Out144[0] }), .Read1(\Level16Load128[0] ), .Read2(
        \Level16Load144[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_31 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanOut({\ScanLink32[31] , 
        \ScanLink32[30] , \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , 
        \ScanLink32[26] , \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , 
        \ScanLink32[22] , \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , 
        \ScanLink32[18] , \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , 
        \ScanLink32[14] , \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , 
        \ScanLink32[10] , \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , 
        \ScanLink32[6] , \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , 
        \ScanLink32[2] , \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load31[0] ), .Out({
        \Level1Out31[31] , \Level1Out31[30] , \Level1Out31[29] , 
        \Level1Out31[28] , \Level1Out31[27] , \Level1Out31[26] , 
        \Level1Out31[25] , \Level1Out31[24] , \Level1Out31[23] , 
        \Level1Out31[22] , \Level1Out31[21] , \Level1Out31[20] , 
        \Level1Out31[19] , \Level1Out31[18] , \Level1Out31[17] , 
        \Level1Out31[16] , \Level1Out31[15] , \Level1Out31[14] , 
        \Level1Out31[13] , \Level1Out31[12] , \Level1Out31[11] , 
        \Level1Out31[10] , \Level1Out31[9] , \Level1Out31[8] , 
        \Level1Out31[7] , \Level1Out31[6] , \Level1Out31[5] , \Level1Out31[4] , 
        \Level1Out31[3] , \Level1Out31[2] , \Level1Out31[1] , \Level1Out31[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_101 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink101[31] , \ScanLink101[30] , 
        \ScanLink101[29] , \ScanLink101[28] , \ScanLink101[27] , 
        \ScanLink101[26] , \ScanLink101[25] , \ScanLink101[24] , 
        \ScanLink101[23] , \ScanLink101[22] , \ScanLink101[21] , 
        \ScanLink101[20] , \ScanLink101[19] , \ScanLink101[18] , 
        \ScanLink101[17] , \ScanLink101[16] , \ScanLink101[15] , 
        \ScanLink101[14] , \ScanLink101[13] , \ScanLink101[12] , 
        \ScanLink101[11] , \ScanLink101[10] , \ScanLink101[9] , 
        \ScanLink101[8] , \ScanLink101[7] , \ScanLink101[6] , \ScanLink101[5] , 
        \ScanLink101[4] , \ScanLink101[3] , \ScanLink101[2] , \ScanLink101[1] , 
        \ScanLink101[0] }), .ScanOut({\ScanLink102[31] , \ScanLink102[30] , 
        \ScanLink102[29] , \ScanLink102[28] , \ScanLink102[27] , 
        \ScanLink102[26] , \ScanLink102[25] , \ScanLink102[24] , 
        \ScanLink102[23] , \ScanLink102[22] , \ScanLink102[21] , 
        \ScanLink102[20] , \ScanLink102[19] , \ScanLink102[18] , 
        \ScanLink102[17] , \ScanLink102[16] , \ScanLink102[15] , 
        \ScanLink102[14] , \ScanLink102[13] , \ScanLink102[12] , 
        \ScanLink102[11] , \ScanLink102[10] , \ScanLink102[9] , 
        \ScanLink102[8] , \ScanLink102[7] , \ScanLink102[6] , \ScanLink102[5] , 
        \ScanLink102[4] , \ScanLink102[3] , \ScanLink102[2] , \ScanLink102[1] , 
        \ScanLink102[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load101[0] ), .Out({\Level1Out101[31] , \Level1Out101[30] , 
        \Level1Out101[29] , \Level1Out101[28] , \Level1Out101[27] , 
        \Level1Out101[26] , \Level1Out101[25] , \Level1Out101[24] , 
        \Level1Out101[23] , \Level1Out101[22] , \Level1Out101[21] , 
        \Level1Out101[20] , \Level1Out101[19] , \Level1Out101[18] , 
        \Level1Out101[17] , \Level1Out101[16] , \Level1Out101[15] , 
        \Level1Out101[14] , \Level1Out101[13] , \Level1Out101[12] , 
        \Level1Out101[11] , \Level1Out101[10] , \Level1Out101[9] , 
        \Level1Out101[8] , \Level1Out101[7] , \Level1Out101[6] , 
        \Level1Out101[5] , \Level1Out101[4] , \Level1Out101[3] , 
        \Level1Out101[2] , \Level1Out101[1] , \Level1Out101[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_126 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink126[31] , \ScanLink126[30] , 
        \ScanLink126[29] , \ScanLink126[28] , \ScanLink126[27] , 
        \ScanLink126[26] , \ScanLink126[25] , \ScanLink126[24] , 
        \ScanLink126[23] , \ScanLink126[22] , \ScanLink126[21] , 
        \ScanLink126[20] , \ScanLink126[19] , \ScanLink126[18] , 
        \ScanLink126[17] , \ScanLink126[16] , \ScanLink126[15] , 
        \ScanLink126[14] , \ScanLink126[13] , \ScanLink126[12] , 
        \ScanLink126[11] , \ScanLink126[10] , \ScanLink126[9] , 
        \ScanLink126[8] , \ScanLink126[7] , \ScanLink126[6] , \ScanLink126[5] , 
        \ScanLink126[4] , \ScanLink126[3] , \ScanLink126[2] , \ScanLink126[1] , 
        \ScanLink126[0] }), .ScanOut({\ScanLink127[31] , \ScanLink127[30] , 
        \ScanLink127[29] , \ScanLink127[28] , \ScanLink127[27] , 
        \ScanLink127[26] , \ScanLink127[25] , \ScanLink127[24] , 
        \ScanLink127[23] , \ScanLink127[22] , \ScanLink127[21] , 
        \ScanLink127[20] , \ScanLink127[19] , \ScanLink127[18] , 
        \ScanLink127[17] , \ScanLink127[16] , \ScanLink127[15] , 
        \ScanLink127[14] , \ScanLink127[13] , \ScanLink127[12] , 
        \ScanLink127[11] , \ScanLink127[10] , \ScanLink127[9] , 
        \ScanLink127[8] , \ScanLink127[7] , \ScanLink127[6] , \ScanLink127[5] , 
        \ScanLink127[4] , \ScanLink127[3] , \ScanLink127[2] , \ScanLink127[1] , 
        \ScanLink127[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load126[0] ), .Out({\Level1Out126[31] , \Level1Out126[30] , 
        \Level1Out126[29] , \Level1Out126[28] , \Level1Out126[27] , 
        \Level1Out126[26] , \Level1Out126[25] , \Level1Out126[24] , 
        \Level1Out126[23] , \Level1Out126[22] , \Level1Out126[21] , 
        \Level1Out126[20] , \Level1Out126[19] , \Level1Out126[18] , 
        \Level1Out126[17] , \Level1Out126[16] , \Level1Out126[15] , 
        \Level1Out126[14] , \Level1Out126[13] , \Level1Out126[12] , 
        \Level1Out126[11] , \Level1Out126[10] , \Level1Out126[9] , 
        \Level1Out126[8] , \Level1Out126[7] , \Level1Out126[6] , 
        \Level1Out126[5] , \Level1Out126[4] , \Level1Out126[3] , 
        \Level1Out126[2] , \Level1Out126[1] , \Level1Out126[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_216 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink216[31] , \ScanLink216[30] , 
        \ScanLink216[29] , \ScanLink216[28] , \ScanLink216[27] , 
        \ScanLink216[26] , \ScanLink216[25] , \ScanLink216[24] , 
        \ScanLink216[23] , \ScanLink216[22] , \ScanLink216[21] , 
        \ScanLink216[20] , \ScanLink216[19] , \ScanLink216[18] , 
        \ScanLink216[17] , \ScanLink216[16] , \ScanLink216[15] , 
        \ScanLink216[14] , \ScanLink216[13] , \ScanLink216[12] , 
        \ScanLink216[11] , \ScanLink216[10] , \ScanLink216[9] , 
        \ScanLink216[8] , \ScanLink216[7] , \ScanLink216[6] , \ScanLink216[5] , 
        \ScanLink216[4] , \ScanLink216[3] , \ScanLink216[2] , \ScanLink216[1] , 
        \ScanLink216[0] }), .ScanOut({\ScanLink217[31] , \ScanLink217[30] , 
        \ScanLink217[29] , \ScanLink217[28] , \ScanLink217[27] , 
        \ScanLink217[26] , \ScanLink217[25] , \ScanLink217[24] , 
        \ScanLink217[23] , \ScanLink217[22] , \ScanLink217[21] , 
        \ScanLink217[20] , \ScanLink217[19] , \ScanLink217[18] , 
        \ScanLink217[17] , \ScanLink217[16] , \ScanLink217[15] , 
        \ScanLink217[14] , \ScanLink217[13] , \ScanLink217[12] , 
        \ScanLink217[11] , \ScanLink217[10] , \ScanLink217[9] , 
        \ScanLink217[8] , \ScanLink217[7] , \ScanLink217[6] , \ScanLink217[5] , 
        \ScanLink217[4] , \ScanLink217[3] , \ScanLink217[2] , \ScanLink217[1] , 
        \ScanLink217[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load216[0] ), .Out({\Level1Out216[31] , \Level1Out216[30] , 
        \Level1Out216[29] , \Level1Out216[28] , \Level1Out216[27] , 
        \Level1Out216[26] , \Level1Out216[25] , \Level1Out216[24] , 
        \Level1Out216[23] , \Level1Out216[22] , \Level1Out216[21] , 
        \Level1Out216[20] , \Level1Out216[19] , \Level1Out216[18] , 
        \Level1Out216[17] , \Level1Out216[16] , \Level1Out216[15] , 
        \Level1Out216[14] , \Level1Out216[13] , \Level1Out216[12] , 
        \Level1Out216[11] , \Level1Out216[10] , \Level1Out216[9] , 
        \Level1Out216[8] , \Level1Out216[7] , \Level1Out216[6] , 
        \Level1Out216[5] , \Level1Out216[4] , \Level1Out216[3] , 
        \Level1Out216[2] , \Level1Out216[1] , \Level1Out216[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_96_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load96[0] ), .Out({\Level16Out96[31] , \Level16Out96[30] , 
        \Level16Out96[29] , \Level16Out96[28] , \Level16Out96[27] , 
        \Level16Out96[26] , \Level16Out96[25] , \Level16Out96[24] , 
        \Level16Out96[23] , \Level16Out96[22] , \Level16Out96[21] , 
        \Level16Out96[20] , \Level16Out96[19] , \Level16Out96[18] , 
        \Level16Out96[17] , \Level16Out96[16] , \Level16Out96[15] , 
        \Level16Out96[14] , \Level16Out96[13] , \Level16Out96[12] , 
        \Level16Out96[11] , \Level16Out96[10] , \Level16Out96[9] , 
        \Level16Out96[8] , \Level16Out96[7] , \Level16Out96[6] , 
        \Level16Out96[5] , \Level16Out96[4] , \Level16Out96[3] , 
        \Level16Out96[2] , \Level16Out96[1] , \Level16Out96[0] }), .In1({
        \Level8Out96[31] , \Level8Out96[30] , \Level8Out96[29] , 
        \Level8Out96[28] , \Level8Out96[27] , \Level8Out96[26] , 
        \Level8Out96[25] , \Level8Out96[24] , \Level8Out96[23] , 
        \Level8Out96[22] , \Level8Out96[21] , \Level8Out96[20] , 
        \Level8Out96[19] , \Level8Out96[18] , \Level8Out96[17] , 
        \Level8Out96[16] , \Level8Out96[15] , \Level8Out96[14] , 
        \Level8Out96[13] , \Level8Out96[12] , \Level8Out96[11] , 
        \Level8Out96[10] , \Level8Out96[9] , \Level8Out96[8] , 
        \Level8Out96[7] , \Level8Out96[6] , \Level8Out96[5] , \Level8Out96[4] , 
        \Level8Out96[3] , \Level8Out96[2] , \Level8Out96[1] , \Level8Out96[0] 
        }), .In2({\Level8Out104[31] , \Level8Out104[30] , \Level8Out104[29] , 
        \Level8Out104[28] , \Level8Out104[27] , \Level8Out104[26] , 
        \Level8Out104[25] , \Level8Out104[24] , \Level8Out104[23] , 
        \Level8Out104[22] , \Level8Out104[21] , \Level8Out104[20] , 
        \Level8Out104[19] , \Level8Out104[18] , \Level8Out104[17] , 
        \Level8Out104[16] , \Level8Out104[15] , \Level8Out104[14] , 
        \Level8Out104[13] , \Level8Out104[12] , \Level8Out104[11] , 
        \Level8Out104[10] , \Level8Out104[9] , \Level8Out104[8] , 
        \Level8Out104[7] , \Level8Out104[6] , \Level8Out104[5] , 
        \Level8Out104[4] , \Level8Out104[3] , \Level8Out104[2] , 
        \Level8Out104[1] , \Level8Out104[0] }), .Read1(\Level8Load96[0] ), 
        .Read2(\Level8Load104[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_113 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink113[31] , \ScanLink113[30] , 
        \ScanLink113[29] , \ScanLink113[28] , \ScanLink113[27] , 
        \ScanLink113[26] , \ScanLink113[25] , \ScanLink113[24] , 
        \ScanLink113[23] , \ScanLink113[22] , \ScanLink113[21] , 
        \ScanLink113[20] , \ScanLink113[19] , \ScanLink113[18] , 
        \ScanLink113[17] , \ScanLink113[16] , \ScanLink113[15] , 
        \ScanLink113[14] , \ScanLink113[13] , \ScanLink113[12] , 
        \ScanLink113[11] , \ScanLink113[10] , \ScanLink113[9] , 
        \ScanLink113[8] , \ScanLink113[7] , \ScanLink113[6] , \ScanLink113[5] , 
        \ScanLink113[4] , \ScanLink113[3] , \ScanLink113[2] , \ScanLink113[1] , 
        \ScanLink113[0] }), .ScanOut({\ScanLink114[31] , \ScanLink114[30] , 
        \ScanLink114[29] , \ScanLink114[28] , \ScanLink114[27] , 
        \ScanLink114[26] , \ScanLink114[25] , \ScanLink114[24] , 
        \ScanLink114[23] , \ScanLink114[22] , \ScanLink114[21] , 
        \ScanLink114[20] , \ScanLink114[19] , \ScanLink114[18] , 
        \ScanLink114[17] , \ScanLink114[16] , \ScanLink114[15] , 
        \ScanLink114[14] , \ScanLink114[13] , \ScanLink114[12] , 
        \ScanLink114[11] , \ScanLink114[10] , \ScanLink114[9] , 
        \ScanLink114[8] , \ScanLink114[7] , \ScanLink114[6] , \ScanLink114[5] , 
        \ScanLink114[4] , \ScanLink114[3] , \ScanLink114[2] , \ScanLink114[1] , 
        \ScanLink114[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load113[0] ), .Out({\Level1Out113[31] , \Level1Out113[30] , 
        \Level1Out113[29] , \Level1Out113[28] , \Level1Out113[27] , 
        \Level1Out113[26] , \Level1Out113[25] , \Level1Out113[24] , 
        \Level1Out113[23] , \Level1Out113[22] , \Level1Out113[21] , 
        \Level1Out113[20] , \Level1Out113[19] , \Level1Out113[18] , 
        \Level1Out113[17] , \Level1Out113[16] , \Level1Out113[15] , 
        \Level1Out113[14] , \Level1Out113[13] , \Level1Out113[12] , 
        \Level1Out113[11] , \Level1Out113[10] , \Level1Out113[9] , 
        \Level1Out113[8] , \Level1Out113[7] , \Level1Out113[6] , 
        \Level1Out113[5] , \Level1Out113[4] , \Level1Out113[3] , 
        \Level1Out113[2] , \Level1Out113[1] , \Level1Out113[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_134 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink134[31] , \ScanLink134[30] , 
        \ScanLink134[29] , \ScanLink134[28] , \ScanLink134[27] , 
        \ScanLink134[26] , \ScanLink134[25] , \ScanLink134[24] , 
        \ScanLink134[23] , \ScanLink134[22] , \ScanLink134[21] , 
        \ScanLink134[20] , \ScanLink134[19] , \ScanLink134[18] , 
        \ScanLink134[17] , \ScanLink134[16] , \ScanLink134[15] , 
        \ScanLink134[14] , \ScanLink134[13] , \ScanLink134[12] , 
        \ScanLink134[11] , \ScanLink134[10] , \ScanLink134[9] , 
        \ScanLink134[8] , \ScanLink134[7] , \ScanLink134[6] , \ScanLink134[5] , 
        \ScanLink134[4] , \ScanLink134[3] , \ScanLink134[2] , \ScanLink134[1] , 
        \ScanLink134[0] }), .ScanOut({\ScanLink135[31] , \ScanLink135[30] , 
        \ScanLink135[29] , \ScanLink135[28] , \ScanLink135[27] , 
        \ScanLink135[26] , \ScanLink135[25] , \ScanLink135[24] , 
        \ScanLink135[23] , \ScanLink135[22] , \ScanLink135[21] , 
        \ScanLink135[20] , \ScanLink135[19] , \ScanLink135[18] , 
        \ScanLink135[17] , \ScanLink135[16] , \ScanLink135[15] , 
        \ScanLink135[14] , \ScanLink135[13] , \ScanLink135[12] , 
        \ScanLink135[11] , \ScanLink135[10] , \ScanLink135[9] , 
        \ScanLink135[8] , \ScanLink135[7] , \ScanLink135[6] , \ScanLink135[5] , 
        \ScanLink135[4] , \ScanLink135[3] , \ScanLink135[2] , \ScanLink135[1] , 
        \ScanLink135[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load134[0] ), .Out({\Level1Out134[31] , \Level1Out134[30] , 
        \Level1Out134[29] , \Level1Out134[28] , \Level1Out134[27] , 
        \Level1Out134[26] , \Level1Out134[25] , \Level1Out134[24] , 
        \Level1Out134[23] , \Level1Out134[22] , \Level1Out134[21] , 
        \Level1Out134[20] , \Level1Out134[19] , \Level1Out134[18] , 
        \Level1Out134[17] , \Level1Out134[16] , \Level1Out134[15] , 
        \Level1Out134[14] , \Level1Out134[13] , \Level1Out134[12] , 
        \Level1Out134[11] , \Level1Out134[10] , \Level1Out134[9] , 
        \Level1Out134[8] , \Level1Out134[7] , \Level1Out134[6] , 
        \Level1Out134[5] , \Level1Out134[4] , \Level1Out134[3] , 
        \Level1Out134[2] , \Level1Out134[1] , \Level1Out134[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_204 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink204[31] , \ScanLink204[30] , 
        \ScanLink204[29] , \ScanLink204[28] , \ScanLink204[27] , 
        \ScanLink204[26] , \ScanLink204[25] , \ScanLink204[24] , 
        \ScanLink204[23] , \ScanLink204[22] , \ScanLink204[21] , 
        \ScanLink204[20] , \ScanLink204[19] , \ScanLink204[18] , 
        \ScanLink204[17] , \ScanLink204[16] , \ScanLink204[15] , 
        \ScanLink204[14] , \ScanLink204[13] , \ScanLink204[12] , 
        \ScanLink204[11] , \ScanLink204[10] , \ScanLink204[9] , 
        \ScanLink204[8] , \ScanLink204[7] , \ScanLink204[6] , \ScanLink204[5] , 
        \ScanLink204[4] , \ScanLink204[3] , \ScanLink204[2] , \ScanLink204[1] , 
        \ScanLink204[0] }), .ScanOut({\ScanLink205[31] , \ScanLink205[30] , 
        \ScanLink205[29] , \ScanLink205[28] , \ScanLink205[27] , 
        \ScanLink205[26] , \ScanLink205[25] , \ScanLink205[24] , 
        \ScanLink205[23] , \ScanLink205[22] , \ScanLink205[21] , 
        \ScanLink205[20] , \ScanLink205[19] , \ScanLink205[18] , 
        \ScanLink205[17] , \ScanLink205[16] , \ScanLink205[15] , 
        \ScanLink205[14] , \ScanLink205[13] , \ScanLink205[12] , 
        \ScanLink205[11] , \ScanLink205[10] , \ScanLink205[9] , 
        \ScanLink205[8] , \ScanLink205[7] , \ScanLink205[6] , \ScanLink205[5] , 
        \ScanLink205[4] , \ScanLink205[3] , \ScanLink205[2] , \ScanLink205[1] , 
        \ScanLink205[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load204[0] ), .Out({\Level1Out204[31] , \Level1Out204[30] , 
        \Level1Out204[29] , \Level1Out204[28] , \Level1Out204[27] , 
        \Level1Out204[26] , \Level1Out204[25] , \Level1Out204[24] , 
        \Level1Out204[23] , \Level1Out204[22] , \Level1Out204[21] , 
        \Level1Out204[20] , \Level1Out204[19] , \Level1Out204[18] , 
        \Level1Out204[17] , \Level1Out204[16] , \Level1Out204[15] , 
        \Level1Out204[14] , \Level1Out204[13] , \Level1Out204[12] , 
        \Level1Out204[11] , \Level1Out204[10] , \Level1Out204[9] , 
        \Level1Out204[8] , \Level1Out204[7] , \Level1Out204[6] , 
        \Level1Out204[5] , \Level1Out204[4] , \Level1Out204[3] , 
        \Level1Out204[2] , \Level1Out204[1] , \Level1Out204[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_231 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink231[31] , \ScanLink231[30] , 
        \ScanLink231[29] , \ScanLink231[28] , \ScanLink231[27] , 
        \ScanLink231[26] , \ScanLink231[25] , \ScanLink231[24] , 
        \ScanLink231[23] , \ScanLink231[22] , \ScanLink231[21] , 
        \ScanLink231[20] , \ScanLink231[19] , \ScanLink231[18] , 
        \ScanLink231[17] , \ScanLink231[16] , \ScanLink231[15] , 
        \ScanLink231[14] , \ScanLink231[13] , \ScanLink231[12] , 
        \ScanLink231[11] , \ScanLink231[10] , \ScanLink231[9] , 
        \ScanLink231[8] , \ScanLink231[7] , \ScanLink231[6] , \ScanLink231[5] , 
        \ScanLink231[4] , \ScanLink231[3] , \ScanLink231[2] , \ScanLink231[1] , 
        \ScanLink231[0] }), .ScanOut({\ScanLink232[31] , \ScanLink232[30] , 
        \ScanLink232[29] , \ScanLink232[28] , \ScanLink232[27] , 
        \ScanLink232[26] , \ScanLink232[25] , \ScanLink232[24] , 
        \ScanLink232[23] , \ScanLink232[22] , \ScanLink232[21] , 
        \ScanLink232[20] , \ScanLink232[19] , \ScanLink232[18] , 
        \ScanLink232[17] , \ScanLink232[16] , \ScanLink232[15] , 
        \ScanLink232[14] , \ScanLink232[13] , \ScanLink232[12] , 
        \ScanLink232[11] , \ScanLink232[10] , \ScanLink232[9] , 
        \ScanLink232[8] , \ScanLink232[7] , \ScanLink232[6] , \ScanLink232[5] , 
        \ScanLink232[4] , \ScanLink232[3] , \ScanLink232[2] , \ScanLink232[1] , 
        \ScanLink232[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load231[0] ), .Out({\Level1Out231[31] , \Level1Out231[30] , 
        \Level1Out231[29] , \Level1Out231[28] , \Level1Out231[27] , 
        \Level1Out231[26] , \Level1Out231[25] , \Level1Out231[24] , 
        \Level1Out231[23] , \Level1Out231[22] , \Level1Out231[21] , 
        \Level1Out231[20] , \Level1Out231[19] , \Level1Out231[18] , 
        \Level1Out231[17] , \Level1Out231[16] , \Level1Out231[15] , 
        \Level1Out231[14] , \Level1Out231[13] , \Level1Out231[12] , 
        \Level1Out231[11] , \Level1Out231[10] , \Level1Out231[9] , 
        \Level1Out231[8] , \Level1Out231[7] , \Level1Out231[6] , 
        \Level1Out231[5] , \Level1Out231[4] , \Level1Out231[3] , 
        \Level1Out231[2] , \Level1Out231[1] , \Level1Out231[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_12_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load12[0] ), .Out({\Level2Out12[31] , \Level2Out12[30] , 
        \Level2Out12[29] , \Level2Out12[28] , \Level2Out12[27] , 
        \Level2Out12[26] , \Level2Out12[25] , \Level2Out12[24] , 
        \Level2Out12[23] , \Level2Out12[22] , \Level2Out12[21] , 
        \Level2Out12[20] , \Level2Out12[19] , \Level2Out12[18] , 
        \Level2Out12[17] , \Level2Out12[16] , \Level2Out12[15] , 
        \Level2Out12[14] , \Level2Out12[13] , \Level2Out12[12] , 
        \Level2Out12[11] , \Level2Out12[10] , \Level2Out12[9] , 
        \Level2Out12[8] , \Level2Out12[7] , \Level2Out12[6] , \Level2Out12[5] , 
        \Level2Out12[4] , \Level2Out12[3] , \Level2Out12[2] , \Level2Out12[1] , 
        \Level2Out12[0] }), .In1({\Level1Out12[31] , \Level1Out12[30] , 
        \Level1Out12[29] , \Level1Out12[28] , \Level1Out12[27] , 
        \Level1Out12[26] , \Level1Out12[25] , \Level1Out12[24] , 
        \Level1Out12[23] , \Level1Out12[22] , \Level1Out12[21] , 
        \Level1Out12[20] , \Level1Out12[19] , \Level1Out12[18] , 
        \Level1Out12[17] , \Level1Out12[16] , \Level1Out12[15] , 
        \Level1Out12[14] , \Level1Out12[13] , \Level1Out12[12] , 
        \Level1Out12[11] , \Level1Out12[10] , \Level1Out12[9] , 
        \Level1Out12[8] , \Level1Out12[7] , \Level1Out12[6] , \Level1Out12[5] , 
        \Level1Out12[4] , \Level1Out12[3] , \Level1Out12[2] , \Level1Out12[1] , 
        \Level1Out12[0] }), .In2({\Level1Out13[31] , \Level1Out13[30] , 
        \Level1Out13[29] , \Level1Out13[28] , \Level1Out13[27] , 
        \Level1Out13[26] , \Level1Out13[25] , \Level1Out13[24] , 
        \Level1Out13[23] , \Level1Out13[22] , \Level1Out13[21] , 
        \Level1Out13[20] , \Level1Out13[19] , \Level1Out13[18] , 
        \Level1Out13[17] , \Level1Out13[16] , \Level1Out13[15] , 
        \Level1Out13[14] , \Level1Out13[13] , \Level1Out13[12] , 
        \Level1Out13[11] , \Level1Out13[10] , \Level1Out13[9] , 
        \Level1Out13[8] , \Level1Out13[7] , \Level1Out13[6] , \Level1Out13[5] , 
        \Level1Out13[4] , \Level1Out13[3] , \Level1Out13[2] , \Level1Out13[1] , 
        \Level1Out13[0] }), .Read1(\Level1Load12[0] ), .Read2(
        \Level1Load13[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_154_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load154[0] ), .Out({\Level2Out154[31] , \Level2Out154[30] , 
        \Level2Out154[29] , \Level2Out154[28] , \Level2Out154[27] , 
        \Level2Out154[26] , \Level2Out154[25] , \Level2Out154[24] , 
        \Level2Out154[23] , \Level2Out154[22] , \Level2Out154[21] , 
        \Level2Out154[20] , \Level2Out154[19] , \Level2Out154[18] , 
        \Level2Out154[17] , \Level2Out154[16] , \Level2Out154[15] , 
        \Level2Out154[14] , \Level2Out154[13] , \Level2Out154[12] , 
        \Level2Out154[11] , \Level2Out154[10] , \Level2Out154[9] , 
        \Level2Out154[8] , \Level2Out154[7] , \Level2Out154[6] , 
        \Level2Out154[5] , \Level2Out154[4] , \Level2Out154[3] , 
        \Level2Out154[2] , \Level2Out154[1] , \Level2Out154[0] }), .In1({
        \Level1Out154[31] , \Level1Out154[30] , \Level1Out154[29] , 
        \Level1Out154[28] , \Level1Out154[27] , \Level1Out154[26] , 
        \Level1Out154[25] , \Level1Out154[24] , \Level1Out154[23] , 
        \Level1Out154[22] , \Level1Out154[21] , \Level1Out154[20] , 
        \Level1Out154[19] , \Level1Out154[18] , \Level1Out154[17] , 
        \Level1Out154[16] , \Level1Out154[15] , \Level1Out154[14] , 
        \Level1Out154[13] , \Level1Out154[12] , \Level1Out154[11] , 
        \Level1Out154[10] , \Level1Out154[9] , \Level1Out154[8] , 
        \Level1Out154[7] , \Level1Out154[6] , \Level1Out154[5] , 
        \Level1Out154[4] , \Level1Out154[3] , \Level1Out154[2] , 
        \Level1Out154[1] , \Level1Out154[0] }), .In2({\Level1Out155[31] , 
        \Level1Out155[30] , \Level1Out155[29] , \Level1Out155[28] , 
        \Level1Out155[27] , \Level1Out155[26] , \Level1Out155[25] , 
        \Level1Out155[24] , \Level1Out155[23] , \Level1Out155[22] , 
        \Level1Out155[21] , \Level1Out155[20] , \Level1Out155[19] , 
        \Level1Out155[18] , \Level1Out155[17] , \Level1Out155[16] , 
        \Level1Out155[15] , \Level1Out155[14] , \Level1Out155[13] , 
        \Level1Out155[12] , \Level1Out155[11] , \Level1Out155[10] , 
        \Level1Out155[9] , \Level1Out155[8] , \Level1Out155[7] , 
        \Level1Out155[6] , \Level1Out155[5] , \Level1Out155[4] , 
        \Level1Out155[3] , \Level1Out155[2] , \Level1Out155[1] , 
        \Level1Out155[0] }), .Read1(\Level1Load154[0] ), .Read2(
        \Level1Load155[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_148_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load148[0] ), .Out({\Level4Out148[31] , \Level4Out148[30] , 
        \Level4Out148[29] , \Level4Out148[28] , \Level4Out148[27] , 
        \Level4Out148[26] , \Level4Out148[25] , \Level4Out148[24] , 
        \Level4Out148[23] , \Level4Out148[22] , \Level4Out148[21] , 
        \Level4Out148[20] , \Level4Out148[19] , \Level4Out148[18] , 
        \Level4Out148[17] , \Level4Out148[16] , \Level4Out148[15] , 
        \Level4Out148[14] , \Level4Out148[13] , \Level4Out148[12] , 
        \Level4Out148[11] , \Level4Out148[10] , \Level4Out148[9] , 
        \Level4Out148[8] , \Level4Out148[7] , \Level4Out148[6] , 
        \Level4Out148[5] , \Level4Out148[4] , \Level4Out148[3] , 
        \Level4Out148[2] , \Level4Out148[1] , \Level4Out148[0] }), .In1({
        \Level2Out148[31] , \Level2Out148[30] , \Level2Out148[29] , 
        \Level2Out148[28] , \Level2Out148[27] , \Level2Out148[26] , 
        \Level2Out148[25] , \Level2Out148[24] , \Level2Out148[23] , 
        \Level2Out148[22] , \Level2Out148[21] , \Level2Out148[20] , 
        \Level2Out148[19] , \Level2Out148[18] , \Level2Out148[17] , 
        \Level2Out148[16] , \Level2Out148[15] , \Level2Out148[14] , 
        \Level2Out148[13] , \Level2Out148[12] , \Level2Out148[11] , 
        \Level2Out148[10] , \Level2Out148[9] , \Level2Out148[8] , 
        \Level2Out148[7] , \Level2Out148[6] , \Level2Out148[5] , 
        \Level2Out148[4] , \Level2Out148[3] , \Level2Out148[2] , 
        \Level2Out148[1] , \Level2Out148[0] }), .In2({\Level2Out150[31] , 
        \Level2Out150[30] , \Level2Out150[29] , \Level2Out150[28] , 
        \Level2Out150[27] , \Level2Out150[26] , \Level2Out150[25] , 
        \Level2Out150[24] , \Level2Out150[23] , \Level2Out150[22] , 
        \Level2Out150[21] , \Level2Out150[20] , \Level2Out150[19] , 
        \Level2Out150[18] , \Level2Out150[17] , \Level2Out150[16] , 
        \Level2Out150[15] , \Level2Out150[14] , \Level2Out150[13] , 
        \Level2Out150[12] , \Level2Out150[11] , \Level2Out150[10] , 
        \Level2Out150[9] , \Level2Out150[8] , \Level2Out150[7] , 
        \Level2Out150[6] , \Level2Out150[5] , \Level2Out150[4] , 
        \Level2Out150[3] , \Level2Out150[2] , \Level2Out150[1] , 
        \Level2Out150[0] }), .Read1(\Level2Load148[0] ), .Read2(
        \Level2Load150[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_223 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink223[31] , \ScanLink223[30] , 
        \ScanLink223[29] , \ScanLink223[28] , \ScanLink223[27] , 
        \ScanLink223[26] , \ScanLink223[25] , \ScanLink223[24] , 
        \ScanLink223[23] , \ScanLink223[22] , \ScanLink223[21] , 
        \ScanLink223[20] , \ScanLink223[19] , \ScanLink223[18] , 
        \ScanLink223[17] , \ScanLink223[16] , \ScanLink223[15] , 
        \ScanLink223[14] , \ScanLink223[13] , \ScanLink223[12] , 
        \ScanLink223[11] , \ScanLink223[10] , \ScanLink223[9] , 
        \ScanLink223[8] , \ScanLink223[7] , \ScanLink223[6] , \ScanLink223[5] , 
        \ScanLink223[4] , \ScanLink223[3] , \ScanLink223[2] , \ScanLink223[1] , 
        \ScanLink223[0] }), .ScanOut({\ScanLink224[31] , \ScanLink224[30] , 
        \ScanLink224[29] , \ScanLink224[28] , \ScanLink224[27] , 
        \ScanLink224[26] , \ScanLink224[25] , \ScanLink224[24] , 
        \ScanLink224[23] , \ScanLink224[22] , \ScanLink224[21] , 
        \ScanLink224[20] , \ScanLink224[19] , \ScanLink224[18] , 
        \ScanLink224[17] , \ScanLink224[16] , \ScanLink224[15] , 
        \ScanLink224[14] , \ScanLink224[13] , \ScanLink224[12] , 
        \ScanLink224[11] , \ScanLink224[10] , \ScanLink224[9] , 
        \ScanLink224[8] , \ScanLink224[7] , \ScanLink224[6] , \ScanLink224[5] , 
        \ScanLink224[4] , \ScanLink224[3] , \ScanLink224[2] , \ScanLink224[1] , 
        \ScanLink224[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load223[0] ), .Out({\Level1Out223[31] , \Level1Out223[30] , 
        \Level1Out223[29] , \Level1Out223[28] , \Level1Out223[27] , 
        \Level1Out223[26] , \Level1Out223[25] , \Level1Out223[24] , 
        \Level1Out223[23] , \Level1Out223[22] , \Level1Out223[21] , 
        \Level1Out223[20] , \Level1Out223[19] , \Level1Out223[18] , 
        \Level1Out223[17] , \Level1Out223[16] , \Level1Out223[15] , 
        \Level1Out223[14] , \Level1Out223[13] , \Level1Out223[12] , 
        \Level1Out223[11] , \Level1Out223[10] , \Level1Out223[9] , 
        \Level1Out223[8] , \Level1Out223[7] , \Level1Out223[6] , 
        \Level1Out223[5] , \Level1Out223[4] , \Level1Out223[3] , 
        \Level1Out223[2] , \Level1Out223[1] , \Level1Out223[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_38_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load38[0] ), .Out({\Level2Out38[31] , \Level2Out38[30] , 
        \Level2Out38[29] , \Level2Out38[28] , \Level2Out38[27] , 
        \Level2Out38[26] , \Level2Out38[25] , \Level2Out38[24] , 
        \Level2Out38[23] , \Level2Out38[22] , \Level2Out38[21] , 
        \Level2Out38[20] , \Level2Out38[19] , \Level2Out38[18] , 
        \Level2Out38[17] , \Level2Out38[16] , \Level2Out38[15] , 
        \Level2Out38[14] , \Level2Out38[13] , \Level2Out38[12] , 
        \Level2Out38[11] , \Level2Out38[10] , \Level2Out38[9] , 
        \Level2Out38[8] , \Level2Out38[7] , \Level2Out38[6] , \Level2Out38[5] , 
        \Level2Out38[4] , \Level2Out38[3] , \Level2Out38[2] , \Level2Out38[1] , 
        \Level2Out38[0] }), .In1({\Level1Out38[31] , \Level1Out38[30] , 
        \Level1Out38[29] , \Level1Out38[28] , \Level1Out38[27] , 
        \Level1Out38[26] , \Level1Out38[25] , \Level1Out38[24] , 
        \Level1Out38[23] , \Level1Out38[22] , \Level1Out38[21] , 
        \Level1Out38[20] , \Level1Out38[19] , \Level1Out38[18] , 
        \Level1Out38[17] , \Level1Out38[16] , \Level1Out38[15] , 
        \Level1Out38[14] , \Level1Out38[13] , \Level1Out38[12] , 
        \Level1Out38[11] , \Level1Out38[10] , \Level1Out38[9] , 
        \Level1Out38[8] , \Level1Out38[7] , \Level1Out38[6] , \Level1Out38[5] , 
        \Level1Out38[4] , \Level1Out38[3] , \Level1Out38[2] , \Level1Out38[1] , 
        \Level1Out38[0] }), .In2({\Level1Out39[31] , \Level1Out39[30] , 
        \Level1Out39[29] , \Level1Out39[28] , \Level1Out39[27] , 
        \Level1Out39[26] , \Level1Out39[25] , \Level1Out39[24] , 
        \Level1Out39[23] , \Level1Out39[22] , \Level1Out39[21] , 
        \Level1Out39[20] , \Level1Out39[19] , \Level1Out39[18] , 
        \Level1Out39[17] , \Level1Out39[16] , \Level1Out39[15] , 
        \Level1Out39[14] , \Level1Out39[13] , \Level1Out39[12] , 
        \Level1Out39[11] , \Level1Out39[10] , \Level1Out39[9] , 
        \Level1Out39[8] , \Level1Out39[7] , \Level1Out39[6] , \Level1Out39[5] , 
        \Level1Out39[4] , \Level1Out39[3] , \Level1Out39[2] , \Level1Out39[1] , 
        \Level1Out39[0] }), .Read1(\Level1Load38[0] ), .Read2(
        \Level1Load39[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load24[0] ), .Out({\Level4Out24[31] , \Level4Out24[30] , 
        \Level4Out24[29] , \Level4Out24[28] , \Level4Out24[27] , 
        \Level4Out24[26] , \Level4Out24[25] , \Level4Out24[24] , 
        \Level4Out24[23] , \Level4Out24[22] , \Level4Out24[21] , 
        \Level4Out24[20] , \Level4Out24[19] , \Level4Out24[18] , 
        \Level4Out24[17] , \Level4Out24[16] , \Level4Out24[15] , 
        \Level4Out24[14] , \Level4Out24[13] , \Level4Out24[12] , 
        \Level4Out24[11] , \Level4Out24[10] , \Level4Out24[9] , 
        \Level4Out24[8] , \Level4Out24[7] , \Level4Out24[6] , \Level4Out24[5] , 
        \Level4Out24[4] , \Level4Out24[3] , \Level4Out24[2] , \Level4Out24[1] , 
        \Level4Out24[0] }), .In1({\Level2Out24[31] , \Level2Out24[30] , 
        \Level2Out24[29] , \Level2Out24[28] , \Level2Out24[27] , 
        \Level2Out24[26] , \Level2Out24[25] , \Level2Out24[24] , 
        \Level2Out24[23] , \Level2Out24[22] , \Level2Out24[21] , 
        \Level2Out24[20] , \Level2Out24[19] , \Level2Out24[18] , 
        \Level2Out24[17] , \Level2Out24[16] , \Level2Out24[15] , 
        \Level2Out24[14] , \Level2Out24[13] , \Level2Out24[12] , 
        \Level2Out24[11] , \Level2Out24[10] , \Level2Out24[9] , 
        \Level2Out24[8] , \Level2Out24[7] , \Level2Out24[6] , \Level2Out24[5] , 
        \Level2Out24[4] , \Level2Out24[3] , \Level2Out24[2] , \Level2Out24[1] , 
        \Level2Out24[0] }), .In2({\Level2Out26[31] , \Level2Out26[30] , 
        \Level2Out26[29] , \Level2Out26[28] , \Level2Out26[27] , 
        \Level2Out26[26] , \Level2Out26[25] , \Level2Out26[24] , 
        \Level2Out26[23] , \Level2Out26[22] , \Level2Out26[21] , 
        \Level2Out26[20] , \Level2Out26[19] , \Level2Out26[18] , 
        \Level2Out26[17] , \Level2Out26[16] , \Level2Out26[15] , 
        \Level2Out26[14] , \Level2Out26[13] , \Level2Out26[12] , 
        \Level2Out26[11] , \Level2Out26[10] , \Level2Out26[9] , 
        \Level2Out26[8] , \Level2Out26[7] , \Level2Out26[6] , \Level2Out26[5] , 
        \Level2Out26[4] , \Level2Out26[3] , \Level2Out26[2] , \Level2Out26[1] , 
        \Level2Out26[0] }), .Read1(\Level2Load24[0] ), .Read2(
        \Level2Load26[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_84_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load84[0] ), .Out({\Level2Out84[31] , \Level2Out84[30] , 
        \Level2Out84[29] , \Level2Out84[28] , \Level2Out84[27] , 
        \Level2Out84[26] , \Level2Out84[25] , \Level2Out84[24] , 
        \Level2Out84[23] , \Level2Out84[22] , \Level2Out84[21] , 
        \Level2Out84[20] , \Level2Out84[19] , \Level2Out84[18] , 
        \Level2Out84[17] , \Level2Out84[16] , \Level2Out84[15] , 
        \Level2Out84[14] , \Level2Out84[13] , \Level2Out84[12] , 
        \Level2Out84[11] , \Level2Out84[10] , \Level2Out84[9] , 
        \Level2Out84[8] , \Level2Out84[7] , \Level2Out84[6] , \Level2Out84[5] , 
        \Level2Out84[4] , \Level2Out84[3] , \Level2Out84[2] , \Level2Out84[1] , 
        \Level2Out84[0] }), .In1({\Level1Out84[31] , \Level1Out84[30] , 
        \Level1Out84[29] , \Level1Out84[28] , \Level1Out84[27] , 
        \Level1Out84[26] , \Level1Out84[25] , \Level1Out84[24] , 
        \Level1Out84[23] , \Level1Out84[22] , \Level1Out84[21] , 
        \Level1Out84[20] , \Level1Out84[19] , \Level1Out84[18] , 
        \Level1Out84[17] , \Level1Out84[16] , \Level1Out84[15] , 
        \Level1Out84[14] , \Level1Out84[13] , \Level1Out84[12] , 
        \Level1Out84[11] , \Level1Out84[10] , \Level1Out84[9] , 
        \Level1Out84[8] , \Level1Out84[7] , \Level1Out84[6] , \Level1Out84[5] , 
        \Level1Out84[4] , \Level1Out84[3] , \Level1Out84[2] , \Level1Out84[1] , 
        \Level1Out84[0] }), .In2({\Level1Out85[31] , \Level1Out85[30] , 
        \Level1Out85[29] , \Level1Out85[28] , \Level1Out85[27] , 
        \Level1Out85[26] , \Level1Out85[25] , \Level1Out85[24] , 
        \Level1Out85[23] , \Level1Out85[22] , \Level1Out85[21] , 
        \Level1Out85[20] , \Level1Out85[19] , \Level1Out85[18] , 
        \Level1Out85[17] , \Level1Out85[16] , \Level1Out85[15] , 
        \Level1Out85[14] , \Level1Out85[13] , \Level1Out85[12] , 
        \Level1Out85[11] , \Level1Out85[10] , \Level1Out85[9] , 
        \Level1Out85[8] , \Level1Out85[7] , \Level1Out85[6] , \Level1Out85[5] , 
        \Level1Out85[4] , \Level1Out85[3] , \Level1Out85[2] , \Level1Out85[1] , 
        \Level1Out85[0] }), .Read1(\Level1Load84[0] ), .Read2(
        \Level1Load85[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_44 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanOut({\ScanLink45[31] , 
        \ScanLink45[30] , \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , 
        \ScanLink45[26] , \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , 
        \ScanLink45[22] , \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , 
        \ScanLink45[18] , \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , 
        \ScanLink45[14] , \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , 
        \ScanLink45[10] , \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , 
        \ScanLink45[6] , \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , 
        \ScanLink45[2] , \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load44[0] ), .Out({
        \Level1Out44[31] , \Level1Out44[30] , \Level1Out44[29] , 
        \Level1Out44[28] , \Level1Out44[27] , \Level1Out44[26] , 
        \Level1Out44[25] , \Level1Out44[24] , \Level1Out44[23] , 
        \Level1Out44[22] , \Level1Out44[21] , \Level1Out44[20] , 
        \Level1Out44[19] , \Level1Out44[18] , \Level1Out44[17] , 
        \Level1Out44[16] , \Level1Out44[15] , \Level1Out44[14] , 
        \Level1Out44[13] , \Level1Out44[12] , \Level1Out44[11] , 
        \Level1Out44[10] , \Level1Out44[9] , \Level1Out44[8] , 
        \Level1Out44[7] , \Level1Out44[6] , \Level1Out44[5] , \Level1Out44[4] , 
        \Level1Out44[3] , \Level1Out44[2] , \Level1Out44[1] , \Level1Out44[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_78 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink78[31] , \ScanLink78[30] , 
        \ScanLink78[29] , \ScanLink78[28] , \ScanLink78[27] , \ScanLink78[26] , 
        \ScanLink78[25] , \ScanLink78[24] , \ScanLink78[23] , \ScanLink78[22] , 
        \ScanLink78[21] , \ScanLink78[20] , \ScanLink78[19] , \ScanLink78[18] , 
        \ScanLink78[17] , \ScanLink78[16] , \ScanLink78[15] , \ScanLink78[14] , 
        \ScanLink78[13] , \ScanLink78[12] , \ScanLink78[11] , \ScanLink78[10] , 
        \ScanLink78[9] , \ScanLink78[8] , \ScanLink78[7] , \ScanLink78[6] , 
        \ScanLink78[5] , \ScanLink78[4] , \ScanLink78[3] , \ScanLink78[2] , 
        \ScanLink78[1] , \ScanLink78[0] }), .ScanOut({\ScanLink79[31] , 
        \ScanLink79[30] , \ScanLink79[29] , \ScanLink79[28] , \ScanLink79[27] , 
        \ScanLink79[26] , \ScanLink79[25] , \ScanLink79[24] , \ScanLink79[23] , 
        \ScanLink79[22] , \ScanLink79[21] , \ScanLink79[20] , \ScanLink79[19] , 
        \ScanLink79[18] , \ScanLink79[17] , \ScanLink79[16] , \ScanLink79[15] , 
        \ScanLink79[14] , \ScanLink79[13] , \ScanLink79[12] , \ScanLink79[11] , 
        \ScanLink79[10] , \ScanLink79[9] , \ScanLink79[8] , \ScanLink79[7] , 
        \ScanLink79[6] , \ScanLink79[5] , \ScanLink79[4] , \ScanLink79[3] , 
        \ScanLink79[2] , \ScanLink79[1] , \ScanLink79[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load78[0] ), .Out({
        \Level1Out78[31] , \Level1Out78[30] , \Level1Out78[29] , 
        \Level1Out78[28] , \Level1Out78[27] , \Level1Out78[26] , 
        \Level1Out78[25] , \Level1Out78[24] , \Level1Out78[23] , 
        \Level1Out78[22] , \Level1Out78[21] , \Level1Out78[20] , 
        \Level1Out78[19] , \Level1Out78[18] , \Level1Out78[17] , 
        \Level1Out78[16] , \Level1Out78[15] , \Level1Out78[14] , 
        \Level1Out78[13] , \Level1Out78[12] , \Level1Out78[11] , 
        \Level1Out78[10] , \Level1Out78[9] , \Level1Out78[8] , 
        \Level1Out78[7] , \Level1Out78[6] , \Level1Out78[5] , \Level1Out78[4] , 
        \Level1Out78[3] , \Level1Out78[2] , \Level1Out78[1] , \Level1Out78[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_198 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink198[31] , \ScanLink198[30] , 
        \ScanLink198[29] , \ScanLink198[28] , \ScanLink198[27] , 
        \ScanLink198[26] , \ScanLink198[25] , \ScanLink198[24] , 
        \ScanLink198[23] , \ScanLink198[22] , \ScanLink198[21] , 
        \ScanLink198[20] , \ScanLink198[19] , \ScanLink198[18] , 
        \ScanLink198[17] , \ScanLink198[16] , \ScanLink198[15] , 
        \ScanLink198[14] , \ScanLink198[13] , \ScanLink198[12] , 
        \ScanLink198[11] , \ScanLink198[10] , \ScanLink198[9] , 
        \ScanLink198[8] , \ScanLink198[7] , \ScanLink198[6] , \ScanLink198[5] , 
        \ScanLink198[4] , \ScanLink198[3] , \ScanLink198[2] , \ScanLink198[1] , 
        \ScanLink198[0] }), .ScanOut({\ScanLink199[31] , \ScanLink199[30] , 
        \ScanLink199[29] , \ScanLink199[28] , \ScanLink199[27] , 
        \ScanLink199[26] , \ScanLink199[25] , \ScanLink199[24] , 
        \ScanLink199[23] , \ScanLink199[22] , \ScanLink199[21] , 
        \ScanLink199[20] , \ScanLink199[19] , \ScanLink199[18] , 
        \ScanLink199[17] , \ScanLink199[16] , \ScanLink199[15] , 
        \ScanLink199[14] , \ScanLink199[13] , \ScanLink199[12] , 
        \ScanLink199[11] , \ScanLink199[10] , \ScanLink199[9] , 
        \ScanLink199[8] , \ScanLink199[7] , \ScanLink199[6] , \ScanLink199[5] , 
        \ScanLink199[4] , \ScanLink199[3] , \ScanLink199[2] , \ScanLink199[1] , 
        \ScanLink199[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load198[0] ), .Out({\Level1Out198[31] , \Level1Out198[30] , 
        \Level1Out198[29] , \Level1Out198[28] , \Level1Out198[27] , 
        \Level1Out198[26] , \Level1Out198[25] , \Level1Out198[24] , 
        \Level1Out198[23] , \Level1Out198[22] , \Level1Out198[21] , 
        \Level1Out198[20] , \Level1Out198[19] , \Level1Out198[18] , 
        \Level1Out198[17] , \Level1Out198[16] , \Level1Out198[15] , 
        \Level1Out198[14] , \Level1Out198[13] , \Level1Out198[12] , 
        \Level1Out198[11] , \Level1Out198[10] , \Level1Out198[9] , 
        \Level1Out198[8] , \Level1Out198[7] , \Level1Out198[6] , 
        \Level1Out198[5] , \Level1Out198[4] , \Level1Out198[3] , 
        \Level1Out198[2] , \Level1Out198[1] , \Level1Out198[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_160_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load160[0] ), .Out({\Level8Out160[31] , \Level8Out160[30] , 
        \Level8Out160[29] , \Level8Out160[28] , \Level8Out160[27] , 
        \Level8Out160[26] , \Level8Out160[25] , \Level8Out160[24] , 
        \Level8Out160[23] , \Level8Out160[22] , \Level8Out160[21] , 
        \Level8Out160[20] , \Level8Out160[19] , \Level8Out160[18] , 
        \Level8Out160[17] , \Level8Out160[16] , \Level8Out160[15] , 
        \Level8Out160[14] , \Level8Out160[13] , \Level8Out160[12] , 
        \Level8Out160[11] , \Level8Out160[10] , \Level8Out160[9] , 
        \Level8Out160[8] , \Level8Out160[7] , \Level8Out160[6] , 
        \Level8Out160[5] , \Level8Out160[4] , \Level8Out160[3] , 
        \Level8Out160[2] , \Level8Out160[1] , \Level8Out160[0] }), .In1({
        \Level4Out160[31] , \Level4Out160[30] , \Level4Out160[29] , 
        \Level4Out160[28] , \Level4Out160[27] , \Level4Out160[26] , 
        \Level4Out160[25] , \Level4Out160[24] , \Level4Out160[23] , 
        \Level4Out160[22] , \Level4Out160[21] , \Level4Out160[20] , 
        \Level4Out160[19] , \Level4Out160[18] , \Level4Out160[17] , 
        \Level4Out160[16] , \Level4Out160[15] , \Level4Out160[14] , 
        \Level4Out160[13] , \Level4Out160[12] , \Level4Out160[11] , 
        \Level4Out160[10] , \Level4Out160[9] , \Level4Out160[8] , 
        \Level4Out160[7] , \Level4Out160[6] , \Level4Out160[5] , 
        \Level4Out160[4] , \Level4Out160[3] , \Level4Out160[2] , 
        \Level4Out160[1] , \Level4Out160[0] }), .In2({\Level4Out164[31] , 
        \Level4Out164[30] , \Level4Out164[29] , \Level4Out164[28] , 
        \Level4Out164[27] , \Level4Out164[26] , \Level4Out164[25] , 
        \Level4Out164[24] , \Level4Out164[23] , \Level4Out164[22] , 
        \Level4Out164[21] , \Level4Out164[20] , \Level4Out164[19] , 
        \Level4Out164[18] , \Level4Out164[17] , \Level4Out164[16] , 
        \Level4Out164[15] , \Level4Out164[14] , \Level4Out164[13] , 
        \Level4Out164[12] , \Level4Out164[11] , \Level4Out164[10] , 
        \Level4Out164[9] , \Level4Out164[8] , \Level4Out164[7] , 
        \Level4Out164[6] , \Level4Out164[5] , \Level4Out164[4] , 
        \Level4Out164[3] , \Level4Out164[2] , \Level4Out164[1] , 
        \Level4Out164[0] }), .Read1(\Level4Load160[0] ), .Read2(
        \Level4Load164[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_141 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink141[31] , \ScanLink141[30] , 
        \ScanLink141[29] , \ScanLink141[28] , \ScanLink141[27] , 
        \ScanLink141[26] , \ScanLink141[25] , \ScanLink141[24] , 
        \ScanLink141[23] , \ScanLink141[22] , \ScanLink141[21] , 
        \ScanLink141[20] , \ScanLink141[19] , \ScanLink141[18] , 
        \ScanLink141[17] , \ScanLink141[16] , \ScanLink141[15] , 
        \ScanLink141[14] , \ScanLink141[13] , \ScanLink141[12] , 
        \ScanLink141[11] , \ScanLink141[10] , \ScanLink141[9] , 
        \ScanLink141[8] , \ScanLink141[7] , \ScanLink141[6] , \ScanLink141[5] , 
        \ScanLink141[4] , \ScanLink141[3] , \ScanLink141[2] , \ScanLink141[1] , 
        \ScanLink141[0] }), .ScanOut({\ScanLink142[31] , \ScanLink142[30] , 
        \ScanLink142[29] , \ScanLink142[28] , \ScanLink142[27] , 
        \ScanLink142[26] , \ScanLink142[25] , \ScanLink142[24] , 
        \ScanLink142[23] , \ScanLink142[22] , \ScanLink142[21] , 
        \ScanLink142[20] , \ScanLink142[19] , \ScanLink142[18] , 
        \ScanLink142[17] , \ScanLink142[16] , \ScanLink142[15] , 
        \ScanLink142[14] , \ScanLink142[13] , \ScanLink142[12] , 
        \ScanLink142[11] , \ScanLink142[10] , \ScanLink142[9] , 
        \ScanLink142[8] , \ScanLink142[7] , \ScanLink142[6] , \ScanLink142[5] , 
        \ScanLink142[4] , \ScanLink142[3] , \ScanLink142[2] , \ScanLink142[1] , 
        \ScanLink142[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load141[0] ), .Out({\Level1Out141[31] , \Level1Out141[30] , 
        \Level1Out141[29] , \Level1Out141[28] , \Level1Out141[27] , 
        \Level1Out141[26] , \Level1Out141[25] , \Level1Out141[24] , 
        \Level1Out141[23] , \Level1Out141[22] , \Level1Out141[21] , 
        \Level1Out141[20] , \Level1Out141[19] , \Level1Out141[18] , 
        \Level1Out141[17] , \Level1Out141[16] , \Level1Out141[15] , 
        \Level1Out141[14] , \Level1Out141[13] , \Level1Out141[12] , 
        \Level1Out141[11] , \Level1Out141[10] , \Level1Out141[9] , 
        \Level1Out141[8] , \Level1Out141[7] , \Level1Out141[6] , 
        \Level1Out141[5] , \Level1Out141[4] , \Level1Out141[3] , 
        \Level1Out141[2] , \Level1Out141[1] , \Level1Out141[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_166 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink166[31] , \ScanLink166[30] , 
        \ScanLink166[29] , \ScanLink166[28] , \ScanLink166[27] , 
        \ScanLink166[26] , \ScanLink166[25] , \ScanLink166[24] , 
        \ScanLink166[23] , \ScanLink166[22] , \ScanLink166[21] , 
        \ScanLink166[20] , \ScanLink166[19] , \ScanLink166[18] , 
        \ScanLink166[17] , \ScanLink166[16] , \ScanLink166[15] , 
        \ScanLink166[14] , \ScanLink166[13] , \ScanLink166[12] , 
        \ScanLink166[11] , \ScanLink166[10] , \ScanLink166[9] , 
        \ScanLink166[8] , \ScanLink166[7] , \ScanLink166[6] , \ScanLink166[5] , 
        \ScanLink166[4] , \ScanLink166[3] , \ScanLink166[2] , \ScanLink166[1] , 
        \ScanLink166[0] }), .ScanOut({\ScanLink167[31] , \ScanLink167[30] , 
        \ScanLink167[29] , \ScanLink167[28] , \ScanLink167[27] , 
        \ScanLink167[26] , \ScanLink167[25] , \ScanLink167[24] , 
        \ScanLink167[23] , \ScanLink167[22] , \ScanLink167[21] , 
        \ScanLink167[20] , \ScanLink167[19] , \ScanLink167[18] , 
        \ScanLink167[17] , \ScanLink167[16] , \ScanLink167[15] , 
        \ScanLink167[14] , \ScanLink167[13] , \ScanLink167[12] , 
        \ScanLink167[11] , \ScanLink167[10] , \ScanLink167[9] , 
        \ScanLink167[8] , \ScanLink167[7] , \ScanLink167[6] , \ScanLink167[5] , 
        \ScanLink167[4] , \ScanLink167[3] , \ScanLink167[2] , \ScanLink167[1] , 
        \ScanLink167[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load166[0] ), .Out({\Level1Out166[31] , \Level1Out166[30] , 
        \Level1Out166[29] , \Level1Out166[28] , \Level1Out166[27] , 
        \Level1Out166[26] , \Level1Out166[25] , \Level1Out166[24] , 
        \Level1Out166[23] , \Level1Out166[22] , \Level1Out166[21] , 
        \Level1Out166[20] , \Level1Out166[19] , \Level1Out166[18] , 
        \Level1Out166[17] , \Level1Out166[16] , \Level1Out166[15] , 
        \Level1Out166[14] , \Level1Out166[13] , \Level1Out166[12] , 
        \Level1Out166[11] , \Level1Out166[10] , \Level1Out166[9] , 
        \Level1Out166[8] , \Level1Out166[7] , \Level1Out166[6] , 
        \Level1Out166[5] , \Level1Out166[4] , \Level1Out166[3] , 
        \Level1Out166[2] , \Level1Out166[1] , \Level1Out166[0] }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_63 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanOut({\ScanLink64[31] , 
        \ScanLink64[30] , \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , 
        \ScanLink64[26] , \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , 
        \ScanLink64[22] , \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , 
        \ScanLink64[18] , \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , 
        \ScanLink64[14] , \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , 
        \ScanLink64[10] , \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , 
        \ScanLink64[6] , \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , 
        \ScanLink64[2] , \ScanLink64[1] , \ScanLink64[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load63[0] ), .Out({
        \Level1Out63[31] , \Level1Out63[30] , \Level1Out63[29] , 
        \Level1Out63[28] , \Level1Out63[27] , \Level1Out63[26] , 
        \Level1Out63[25] , \Level1Out63[24] , \Level1Out63[23] , 
        \Level1Out63[22] , \Level1Out63[21] , \Level1Out63[20] , 
        \Level1Out63[19] , \Level1Out63[18] , \Level1Out63[17] , 
        \Level1Out63[16] , \Level1Out63[15] , \Level1Out63[14] , 
        \Level1Out63[13] , \Level1Out63[12] , \Level1Out63[11] , 
        \Level1Out63[10] , \Level1Out63[9] , \Level1Out63[8] , 
        \Level1Out63[7] , \Level1Out63[6] , \Level1Out63[5] , \Level1Out63[4] , 
        \Level1Out63[3] , \Level1Out63[2] , \Level1Out63[1] , \Level1Out63[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_86 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink86[31] , \ScanLink86[30] , 
        \ScanLink86[29] , \ScanLink86[28] , \ScanLink86[27] , \ScanLink86[26] , 
        \ScanLink86[25] , \ScanLink86[24] , \ScanLink86[23] , \ScanLink86[22] , 
        \ScanLink86[21] , \ScanLink86[20] , \ScanLink86[19] , \ScanLink86[18] , 
        \ScanLink86[17] , \ScanLink86[16] , \ScanLink86[15] , \ScanLink86[14] , 
        \ScanLink86[13] , \ScanLink86[12] , \ScanLink86[11] , \ScanLink86[10] , 
        \ScanLink86[9] , \ScanLink86[8] , \ScanLink86[7] , \ScanLink86[6] , 
        \ScanLink86[5] , \ScanLink86[4] , \ScanLink86[3] , \ScanLink86[2] , 
        \ScanLink86[1] , \ScanLink86[0] }), .ScanOut({\ScanLink87[31] , 
        \ScanLink87[30] , \ScanLink87[29] , \ScanLink87[28] , \ScanLink87[27] , 
        \ScanLink87[26] , \ScanLink87[25] , \ScanLink87[24] , \ScanLink87[23] , 
        \ScanLink87[22] , \ScanLink87[21] , \ScanLink87[20] , \ScanLink87[19] , 
        \ScanLink87[18] , \ScanLink87[17] , \ScanLink87[16] , \ScanLink87[15] , 
        \ScanLink87[14] , \ScanLink87[13] , \ScanLink87[12] , \ScanLink87[11] , 
        \ScanLink87[10] , \ScanLink87[9] , \ScanLink87[8] , \ScanLink87[7] , 
        \ScanLink87[6] , \ScanLink87[5] , \ScanLink87[4] , \ScanLink87[3] , 
        \ScanLink87[2] , \ScanLink87[1] , \ScanLink87[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load86[0] ), .Out({
        \Level1Out86[31] , \Level1Out86[30] , \Level1Out86[29] , 
        \Level1Out86[28] , \Level1Out86[27] , \Level1Out86[26] , 
        \Level1Out86[25] , \Level1Out86[24] , \Level1Out86[23] , 
        \Level1Out86[22] , \Level1Out86[21] , \Level1Out86[20] , 
        \Level1Out86[19] , \Level1Out86[18] , \Level1Out86[17] , 
        \Level1Out86[16] , \Level1Out86[15] , \Level1Out86[14] , 
        \Level1Out86[13] , \Level1Out86[12] , \Level1Out86[11] , 
        \Level1Out86[10] , \Level1Out86[9] , \Level1Out86[8] , 
        \Level1Out86[7] , \Level1Out86[6] , \Level1Out86[5] , \Level1Out86[4] , 
        \Level1Out86[3] , \Level1Out86[2] , \Level1Out86[1] , \Level1Out86[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_183 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink183[31] , \ScanLink183[30] , 
        \ScanLink183[29] , \ScanLink183[28] , \ScanLink183[27] , 
        \ScanLink183[26] , \ScanLink183[25] , \ScanLink183[24] , 
        \ScanLink183[23] , \ScanLink183[22] , \ScanLink183[21] , 
        \ScanLink183[20] , \ScanLink183[19] , \ScanLink183[18] , 
        \ScanLink183[17] , \ScanLink183[16] , \ScanLink183[15] , 
        \ScanLink183[14] , \ScanLink183[13] , \ScanLink183[12] , 
        \ScanLink183[11] , \ScanLink183[10] , \ScanLink183[9] , 
        \ScanLink183[8] , \ScanLink183[7] , \ScanLink183[6] , \ScanLink183[5] , 
        \ScanLink183[4] , \ScanLink183[3] , \ScanLink183[2] , \ScanLink183[1] , 
        \ScanLink183[0] }), .ScanOut({\ScanLink184[31] , \ScanLink184[30] , 
        \ScanLink184[29] , \ScanLink184[28] , \ScanLink184[27] , 
        \ScanLink184[26] , \ScanLink184[25] , \ScanLink184[24] , 
        \ScanLink184[23] , \ScanLink184[22] , \ScanLink184[21] , 
        \ScanLink184[20] , \ScanLink184[19] , \ScanLink184[18] , 
        \ScanLink184[17] , \ScanLink184[16] , \ScanLink184[15] , 
        \ScanLink184[14] , \ScanLink184[13] , \ScanLink184[12] , 
        \ScanLink184[11] , \ScanLink184[10] , \ScanLink184[9] , 
        \ScanLink184[8] , \ScanLink184[7] , \ScanLink184[6] , \ScanLink184[5] , 
        \ScanLink184[4] , \ScanLink184[3] , \ScanLink184[2] , \ScanLink184[1] , 
        \ScanLink184[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b1), .Load(
        \Level1Load183[0] ), .Out({\Level1Out183[31] , \Level1Out183[30] , 
        \Level1Out183[29] , \Level1Out183[28] , \Level1Out183[27] , 
        \Level1Out183[26] , \Level1Out183[25] , \Level1Out183[24] , 
        \Level1Out183[23] , \Level1Out183[22] , \Level1Out183[21] , 
        \Level1Out183[20] , \Level1Out183[19] , \Level1Out183[18] , 
        \Level1Out183[17] , \Level1Out183[16] , \Level1Out183[15] , 
        \Level1Out183[14] , \Level1Out183[13] , \Level1Out183[12] , 
        \Level1Out183[11] , \Level1Out183[10] , \Level1Out183[9] , 
        \Level1Out183[8] , \Level1Out183[7] , \Level1Out183[6] , 
        \Level1Out183[5] , \Level1Out183[4] , \Level1Out183[3] , 
        \Level1Out183[2] , \Level1Out183[1] , \Level1Out183[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_166_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load166[0] ), .Out({\Level2Out166[31] , \Level2Out166[30] , 
        \Level2Out166[29] , \Level2Out166[28] , \Level2Out166[27] , 
        \Level2Out166[26] , \Level2Out166[25] , \Level2Out166[24] , 
        \Level2Out166[23] , \Level2Out166[22] , \Level2Out166[21] , 
        \Level2Out166[20] , \Level2Out166[19] , \Level2Out166[18] , 
        \Level2Out166[17] , \Level2Out166[16] , \Level2Out166[15] , 
        \Level2Out166[14] , \Level2Out166[13] , \Level2Out166[12] , 
        \Level2Out166[11] , \Level2Out166[10] , \Level2Out166[9] , 
        \Level2Out166[8] , \Level2Out166[7] , \Level2Out166[6] , 
        \Level2Out166[5] , \Level2Out166[4] , \Level2Out166[3] , 
        \Level2Out166[2] , \Level2Out166[1] , \Level2Out166[0] }), .In1({
        \Level1Out166[31] , \Level1Out166[30] , \Level1Out166[29] , 
        \Level1Out166[28] , \Level1Out166[27] , \Level1Out166[26] , 
        \Level1Out166[25] , \Level1Out166[24] , \Level1Out166[23] , 
        \Level1Out166[22] , \Level1Out166[21] , \Level1Out166[20] , 
        \Level1Out166[19] , \Level1Out166[18] , \Level1Out166[17] , 
        \Level1Out166[16] , \Level1Out166[15] , \Level1Out166[14] , 
        \Level1Out166[13] , \Level1Out166[12] , \Level1Out166[11] , 
        \Level1Out166[10] , \Level1Out166[9] , \Level1Out166[8] , 
        \Level1Out166[7] , \Level1Out166[6] , \Level1Out166[5] , 
        \Level1Out166[4] , \Level1Out166[3] , \Level1Out166[2] , 
        \Level1Out166[1] , \Level1Out166[0] }), .In2({\Level1Out167[31] , 
        \Level1Out167[30] , \Level1Out167[29] , \Level1Out167[28] , 
        \Level1Out167[27] , \Level1Out167[26] , \Level1Out167[25] , 
        \Level1Out167[24] , \Level1Out167[23] , \Level1Out167[22] , 
        \Level1Out167[21] , \Level1Out167[20] , \Level1Out167[19] , 
        \Level1Out167[18] , \Level1Out167[17] , \Level1Out167[16] , 
        \Level1Out167[15] , \Level1Out167[14] , \Level1Out167[13] , 
        \Level1Out167[12] , \Level1Out167[11] , \Level1Out167[10] , 
        \Level1Out167[9] , \Level1Out167[8] , \Level1Out167[7] , 
        \Level1Out167[6] , \Level1Out167[5] , \Level1Out167[4] , 
        \Level1Out167[3] , \Level1Out167[2] , \Level1Out167[1] , 
        \Level1Out167[0] }), .Read1(\Level1Load166[0] ), .Read2(
        \Level1Load167[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load16[0] ), .Out({\Level4Out16[31] , \Level4Out16[30] , 
        \Level4Out16[29] , \Level4Out16[28] , \Level4Out16[27] , 
        \Level4Out16[26] , \Level4Out16[25] , \Level4Out16[24] , 
        \Level4Out16[23] , \Level4Out16[22] , \Level4Out16[21] , 
        \Level4Out16[20] , \Level4Out16[19] , \Level4Out16[18] , 
        \Level4Out16[17] , \Level4Out16[16] , \Level4Out16[15] , 
        \Level4Out16[14] , \Level4Out16[13] , \Level4Out16[12] , 
        \Level4Out16[11] , \Level4Out16[10] , \Level4Out16[9] , 
        \Level4Out16[8] , \Level4Out16[7] , \Level4Out16[6] , \Level4Out16[5] , 
        \Level4Out16[4] , \Level4Out16[3] , \Level4Out16[2] , \Level4Out16[1] , 
        \Level4Out16[0] }), .In1({\Level2Out16[31] , \Level2Out16[30] , 
        \Level2Out16[29] , \Level2Out16[28] , \Level2Out16[27] , 
        \Level2Out16[26] , \Level2Out16[25] , \Level2Out16[24] , 
        \Level2Out16[23] , \Level2Out16[22] , \Level2Out16[21] , 
        \Level2Out16[20] , \Level2Out16[19] , \Level2Out16[18] , 
        \Level2Out16[17] , \Level2Out16[16] , \Level2Out16[15] , 
        \Level2Out16[14] , \Level2Out16[13] , \Level2Out16[12] , 
        \Level2Out16[11] , \Level2Out16[10] , \Level2Out16[9] , 
        \Level2Out16[8] , \Level2Out16[7] , \Level2Out16[6] , \Level2Out16[5] , 
        \Level2Out16[4] , \Level2Out16[3] , \Level2Out16[2] , \Level2Out16[1] , 
        \Level2Out16[0] }), .In2({\Level2Out18[31] , \Level2Out18[30] , 
        \Level2Out18[29] , \Level2Out18[28] , \Level2Out18[27] , 
        \Level2Out18[26] , \Level2Out18[25] , \Level2Out18[24] , 
        \Level2Out18[23] , \Level2Out18[22] , \Level2Out18[21] , 
        \Level2Out18[20] , \Level2Out18[19] , \Level2Out18[18] , 
        \Level2Out18[17] , \Level2Out18[16] , \Level2Out18[15] , 
        \Level2Out18[14] , \Level2Out18[13] , \Level2Out18[12] , 
        \Level2Out18[11] , \Level2Out18[10] , \Level2Out18[9] , 
        \Level2Out18[8] , \Level2Out18[7] , \Level2Out18[6] , \Level2Out18[5] , 
        \Level2Out18[4] , \Level2Out18[3] , \Level2Out18[2] , \Level2Out18[1] , 
        \Level2Out18[0] }), .Read1(\Level2Load16[0] ), .Read2(
        \Level2Load18[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_238 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink238[31] , \ScanLink238[30] , 
        \ScanLink238[29] , \ScanLink238[28] , \ScanLink238[27] , 
        \ScanLink238[26] , \ScanLink238[25] , \ScanLink238[24] , 
        \ScanLink238[23] , \ScanLink238[22] , \ScanLink238[21] , 
        \ScanLink238[20] , \ScanLink238[19] , \ScanLink238[18] , 
        \ScanLink238[17] , \ScanLink238[16] , \ScanLink238[15] , 
        \ScanLink238[14] , \ScanLink238[13] , \ScanLink238[12] , 
        \ScanLink238[11] , \ScanLink238[10] , \ScanLink238[9] , 
        \ScanLink238[8] , \ScanLink238[7] , \ScanLink238[6] , \ScanLink238[5] , 
        \ScanLink238[4] , \ScanLink238[3] , \ScanLink238[2] , \ScanLink238[1] , 
        \ScanLink238[0] }), .ScanOut({\ScanLink239[31] , \ScanLink239[30] , 
        \ScanLink239[29] , \ScanLink239[28] , \ScanLink239[27] , 
        \ScanLink239[26] , \ScanLink239[25] , \ScanLink239[24] , 
        \ScanLink239[23] , \ScanLink239[22] , \ScanLink239[21] , 
        \ScanLink239[20] , \ScanLink239[19] , \ScanLink239[18] , 
        \ScanLink239[17] , \ScanLink239[16] , \ScanLink239[15] , 
        \ScanLink239[14] , \ScanLink239[13] , \ScanLink239[12] , 
        \ScanLink239[11] , \ScanLink239[10] , \ScanLink239[9] , 
        \ScanLink239[8] , \ScanLink239[7] , \ScanLink239[6] , \ScanLink239[5] , 
        \ScanLink239[4] , \ScanLink239[3] , \ScanLink239[2] , \ScanLink239[1] , 
        \ScanLink239[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load238[0] ), .Out({\Level1Out238[31] , \Level1Out238[30] , 
        \Level1Out238[29] , \Level1Out238[28] , \Level1Out238[27] , 
        \Level1Out238[26] , \Level1Out238[25] , \Level1Out238[24] , 
        \Level1Out238[23] , \Level1Out238[22] , \Level1Out238[21] , 
        \Level1Out238[20] , \Level1Out238[19] , \Level1Out238[18] , 
        \Level1Out238[17] , \Level1Out238[16] , \Level1Out238[15] , 
        \Level1Out238[14] , \Level1Out238[13] , \Level1Out238[12] , 
        \Level1Out238[11] , \Level1Out238[10] , \Level1Out238[9] , 
        \Level1Out238[8] , \Level1Out238[7] , \Level1Out238[6] , 
        \Level1Out238[5] , \Level1Out238[4] , \Level1Out238[3] , 
        \Level1Out238[2] , \Level1Out238[1] , \Level1Out238[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_20_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load20[0] ), .Out({\Level2Out20[31] , \Level2Out20[30] , 
        \Level2Out20[29] , \Level2Out20[28] , \Level2Out20[27] , 
        \Level2Out20[26] , \Level2Out20[25] , \Level2Out20[24] , 
        \Level2Out20[23] , \Level2Out20[22] , \Level2Out20[21] , 
        \Level2Out20[20] , \Level2Out20[19] , \Level2Out20[18] , 
        \Level2Out20[17] , \Level2Out20[16] , \Level2Out20[15] , 
        \Level2Out20[14] , \Level2Out20[13] , \Level2Out20[12] , 
        \Level2Out20[11] , \Level2Out20[10] , \Level2Out20[9] , 
        \Level2Out20[8] , \Level2Out20[7] , \Level2Out20[6] , \Level2Out20[5] , 
        \Level2Out20[4] , \Level2Out20[3] , \Level2Out20[2] , \Level2Out20[1] , 
        \Level2Out20[0] }), .In1({\Level1Out20[31] , \Level1Out20[30] , 
        \Level1Out20[29] , \Level1Out20[28] , \Level1Out20[27] , 
        \Level1Out20[26] , \Level1Out20[25] , \Level1Out20[24] , 
        \Level1Out20[23] , \Level1Out20[22] , \Level1Out20[21] , 
        \Level1Out20[20] , \Level1Out20[19] , \Level1Out20[18] , 
        \Level1Out20[17] , \Level1Out20[16] , \Level1Out20[15] , 
        \Level1Out20[14] , \Level1Out20[13] , \Level1Out20[12] , 
        \Level1Out20[11] , \Level1Out20[10] , \Level1Out20[9] , 
        \Level1Out20[8] , \Level1Out20[7] , \Level1Out20[6] , \Level1Out20[5] , 
        \Level1Out20[4] , \Level1Out20[3] , \Level1Out20[2] , \Level1Out20[1] , 
        \Level1Out20[0] }), .In2({\Level1Out21[31] , \Level1Out21[30] , 
        \Level1Out21[29] , \Level1Out21[28] , \Level1Out21[27] , 
        \Level1Out21[26] , \Level1Out21[25] , \Level1Out21[24] , 
        \Level1Out21[23] , \Level1Out21[22] , \Level1Out21[21] , 
        \Level1Out21[20] , \Level1Out21[19] , \Level1Out21[18] , 
        \Level1Out21[17] , \Level1Out21[16] , \Level1Out21[15] , 
        \Level1Out21[14] , \Level1Out21[13] , \Level1Out21[12] , 
        \Level1Out21[11] , \Level1Out21[10] , \Level1Out21[9] , 
        \Level1Out21[8] , \Level1Out21[7] , \Level1Out21[6] , \Level1Out21[5] , 
        \Level1Out21[4] , \Level1Out21[3] , \Level1Out21[2] , \Level1Out21[1] , 
        \Level1Out21[0] }), .Read1(\Level1Load20[0] ), .Read2(
        \Level1Load21[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_80_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load80[0] ), .Out({\Level16Out80[31] , \Level16Out80[30] , 
        \Level16Out80[29] , \Level16Out80[28] , \Level16Out80[27] , 
        \Level16Out80[26] , \Level16Out80[25] , \Level16Out80[24] , 
        \Level16Out80[23] , \Level16Out80[22] , \Level16Out80[21] , 
        \Level16Out80[20] , \Level16Out80[19] , \Level16Out80[18] , 
        \Level16Out80[17] , \Level16Out80[16] , \Level16Out80[15] , 
        \Level16Out80[14] , \Level16Out80[13] , \Level16Out80[12] , 
        \Level16Out80[11] , \Level16Out80[10] , \Level16Out80[9] , 
        \Level16Out80[8] , \Level16Out80[7] , \Level16Out80[6] , 
        \Level16Out80[5] , \Level16Out80[4] , \Level16Out80[3] , 
        \Level16Out80[2] , \Level16Out80[1] , \Level16Out80[0] }), .In1({
        \Level8Out80[31] , \Level8Out80[30] , \Level8Out80[29] , 
        \Level8Out80[28] , \Level8Out80[27] , \Level8Out80[26] , 
        \Level8Out80[25] , \Level8Out80[24] , \Level8Out80[23] , 
        \Level8Out80[22] , \Level8Out80[21] , \Level8Out80[20] , 
        \Level8Out80[19] , \Level8Out80[18] , \Level8Out80[17] , 
        \Level8Out80[16] , \Level8Out80[15] , \Level8Out80[14] , 
        \Level8Out80[13] , \Level8Out80[12] , \Level8Out80[11] , 
        \Level8Out80[10] , \Level8Out80[9] , \Level8Out80[8] , 
        \Level8Out80[7] , \Level8Out80[6] , \Level8Out80[5] , \Level8Out80[4] , 
        \Level8Out80[3] , \Level8Out80[2] , \Level8Out80[1] , \Level8Out80[0] 
        }), .In2({\Level8Out88[31] , \Level8Out88[30] , \Level8Out88[29] , 
        \Level8Out88[28] , \Level8Out88[27] , \Level8Out88[26] , 
        \Level8Out88[25] , \Level8Out88[24] , \Level8Out88[23] , 
        \Level8Out88[22] , \Level8Out88[21] , \Level8Out88[20] , 
        \Level8Out88[19] , \Level8Out88[18] , \Level8Out88[17] , 
        \Level8Out88[16] , \Level8Out88[15] , \Level8Out88[14] , 
        \Level8Out88[13] , \Level8Out88[12] , \Level8Out88[11] , 
        \Level8Out88[10] , \Level8Out88[9] , \Level8Out88[8] , 
        \Level8Out88[7] , \Level8Out88[6] , \Level8Out88[5] , \Level8Out88[4] , 
        \Level8Out88[3] , \Level8Out88[2] , \Level8Out88[1] , \Level8Out88[0] 
        }), .Read1(\Level8Load80[0] ), .Read2(\Level8Load88[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_252_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load252[0] ), .Out({\Level2Out252[31] , \Level2Out252[30] , 
        \Level2Out252[29] , \Level2Out252[28] , \Level2Out252[27] , 
        \Level2Out252[26] , \Level2Out252[25] , \Level2Out252[24] , 
        \Level2Out252[23] , \Level2Out252[22] , \Level2Out252[21] , 
        \Level2Out252[20] , \Level2Out252[19] , \Level2Out252[18] , 
        \Level2Out252[17] , \Level2Out252[16] , \Level2Out252[15] , 
        \Level2Out252[14] , \Level2Out252[13] , \Level2Out252[12] , 
        \Level2Out252[11] , \Level2Out252[10] , \Level2Out252[9] , 
        \Level2Out252[8] , \Level2Out252[7] , \Level2Out252[6] , 
        \Level2Out252[5] , \Level2Out252[4] , \Level2Out252[3] , 
        \Level2Out252[2] , \Level2Out252[1] , \Level2Out252[0] }), .In1({
        \Level1Out252[31] , \Level1Out252[30] , \Level1Out252[29] , 
        \Level1Out252[28] , \Level1Out252[27] , \Level1Out252[26] , 
        \Level1Out252[25] , \Level1Out252[24] , \Level1Out252[23] , 
        \Level1Out252[22] , \Level1Out252[21] , \Level1Out252[20] , 
        \Level1Out252[19] , \Level1Out252[18] , \Level1Out252[17] , 
        \Level1Out252[16] , \Level1Out252[15] , \Level1Out252[14] , 
        \Level1Out252[13] , \Level1Out252[12] , \Level1Out252[11] , 
        \Level1Out252[10] , \Level1Out252[9] , \Level1Out252[8] , 
        \Level1Out252[7] , \Level1Out252[6] , \Level1Out252[5] , 
        \Level1Out252[4] , \Level1Out252[3] , \Level1Out252[2] , 
        \Level1Out252[1] , \Level1Out252[0] }), .In2({\Level1Out253[31] , 
        \Level1Out253[30] , \Level1Out253[29] , \Level1Out253[28] , 
        \Level1Out253[27] , \Level1Out253[26] , \Level1Out253[25] , 
        \Level1Out253[24] , \Level1Out253[23] , \Level1Out253[22] , 
        \Level1Out253[21] , \Level1Out253[20] , \Level1Out253[19] , 
        \Level1Out253[18] , \Level1Out253[17] , \Level1Out253[16] , 
        \Level1Out253[15] , \Level1Out253[14] , \Level1Out253[13] , 
        \Level1Out253[12] , \Level1Out253[11] , \Level1Out253[10] , 
        \Level1Out253[9] , \Level1Out253[8] , \Level1Out253[7] , 
        \Level1Out253[6] , \Level1Out253[5] , \Level1Out253[4] , 
        \Level1Out253[3] , \Level1Out253[2] , \Level1Out253[1] , 
        \Level1Out253[0] }), .Read1(\Level1Load252[0] ), .Read2(
        \Level1Load253[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_80_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load80[0] ), .Out({\Level4Out80[31] , \Level4Out80[30] , 
        \Level4Out80[29] , \Level4Out80[28] , \Level4Out80[27] , 
        \Level4Out80[26] , \Level4Out80[25] , \Level4Out80[24] , 
        \Level4Out80[23] , \Level4Out80[22] , \Level4Out80[21] , 
        \Level4Out80[20] , \Level4Out80[19] , \Level4Out80[18] , 
        \Level4Out80[17] , \Level4Out80[16] , \Level4Out80[15] , 
        \Level4Out80[14] , \Level4Out80[13] , \Level4Out80[12] , 
        \Level4Out80[11] , \Level4Out80[10] , \Level4Out80[9] , 
        \Level4Out80[8] , \Level4Out80[7] , \Level4Out80[6] , \Level4Out80[5] , 
        \Level4Out80[4] , \Level4Out80[3] , \Level4Out80[2] , \Level4Out80[1] , 
        \Level4Out80[0] }), .In1({\Level2Out80[31] , \Level2Out80[30] , 
        \Level2Out80[29] , \Level2Out80[28] , \Level2Out80[27] , 
        \Level2Out80[26] , \Level2Out80[25] , \Level2Out80[24] , 
        \Level2Out80[23] , \Level2Out80[22] , \Level2Out80[21] , 
        \Level2Out80[20] , \Level2Out80[19] , \Level2Out80[18] , 
        \Level2Out80[17] , \Level2Out80[16] , \Level2Out80[15] , 
        \Level2Out80[14] , \Level2Out80[13] , \Level2Out80[12] , 
        \Level2Out80[11] , \Level2Out80[10] , \Level2Out80[9] , 
        \Level2Out80[8] , \Level2Out80[7] , \Level2Out80[6] , \Level2Out80[5] , 
        \Level2Out80[4] , \Level2Out80[3] , \Level2Out80[2] , \Level2Out80[1] , 
        \Level2Out80[0] }), .In2({\Level2Out82[31] , \Level2Out82[30] , 
        \Level2Out82[29] , \Level2Out82[28] , \Level2Out82[27] , 
        \Level2Out82[26] , \Level2Out82[25] , \Level2Out82[24] , 
        \Level2Out82[23] , \Level2Out82[22] , \Level2Out82[21] , 
        \Level2Out82[20] , \Level2Out82[19] , \Level2Out82[18] , 
        \Level2Out82[17] , \Level2Out82[16] , \Level2Out82[15] , 
        \Level2Out82[14] , \Level2Out82[13] , \Level2Out82[12] , 
        \Level2Out82[11] , \Level2Out82[10] , \Level2Out82[9] , 
        \Level2Out82[8] , \Level2Out82[7] , \Level2Out82[6] , \Level2Out82[5] , 
        \Level2Out82[4] , \Level2Out82[3] , \Level2Out82[2] , \Level2Out82[1] , 
        \Level2Out82[0] }), .Read1(\Level2Load80[0] ), .Read2(
        \Level2Load82[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_108 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink108[31] , \ScanLink108[30] , 
        \ScanLink108[29] , \ScanLink108[28] , \ScanLink108[27] , 
        \ScanLink108[26] , \ScanLink108[25] , \ScanLink108[24] , 
        \ScanLink108[23] , \ScanLink108[22] , \ScanLink108[21] , 
        \ScanLink108[20] , \ScanLink108[19] , \ScanLink108[18] , 
        \ScanLink108[17] , \ScanLink108[16] , \ScanLink108[15] , 
        \ScanLink108[14] , \ScanLink108[13] , \ScanLink108[12] , 
        \ScanLink108[11] , \ScanLink108[10] , \ScanLink108[9] , 
        \ScanLink108[8] , \ScanLink108[7] , \ScanLink108[6] , \ScanLink108[5] , 
        \ScanLink108[4] , \ScanLink108[3] , \ScanLink108[2] , \ScanLink108[1] , 
        \ScanLink108[0] }), .ScanOut({\ScanLink109[31] , \ScanLink109[30] , 
        \ScanLink109[29] , \ScanLink109[28] , \ScanLink109[27] , 
        \ScanLink109[26] , \ScanLink109[25] , \ScanLink109[24] , 
        \ScanLink109[23] , \ScanLink109[22] , \ScanLink109[21] , 
        \ScanLink109[20] , \ScanLink109[19] , \ScanLink109[18] , 
        \ScanLink109[17] , \ScanLink109[16] , \ScanLink109[15] , 
        \ScanLink109[14] , \ScanLink109[13] , \ScanLink109[12] , 
        \ScanLink109[11] , \ScanLink109[10] , \ScanLink109[9] , 
        \ScanLink109[8] , \ScanLink109[7] , \ScanLink109[6] , \ScanLink109[5] , 
        \ScanLink109[4] , \ScanLink109[3] , \ScanLink109[2] , \ScanLink109[1] , 
        \ScanLink109[0] }), .ScanEnable(\ScanEnable[0] ), .Id(1'b0), .Load(
        \Level1Load108[0] ), .Out({\Level1Out108[31] , \Level1Out108[30] , 
        \Level1Out108[29] , \Level1Out108[28] , \Level1Out108[27] , 
        \Level1Out108[26] , \Level1Out108[25] , \Level1Out108[24] , 
        \Level1Out108[23] , \Level1Out108[22] , \Level1Out108[21] , 
        \Level1Out108[20] , \Level1Out108[19] , \Level1Out108[18] , 
        \Level1Out108[17] , \Level1Out108[16] , \Level1Out108[15] , 
        \Level1Out108[14] , \Level1Out108[13] , \Level1Out108[12] , 
        \Level1Out108[11] , \Level1Out108[10] , \Level1Out108[9] , 
        \Level1Out108[8] , \Level1Out108[7] , \Level1Out108[6] , 
        \Level1Out108[5] , \Level1Out108[4] , \Level1Out108[3] , 
        \Level1Out108[2] , \Level1Out108[1] , \Level1Out108[0] }) );
    Merge_Node_DWIDTH32 U_Merge_Node_152_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load152[0] ), .Out({\Level8Out152[31] , \Level8Out152[30] , 
        \Level8Out152[29] , \Level8Out152[28] , \Level8Out152[27] , 
        \Level8Out152[26] , \Level8Out152[25] , \Level8Out152[24] , 
        \Level8Out152[23] , \Level8Out152[22] , \Level8Out152[21] , 
        \Level8Out152[20] , \Level8Out152[19] , \Level8Out152[18] , 
        \Level8Out152[17] , \Level8Out152[16] , \Level8Out152[15] , 
        \Level8Out152[14] , \Level8Out152[13] , \Level8Out152[12] , 
        \Level8Out152[11] , \Level8Out152[10] , \Level8Out152[9] , 
        \Level8Out152[8] , \Level8Out152[7] , \Level8Out152[6] , 
        \Level8Out152[5] , \Level8Out152[4] , \Level8Out152[3] , 
        \Level8Out152[2] , \Level8Out152[1] , \Level8Out152[0] }), .In1({
        \Level4Out152[31] , \Level4Out152[30] , \Level4Out152[29] , 
        \Level4Out152[28] , \Level4Out152[27] , \Level4Out152[26] , 
        \Level4Out152[25] , \Level4Out152[24] , \Level4Out152[23] , 
        \Level4Out152[22] , \Level4Out152[21] , \Level4Out152[20] , 
        \Level4Out152[19] , \Level4Out152[18] , \Level4Out152[17] , 
        \Level4Out152[16] , \Level4Out152[15] , \Level4Out152[14] , 
        \Level4Out152[13] , \Level4Out152[12] , \Level4Out152[11] , 
        \Level4Out152[10] , \Level4Out152[9] , \Level4Out152[8] , 
        \Level4Out152[7] , \Level4Out152[6] , \Level4Out152[5] , 
        \Level4Out152[4] , \Level4Out152[3] , \Level4Out152[2] , 
        \Level4Out152[1] , \Level4Out152[0] }), .In2({\Level4Out156[31] , 
        \Level4Out156[30] , \Level4Out156[29] , \Level4Out156[28] , 
        \Level4Out156[27] , \Level4Out156[26] , \Level4Out156[25] , 
        \Level4Out156[24] , \Level4Out156[23] , \Level4Out156[22] , 
        \Level4Out156[21] , \Level4Out156[20] , \Level4Out156[19] , 
        \Level4Out156[18] , \Level4Out156[17] , \Level4Out156[16] , 
        \Level4Out156[15] , \Level4Out156[14] , \Level4Out156[13] , 
        \Level4Out156[12] , \Level4Out156[11] , \Level4Out156[10] , 
        \Level4Out156[9] , \Level4Out156[8] , \Level4Out156[7] , 
        \Level4Out156[6] , \Level4Out156[5] , \Level4Out156[4] , 
        \Level4Out156[3] , \Level4Out156[2] , \Level4Out156[1] , 
        \Level4Out156[0] }), .Read1(\Level4Load152[0] ), .Read2(
        \Level4Load156[0] ) );
endmodule

