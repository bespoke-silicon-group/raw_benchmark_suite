/*
 * $Header: /projects/raw/cvsroot/benchmark/include/common/main_trailer.v,v 1.2 1997/08/09 05:56:14 jbabb Exp $
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
