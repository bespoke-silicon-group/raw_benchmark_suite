
module NORMALIZE_SIZE8_DW01_dec_8_0 ( A, SUM );
input  [7:0] A;
output [7:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n11, n10;
    VMW_AO21 U3 ( .A(n5), .B(A[5]), .C(n6), .Z(SUM[5]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n7), .Z(SUM[1]) );
    VMW_OAI21 U6 ( .A(n10), .B(n11), .C(n5), .Z(SUM[4]) );
    VMW_NOR2 U14 ( .A(n5), .B(A[5]), .Z(n6) );
    VMW_INV U7 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO21 U8 ( .A(n9), .B(A[3]), .C(n10), .Z(SUM[3]) );
    VMW_NAND2 U13 ( .A(n10), .B(n11), .Z(n5) );
    VMW_NOR2 U9 ( .A(A[6]), .B(n13), .Z(n12) );
    VMW_NOR2 U12 ( .A(n9), .B(A[3]), .Z(n10) );
    VMW_XOR2 U15 ( .A(A[7]), .B(n12), .Z(SUM[7]) );
    VMW_INV U17 ( .A(A[2]), .Z(n8) );
    VMW_NOR2 U10 ( .A(A[0]), .B(A[1]), .Z(n7) );
    VMW_NAND2 U11 ( .A(n7), .B(n8), .Z(n9) );
    VMW_INV U19 ( .A(n6), .Z(n13) );
    VMW_OAI21 U4 ( .A(n7), .B(n8), .C(n9), .Z(SUM[2]) );
    VMW_INV U18 ( .A(A[4]), .Z(n11) );
    VMW_MUX2I U16 ( .A(n13), .B(n6), .S(A[6]), .Z(SUM[6]) );
endmodule


module NORMALIZE_SIZE8 ( a, b );
input  [8:0] a;
output [8:0] b;
    wire \b99[4] , n182, \b99[6] , n176, \b99[2] , n178, n181, n179, \b99[3] , 
        n177, \b99[7] , \b99[5] , \b99[8] , \b99[1] , n180;
    VMW_NOR4 U22 ( .A(a[3]), .B(a[4]), .C(n176), .D(n177), .Z(b[8]) );
    VMW_AO22 U26 ( .A(\b99[5] ), .B(n178), .C(a[4]), .D(n179), .Z(b[4]) );
    VMW_AO22 U28 ( .A(\b99[3] ), .B(n178), .C(a[2]), .D(n179), .Z(b[2]) );
    VMW_OR4 U33 ( .A(a[4]), .B(a[5]), .C(a[6]), .D(a[7]), .Z(n181) );
    VMW_OR4 U34 ( .A(a[0]), .B(a[1]), .C(a[2]), .D(a[3]), .Z(n182) );
    VMW_AO22 U27 ( .A(\b99[4] ), .B(n178), .C(a[3]), .D(n179), .Z(b[3]) );
    VMW_OAI21 U35 ( .A(n181), .B(n182), .C(a[8]), .Z(n179) );
    NORMALIZE_SIZE8_DW01_dec_8_0 sub_217 ( .A(a[7:0]), .SUM({\b99[8] , 
        \b99[7] , \b99[6] , \b99[5] , \b99[4] , \b99[3] , \b99[2] , \b99[1] })
         );
    VMW_AO22 U29 ( .A(\b99[2] ), .B(n178), .C(a[1]), .D(n179), .Z(b[1]) );
    VMW_OR4 U32 ( .A(n180), .B(a[0]), .C(a[1]), .D(a[2]), .Z(n177) );
    VMW_AO22 U23 ( .A(\b99[8] ), .B(n178), .C(a[7]), .D(n179), .Z(b[7]) );
    VMW_AO22 U24 ( .A(\b99[7] ), .B(n178), .C(a[6]), .D(n179), .Z(b[6]) );
    VMW_AO22 U25 ( .A(\b99[6] ), .B(n178), .C(a[5]), .D(n179), .Z(b[5]) );
    VMW_AO22 U30 ( .A(\b99[1] ), .B(n178), .C(a[0]), .D(n179), .Z(b[0]) );
    VMW_INV U37 ( .A(a[8]), .Z(n180) );
    VMW_INV U36 ( .A(n179), .Z(n178) );
    VMW_OR3 U31 ( .A(a[5]), .B(a[7]), .C(a[6]), .Z(n176) );
endmodule


module ADD_NN_SIZE8_DW01_add_8_0 ( A, B, CI, SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_AND2 U1 ( .A(A[0]), .B(B[0]), .Z(\carry[1] ) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_XOR2 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module ADD_NN_SIZE8 ( a, b, c );
input  [8:0] a;
input  [8:0] b;
output [8:0] c;
    wire \arr[8] , \arr[7] , \arr[3] , \arr[5] , \arr[6] , \arr[4] , \arr[1] , 
        \arr[0] , n56, \arr[2] , n58, n59, n57;
    NORMALIZE_SIZE8 norm ( .a({\arr[8] , \arr[7] , \arr[6] , \arr[5] , 
        \arr[4] , \arr[3] , \arr[2] , \arr[1] , \arr[0] }), .b(c) );
    VMW_INV U6 ( .A(n58), .Z(n57) );
    ADD_NN_SIZE8_DW01_add_8_0 add_234 ( .A(a[7:0]), .B(b[7:0]), .CI(n59), 
        .SUM({\arr[7] , \arr[6] , \arr[5] , \arr[4] , \arr[3] , \arr[2] , 
        \arr[1] , \arr[0] }) );
    VMW_PULLDOWN U2 ( .Z(n59) );
    VMW_INV U5 ( .A(\arr[7] ), .Z(n56) );
    VMW_AO21 U3 ( .A(n56), .B(b[7]), .C(n57), .Z(\arr[8] ) );
    VMW_OAI21 U4 ( .A(b[7]), .B(n56), .C(a[7]), .Z(n58) );
endmodule


module ADD_MINUS_1_SIZE8_DW01_dec_8_0 ( A, SUM );
input  [7:0] A;
output [7:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n11, n10;
    VMW_AO21 U3 ( .A(n5), .B(A[5]), .C(n6), .Z(SUM[5]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n7), .Z(SUM[1]) );
    VMW_OAI21 U6 ( .A(n10), .B(n11), .C(n5), .Z(SUM[4]) );
    VMW_NOR2 U14 ( .A(n5), .B(A[5]), .Z(n6) );
    VMW_INV U7 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO21 U8 ( .A(n9), .B(A[3]), .C(n10), .Z(SUM[3]) );
    VMW_NAND2 U13 ( .A(n10), .B(n11), .Z(n5) );
    VMW_NOR2 U9 ( .A(A[6]), .B(n13), .Z(n12) );
    VMW_NOR2 U12 ( .A(n9), .B(A[3]), .Z(n10) );
    VMW_XOR2 U15 ( .A(A[7]), .B(n12), .Z(SUM[7]) );
    VMW_INV U17 ( .A(A[2]), .Z(n8) );
    VMW_NOR2 U10 ( .A(A[0]), .B(A[1]), .Z(n7) );
    VMW_NAND2 U11 ( .A(n7), .B(n8), .Z(n9) );
    VMW_INV U19 ( .A(n6), .Z(n13) );
    VMW_OAI21 U4 ( .A(n7), .B(n8), .C(n9), .Z(SUM[2]) );
    VMW_INV U18 ( .A(A[4]), .Z(n11) );
    VMW_MUX2I U16 ( .A(n13), .B(n6), .S(A[6]), .Z(SUM[6]) );
endmodule


module ADD_MINUS_1_SIZE8 ( a, b );
input  [8:0] a;
output [8:0] b;
    wire n158, \c82[7] , \c82[3] , \c82[8] , \c82[1] , \c82[5] , n159, 
        \c82[4] , \c82[2] , \c82[6] ;
    VMW_NOR4 U20 ( .A(n158), .B(n159), .C(a[5]), .D(a[4]), .Z(b[8]) );
    VMW_OR2 U21 ( .A(\c82[8] ), .B(a[8]), .Z(b[7]) );
    VMW_OR2 U26 ( .A(\c82[3] ), .B(a[8]), .Z(b[2]) );
    VMW_OR2 U28 ( .A(\c82[1] ), .B(a[8]), .Z(b[0]) );
    VMW_OR2 U27 ( .A(\c82[2] ), .B(a[8]), .Z(b[1]) );
    ADD_MINUS_1_SIZE8_DW01_dec_8_0 sub_199 ( .A(a[7:0]), .SUM({\c82[8] , 
        \c82[7] , \c82[6] , \c82[5] , \c82[4] , \c82[3] , \c82[2] , \c82[1] })
         );
    VMW_OR2 U22 ( .A(\c82[7] ), .B(a[8]), .Z(b[6]) );
    VMW_OR3 U29 ( .A(a[8]), .B(a[7]), .C(a[6]), .Z(n159) );
    VMW_OR2 U23 ( .A(\c82[6] ), .B(a[8]), .Z(b[5]) );
    VMW_OR2 U24 ( .A(\c82[5] ), .B(a[8]), .Z(b[4]) );
    VMW_OR2 U25 ( .A(\c82[4] ), .B(a[8]), .Z(b[3]) );
    VMW_OR4 U30 ( .A(a[1]), .B(a[0]), .C(a[3]), .D(a[2]), .Z(n158) );
endmodule


module ADD_SIZE8 ( a, b, c );
input  [8:0] a;
input  [8:0] b;
output [8:0] c;
    wire \sum1[6] , n97, \sum2[5] , \sum2[8] , \sum1[2] , \sum2[1] , \sum1[0] , 
        \sum2[3] , n99, \sum1[4] , \sum2[7] , \sum3[8] , \sum3[7] , \sum3[3] , 
        n90, n98, \sum3[5] , n91, n96, \sum3[6] , \sum3[4] , \sum3[1] , 
        \sum3[0] , n94, \sum3[2] , n93, \sum1[5] , \sum1[1] , \sum2[6] , 
        \sum2[2] , n92, \sum1[8] , n89, n95, \sum1[7] , \sum1[3] , \sum2[4] , 
        \sum2[0] ;
    ADD_NN_SIZE8 add_nn ( .a(a), .b(b), .c({\sum1[8] , \sum1[7] , \sum1[6] , 
        \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }) );
    ADD_MINUS_1_SIZE8 am2 ( .a(b), .b({\sum3[8] , \sum3[7] , \sum3[6] , 
        \sum3[5] , \sum3[4] , \sum3[3] , \sum3[2] , \sum3[1] , \sum3[0] }) );
    VMW_AO21 U20 ( .A(\sum1[5] ), .B(n89), .C(n93), .Z(c[5]) );
    VMW_AO21 U21 ( .A(\sum1[4] ), .B(n89), .C(n94), .Z(c[4]) );
    VMW_NOR2 U26 ( .A(n89), .B(a[8]), .Z(n99) );
    VMW_AO22 U28 ( .A(\sum3[8] ), .B(a[8]), .C(\sum2[8] ), .D(n99), .Z(n90) );
    VMW_AO22 U33 ( .A(\sum3[3] ), .B(a[8]), .C(\sum2[3] ), .D(n99), .Z(n95) );
    VMW_AO22 U34 ( .A(\sum3[2] ), .B(a[8]), .C(\sum2[2] ), .D(n99), .Z(n96) );
    VMW_NOR2 U27 ( .A(a[8]), .B(b[8]), .Z(n89) );
    VMW_AO22 U35 ( .A(\sum3[1] ), .B(a[8]), .C(\sum2[1] ), .D(n99), .Z(n97) );
    VMW_AO22 U29 ( .A(\sum3[7] ), .B(a[8]), .C(\sum2[7] ), .D(n99), .Z(n91) );
    VMW_AO21 U17 ( .A(n89), .B(\sum1[8] ), .C(n90), .Z(c[8]) );
    VMW_AO21 U22 ( .A(\sum1[3] ), .B(n89), .C(n95), .Z(c[3]) );
    VMW_AO22 U32 ( .A(\sum3[4] ), .B(a[8]), .C(\sum2[4] ), .D(n99), .Z(n94) );
    VMW_AO22 U30 ( .A(\sum3[6] ), .B(a[8]), .C(\sum2[6] ), .D(n99), .Z(n92) );
    VMW_AO21 U18 ( .A(\sum1[7] ), .B(n89), .C(n91), .Z(c[7]) );
    VMW_AO21 U19 ( .A(\sum1[6] ), .B(n89), .C(n92), .Z(c[6]) );
    VMW_AO21 U25 ( .A(\sum1[0] ), .B(n89), .C(n98), .Z(c[0]) );
    VMW_AO22 U36 ( .A(\sum3[0] ), .B(a[8]), .C(\sum2[0] ), .D(n99), .Z(n98) );
    VMW_AO21 U23 ( .A(\sum1[2] ), .B(n89), .C(n96), .Z(c[2]) );
    VMW_AO21 U24 ( .A(\sum1[1] ), .B(n89), .C(n97), .Z(c[1]) );
    ADD_MINUS_1_SIZE8 am1 ( .a(a), .b({\sum2[8] , \sum2[7] , \sum2[6] , 
        \sum2[5] , \sum2[4] , \sum2[3] , \sum2[2] , \sum2[1] , \sum2[0] }) );
    VMW_AO22 U31 ( .A(\sum3[5] ), .B(a[8]), .C(\sum2[5] ), .D(n99), .Z(n93) );
endmodule


module NEGATE_SIZE8_DW01_sub_9_0 ( A, B, CI, DIFF, CO );
input  [8:0] A;
input  [8:0] B;
output [8:0] DIFF;
input  CI;
output CO;
    wire \carry[8] , \B_not[8] , \B_not[7] , \carry[4] , \B_not[3] , 
        \carry[6] , \B_not[5] , \carry[2] , \carry[7] , \B_not[4] , \carry[3] , 
        \B_not[6] , \carry[5] , \B_not[2] ;
    VMW_XNOR2 U3 ( .A(\carry[8] ), .B(\B_not[8] ), .Z(DIFF[8]) );
    VMW_XOR2 U5 ( .A(\carry[7] ), .B(\B_not[7] ), .Z(DIFF[7]) );
    VMW_AND2 U6 ( .A(\carry[6] ), .B(\B_not[6] ), .Z(\carry[7] ) );
    VMW_AND2 U14 ( .A(\carry[2] ), .B(\B_not[2] ), .Z(\carry[3] ) );
    VMW_INV U21 ( .A(B[7]), .Z(\B_not[7] ) );
    VMW_XOR2 U7 ( .A(\carry[6] ), .B(\B_not[6] ), .Z(DIFF[6]) );
    VMW_AND2 U8 ( .A(\carry[5] ), .B(\B_not[5] ), .Z(\carry[6] ) );
    VMW_XOR2 U13 ( .A(\carry[3] ), .B(\B_not[3] ), .Z(DIFF[3]) );
    VMW_XOR2 U9 ( .A(\carry[5] ), .B(\B_not[5] ), .Z(DIFF[5]) );
    VMW_AND2 U12 ( .A(\carry[3] ), .B(\B_not[3] ), .Z(\carry[4] ) );
    VMW_INV U20 ( .A(B[2]), .Z(\B_not[2] ) );
    VMW_XOR2 U15 ( .A(\carry[2] ), .B(\B_not[2] ), .Z(DIFF[2]) );
    VMW_INV U17 ( .A(B[4]), .Z(\B_not[4] ) );
    VMW_INV U22 ( .A(B[6]), .Z(\B_not[6] ) );
    VMW_AND2 U10 ( .A(\carry[4] ), .B(\B_not[4] ), .Z(\carry[5] ) );
    VMW_XOR2 U11 ( .A(\carry[4] ), .B(\B_not[4] ), .Z(DIFF[4]) );
    VMW_INV U19 ( .A(B[5]), .Z(\B_not[5] ) );
    VMW_INV U25 ( .A(B[1]), .Z(\carry[2] ) );
    VMW_AND2 U4 ( .A(\carry[7] ), .B(\B_not[7] ), .Z(\carry[8] ) );
    VMW_INV U18 ( .A(B[3]), .Z(\B_not[3] ) );
    VMW_INV U23 ( .A(B[0]), .Z(DIFF[0]) );
    VMW_INV U24 ( .A(B[8]), .Z(\B_not[8] ) );
    VMW_INV U16 ( .A(\carry[2] ), .Z(DIFF[1]) );
endmodule


module NEGATE_SIZE8 ( a, b );
input  [8:0] a;
output [8:0] b;
    wire n239, \c164[8] , \c164[1] , \ozzo[1] , \ozzo[0] , \c164[7] , 
        \c164[3] , n236, n237, n238, \c164[9] , n234, n235, \c164[6] , 
        \n135[28] , \c164[2] , \c164[4] ;
    VMW_PULLDOWN U51 ( .Z(n239) );
    VMW_PULLDOWN U52 ( .Z(\ozzo[1] ) );
    VMW_PULLUP U53 ( .Z(\ozzo[0] ) );
    VMW_AO22 U54 ( .A(\c164[9] ), .B(n234), .C(n235), .D(a[0]), .Z(b[8]) );
    VMW_AND2 U61 ( .A(\c164[2] ), .B(n234), .Z(b[1]) );
    NEGATE_SIZE8_DW01_sub_9_0 sub_276 ( .A({\ozzo[0] , \ozzo[1] , \ozzo[1] , 
        \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[1] , \ozzo[0] }), 
        .B(a), .CI(n239), .DIFF({\c164[9] , \c164[8] , \c164[7] , \c164[6] , 
        \n135[28] , \c164[4] , \c164[3] , \c164[2] , \c164[1] }) );
    VMW_NOR2 U66 ( .A(n236), .B(a[8]), .Z(n235) );
    VMW_INV U67 ( .A(n237), .Z(n236) );
    VMW_AND2 U55 ( .A(\c164[8] ), .B(n234), .Z(b[7]) );
    VMW_AND2 U57 ( .A(\c164[6] ), .B(n234), .Z(b[5]) );
    VMW_AND2 U60 ( .A(\c164[3] ), .B(n234), .Z(b[2]) );
    VMW_AND2 U58 ( .A(\n135[28] ), .B(n234), .Z(b[4]) );
    VMW_AND2 U59 ( .A(\c164[4] ), .B(n234), .Z(b[3]) );
    VMW_AO21 U62 ( .A(\c164[1] ), .B(n236), .C(a[8]), .Z(b[0]) );
    VMW_OR4 U65 ( .A(a[3]), .B(a[4]), .C(a[1]), .D(a[2]), .Z(n238) );
    VMW_NOR2 U64 ( .A(a[8]), .B(n237), .Z(n234) );
    VMW_AND2 U56 ( .A(\c164[7] ), .B(n234), .Z(b[6]) );
    VMW_NOR4 U63 ( .A(a[5]), .B(a[7]), .C(a[6]), .D(n238), .Z(n237) );
endmodule


module SHIFT_UP_SIZE8_s17 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[2] , Logic0, 
        \nb2[5] , \nb2[8] , \nb2[1] , \sum1[0] , \nb2[3] , \nb2[7] , \nb2[6] , 
        \sum1[1] , \nb2[2] , \sum1[7] , \sum1[3] , \nb2[4] , \nb2[0] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({\sum1[8] , 
        \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , \sum1[2] , 
        \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U10 ( .Z(Logic0) );
endmodule


module COMBINATIONAL_SIZE8_s17 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \b[2] , \t2[5] , \t1[6] , \b[0] , \b[4] , \t2[1] , \t1[2] , \t2[8] , 
        \b[5] , \b[6] , \a[3]1 , \t2[3] , \t1[0] , \a[8]1 , \a[2]1 , \t2[7] , 
        \t1[4] , \a[7]1 , \a[6]1 , \a[5]1 , \a[4]1 , \b[8] , \b[3] , \b[7] , 
        \t2[6] , \t1[5] , \t1[8] , \t2[2] , \t1[1] , \t2[0] , \t1[3] , \a[1]1 , 
        \b[1] , \t1[7] , \t2[4] , \a[0]1 ;
    assign \a[8]1  = a[8];
    assign \a[7]1  = a[7];
    assign \a[6]1  = a[6];
    assign \a[5]1  = a[5];
    assign \a[4]1  = a[4];
    assign \a[3]1  = a[3];
    assign \a[2]1  = a[2];
    assign \a[1]1  = a[1];
    assign \a[0]1  = a[0];
    assign \b[8]  = b[8];
    assign \b[7]  = b[7];
    assign \b[6]  = b[6];
    assign \b[5]  = b[5];
    assign \b[4]  = b[4];
    assign \b[3]  = b[3];
    assign \b[2]  = b[2];
    assign \b[1]  = b[1];
    assign \b[0]  = b[0];
    assign x[8] = \a[8]1 ;
    assign x[7] = \a[7]1 ;
    assign x[6] = \a[6]1 ;
    assign x[5] = \a[5]1 ;
    assign x[4] = \a[4]1 ;
    assign x[3] = \a[3]1 ;
    assign x[2] = \a[2]1 ;
    assign x[1] = \a[1]1 ;
    assign x[0] = \a[0]1 ;
    assign y[8] = \b[8] ;
    assign y[7] = \b[7] ;
    assign y[6] = \b[6] ;
    assign y[5] = \b[5] ;
    assign y[4] = \b[4] ;
    assign y[3] = \b[3] ;
    assign y[2] = \b[2] ;
    assign y[1] = \b[1] ;
    assign y[0] = \b[0] ;
    ADD_SIZE8 add2 ( .a({\a[8]1 , \a[7]1 , \a[6]1 , \a[5]1 , \a[4]1 , \a[3]1 , 
        \a[2]1 , \a[1]1 , \a[0]1 }), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , 
        \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    ADD_SIZE8 add1 ( .a({\a[8]1 , \a[7]1 , \a[6]1 , \a[5]1 , \a[4]1 , \a[3]1 , 
        \a[2]1 , \a[1]1 , \a[0]1 }), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    SHIFT_UP_SIZE8_s17 shift ( .a({\b[8] , \b[7] , \b[6] , \b[5] , \b[4] , 
        \b[3] , \b[2] , \b[1] , \b[0] }), .c({\t1[8] , \t1[7] , \t1[6] , 
        \t1[5] , \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s17 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s0 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \a[8] , \a[7] , \sum1[6] , \b1[5] , \nb2[5] , \a[3] , \nb2[8] , 
        \b1[8] , \b1[1] , \a[1] , \sum1[2] , \nb2[1] , \sum1[0] , \nb2[3] , 
        \b1[3] , \a[6] , \a[5] , \a[4] , \nb2[7] , \sum1[4] , \b1[7] , n166, 
        \a[2] , \a[0] , \sum1[5] , \nb2[6] , \sum1[1] , \b1[6] , \nb2[2] , 
        \sum1[8] , \b1[2] , Logic01, \b1[0] , \nb2[0] , \sum1[3] , \sum1[7] , 
        \nb2[4] , \b1[4] ;
    assign \a[8]  = a[8];
    assign \a[7]  = a[7];
    assign \a[6]  = a[6];
    assign \a[5]  = a[5];
    assign \a[4]  = a[4];
    assign \a[3]  = a[3];
    assign \a[2]  = a[2];
    assign \a[1]  = a[1];
    assign \a[0]  = a[0];
    assign c[8] = \a[8] ;
    assign c[7] = \a[7] ;
    assign c[6] = \a[6] ;
    assign c[5] = \a[5] ;
    assign c[4] = \a[4] ;
    assign c[3] = \a[3] ;
    assign c[2] = \a[2] ;
    assign c[1] = \a[1] ;
    assign c[0] = \a[0] ;
    VMW_AND2 U21 ( .A(\a[1] ), .B(n166), .Z(\b1[1] ) );
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01, Logic01, Logic01, Logic01}) );
    VMW_PULLDOWN U13 ( .Z(\b1[8] ) );
    VMW_PULLDOWN U14 ( .Z(Logic01) );
    VMW_AND2 U15 ( .A(\a[7] ), .B(n166), .Z(\b1[7] ) );
    VMW_AND2 U20 ( .A(\a[2] ), .B(n166), .Z(\b1[2] ) );
    NEGATE_SIZE8 negate ( .a({Logic01, Logic01, Logic01, Logic01, Logic01, 
        Logic01, Logic01, Logic01, Logic01}), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_AND2 U17 ( .A(\a[5] ), .B(n166), .Z(\b1[5] ) );
    VMW_AND2 U22 ( .A(\a[0] ), .B(n166), .Z(\b1[0] ) );
    VMW_AND2 U16 ( .A(\a[6] ), .B(n166), .Z(\b1[6] ) );
    VMW_AND2 U18 ( .A(\a[4] ), .B(n166), .Z(\b1[4] ) );
    VMW_AND2 U19 ( .A(\a[3] ), .B(n166), .Z(\b1[3] ) );
    VMW_INV U23 ( .A(\a[8] ), .Z(n166) );
endmodule


module COMBINATIONAL_SIZE8_s0 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s0 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s0 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s4 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , \nb2[6] , \sum1[1] , \b1[6] , 
        \nb2[2] , \b1[2] , n170, \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[2] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n170), .Z(\b1[5] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[3] ) );
    VMW_AND2 U20 ( .A(a[2]), .B(n170), .Z(\b1[6] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[1] ) );
    VMW_AND2 U22 ( .A(a[0]), .B(n170), .Z(\b1[4] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[8] ) );
    VMW_PULLDOWN U18 ( .Z(Logic0) );
    VMW_AND2 U19 ( .A(a[3]), .B(n170), .Z(\b1[7] ) );
    VMW_INV U23 ( .A(a[8]), .Z(n170) );
endmodule


module COMBINATIONAL_SIZE8_s4 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s4 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comright[6] , n438, \comleft[5] , n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s4 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s2 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , n168, \nb2[6] , \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[8] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n168), .Z(\b1[3] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[1] ) );
    VMW_AND2 U20 ( .A(a[2]), .B(n168), .Z(\b1[4] ) );
    VMW_AND2 U17 ( .A(a[5]), .B(n168), .Z(\b1[7] ) );
    VMW_AND2 U22 ( .A(a[0]), .B(n168), .Z(\b1[2] ) );
    VMW_PULLDOWN U16 ( .Z(Logic0) );
    VMW_AND2 U18 ( .A(a[4]), .B(n168), .Z(\b1[6] ) );
    VMW_AND2 U19 ( .A(a[3]), .B(n168), .Z(\b1[5] ) );
    VMW_INV U23 ( .A(a[8]), .Z(n168) );
endmodule


module COMBINATIONAL_SIZE8_s2 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s2 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s2_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s2 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s6 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , n172, \nb2[6] , \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n172), .Z(\b1[7] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(\b1[5] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[8] ) );
    VMW_AND2 U22 ( .A(a[0]), .B(n172), .Z(\b1[6] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U19 ( .Z(Logic0) );
    VMW_INV U23 ( .A(a[8]), .Z(n172) );
endmodule


module COMBINATIONAL_SIZE8_s6 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s6 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s6_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s6 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s1 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , n167, 
        \sum1[0] , \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , \nb2[6] , \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[8] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n167), .Z(\b1[2] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(Logic0) );
    VMW_AND2 U20 ( .A(a[2]), .B(n167), .Z(\b1[3] ) );
    VMW_AND2 U17 ( .A(a[5]), .B(n167), .Z(\b1[6] ) );
    VMW_AND2 U22 ( .A(a[0]), .B(n167), .Z(\b1[1] ) );
    VMW_AND2 U16 ( .A(a[6]), .B(n167), .Z(\b1[7] ) );
    VMW_AND2 U18 ( .A(a[4]), .B(n167), .Z(\b1[5] ) );
    VMW_AND2 U19 ( .A(a[3]), .B(n167), .Z(\b1[4] ) );
    VMW_INV U23 ( .A(a[8]), .Z(n167) );
endmodule


module COMBINATIONAL_SIZE8_s1 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s1 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[4] , \outleft[0] , \ScanReg[2] , 
        n467, n440, n475, n449, n452, \outleft[6] , \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s1 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s3 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , n169, \b1[7] , \nb2[6] , \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[2] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n169), .Z(\b1[4] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[8] ) );
    VMW_AND2 U20 ( .A(a[2]), .B(n169), .Z(\b1[5] ) );
    VMW_PULLDOWN U17 ( .Z(Logic0) );
    VMW_AND2 U22 ( .A(a[0]), .B(n169), .Z(\b1[3] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[1] ) );
    VMW_AND2 U18 ( .A(a[4]), .B(n169), .Z(\b1[7] ) );
    VMW_AND2 U19 ( .A(a[3]), .B(n169), .Z(\b1[6] ) );
    VMW_INV U23 ( .A(a[8]), .Z(n169) );
endmodule


module COMBINATIONAL_SIZE8_s3 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s3 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s3_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s3 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s5 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , \nb2[6] , n171, \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_AND2 U21 ( .A(a[1]), .B(n171), .Z(\b1[6] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_AND2 U20 ( .A(a[2]), .B(n171), .Z(\b1[7] ) );
    VMW_PULLDOWN U17 ( .Z(\b1[8] ) );
    VMW_AND2 U22 ( .A(a[0]), .B(n171), .Z(\b1[5] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[3] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[1] ) );
    VMW_PULLDOWN U19 ( .Z(Logic0) );
    VMW_INV U23 ( .A(a[8]), .Z(n171) );
endmodule


module COMBINATIONAL_SIZE8_s5 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s5 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s5_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[0] , \ScanReg[2] , n467, n440, 
        n475, n449, n452, \outleft[6] , \outleft[4] , \ScanReg[4] , 
        \ScanReg[6] , n469, \outleft[2] , n472, n455, n429, n460, n447, n432, 
        \outleft[3] , \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , 
        n462, n445, n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, 
        \ScanReg[3] , n477, n450, n436, n443, \comleft[7] , n464, 
        \comright[4] , \comleft[3] , \comright[0] , n476, n451, \comleft[1] , 
        \comright[2] , n471, n456, \comleft[8] , \comleft[5] , \comright[6] , 
        n438, n463, n444, n478, n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s5 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module SHIFT_UP_SIZE8_s7 ( a, c );
input  [8:0] a;
output [8:0] c;
    wire \sum1[8] , \sum1[6] , \b1[5] , \sum1[5] , \sum1[4] , \sum1[2] , 
        Logic0, \nb2[5] , \nb2[8] , \nb2[1] , \b1[8] , \b1[1] , \sum1[0] , 
        \nb2[3] , \b1[3] , \nb2[7] , \b1[7] , n173, \nb2[6] , \sum1[1] , 
        \b1[6] , \nb2[2] , \b1[2] , \sum1[7] , \sum1[3] , \b1[0] , \nb2[4] , 
        \nb2[0] , \b1[4] ;
    ADD_SIZE8 add2 ( .a({\sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , 
        \sum1[3] , \sum1[2] , \sum1[1] , \sum1[0] }), .b({Logic0, Logic0, 
        Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, Logic0}), .c(c) );
    VMW_PULLDOWN U13 ( .Z(\b1[4] ) );
    VMW_PULLDOWN U14 ( .Z(\b1[0] ) );
    VMW_PULLDOWN U21 ( .Z(\b1[5] ) );
    NEGATE_SIZE8 negate ( .a({Logic0, Logic0, Logic0, Logic0, Logic0, Logic0, 
        Logic0, Logic0, Logic0}), .b({\nb2[8] , \nb2[7] , \nb2[6] , \nb2[5] , 
        \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }) );
    ADD_SIZE8 add1 ( .a({\b1[8] , \b1[7] , \b1[6] , \b1[5] , \b1[4] , \b1[3] , 
        \b1[2] , \b1[1] , \b1[0] }), .b({\nb2[8] , \nb2[7] , \nb2[6] , 
        \nb2[5] , \nb2[4] , \nb2[3] , \nb2[2] , \nb2[1] , \nb2[0] }), .c({
        \sum1[8] , \sum1[7] , \sum1[6] , \sum1[5] , \sum1[4] , \sum1[3] , 
        \sum1[2] , \sum1[1] , \sum1[0] }) );
    VMW_PULLDOWN U15 ( .Z(\b1[2] ) );
    VMW_PULLDOWN U20 ( .Z(Logic0) );
    VMW_PULLDOWN U17 ( .Z(\b1[3] ) );
    VMW_NOR2 U22 ( .A(n173), .B(a[8]), .Z(\b1[7] ) );
    VMW_PULLDOWN U16 ( .Z(\b1[6] ) );
    VMW_PULLDOWN U18 ( .Z(\b1[8] ) );
    VMW_PULLDOWN U19 ( .Z(\b1[1] ) );
    VMW_INV U23 ( .A(a[0]), .Z(n173) );
endmodule


module COMBINATIONAL_SIZE8_s7 ( a, b, x, y );
input  [8:0] a;
output [8:0] y;
input  [8:0] b;
output [8:0] x;
    wire \t2[5] , \t1[6] , \t4[2] , \t2[1] , \t1[2] , \t2[8] , \t4[6] , 
        \t4[4] , \t2[3] , \t1[0] , \t2[7] , \t4[0] , \t1[4] , \t3[3] , n154, 
        \t3[7] , \t3[5] , \t3[1] , n153, \t3[4] , \t3[0] , \t3[6] , \t3[2] , 
        \t2[6] , \t4[1] , \t1[5] , \t4[5] , \t1[8] , \t2[2] , \t2[0] , \t1[3] , 
        \t1[1] , \t2[4] , \t4[7] , \t4[3] , \t1[7] ;
    ADD_SIZE8 add2 ( .a(a), .b({\t2[8] , \t2[7] , \t2[6] , \t2[5] , \t2[4] , 
        \t2[3] , \t2[2] , \t2[1] , \t2[0] }), .c({y[8], \t4[7] , \t4[6] , 
        \t4[5] , \t4[4] , \t4[3] , \t4[2] , \t4[1] , \t4[0] }) );
    VMW_AND2 U21 ( .A(\t3[6] ), .B(n153), .Z(x[6]) );
    VMW_AND2 U26 ( .A(\t3[1] ), .B(n153), .Z(x[1]) );
    VMW_AND2 U28 ( .A(\t4[7] ), .B(n154), .Z(y[7]) );
    VMW_AND2 U33 ( .A(\t4[2] ), .B(n154), .Z(y[2]) );
    VMW_AND2 U34 ( .A(\t4[1] ), .B(n154), .Z(y[1]) );
    ADD_SIZE8 add1 ( .a(a), .b({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .c({x[8], \t3[7] , \t3[6] , 
        \t3[5] , \t3[4] , \t3[3] , \t3[2] , \t3[1] , \t3[0] }) );
    VMW_AND2 U20 ( .A(\t3[7] ), .B(n153), .Z(x[7]) );
    VMW_AND2 U27 ( .A(\t3[0] ), .B(n153), .Z(x[0]) );
    VMW_AND2 U35 ( .A(\t4[0] ), .B(n154), .Z(y[0]) );
    VMW_AND2 U22 ( .A(\t3[5] ), .B(n153), .Z(x[5]) );
    VMW_AND2 U29 ( .A(\t4[6] ), .B(n154), .Z(y[6]) );
    VMW_AND2 U32 ( .A(\t4[3] ), .B(n154), .Z(y[3]) );
    VMW_AND2 U30 ( .A(\t4[5] ), .B(n154), .Z(y[5]) );
    VMW_INV U37 ( .A(x[8]), .Z(n153) );
    SHIFT_UP_SIZE8_s7 shift ( .a(b), .c({\t1[8] , \t1[7] , \t1[6] , \t1[5] , 
        \t1[4] , \t1[3] , \t1[2] , \t1[1] , \t1[0] }) );
    VMW_AND2 U25 ( .A(\t3[2] ), .B(n153), .Z(x[2]) );
    VMW_INV U36 ( .A(y[8]), .Z(n154) );
    NEGATE_SIZE8 neg ( .a({\t1[8] , \t1[7] , \t1[6] , \t1[5] , \t1[4] , 
        \t1[3] , \t1[2] , \t1[1] , \t1[0] }), .b({\t2[8] , \t2[7] , \t2[6] , 
        \t2[5] , \t2[4] , \t2[3] , \t2[2] , \t2[1] , \t2[0] }) );
    VMW_AND2 U23 ( .A(\t3[4] ), .B(n153), .Z(x[4]) );
    VMW_AND2 U24 ( .A(\t3[3] ), .B(n153), .Z(x[3]) );
    VMW_AND2 U31 ( .A(\t4[4] ), .B(n154), .Z(y[4]) );
endmodule


module FFT_Node_SIZE8_IDWIDTH1_s7_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, Idl, Idr, Ids, Enable, inleft, 
    inright, outleft, outright );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Idl;
input  [0:0] Ids;
output [8:0] outleft;
input  [7:0] ScanIn;
input  [0:0] Idr;
input  [8:0] inleft;
input  [8:0] inright;
output [7:0] ScanOut;
output [8:0] outright;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \outleft[7] , n448, n468, \comright[7] , \comleft[4] , n473, n454, 
        n433, \comleft[0] , \comright[3] , n461, n446, \comright[8] , n466, 
        n441, \comright[1] , \comleft[2] , n434, \comleft[6] , n474, 
        \comright[5] , n453, n435, \outleft[6] , \outleft[4] , \outleft[0] , 
        \ScanReg[2] , n467, n440, n475, n449, n452, \ScanReg[4] , \ScanReg[6] , 
        n469, \outleft[2] , n472, n455, n429, n460, n447, n432, \outleft[3] , 
        \ScanReg[5] , n470, n439, n457, n430, n458, \outleft[5] , n462, n445, 
        n465, n442, n459, \outleft[1] , \ScanReg[7] , n437, \ScanReg[3] , n477, 
        n450, n436, n443, \comleft[7] , n464, \comright[4] , \comleft[3] , 
        \comright[0] , n476, n451, \comleft[1] , \comright[2] , n471, n456, 
        \comleft[8] , \comleft[5] , \comright[6] , n438, n463, n444, n478, 
        n431;
    assign ScanOut[7] = \outleft[7] ;
    assign ScanOut[6] = \outleft[6] ;
    assign ScanOut[5] = \outleft[5] ;
    assign ScanOut[4] = \outleft[4] ;
    assign ScanOut[3] = \outleft[3] ;
    assign ScanOut[2] = \outleft[2] ;
    assign ScanOut[1] = \outleft[1] ;
    assign ScanOut[0] = \outleft[0] ;
    assign outleft[7] = \outleft[7] ;
    assign outleft[6] = \outleft[6] ;
    assign outleft[5] = \outleft[5] ;
    assign outleft[4] = \outleft[4] ;
    assign outleft[3] = \outleft[3] ;
    assign outleft[2] = \outleft[2] ;
    assign outleft[1] = \outleft[1] ;
    assign outleft[0] = \outleft[0] ;
    VMW_AO22 U54 ( .A(ScanIn[3]), .B(n429), .C(\ScanReg[3] ), .D(n430), .Z(
        n477) );
    VMW_AO21 U73 ( .A(\outleft[5] ), .B(n431), .C(n446), .Z(n458) );
    VMW_AO21 U68 ( .A(\outleft[0] ), .B(n431), .C(n441), .Z(n463) );
    VMW_AO22 U96 ( .A(outright[4]), .B(n454), .C(\comleft[4] ), .D(n452), .Z(
        n445) );
    VMW_FD \outright_reg[0]  ( .D(n472), .CP(Clk), .Q(outright[0]) );
    VMW_FD \outleft_reg[4]  ( .D(n459), .CP(Clk), .Q(\outleft[4] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(n475), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_AO22 U53 ( .A(ScanIn[2]), .B(n429), .C(\ScanReg[2] ), .D(n430), .Z(
        n478) );
    VMW_AO21 U61 ( .A(outright[2]), .B(n431), .C(n434), .Z(n470) );
    VMW_AO22 U84 ( .A(\ScanReg[7] ), .B(n454), .C(\comright[7] ), .D(n452), 
        .Z(n439) );
    VMW_FD \outleft_reg[0]  ( .D(n463), .CP(Clk), .Q(\outleft[0] ) );
    VMW_FD \outright_reg[4]  ( .D(n468), .CP(Clk), .Q(outright[4]) );
    VMW_AO21 U66 ( .A(outright[7]), .B(n431), .C(n439), .Z(n465) );
    VMW_INV U101 ( .A(ScanEnable), .Z(n453) );
    VMW_AO22 U83 ( .A(ScanIn[1]), .B(n454), .C(\comright[8] ), .D(n452), .Z(
        n440) );
    VMW_AO22 U91 ( .A(outleft[8]), .B(n454), .C(\comright[0] ), .D(n452), .Z(
        n432) );
    VMW_AO22 U98 ( .A(outright[2]), .B(n454), .C(\comleft[2] ), .D(n452), .Z(
        n443) );
    VMW_FD \outleft_reg[2]  ( .D(n461), .CP(Clk), .Q(\outleft[2] ) );
    VMW_FD \outright_reg[6]  ( .D(n466), .CP(Clk), .Q(outright[6]) );
    VMW_FD \ScanReg_reg[3]  ( .D(n477), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_FD \outleft_reg[6]  ( .D(n457), .CP(Clk), .Q(\outleft[6] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(n473), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_AO21 U74 ( .A(\outleft[6] ), .B(n431), .C(n447), .Z(n457) );
    VMW_AO22 U99 ( .A(outright[1]), .B(n454), .C(\comleft[1] ), .D(n452), .Z(
        n442) );
    VMW_FD \outright_reg[2]  ( .D(n470), .CP(Clk), .Q(outright[2]) );
    VMW_AO22 U55 ( .A(ScanIn[4]), .B(n429), .C(\ScanReg[4] ), .D(n430), .Z(
        n476) );
    VMW_AO21 U67 ( .A(outright[8]), .B(n431), .C(n440), .Z(n464) );
    VMW_NOR2 U82 ( .A(n453), .B(Reset), .Z(n429) );
    VMW_AO21 U69 ( .A(\outleft[1] ), .B(n431), .C(n442), .Z(n462) );
    VMW_AO21 U75 ( .A(\outleft[7] ), .B(n431), .C(n448), .Z(n456) );
    VMW_AO22 U90 ( .A(outright[8]), .B(n454), .C(\comright[1] ), .D(n452), .Z(
        n433) );
    VMW_AO21 U72 ( .A(\outleft[4] ), .B(n431), .C(n445), .Z(n459) );
    VMW_AO22 U97 ( .A(outright[3]), .B(n454), .C(\comleft[3] ), .D(n452), .Z(
        n444) );
    VMW_AO21 U60 ( .A(outright[1]), .B(n431), .C(n433), .Z(n471) );
    VMW_AO22 U85 ( .A(\ScanReg[6] ), .B(n454), .C(\comright[6] ), .D(n452), 
        .Z(n438) );
    VMW_AO22 U100 ( .A(outright[0]), .B(n454), .C(\comleft[0] ), .D(n452), .Z(
        n441) );
    COMBINATIONAL_SIZE8_s7 com ( .a(inleft), .b(inright), .x({\comleft[8] , 
        \comleft[7] , \comleft[6] , \comleft[5] , \comleft[4] , \comleft[3] , 
        \comleft[2] , \comleft[1] , \comleft[0] }), .y({\comright[8] , 
        \comright[7] , \comright[6] , \comright[5] , \comright[4] , 
        \comright[3] , \comright[2] , \comright[1] , \comright[0] }) );
    VMW_AO22 U57 ( .A(ScanIn[6]), .B(n429), .C(\ScanReg[6] ), .D(n430), .Z(
        n474) );
    VMW_AO21 U62 ( .A(outright[3]), .B(n431), .C(n435), .Z(n469) );
    VMW_AO21 U70 ( .A(\outleft[2] ), .B(n431), .C(n443), .Z(n461) );
    VMW_AND2 U79 ( .A(n453), .B(n451), .Z(n452) );
    VMW_AO22 U95 ( .A(outright[5]), .B(n454), .C(\comleft[5] ), .D(n452), .Z(
        n446) );
    VMW_AO22 U87 ( .A(\ScanReg[4] ), .B(n454), .C(\comright[4] ), .D(n452), 
        .Z(n436) );
    VMW_AO21 U65 ( .A(outright[6]), .B(n431), .C(n438), .Z(n466) );
    VMW_INV U102 ( .A(n450), .Z(n430) );
    VMW_AO22 U56 ( .A(ScanIn[5]), .B(n429), .C(\ScanReg[5] ), .D(n430), .Z(
        n475) );
    VMW_AO22 U58 ( .A(ScanIn[7]), .B(n429), .C(\ScanReg[7] ), .D(n430), .Z(
        n473) );
    VMW_AO21 U59 ( .A(outright[0]), .B(n431), .C(n432), .Z(n472) );
    VMW_AND2 U80 ( .A(n451), .B(ScanEnable), .Z(n454) );
    VMW_OR2 U77 ( .A(ScanEnable), .B(Reset), .Z(n450) );
    VMW_AO22 U89 ( .A(\ScanReg[2] ), .B(n454), .C(\comright[2] ), .D(n452), 
        .Z(n434) );
    VMW_AO22 U92 ( .A(ScanIn[0]), .B(n454), .C(\comleft[8] ), .D(n452), .Z(
        n449) );
    VMW_FD \outleft_reg[7]  ( .D(n456), .CP(Clk), .Q(\outleft[7] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(n474), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_AO21 U64 ( .A(outright[5]), .B(n431), .C(n437), .Z(n467) );
    VMW_NOR2 U81 ( .A(Enable), .B(n450), .Z(n431) );
    VMW_AO21 U76 ( .A(outleft[8]), .B(n431), .C(n449), .Z(n455) );
    VMW_FD \outright_reg[3]  ( .D(n469), .CP(Clk), .Q(outright[3]) );
    VMW_AO22 U88 ( .A(\ScanReg[3] ), .B(n454), .C(\comright[3] ), .D(n452), 
        .Z(n435) );
    VMW_AO22 U93 ( .A(outright[7]), .B(n454), .C(\comleft[7] ), .D(n452), .Z(
        n448) );
    VMW_FD \ScanReg_reg[2]  ( .D(n478), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_FD \outleft_reg[3]  ( .D(n460), .CP(Clk), .Q(\outleft[3] ) );
    VMW_AO22 U94 ( .A(outright[6]), .B(n454), .C(\comleft[6] ), .D(n452), .Z(
        n447) );
    VMW_FD \outleft_reg[8]  ( .D(n455), .CP(Clk), .Q(outleft[8]) );
    VMW_FD \outright_reg[7]  ( .D(n465), .CP(Clk), .Q(outright[7]) );
    VMW_FD \outright_reg[5]  ( .D(n467), .CP(Clk), .Q(outright[5]) );
    VMW_FD \outleft_reg[1]  ( .D(n462), .CP(Clk), .Q(\outleft[1] ) );
    VMW_AO21 U63 ( .A(outright[4]), .B(n431), .C(n436), .Z(n468) );
    VMW_AO21 U71 ( .A(\outleft[3] ), .B(n431), .C(n444), .Z(n460) );
    VMW_NOR2 U78 ( .A(Reset), .B(n431), .Z(n451) );
    VMW_AO22 U86 ( .A(\ScanReg[5] ), .B(n454), .C(\comright[5] ), .D(n452), 
        .Z(n437) );
    VMW_FD \outright_reg[1]  ( .D(n471), .CP(Clk), .Q(outright[1]) );
    VMW_FD \outleft_reg[5]  ( .D(n458), .CP(Clk), .Q(\outleft[5] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(n476), .CP(Clk), .Q(\ScanReg[4] ) );
    VMW_FD \outright_reg[8]  ( .D(n464), .CP(Clk), .Q(outright[8]) );
endmodule


module FFT_Control_SIZE8_IDWIDTH1_SCAN1_DW01_dec_32_0 ( A, SUM );
input  [31:0] A;
output [31:0] SUM;
    wire n20, n15, n32, n29, n9, n47, n7, n12, n40, n35, n27, n49, n13, n34, 
        n41, n6, n26, n48, n21, n8, n46, n28, n33, n14, n38, n23, n16, n31, 
        n43, n44, n36, n11, n24, n18, n10, n37, n42, n5, n19, n25, n22, n39, 
        n45, n17, n30;
    VMW_INV U3 ( .A(A[0]), .Z(SUM[0]) );
    VMW_OAI21 U5 ( .A(n8), .B(n9), .C(n10), .Z(SUM[20]) );
    VMW_OAI21 U6 ( .A(n11), .B(n12), .C(n13), .Z(SUM[2]) );
    VMW_AO21 U14 ( .A(n25), .B(A[17]), .C(n14), .Z(SUM[17]) );
    VMW_AO21 U21 ( .A(n33), .B(A[29]), .C(n34), .Z(SUM[29]) );
    VMW_NOR2 U54 ( .A(n10), .B(A[21]), .Z(n41) );
    VMW_INV U73 ( .A(A[4]), .Z(n35) );
    VMW_INV U68 ( .A(A[2]), .Z(n12) );
    VMW_AO21 U28 ( .A(n36), .B(A[5]), .C(n43), .Z(SUM[5]) );
    VMW_NOR2 U33 ( .A(A[30]), .B(n49), .Z(n48) );
    VMW_OAI21 U7 ( .A(n14), .B(n15), .C(n16), .Z(SUM[18]) );
    VMW_AO21 U8 ( .A(n17), .B(A[25]), .C(n18), .Z(SUM[25]) );
    VMW_AO21 U13 ( .A(n13), .B(A[3]), .C(n24), .Z(SUM[3]) );
    VMW_NOR2 U34 ( .A(A[1]), .B(A[0]), .Z(n11) );
    VMW_NAND2 U41 ( .A(n39), .B(n46), .Z(n30) );
    VMW_NOR2 U46 ( .A(n7), .B(A[13]), .Z(n22) );
    VMW_NAND2 U61 ( .A(n47), .B(n45), .Z(n33) );
    VMW_INV U66 ( .A(A[12]), .Z(n6) );
    VMW_OAI21 U26 ( .A(n41), .B(n42), .C(n28), .Z(SUM[22]) );
    VMW_NOR2 U48 ( .A(n19), .B(A[15]), .Z(n20) );
    VMW_AO21 U9 ( .A(n19), .B(A[15]), .C(n20), .Z(SUM[15]) );
    VMW_AO21 U12 ( .A(A[0]), .B(A[1]), .C(n11), .Z(SUM[1]) );
    VMW_NAND2 U35 ( .A(n11), .B(n12), .Z(n13) );
    VMW_NAND2 U53 ( .A(n9), .B(n8), .Z(n10) );
    VMW_INV U74 ( .A(A[16]), .Z(n37) );
    VMW_AO21 U27 ( .A(n10), .B(A[21]), .C(n41), .Z(SUM[21]) );
    VMW_NOR2 U40 ( .A(A[7]), .B(n38), .Z(n39) );
    VMW_NOR2 U52 ( .A(n16), .B(A[19]), .Z(n8) );
    VMW_INV U67 ( .A(A[20]), .Z(n9) );
    VMW_INV U75 ( .A(A[10]), .Z(n40) );
    VMW_OAI21 U20 ( .A(n29), .B(n32), .C(n17), .Z(SUM[24]) );
    VMW_NAND2 U49 ( .A(n37), .B(n20), .Z(n25) );
    VMW_INV U69 ( .A(A[18]), .Z(n15) );
    VMW_OAI21 U29 ( .A(n43), .B(n44), .C(n38), .Z(SUM[6]) );
    VMW_NAND2 U47 ( .A(n23), .B(n22), .Z(n19) );
    VMW_NAND2 U55 ( .A(n42), .B(n41), .Z(n28) );
    VMW_INV U72 ( .A(A[24]), .Z(n32) );
    VMW_NOR2 U60 ( .A(n27), .B(A[27]), .Z(n45) );
    VMW_OAI21 U15 ( .A(n18), .B(n26), .C(n27), .Z(SUM[26]) );
    VMW_AO21 U17 ( .A(n28), .B(A[23]), .C(n29), .Z(SUM[23]) );
    VMW_OAI21 U22 ( .A(n24), .B(n35), .C(n36), .Z(SUM[4]) );
    VMW_OAI21 U32 ( .A(n45), .B(n47), .C(n33), .Z(SUM[28]) );
    VMW_NAND2 U39 ( .A(n43), .B(n44), .Z(n38) );
    VMW_NAND2 U57 ( .A(n32), .B(n29), .Z(n17) );
    VMW_INV U70 ( .A(A[14]), .Z(n23) );
    VMW_AO21 U30 ( .A(n27), .B(A[27]), .C(n45), .Z(SUM[27]) );
    VMW_INV U79 ( .A(A[28]), .Z(n47) );
    VMW_AO21 U10 ( .A(n21), .B(A[11]), .C(n5), .Z(SUM[11]) );
    VMW_NOR2 U42 ( .A(n30), .B(A[9]), .Z(n31) );
    VMW_NAND2 U45 ( .A(n6), .B(n5), .Z(n7) );
    VMW_OR2 U62 ( .A(n33), .B(A[29]), .Z(n49) );
    VMW_INV U65 ( .A(n49), .Z(n34) );
    VMW_OAI21 U11 ( .A(n22), .B(n23), .C(n19), .Z(SUM[14]) );
    VMW_AO21 U19 ( .A(n30), .B(A[9]), .C(n31), .Z(SUM[9]) );
    VMW_OAI21 U25 ( .A(n31), .B(n40), .C(n21), .Z(SUM[10]) );
    VMW_NAND2 U37 ( .A(n24), .B(n35), .Z(n36) );
    VMW_NAND2 U59 ( .A(n26), .B(n18), .Z(n27) );
    VMW_NOR2 U50 ( .A(n25), .B(A[17]), .Z(n14) );
    VMW_INV U77 ( .A(A[6]), .Z(n44) );
    VMW_NOR2 U58 ( .A(n17), .B(A[25]), .Z(n18) );
    VMW_NOR2 U36 ( .A(n13), .B(A[3]), .Z(n24) );
    VMW_OAI21 U4 ( .A(n5), .B(n6), .C(n7), .Z(SUM[12]) );
    VMW_AO21 U18 ( .A(n7), .B(A[13]), .C(n22), .Z(SUM[13]) );
    VMW_NAND2 U43 ( .A(n40), .B(n31), .Z(n21) );
    VMW_MUX2I U64 ( .A(n49), .B(n34), .S(A[30]), .Z(SUM[30]) );
    VMW_NAND2 U51 ( .A(n15), .B(n14), .Z(n16) );
    VMW_INV U76 ( .A(A[22]), .Z(n42) );
    VMW_OAI21 U23 ( .A(n20), .B(n37), .C(n25), .Z(SUM[16]) );
    VMW_AO21 U24 ( .A(n38), .B(A[7]), .C(n39), .Z(SUM[7]) );
    VMW_NOR2 U38 ( .A(n36), .B(A[5]), .Z(n43) );
    VMW_NOR2 U44 ( .A(n21), .B(A[11]), .Z(n5) );
    VMW_NOR2 U56 ( .A(n28), .B(A[23]), .Z(n29) );
    VMW_INV U71 ( .A(A[26]), .Z(n26) );
    VMW_XOR2 U63 ( .A(A[31]), .B(n48), .Z(SUM[31]) );
    VMW_AO21 U16 ( .A(n16), .B(A[19]), .C(n8), .Z(SUM[19]) );
    VMW_OAI21 U31 ( .A(n39), .B(n46), .C(n30), .Z(SUM[8]) );
    VMW_INV U78 ( .A(A[8]), .Z(n46) );
endmodule


module FFT_Control_SIZE8_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, 
    DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] ScanIn;
output [7:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire \DataIn[4] , n317, \count241[28] , n330, \count[17] , \count[24] , 
        \count[2] , \DataIn[0] , n362, \count241[12] , \count241[21] , n345, 
        n370, n339, \count[20] , \count[13] , \count[6] , n357, \count241[16] , 
        \count241[25] , n295, n305, n322, \DataIn[6] , \DataIn[2] , n302, n292, 
        \count[29] , \count[30] , n325, \count241[14] , \count241[27] , 
        \count[18] , n350, \n239[1] , n289, \count[11] , \count[4] , 
        \count[22] , n319, n342, \count241[10] , \count241[23] , \count[9] , 
        n365, n359, \count[15] , \count[0] , \count[26] , \count241[19] , n310, 
        n337, \count241[1] , n351, n318, \ScanReg[2] , n293, n324, n303, 
        \count241[8] , n336, n311, \count241[5] , n358, n364, n343, 
        \ScanReg[6] , \ScanReg[4] , \count241[7] , n363, n344, n316, n294, 
        n331, n323, n304, \ScanReg[0] , n356, \count241[3] , n338, n333, n314, 
        n361, n346, \ScanReg[1] , \count241[2] , n328, \ScanReg[5] , n354, 
        n368, \count241[6] , n296, n321, n306, \ScanReg[7] , n291, n301, 
        \count241[4] , n326, n353, n348, \count241[0] , n366, n308, n298, n341, 
        \DataIn[7] , \count241[9] , n334, n313, \ScanReg[3] , \count241[11] , 
        \count241[22] , \count[8] , n352, \count[14] , \count[1] , n349, 
        \count[27] , \DataIn[3] , n300, n290, \count241[18] , n312, n327, 
        \count241[15] , \count241[26] , n335, \count[19] , n340, n367, 
        \DataIn[1] , \count[10] , \count[5] , \count[23] , n299, n309, n360, 
        n347, n329, \count[12] , \count[7] , \count[21] , \count241[17] , 
        \count241[24] , \DataIn[5] , n332, \count[28] , n315, \count[31] , 
        n369, \count241[29] , n320, \count241[30] , n297, n307, \count[16] , 
        \count[3] , \count[25] , n355, \count241[20] , \count241[13] ;
    tri \DataOut[27]1 , \DataOut[14]1 , \DataOut[26]1 , \DataOut[15]1 , 
        \DataOut[31] , \DataOut[18]1 , \DataOut[0]1 , \DataOut[19]1 , 
        \DataOut[1]1 , \DataOut[23]1 , \DataOut[22]1 , \DataOut[11]1 , 
        \DataOut[10]1 , \DataOut[9]1 , \DataOut[8]1 , \DataOut[5]1 , 
        \DataOut[4]1 , \DataOut[21]1 , \DataOut[20]1 , \DataOut[13]1 , 
        \DataOut[12]1 , \DataOut[7]1 , \DataOut[6]1 , \DataOut[25]1 , 
        \DataOut[16]1 , \DataOut[24]1 , \DataOut[17]1 , \DataOut[29]1 , 
        \DataOut[30]1 , \DataOut[2]1 , \DataOut[28]1 , \DataOut[3]1 ;
    assign \DataIn[7]  = DataIn[7];
    assign \DataIn[6]  = DataIn[6];
    assign \DataIn[5]  = DataIn[5];
    assign \DataIn[4]  = DataIn[4];
    assign \DataIn[3]  = DataIn[3];
    assign \DataIn[2]  = DataIn[2];
    assign \DataIn[1]  = DataIn[1];
    assign \DataIn[0]  = DataIn[0];
    assign DataOut[31] = \DataOut[31] ;
    assign DataOut[30] = \DataOut[30]1 ;
    assign DataOut[29] = \DataOut[29]1 ;
    assign DataOut[28] = \DataOut[28]1 ;
    assign DataOut[27] = \DataOut[27]1 ;
    assign DataOut[26] = \DataOut[26]1 ;
    assign DataOut[25] = \DataOut[25]1 ;
    assign DataOut[24] = \DataOut[24]1 ;
    assign DataOut[23] = \DataOut[23]1 ;
    assign DataOut[22] = \DataOut[22]1 ;
    assign DataOut[21] = \DataOut[21]1 ;
    assign DataOut[20] = \DataOut[20]1 ;
    assign DataOut[19] = \DataOut[19]1 ;
    assign DataOut[18] = \DataOut[18]1 ;
    assign DataOut[17] = \DataOut[17]1 ;
    assign DataOut[16] = \DataOut[16]1 ;
    assign DataOut[15] = \DataOut[15]1 ;
    assign DataOut[14] = \DataOut[14]1 ;
    assign DataOut[13] = \DataOut[13]1 ;
    assign DataOut[12] = \DataOut[12]1 ;
    assign DataOut[11] = \DataOut[11]1 ;
    assign DataOut[10] = \DataOut[10]1 ;
    assign DataOut[9] = \DataOut[9]1 ;
    assign DataOut[8] = \DataOut[8]1 ;
    assign DataOut[7] = \DataOut[7]1 ;
    assign DataOut[6] = \DataOut[6]1 ;
    assign DataOut[5] = \DataOut[5]1 ;
    assign DataOut[4] = \DataOut[4]1 ;
    assign DataOut[3] = \DataOut[3]1 ;
    assign DataOut[2] = \DataOut[2]1 ;
    assign DataOut[1] = \DataOut[1]1 ;
    assign DataOut[0] = \DataOut[0]1 ;
    assign ScanOut[7] = \DataIn[7] ;
    assign ScanOut[6] = \DataIn[6] ;
    assign ScanOut[5] = \DataIn[5] ;
    assign ScanOut[4] = \DataIn[4] ;
    assign ScanOut[3] = \DataIn[3] ;
    assign ScanOut[2] = \DataIn[2] ;
    assign ScanOut[1] = \DataIn[1] ;
    assign ScanOut[0] = \DataIn[0] ;
    VMW_AO22 U54 ( .A(DataIn[8]), .B(n295), .C(\count241[8] ), .D(n296), .Z(
        n362) );
    VMW_AO22 U73 ( .A(DataIn[27]), .B(n295), .C(\count241[27] ), .D(n296), .Z(
        n343) );
    VMW_AO22 U113 ( .A(\ScanReg[2] ), .B(n298), .C(\count[2] ), .D(n297), .Z(
        n322) );
    VMW_BUFIZ U134 ( .A(n312), .E(n311), .Z(\DataOut[4]1 ) );
    VMW_AO22 U68 ( .A(DataIn[22]), .B(n295), .C(\count241[22] ), .D(n296), .Z(
        n348) );
    VMW_AND2 U96 ( .A(n297), .B(\count[14] ), .Z(n314) );
    VMW_AO22 U108 ( .A(\ScanReg[7] ), .B(n298), .C(\count[7] ), .D(n297), .Z(
        n330) );
    VMW_BUFIZ U141 ( .A(n319), .E(n311), .Z(\DataOut[31] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n364), .CP(Clk), .Q(\count[6] ) );
    VMW_AO22 U46 ( .A(\DataIn[0] ), .B(n295), .C(\count241[0] ), .D(n296), .Z(
        n370) );
    VMW_AO22 U61 ( .A(DataIn[15]), .B(n295), .C(\count241[15] ), .D(n296), .Z(
        n355) );
    VMW_AND2 U84 ( .A(n297), .B(\count[17] ), .Z(n329) );
    VMW_BUFIZ U148 ( .A(n326), .E(n311), .Z(\DataOut[20]1 ) );
    VMW_BUFIZ U153 ( .A(n331), .E(n311), .Z(\DataOut[5]1 ) );
    VMW_FD \count_reg[2]  ( .D(n368), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U101 ( .A(n297), .B(\count[19] ), .Z(n307) );
    VMW_INV U126 ( .A(n289), .Z(Enable) );
    VMW_AO22 U48 ( .A(\DataIn[2] ), .B(n295), .C(\count241[2] ), .D(n296), .Z(
        n368) );
    VMW_AO22 U66 ( .A(DataIn[20]), .B(n295), .C(\count241[20] ), .D(n296), .Z(
        n350) );
    VMW_OAI21 U106 ( .A(RD), .B(WR), .C(n301), .Z(n300) );
    VMW_NOR4 U121 ( .A(\count[12] ), .B(\count[13] ), .C(\count[14] ), .D(
        \count[15] ), .Z(n293) );
    VMW_AND2 U83 ( .A(n297), .B(\count[26] ), .Z(n332) );
    VMW_FD \count_reg[0]  ( .D(n370), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U98 ( .A(n297), .B(\count[9] ), .Z(n310) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_INV U128 ( .A(n300), .Z(ScanEnable) );
    VMW_BUFIZ U154 ( .A(n332), .E(n311), .Z(\DataOut[26]1 ) );
    VMW_FD \count_reg[9]  ( .D(n361), .CP(Clk), .Q(\count[9] ) );
    VMW_FD \count_reg[4]  ( .D(n366), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    FFT_Control_SIZE8_IDWIDTH1_SCAN1_DW01_dec_32_0 sub_183 ( .A({\count[31] , 
        \count[30] , \count[29] , \count[28] , \count[27] , \count[26] , 
        \count[25] , \count[24] , \count[23] , \count[22] , \count[21] , 
        \count[20] , \count[19] , \count[18] , \count[17] , \count[16] , 
        \count[15] , \count[14] , \count[13] , \count[12] , \count[11] , 
        \count[10] , \count[9] , \count[8] , \count[7] , \count[6] , 
        \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , \count[0] 
        }), .SUM({\n239[1] , \count241[30] , \count241[29] , \count241[28] , 
        \count241[27] , \count241[26] , \count241[25] , \count241[24] , 
        \count241[23] , \count241[22] , \count241[21] , \count241[20] , 
        \count241[19] , \count241[18] , \count241[17] , \count241[16] , 
        \count241[15] , \count241[14] , \count241[13] , \count241[12] , 
        \count241[11] , \count241[10] , \count241[9] , \count241[8] , 
        \count241[7] , \count241[6] , \count241[5] , \count241[4] , 
        \count241[3] , \count241[2] , \count241[1] , \count241[0] }) );
    VMW_AO22 U53 ( .A(\DataIn[7] ), .B(n295), .C(\count241[7] ), .D(n296), .Z(
        n363) );
    VMW_AND2 U91 ( .A(n297), .B(\count[21] ), .Z(n320) );
    VMW_BUFIZ U146 ( .A(n324), .E(n311), .Z(\DataOut[30]1 ) );
    VMW_AO22 U74 ( .A(DataIn[28]), .B(n295), .C(\count241[28] ), .D(n296), .Z(
        n342) );
    VMW_AO22 U114 ( .A(\ScanReg[1] ), .B(n298), .C(\count[1] ), .D(n297), .Z(
        n337) );
    VMW_BUFIZ U133 ( .A(n310), .E(n311), .Z(\DataOut[9]1 ) );
    VMW_AO21 U99 ( .A(RD), .B(ScanEnable), .C(n297), .Z(n311) );
    VMW_BUFIZ U155 ( .A(n333), .E(n311), .Z(\DataOut[15]1 ) );
    VMW_FD \count_reg[22]  ( .D(n348), .CP(Clk), .Q(\count[22] ) );
    VMW_FD \count_reg[11]  ( .D(n359), .CP(Clk), .Q(\count[11] ) );
    VMW_AO22 U47 ( .A(\DataIn[1] ), .B(n295), .C(\count241[1] ), .D(n296), .Z(
        n369) );
    VMW_AO22 U49 ( .A(\DataIn[3] ), .B(n295), .C(\count241[3] ), .D(n296), .Z(
        n367) );
    VMW_AO22 U52 ( .A(\DataIn[6] ), .B(n295), .C(\count241[6] ), .D(n296), .Z(
        n364) );
    VMW_AO22 U67 ( .A(DataIn[21]), .B(n295), .C(\count241[21] ), .D(n296), .Z(
        n349) );
    VMW_AND2 U82 ( .A(n297), .B(\count[15] ), .Z(n333) );
    VMW_FD \count_reg[18]  ( .D(n352), .CP(Clk), .Q(\count[18] ) );
    VMW_XNOR2 U107 ( .A(Addr[0]), .B(ScanId), .Z(n301) );
    VMW_AND4 U120 ( .A(n305), .B(n304), .C(n303), .D(n302), .Z(n294) );
    VMW_AO22 U75 ( .A(DataIn[29]), .B(n295), .C(\count241[29] ), .D(n296), .Z(
        n341) );
    VMW_AO22 U115 ( .A(\ScanReg[0] ), .B(n298), .C(\count[0] ), .D(n297), .Z(
        n309) );
    VMW_BUFIZ U132 ( .A(n309), .E(n311), .Z(\DataOut[0]1 ) );
    VMW_FD \count_reg[15]  ( .D(n355), .CP(Clk), .Q(\count[15] ) );
    VMW_FD \count_reg[26]  ( .D(n344), .CP(Clk), .Q(\count[26] ) );
    VMW_AND2 U90 ( .A(n297), .B(\count[28] ), .Z(n321) );
    VMW_BUFIZ U129 ( .A(n306), .E(n311), .Z(\DataOut[23]1 ) );
    VMW_BUFIZ U147 ( .A(n325), .E(n311), .Z(\DataOut[29]1 ) );
    VMW_BUFIZ U160 ( .A(n338), .E(n311), .Z(\DataOut[8]1 ) );
    VMW_AO22 U55 ( .A(DataIn[9]), .B(n295), .C(\count241[9] ), .D(n296), .Z(
        n361) );
    VMW_AO22 U69 ( .A(DataIn[23]), .B(n295), .C(\count241[23] ), .D(n296), .Z(
        n347) );
    VMW_AO22 U109 ( .A(\ScanReg[6] ), .B(n298), .C(\count[6] ), .D(n297), .Z(
        n318) );
    VMW_AO22 U72 ( .A(DataIn[26]), .B(n295), .C(\count241[26] ), .D(n296), .Z(
        n344) );
    VMW_AND2 U97 ( .A(n297), .B(\count[27] ), .Z(n313) );
    VMW_BUFIZ U140 ( .A(n318), .E(n311), .Z(\DataOut[6]1 ) );
    VMW_FD \count_reg[17]  ( .D(n353), .CP(Clk), .Q(\count[17] ) );
    VMW_AO22 U112 ( .A(\ScanReg[3] ), .B(n298), .C(\count[3] ), .D(n297), .Z(
        n327) );
    VMW_FD \count_reg[24]  ( .D(n346), .CP(Clk), .Q(\count[24] ) );
    VMW_BUFIZ U135 ( .A(n313), .E(n311), .Z(\DataOut[27]1 ) );
    VMW_AO22 U60 ( .A(DataIn[14]), .B(n295), .C(\count241[14] ), .D(n296), .Z(
        n356) );
    VMW_AND2 U100 ( .A(n297), .B(\count[10] ), .Z(n308) );
    VMW_INV U127 ( .A(WR), .Z(n299) );
    VMW_AND2 U85 ( .A(n297), .B(\count[24] ), .Z(n328) );
    VMW_BUFIZ U149 ( .A(n327), .E(n311), .Z(\DataOut[3]1 ) );
    VMW_FD \count_reg[30]  ( .D(n340), .CP(Clk), .Q(\count[30] ) );
    VMW_FD \count_reg[29]  ( .D(n341), .CP(Clk), .Q(\count[29] ) );
    VMW_BUFIZ U152 ( .A(n330), .E(n311), .Z(\DataOut[7]1 ) );
    VMW_FD \count_reg[20]  ( .D(n350), .CP(Clk), .Q(\count[20] ) );
    VMW_FD \count_reg[13]  ( .D(n357), .CP(Clk), .Q(\count[13] ) );
    VMW_AND5 U45 ( .A(n290), .B(n291), .C(n292), .D(n293), .E(n294), .Z(n289)
         );
    VMW_AO22 U57 ( .A(DataIn[11]), .B(n295), .C(\count241[11] ), .D(n296), .Z(
        n359) );
    VMW_BUFIZ U137 ( .A(n315), .E(n311), .Z(\DataOut[25]1 ) );
    VMW_AO22 U70 ( .A(DataIn[24]), .B(n295), .C(\count241[24] ), .D(n296), .Z(
        n346) );
    VMW_AND2 U79 ( .A(n297), .B(\count[11] ), .Z(n336) );
    VMW_AND2 U95 ( .A(n297), .B(\count[25] ), .Z(n315) );
    VMW_AO22 U110 ( .A(\ScanReg[5] ), .B(n298), .C(\count[5] ), .D(n297), .Z(
        n331) );
    VMW_BUFIZ U159 ( .A(n337), .E(n311), .Z(\DataOut[1]1 ) );
    VMW_NOR4 U119 ( .A(\count[16] ), .B(\count[17] ), .C(\count[18] ), .D(
        \count[19] ), .Z(n305) );
    VMW_BUFIZ U142 ( .A(n320), .E(n311), .Z(\DataOut[21]1 ) );
    VMW_FD \count_reg[31]  ( .D(n339), .CP(Clk), .Q(\count[31] ) );
    VMW_FD \count_reg[28]  ( .D(n342), .CP(Clk), .Q(\count[28] ) );
    VMW_FD \count_reg[21]  ( .D(n349), .CP(Clk), .Q(\count[21] ) );
    VMW_FD \count_reg[12]  ( .D(n358), .CP(Clk), .Q(\count[12] ) );
    VMW_AND2 U87 ( .A(n297), .B(\count[29] ), .Z(n325) );
    VMW_BUFIZ U150 ( .A(n328), .E(n311), .Z(\DataOut[24]1 ) );
    VMW_INV U125 ( .A(n297), .Z(n298) );
    VMW_AO22 U50 ( .A(\DataIn[4] ), .B(n295), .C(\count241[4] ), .D(n296), .Z(
        n366) );
    VMW_AO22 U59 ( .A(DataIn[13]), .B(n295), .C(\count241[13] ), .D(n296), .Z(
        n357) );
    VMW_AO22 U62 ( .A(DataIn[16]), .B(n295), .C(\count241[16] ), .D(n296), .Z(
        n354) );
    VMW_AO22 U65 ( .A(DataIn[19]), .B(n295), .C(\count241[19] ), .D(n296), .Z(
        n351) );
    VMW_AND2 U102 ( .A(n297), .B(\count[23] ), .Z(n306) );
    VMW_FD \count_reg[25]  ( .D(n345), .CP(Clk), .Q(\count[25] ) );
    VMW_FD \count_reg[16]  ( .D(n354), .CP(Clk), .Q(\count[16] ) );
    VMW_NOR3 U105 ( .A(n298), .B(Reset), .C(n299), .Z(n295) );
    VMW_AND2 U80 ( .A(n297), .B(\count[22] ), .Z(n335) );
    VMW_NOR4 U122 ( .A(\count[8] ), .B(\count[9] ), .C(\count[10] ), .D(
        \count[11] ), .Z(n292) );
    VMW_FD \count_reg[14]  ( .D(n356), .CP(Clk), .Q(\count[14] ) );
    VMW_FD \count_reg[27]  ( .D(n343), .CP(Clk), .Q(\count[27] ) );
    VMW_BUFIZ U139 ( .A(n317), .E(n311), .Z(\DataOut[12]1 ) );
    VMW_BUFIZ U157 ( .A(n335), .E(n311), .Z(\DataOut[22]1 ) );
    VMW_AO22 U77 ( .A(DataIn[31]), .B(n295), .C(\n239[1] ), .D(n296), .Z(n339)
         );
    VMW_AND2 U89 ( .A(n297), .B(\count[13] ), .Z(n323) );
    VMW_AND2 U92 ( .A(n297), .B(\count[31] ), .Z(n319) );
    VMW_BUFIZ U145 ( .A(n323), .E(n311), .Z(\DataOut[13]1 ) );
    VMW_FD \count_reg[23]  ( .D(n347), .CP(Clk), .Q(\count[23] ) );
    VMW_FD \count_reg[10]  ( .D(n360), .CP(Clk), .Q(\count[10] ) );
    VMW_NOR4 U117 ( .A(\count[24] ), .B(\count[25] ), .C(\count[26] ), .D(
        \count[27] ), .Z(n303) );
    VMW_FD \count_reg[19]  ( .D(n351), .CP(Clk), .Q(\count[19] ) );
    VMW_AO22 U51 ( .A(\DataIn[5] ), .B(n295), .C(\count241[5] ), .D(n296), .Z(
        n365) );
    VMW_AO22 U58 ( .A(DataIn[12]), .B(n295), .C(\count241[12] ), .D(n296), .Z(
        n358) );
    VMW_BUFIZ U130 ( .A(n307), .E(n311), .Z(\DataOut[19]1 ) );
    VMW_BUFIZ U138 ( .A(n316), .E(n311), .Z(\DataOut[16]1 ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n365), .CP(Clk), .Q(\count[5] ) );
    VMW_AO22 U64 ( .A(DataIn[18]), .B(n295), .C(\count241[18] ), .D(n296), .Z(
        n352) );
    VMW_AND2 U81 ( .A(n297), .B(\count[18] ), .Z(n334) );
    VMW_BUFIZ U156 ( .A(n334), .E(n311), .Z(\DataOut[18]1 ) );
    VMW_AOI211 U104 ( .A(n297), .B(WR), .C(n289), .D(Reset), .Z(n296) );
    VMW_AO22 U76 ( .A(DataIn[30]), .B(n295), .C(\count241[30] ), .D(n296), .Z(
        n340) );
    VMW_NOR4 U116 ( .A(\count[28] ), .B(\count[29] ), .C(\count[30] ), .D(
        \count[31] ), .Z(n302) );
    VMW_NOR4 U123 ( .A(\count[4] ), .B(\count[5] ), .C(\count[6] ), .D(
        \count[7] ), .Z(n291) );
    VMW_AO22 U56 ( .A(DataIn[10]), .B(n295), .C(\count241[10] ), .D(n296), .Z(
        n360) );
    VMW_AND2 U88 ( .A(n297), .B(\count[30] ), .Z(n324) );
    VMW_AND2 U93 ( .A(n297), .B(\count[12] ), .Z(n317) );
    VMW_BUFIZ U131 ( .A(n308), .E(n311), .Z(\DataOut[10]1 ) );
    VMW_FD \count_reg[1]  ( .D(n369), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(n297), .B(\count[16] ), .Z(n316) );
    VMW_BUFIZ U143 ( .A(n321), .E(n311), .Z(\DataOut[28]1 ) );
    VMW_BUFIZ U144 ( .A(n322), .E(n311), .Z(\DataOut[2]1 ) );
    VMW_FD \count_reg[8]  ( .D(n362), .CP(Clk), .Q(\count[8] ) );
    VMW_BUFIZ U158 ( .A(n336), .E(n311), .Z(\DataOut[11]1 ) );
    VMW_FD \count_reg[3]  ( .D(n367), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n314), .E(n311), .Z(\DataOut[14]1 ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AO22 U63 ( .A(DataIn[17]), .B(n295), .C(\count241[17] ), .D(n296), .Z(
        n353) );
    VMW_AO22 U71 ( .A(DataIn[25]), .B(n295), .C(\count241[25] ), .D(n296), .Z(
        n345) );
    VMW_AO22 U111 ( .A(\ScanReg[4] ), .B(n298), .C(\count[4] ), .D(n297), .Z(
        n312) );
    VMW_NOR4 U124 ( .A(\count[0] ), .B(\count[1] ), .C(\count[2] ), .D(
        \count[3] ), .Z(n290) );
    VMW_AND2 U78 ( .A(n297), .B(\count[8] ), .Z(n338) );
    VMW_AND2 U86 ( .A(n297), .B(\count[20] ), .Z(n326) );
    VMW_XNOR2 U103 ( .A(Addr[0]), .B(Id), .Z(n297) );
    VMW_NOR4 U118 ( .A(\count[20] ), .B(\count[21] ), .C(\count[22] ), .D(
        \count[23] ), .Z(n304) );
    VMW_BUFIZ U151 ( .A(n329), .E(n311), .Z(\DataOut[17]1 ) );
    VMW_FD \count_reg[7]  ( .D(n363), .CP(Clk), .Q(\count[7] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nLeftOut_20[8] , \nRightOut_30[7] , \nRightOut_4[1] , 
        \nLeftOut_5[3] , \nLeftOut_8[6] , \nRightOut_9[4] , \nLeftOut_25[5] , 
        \nRightOut_33[4] , \nLeftOut_26[6] , \ScanLink9[6] , \nLeftOut_14[4] , 
        \nRightOut_14[1] , \nRightOut_17[2] , \nRightOut_28[5] , 
        \ScanLink15[7] , \ScanLink16[4] , \nLeftOut_17[7] , \nLeftOut_19[1] , 
        \nRightOut_19[4] , \nLeftOut_6[0] , \nRightOut_25[0] , 
        \nLeftOut_30[2] , \nLeftOut_33[1] , \nRightOut_26[3] , \nLeftOut_0[7] , 
        \nLeftOut_3[4] , \ScanLink4[3] , \nRightOut_4[8] , \ScanLink7[0] , 
        \nRightOut_7[2] , \nLeftOut_11[0] , \nLeftOut_28[0] , \nLeftOut_12[3] , 
        \nLeftOut_36[5] , \nLeftOut_35[6] , \nRightOut_38[6] , \ScanLink1[7] , 
        \nRightOut_1[5] , \ScanLink2[4] , \nRightOut_2[6] , \nLeftOut_33[8] , 
        \nLeftOut_19[8] , \nLeftOut_20[1] , \nRightOut_20[4] , 
        \nRightOut_23[7] , \nLeftOut_23[2] , \nRightOut_35[3] , 
        \nRightOut_36[0] , \nLeftOut_38[3] , \ScanLink7[4] , \nRightOut_7[6] , 
        \nRightOut_11[5] , \nRightOut_14[8] , \ScanLink10[3] , \ScanLink13[0] , 
        \nRightOut_12[6] , \nRightOut_25[4] , \nRightOut_26[7] , 
        \nLeftOut_28[4] , \ScanLink4[7] , \nRightOut_4[5] , \nLeftOut_36[8] , 
        \ScanEnable[0] , \nRightOut_1[8] , \nLeftOut_5[7] , \nLeftOut_6[4] , 
        \nLeftOut_33[5] , \nRightOut_11[8] , \nLeftOut_14[0] , 
        \nLeftOut_30[6] , \nRightOut_14[5] , \nLeftOut_17[3] , 
        \nRightOut_19[0] , \nRightOut_17[6] , \nLeftOut_19[5] , 
        \ScanLink15[3] , \ScanLink16[0] , \nRightOut_9[0] , \nLeftOut_25[1] , 
        \nLeftOut_26[2] , \ScanLink9[2] , \nRightOut_28[1] , \nLeftOut_8[2] , 
        \nRightOut_33[0] , \nRightOut_11[1] , \nRightOut_12[2] , 
        \nRightOut_30[3] , \ScanLink10[7] , \ScanLink13[4] , \ScanLink1[3] , 
        \nLeftOut_20[5] , \nLeftOut_23[6] , \nLeftOut_25[8] , 
        \nRightOut_28[8] , \nRightOut_35[7] , \nRightOut_36[4] , 
        \nLeftOut_38[7] , \nRightOut_1[1] , \ScanLink2[0] , \nRightOut_2[2] , 
        \nRightOut_20[0] , \nRightOut_23[3] , \nLeftOut_35[2] , 
        \nLeftOut_0[3] , \nLeftOut_36[1] , \nLeftOut_0[1] , \ScanLink1[1] , 
        \ScanLink2[2] , \nRightOut_2[0] , \nLeftOut_3[0] , \nRightOut_38[2] , 
        \nLeftOut_11[4] , \nLeftOut_12[7] , \nRightOut_1[3] , \nLeftOut_3[2] , 
        \nRightOut_20[2] , \nRightOut_23[1] , \nLeftOut_35[0] , 
        \nLeftOut_36[3] , \nRightOut_38[0] , \nLeftOut_11[6] , 
        \nRightOut_11[3] , \nLeftOut_12[5] , \nLeftOut_17[8] , 
        \nRightOut_12[0] , \nRightOut_30[8] , \ScanLink10[5] , \ScanLink13[6] , 
        \nRightOut_9[2] , \nRightOut_14[7] , \nRightOut_17[4] , 
        \nLeftOut_20[7] , \nLeftOut_23[4] , \nRightOut_35[5] , 
        \nRightOut_36[6] , \nLeftOut_38[5] , \nLeftOut_19[7] , 
        \nLeftOut_25[3] , \ScanLink15[1] , \ScanLink16[2] , \nLeftOut_26[0] , 
        \nRightOut_28[3] , \ScanLink9[0] , \nRightOut_30[1] , \nLeftOut_0[8] , 
        \nLeftOut_8[0] , \nRightOut_25[6] , \nRightOut_33[2] , 
        \nRightOut_26[5] , \ScanLink4[5] , \nRightOut_4[7] , \nLeftOut_5[5] , 
        \ScanLink7[6] , \nRightOut_7[4] , \nLeftOut_28[6] , \nLeftOut_6[6] , 
        \nRightOut_23[8] , \nLeftOut_14[2] , \nLeftOut_17[1] , 
        \nLeftOut_30[4] , \nLeftOut_33[7] , \nRightOut_19[2] , 
        \nLeftOut_20[3] , \nRightOut_35[1] , \nRightOut_36[2] , 
        \nLeftOut_38[1] , \nLeftOut_23[0] , \ScanLink10[1] , \ScanLink13[2] , 
        \nLeftOut_0[5] , \nLeftOut_11[2] , \nRightOut_11[7] , 
        \nRightOut_12[4] , \nLeftOut_12[1] , \nLeftOut_35[4] , 
        \nLeftOut_36[7] , \ScanLink1[5] , \nRightOut_1[7] , \nLeftOut_3[6] , 
        \nRightOut_26[8] , \nRightOut_38[4] , \ScanLink2[6] , \nRightOut_2[4] , 
        \nRightOut_4[3] , \nLeftOut_5[8] , \nRightOut_20[6] , \nLeftOut_5[1] , 
        \nLeftOut_6[2] , \nLeftOut_12[8] , \nRightOut_23[5] , \nLeftOut_14[6] , 
        \nLeftOut_17[5] , \nRightOut_19[6] , \ScanLink7[2] , \nRightOut_25[2] , 
        \nRightOut_26[1] , \nLeftOut_30[0] , \nLeftOut_33[3] , 
        \nLeftOut_28[2] , \nRightOut_7[0] , \ScanLink4[1] , \nLeftOut_8[4] , 
        \nRightOut_33[6] , \nRightOut_9[6] , \nRightOut_30[5] , \ScanLink9[4] , 
        \nRightOut_10[3] , \nRightOut_13[0] , \nRightOut_14[3] , 
        \nLeftOut_25[7] , \nLeftOut_26[4] , \nRightOut_28[7] , 
        \nRightOut_35[8] , \nLeftOut_38[8] , \ScanLink15[5] , \ScanLink16[6] , 
        \nRightOut_17[0] , \nLeftOut_19[3] , \nLeftOut_21[7] , \ScanLink11[5] , 
        \ScanLink12[6] , \nLeftOut_22[4] , \nRightOut_31[8] , 
        \nRightOut_34[5] , \nLeftOut_39[5] , \nRightOut_0[3] , \ScanLink0[1] , 
        \nRightOut_21[2] , \nRightOut_37[6] , \nRightOut_22[1] , 
        \nLeftOut_1[1] , \ScanLink3[2] , \nRightOut_3[0] , \nLeftOut_2[2] , 
        \nLeftOut_34[0] , \nRightOut_39[0] , \nLeftOut_37[3] , 
        \nLeftOut_10[6] , \nLeftOut_13[5] , \nLeftOut_1[8] , \ScanLink5[5] , 
        \ScanLink6[6] , \nRightOut_6[4] , \nLeftOut_16[8] , \nLeftOut_29[6] , 
        \nRightOut_5[7] , \nLeftOut_4[5] , \nLeftOut_7[6] , \nRightOut_24[6] , 
        \nRightOut_27[5] , \nLeftOut_31[4] , \nLeftOut_32[7] , 
        \nLeftOut_15[2] , \nRightOut_18[2] , \nRightOut_22[8] , 
        \nLeftOut_16[1] , \ScanLink8[0] , \nRightOut_8[2] , \nRightOut_15[7] , 
        \nLeftOut_18[7] , \nRightOut_16[4] , \nLeftOut_27[0] , 
        \nRightOut_29[3] , \ScanLink14[1] , \nLeftOut_9[0] , \nLeftOut_24[3] , 
        \nLeftOut_10[2] , \nRightOut_31[1] , \nRightOut_32[2] , 
        \nLeftOut_13[1] , \nRightOut_0[7] , \nLeftOut_1[5] , \nLeftOut_2[6] , 
        \nRightOut_39[4] , \ScanLink3[6] , \nLeftOut_4[8] , \nRightOut_27[8] , 
        \nLeftOut_34[4] , \nLeftOut_37[7] , \nRightOut_21[6] , 
        \nRightOut_22[5] , \nRightOut_3[4] , \ScanLink0[5] , \nRightOut_37[2] , 
        \nLeftOut_39[1] , \ScanLink8[4] , \nLeftOut_9[4] , \nRightOut_10[7] , 
        \nLeftOut_21[3] , \nLeftOut_22[0] , \nRightOut_34[1] , \ScanLink11[1] , 
        \ScanLink12[2] , \nRightOut_13[4] , \nRightOut_31[5] , 
        \nRightOut_32[6] , \nLeftOut_24[7] , \nRightOut_29[7] , 
        \nRightOut_34[8] , \nLeftOut_39[8] , \nRightOut_8[6] , 
        \nRightOut_15[3] , \nRightOut_16[0] , \nLeftOut_18[3] , 
        \nLeftOut_27[4] , \ScanLink14[5] , \nLeftOut_13[8] , \nLeftOut_15[6] , 
        \nLeftOut_16[5] , \nRightOut_18[6] , \nLeftOut_31[0] , \nLeftOut_4[1] , 
        \nLeftOut_32[3] , \ScanLink5[1] , \nRightOut_5[3] , \nLeftOut_7[2] , 
        \ScanLink6[2] , \nLeftOut_29[2] , \nRightOut_6[0] , \nRightOut_24[2] , 
        \nRightOut_27[1] , \nLeftOut_4[3] , \nLeftOut_7[0] , \nLeftOut_15[4] , 
        \nRightOut_18[4] , \nLeftOut_16[7] , \nLeftOut_31[2] , 
        \nLeftOut_32[1] , \ScanLink5[3] , \nRightOut_5[1] , \ScanLink6[0] , 
        \nRightOut_6[2] , \nLeftOut_29[0] , \nLeftOut_9[6] , \nRightOut_24[0] , 
        \nRightOut_27[3] , \nLeftOut_21[8] , \nRightOut_31[7] , 
        \nRightOut_32[4] , \nRightOut_29[5] , \ScanLink8[6] , \nLeftOut_27[6] , 
        \nRightOut_8[4] , \nRightOut_15[1] , \nLeftOut_18[1] , 
        \nLeftOut_24[5] , \ScanLink14[7] , \nRightOut_16[2] , 
        \nRightOut_34[3] , \nLeftOut_39[3] , \nLeftOut_21[1] , 
        \nRightOut_37[0] , \nLeftOut_22[2] , \nRightOut_10[5] , 
        \nRightOut_13[6] , \nRightOut_15[8] , \ScanLink11[3] , 
        \nLeftOut_18[8] , \ScanLink12[0] , \nLeftOut_10[0] , \nLeftOut_13[3] , 
        \nRightOut_0[8] , \nRightOut_0[5] , \nLeftOut_1[7] , \nLeftOut_2[4] , 
        \nRightOut_5[8] , \nLeftOut_34[6] , \nRightOut_39[6] , 
        \nLeftOut_37[5] , \nRightOut_21[4] , \nRightOut_22[7] , 
        \nLeftOut_32[8] , \ScanLink0[7] , \ScanLink3[4] , \nRightOut_3[6] , 
        \ScanLink5[7] , \ScanLink8[2] , \nRightOut_8[0] , \nRightOut_10[8] , 
        \nRightOut_15[5] , \nRightOut_16[6] , \nLeftOut_18[5] , 
        \ScanLink14[3] , \nLeftOut_24[1] , \nRightOut_29[1] , \nLeftOut_9[2] , 
        \nLeftOut_27[2] , \nRightOut_31[3] , \nRightOut_32[0] , 
        \nRightOut_5[5] , \nLeftOut_37[8] , \ScanLink6[4] , \nRightOut_6[6] , 
        \nLeftOut_29[4] , \nRightOut_24[4] , \nRightOut_27[7] , 
        \nLeftOut_31[6] , \nLeftOut_32[5] , \nLeftOut_4[7] , \nLeftOut_7[4] , 
        \nLeftOut_15[0] , \nLeftOut_16[3] , \nRightOut_18[0] , 
        \nRightOut_0[1] , \ScanLink0[3] , \ScanLink3[0] , \nRightOut_3[2] , 
        \nRightOut_21[0] , \nRightOut_22[3] , \nLeftOut_1[3] , \nLeftOut_2[0] , 
        \nRightOut_39[2] , \nLeftOut_34[2] , \nLeftOut_37[1] , 
        \nLeftOut_10[4] , \nLeftOut_13[7] , \nRightOut_10[1] , 
        \nRightOut_13[2] , \nLeftOut_21[5] , \nLeftOut_22[6] , \ScanLink11[7] , 
        \ScanLink12[4] , \nLeftOut_24[8] , \nRightOut_37[4] , \nLeftOut_39[7] , 
        \nLeftOut_2[8] , \nLeftOut_4[6] , \nLeftOut_7[5] , \ScanLink8[3] , 
        \nLeftOut_9[3] , \nRightOut_15[4] , \nLeftOut_18[4] , 
        \nRightOut_29[8] , \nRightOut_34[7] , \ScanLink14[2] , 
        \nRightOut_16[7] , \nRightOut_32[1] , \nRightOut_29[0] , 
        \nRightOut_31[2] , \nRightOut_8[1] , \nLeftOut_24[0] , 
        \nLeftOut_27[3] , \nLeftOut_31[7] , \nLeftOut_32[4] , 
        \nRightOut_21[8] , \ScanLink5[6] , \nRightOut_5[4] , \ScanLink6[5] , 
        \nLeftOut_29[5] , \nRightOut_6[7] , \nRightOut_27[6] , 
        \nRightOut_24[5] , \nRightOut_0[0] , \nLeftOut_1[2] , \nLeftOut_15[1] , 
        \nRightOut_18[1] , \nLeftOut_16[2] , \nLeftOut_2[1] , 
        \nRightOut_39[3] , \nRightOut_21[1] , \nLeftOut_34[3] , 
        \nLeftOut_37[0] , \nRightOut_22[2] , \ScanLink0[2] , \ScanLink3[1] , 
        \nRightOut_3[3] , \nLeftOut_13[6] , \nLeftOut_15[8] , 
        \nRightOut_18[8] , \nLeftOut_10[5] , \nRightOut_8[8] , 
        \nRightOut_10[0] , \nRightOut_13[3] , \ScanLink11[6] , \ScanLink12[5] , 
        \nRightOut_34[6] , \nLeftOut_39[6] , \nLeftOut_10[8] , 
        \nLeftOut_15[5] , \nLeftOut_16[6] , \nRightOut_18[5] , 
        \nLeftOut_21[4] , \nRightOut_37[5] , \nLeftOut_22[7] , 
        \nRightOut_32[8] , \nLeftOut_4[2] , \ScanLink5[2] , \nRightOut_5[0] , 
        \ScanLink6[1] , \nRightOut_6[3] , \nRightOut_24[1] , \nLeftOut_29[1] , 
        \nRightOut_27[2] , \nLeftOut_31[3] , \nLeftOut_32[0] , \nLeftOut_7[1] , 
        \nRightOut_29[4] , \nRightOut_37[8] , \ScanLink8[7] , \nRightOut_8[5] , 
        \nLeftOut_24[4] , \nLeftOut_27[7] , \nLeftOut_9[7] , \nRightOut_31[6] , 
        \nRightOut_15[0] , \nRightOut_16[3] , \nLeftOut_18[0] , 
        \nRightOut_32[5] , \nLeftOut_21[0] , \nLeftOut_22[3] , \ScanLink14[6] , 
        \nRightOut_37[1] , \nLeftOut_39[2] , \nLeftOut_10[1] , 
        \nRightOut_10[4] , \nRightOut_34[2] , \nRightOut_13[7] , 
        \ScanLink11[2] , \ScanLink12[1] , \nLeftOut_13[2] , \nRightOut_0[4] , 
        \ScanLink0[6] , \ScanLink3[5] , \nRightOut_3[7] , \nLeftOut_7[8] , 
        \nRightOut_22[6] , \nRightOut_21[5] , \nLeftOut_1[6] , \nLeftOut_2[5] , 
        \nRightOut_24[8] , \nRightOut_39[7] , \nLeftOut_13[0] , 
        \nLeftOut_29[8] , \nLeftOut_34[7] , \nLeftOut_37[4] , \nLeftOut_10[3] , 
        \nRightOut_0[6] , \ScanLink0[4] , \nRightOut_21[7] , \nRightOut_22[4] , 
        \nLeftOut_1[4] , \ScanLink3[7] , \nRightOut_3[5] , \nLeftOut_31[8] , 
        \nLeftOut_2[7] , \nRightOut_39[5] , \nRightOut_6[8] , \nLeftOut_21[2] , 
        \nLeftOut_34[5] , \nLeftOut_37[6] , \nLeftOut_22[1] , 
        \nRightOut_34[0] , \nLeftOut_39[0] , \ScanLink8[5] , \nRightOut_8[7] , 
        \nRightOut_10[6] , \nRightOut_13[5] , \nRightOut_37[3] , 
        \nRightOut_16[8] , \ScanLink11[0] , \ScanLink12[3] , \nRightOut_29[6] , 
        \nLeftOut_9[5] , \nLeftOut_24[6] , \nLeftOut_27[5] , \nRightOut_32[7] , 
        \nRightOut_15[2] , \nLeftOut_18[2] , \nLeftOut_22[8] , 
        \nRightOut_31[4] , \nRightOut_16[1] , \ScanLink14[4] , 
        \nLeftOut_15[7] , \nRightOut_18[7] , \nLeftOut_16[4] , \nLeftOut_4[0] , 
        \ScanLink5[0] , \ScanLink6[3] , \nRightOut_6[1] , \nLeftOut_29[3] , 
        \nRightOut_5[2] , \nLeftOut_7[3] , \nRightOut_24[3] , 
        \nRightOut_27[0] , \nLeftOut_31[1] , \nLeftOut_32[2] , 
        \nRightOut_10[2] , \ScanLink11[4] , \ScanLink12[7] , \nRightOut_13[1] , 
        \nLeftOut_27[8] , \nLeftOut_39[4] , \nRightOut_37[7] , 
        \nRightOut_0[2] , \nLeftOut_1[0] , \nLeftOut_2[3] , \nLeftOut_9[8] , 
        \nLeftOut_21[6] , \nLeftOut_22[5] , \nRightOut_34[4] , 
        \nRightOut_39[1] , \ScanLink3[3] , \nRightOut_21[3] , 
        \nRightOut_22[0] , \nLeftOut_34[1] , \nLeftOut_37[2] , 
        \nRightOut_3[1] , \ScanLink0[0] , \nLeftOut_10[7] , \nLeftOut_13[4] , 
        \nRightOut_3[8] , \nLeftOut_4[4] , \nLeftOut_31[5] , \nLeftOut_32[6] , 
        \ScanLink5[4] , \nRightOut_5[6] , \nLeftOut_7[7] , \ScanLink6[7] , 
        \nRightOut_6[5] , \nRightOut_24[7] , \nLeftOut_29[7] , 
        \nLeftOut_34[8] , \nRightOut_27[4] , \nRightOut_39[8] , \ScanLink8[1] , 
        \nLeftOut_9[1] , \nRightOut_13[8] , \nLeftOut_15[3] , \nLeftOut_16[0] , 
        \nRightOut_18[3] , \ScanLink14[0] , \nRightOut_15[6] , 
        \nRightOut_16[5] , \nLeftOut_18[6] , \nRightOut_31[0] , 
        \nLeftOut_24[2] , \nRightOut_29[2] , \nRightOut_32[3] , 
        \nLeftOut_27[1] , \nRightOut_8[3] , \nRightOut_11[6] , 
        \nLeftOut_20[2] , \nLeftOut_23[1] , \nRightOut_35[0] , 
        \nRightOut_36[3] , \nLeftOut_38[0] , \nRightOut_12[5] , 
        \ScanLink13[3] , \nLeftOut_0[4] , \ScanLink1[4] , \ScanLink2[7] , 
        \nRightOut_2[5] , \nLeftOut_11[3] , \nRightOut_17[8] , \ScanLink10[0] , 
        \nLeftOut_12[0] , \nLeftOut_30[8] , \nRightOut_1[6] , \nLeftOut_3[7] , 
        \nRightOut_7[8] , \nRightOut_20[7] , \nRightOut_23[4] , 
        \nLeftOut_36[6] , \nLeftOut_35[5] , \nRightOut_38[5] , \ScanLink4[0] , 
        \nLeftOut_14[7] , \nLeftOut_17[4] , \nRightOut_19[7] , 
        \nRightOut_25[3] , \nRightOut_26[0] , \nRightOut_4[2] , 
        \nLeftOut_5[0] , \ScanLink7[3] , \nRightOut_7[1] , \nLeftOut_28[3] , 
        \nLeftOut_6[3] , \nRightOut_9[7] , \nLeftOut_25[6] , \nLeftOut_30[1] , 
        \nLeftOut_33[2] , \nLeftOut_23[8] , \nLeftOut_26[5] , \ScanLink9[5] , 
        \nRightOut_28[6] , \nLeftOut_0[0] , \nLeftOut_8[5] , \nRightOut_30[4] , 
        \nRightOut_33[7] , \nRightOut_14[2] , \nRightOut_17[1] , 
        \nLeftOut_19[2] , \nLeftOut_35[1] , \ScanLink15[4] , \ScanLink16[7] , 
        \nLeftOut_36[2] , \ScanLink1[0] , \nRightOut_1[2] , \nLeftOut_3[3] , 
        \nRightOut_38[1] , \ScanLink2[3] , \nRightOut_2[1] , \nLeftOut_11[7] , 
        \nLeftOut_12[4] , \nRightOut_20[3] , \nRightOut_23[0] , 
        \ScanLink10[4] , \ScanLink13[7] , \nLeftOut_8[8] , \nRightOut_11[2] , 
        \nRightOut_12[1] , \nLeftOut_26[8] , \nRightOut_35[4] , 
        \nRightOut_36[7] , \nLeftOut_38[4] , \nLeftOut_20[6] , 
        \nRightOut_12[8] , \nLeftOut_23[5] , \ScanLink16[3] , 
        \nRightOut_14[6] , \ScanLink15[0] , \nRightOut_17[5] , 
        \nLeftOut_19[6] , \nLeftOut_8[1] , \nRightOut_30[0] , 
        \nRightOut_33[3] , \nRightOut_2[8] , \nLeftOut_5[4] , \nLeftOut_6[7] , 
        \nRightOut_9[3] , \nLeftOut_26[1] , \ScanLink9[1] , \nLeftOut_25[2] , 
        \nRightOut_28[2] , \nLeftOut_33[6] , \ScanLink4[4] , \nRightOut_4[6] , 
        \ScanLink7[7] , \nRightOut_25[7] , \nRightOut_26[4] , \nLeftOut_30[5] , 
        \nRightOut_38[8] , \nRightOut_7[5] , \nLeftOut_28[7] , 
        \nLeftOut_35[8] , \nLeftOut_3[8] , \nLeftOut_5[6] , \nLeftOut_14[3] , 
        \nLeftOut_17[0] , \nRightOut_19[3] , \nLeftOut_6[5] , 
        \nRightOut_20[8] , \nLeftOut_30[7] , \nLeftOut_33[4] , \ScanLink4[6] , 
        \nRightOut_4[4] , \nRightOut_25[5] , \nRightOut_26[6] , \ScanLink7[5] , 
        \nLeftOut_28[5] , \nRightOut_7[7] , \nLeftOut_14[1] , \nLeftOut_17[2] , 
        \nRightOut_14[4] , \nRightOut_17[7] , \nRightOut_19[1] , 
        \ScanLink15[2] , \ScanLink16[1] , \nLeftOut_19[4] , \nLeftOut_8[3] , 
        \nRightOut_30[2] , \nRightOut_33[1] , \nRightOut_9[8] , 
        \nRightOut_9[1] , \nLeftOut_25[0] , \ScanLink9[3] , \nRightOut_11[0] , 
        \nLeftOut_26[3] , \nRightOut_28[0] , \ScanLink10[6] , \ScanLink13[5] , 
        \nRightOut_12[3] , \nRightOut_35[6] , \nRightOut_36[5] , 
        \nLeftOut_38[6] , \nLeftOut_20[4] , \nLeftOut_23[7] , 
        \nRightOut_33[8] , \nLeftOut_36[0] , \nEnable[0] , \nLeftOut_0[2] , 
        \nLeftOut_3[1] , \nLeftOut_35[3] , \nRightOut_38[3] , \ScanLink1[2] , 
        \nRightOut_1[0] , \ScanLink2[1] , \nRightOut_2[3] , \nRightOut_20[1] , 
        \nRightOut_23[2] , \nRightOut_9[5] , \nLeftOut_11[5] , 
        \nLeftOut_14[8] , \nRightOut_19[8] , \nLeftOut_12[6] , 
        \nLeftOut_26[7] , \nLeftOut_25[4] , \ScanLink9[7] , \nRightOut_28[4] , 
        \nRightOut_36[8] , \nLeftOut_8[7] , \nRightOut_30[6] , 
        \nRightOut_33[5] , \ScanLink4[2] , \ScanLink7[1] , \nRightOut_7[3] , 
        \nLeftOut_11[8] , \nLeftOut_14[5] , \nRightOut_14[0] , 
        \nRightOut_17[3] , \nLeftOut_19[0] , \ScanLink15[6] , \ScanLink16[5] , 
        \nLeftOut_17[6] , \nRightOut_19[5] , \nRightOut_25[1] , 
        \nRightOut_26[2] , \nLeftOut_28[1] , \nLeftOut_0[6] , \ScanLink1[6] , 
        \nRightOut_4[0] , \nLeftOut_5[2] , \nLeftOut_6[1] , \nLeftOut_11[1] , 
        \nLeftOut_12[2] , \nLeftOut_30[3] , \nLeftOut_33[0] , \nRightOut_1[4] , 
        \ScanLink2[5] , \nRightOut_2[7] , \nLeftOut_6[8] , \nRightOut_20[5] , 
        \nRightOut_23[6] , \nLeftOut_28[8] , \nLeftOut_35[7] , 
        \nLeftOut_36[4] , \nLeftOut_3[5] , \nRightOut_11[4] , 
        \nRightOut_12[7] , \nLeftOut_20[0] , \nRightOut_25[8] , 
        \nRightOut_38[7] , \nLeftOut_23[3] , \nRightOut_35[2] , 
        \nRightOut_36[1] , \nLeftOut_38[2] , \ScanLink10[2] , \ScanLink13[1] ;
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink4[7] , \ScanLink4[6] , \ScanLink4[5] , 
        \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , \ScanLink4[1] , 
        \ScanLink4[0] }), .ScanOut({\ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_4[8] , \nLeftOut_4[7] , \nLeftOut_4[6] , \nLeftOut_4[5] , 
        \nLeftOut_4[4] , \nLeftOut_4[3] , \nLeftOut_4[2] , \nLeftOut_4[1] , 
        \nLeftOut_4[0] }), .inright({\nRightOut_4[8] , \nRightOut_4[7] , 
        \nRightOut_4[6] , \nRightOut_4[5] , \nRightOut_4[4] , \nRightOut_4[3] , 
        \nRightOut_4[2] , \nRightOut_4[1] , \nRightOut_4[0] }), .outleft({
        \nLeftOut_4[8] , \nLeftOut_4[7] , \nLeftOut_4[6] , \nLeftOut_4[5] , 
        \nLeftOut_4[4] , \nLeftOut_4[3] , \nLeftOut_4[2] , \nLeftOut_4[1] , 
        \nLeftOut_4[0] }), .outright({\nRightOut_4[8] , \nRightOut_4[7] , 
        \nRightOut_4[6] , \nRightOut_4[5] , \nRightOut_4[4] , \nRightOut_4[3] , 
        \nRightOut_4[2] , \nRightOut_4[1] , \nRightOut_4[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_2[8] , \nLeftOut_2[7] , 
        \nLeftOut_2[6] , \nLeftOut_2[5] , \nLeftOut_2[4] , \nLeftOut_2[3] , 
        \nLeftOut_2[2] , \nLeftOut_2[1] , \nLeftOut_2[0] }), .inright({
        \nRightOut_2[8] , \nRightOut_2[7] , \nRightOut_2[6] , \nRightOut_2[5] , 
        \nRightOut_2[4] , \nRightOut_2[3] , \nRightOut_2[2] , \nRightOut_2[1] , 
        \nRightOut_2[0] }), .outleft({\nLeftOut_10[8] , \nLeftOut_10[7] , 
        \nLeftOut_10[6] , \nLeftOut_10[5] , \nLeftOut_10[4] , \nLeftOut_10[3] , 
        \nLeftOut_10[2] , \nLeftOut_10[1] , \nLeftOut_10[0] }), .outright({
        \nRightOut_10[8] , \nRightOut_10[7] , \nRightOut_10[6] , 
        \nRightOut_10[5] , \nRightOut_10[4] , \nRightOut_10[3] , 
        \nRightOut_10[2] , \nRightOut_10[1] , \nRightOut_10[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s5_SCAN1 node_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_25[8] , \nRightOut_25[7] , 
        \nRightOut_25[6] , \nRightOut_25[5] , \nRightOut_25[4] , 
        \nRightOut_25[3] , \nRightOut_25[2] , \nRightOut_25[1] , 
        \nRightOut_25[0] }), .inright({\nRightOut_29[8] , \nRightOut_29[7] , 
        \nRightOut_29[6] , \nRightOut_29[5] , \nRightOut_29[4] , 
        \nRightOut_29[3] , \nRightOut_29[2] , \nRightOut_29[1] , 
        \nRightOut_29[0] }), .outleft({\nLeftOut_37[8] , \nLeftOut_37[7] , 
        \nLeftOut_37[6] , \nLeftOut_37[5] , \nLeftOut_37[4] , \nLeftOut_37[3] , 
        \nLeftOut_37[2] , \nLeftOut_37[1] , \nLeftOut_37[0] }), .outright({
        \nRightOut_37[8] , \nRightOut_37[7] , \nRightOut_37[6] , 
        \nRightOut_37[5] , \nRightOut_37[4] , \nRightOut_37[3] , 
        \nRightOut_37[2] , \nRightOut_37[1] , \nRightOut_37[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink10[7] , \ScanLink10[6] , \ScanLink10[5] , 
        \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , \ScanLink10[1] , 
        \ScanLink10[0] }), .ScanOut({\ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_36[8] , \nLeftOut_36[7] , \nLeftOut_36[6] , \nLeftOut_36[5] , 
        \nLeftOut_36[4] , \nLeftOut_36[3] , \nLeftOut_36[2] , \nLeftOut_36[1] , 
        \nLeftOut_36[0] }), .inright({\nLeftOut_37[8] , \nLeftOut_37[7] , 
        \nLeftOut_37[6] , \nLeftOut_37[5] , \nLeftOut_37[4] , \nLeftOut_37[3] , 
        \nLeftOut_37[2] , \nLeftOut_37[1] , \nLeftOut_37[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink0[7] , \ScanLink0[6] , \ScanLink0[5] , 
        \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , \ScanLink0[1] , 
        \ScanLink0[0] }), .ScanOut({\ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_0[8] , \nLeftOut_0[7] , \nLeftOut_0[6] , \nLeftOut_0[5] , 
        \nLeftOut_0[4] , \nLeftOut_0[3] , \nLeftOut_0[2] , \nLeftOut_0[1] , 
        \nLeftOut_0[0] }), .inright({\nRightOut_0[8] , \nRightOut_0[7] , 
        \nRightOut_0[6] , \nRightOut_0[5] , \nRightOut_0[4] , \nRightOut_0[3] , 
        \nRightOut_0[2] , \nRightOut_0[1] , \nRightOut_0[0] }), .outleft({
        \nLeftOut_0[8] , \nLeftOut_0[7] , \nLeftOut_0[6] , \nLeftOut_0[5] , 
        \nLeftOut_0[4] , \nLeftOut_0[3] , \nLeftOut_0[2] , \nLeftOut_0[1] , 
        \nLeftOut_0[0] }), .outright({\nRightOut_0[8] , \nRightOut_0[7] , 
        \nRightOut_0[6] , \nRightOut_0[5] , \nRightOut_0[4] , \nRightOut_0[3] , 
        \nRightOut_0[2] , \nRightOut_0[1] , \nRightOut_0[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink2[7] , \ScanLink2[6] , \ScanLink2[5] , 
        \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , \ScanLink2[1] , 
        \ScanLink2[0] }), .ScanOut({\ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_2[8] , \nLeftOut_2[7] , \nLeftOut_2[6] , \nLeftOut_2[5] , 
        \nLeftOut_2[4] , \nLeftOut_2[3] , \nLeftOut_2[2] , \nLeftOut_2[1] , 
        \nLeftOut_2[0] }), .inright({\nRightOut_2[8] , \nRightOut_2[7] , 
        \nRightOut_2[6] , \nRightOut_2[5] , \nRightOut_2[4] , \nRightOut_2[3] , 
        \nRightOut_2[2] , \nRightOut_2[1] , \nRightOut_2[0] }), .outleft({
        \nLeftOut_2[8] , \nLeftOut_2[7] , \nLeftOut_2[6] , \nLeftOut_2[5] , 
        \nLeftOut_2[4] , \nLeftOut_2[3] , \nLeftOut_2[2] , \nLeftOut_2[1] , 
        \nLeftOut_2[0] }), .outright({\nRightOut_2[8] , \nRightOut_2[7] , 
        \nRightOut_2[6] , \nRightOut_2[5] , \nRightOut_2[4] , \nRightOut_2[3] , 
        \nRightOut_2[2] , \nRightOut_2[1] , \nRightOut_2[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink3[7] , \ScanLink3[6] , \ScanLink3[5] , 
        \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , \ScanLink3[1] , 
        \ScanLink3[0] }), .ScanOut({\ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_3[8] , \nLeftOut_3[7] , \nLeftOut_3[6] , \nLeftOut_3[5] , 
        \nLeftOut_3[4] , \nLeftOut_3[3] , \nLeftOut_3[2] , \nLeftOut_3[1] , 
        \nLeftOut_3[0] }), .inright({\nRightOut_3[8] , \nRightOut_3[7] , 
        \nRightOut_3[6] , \nRightOut_3[5] , \nRightOut_3[4] , \nRightOut_3[3] , 
        \nRightOut_3[2] , \nRightOut_3[1] , \nRightOut_3[0] }), .outleft({
        \nLeftOut_3[8] , \nLeftOut_3[7] , \nLeftOut_3[6] , \nLeftOut_3[5] , 
        \nLeftOut_3[4] , \nLeftOut_3[3] , \nLeftOut_3[2] , \nLeftOut_3[1] , 
        \nLeftOut_3[0] }), .outright({\nRightOut_3[8] , \nRightOut_3[7] , 
        \nRightOut_3[6] , \nRightOut_3[5] , \nRightOut_3[4] , \nRightOut_3[3] , 
        \nRightOut_3[2] , \nRightOut_3[1] , \nRightOut_3[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_10[8] , \nRightOut_10[7] , 
        \nRightOut_10[6] , \nRightOut_10[5] , \nRightOut_10[4] , 
        \nRightOut_10[3] , \nRightOut_10[2] , \nRightOut_10[1] , 
        \nRightOut_10[0] }), .inright({\nRightOut_11[8] , \nRightOut_11[7] , 
        \nRightOut_11[6] , \nRightOut_11[5] , \nRightOut_11[4] , 
        \nRightOut_11[3] , \nRightOut_11[2] , \nRightOut_11[1] , 
        \nRightOut_11[0] }), .outleft({\nLeftOut_19[8] , \nLeftOut_19[7] , 
        \nLeftOut_19[6] , \nLeftOut_19[5] , \nLeftOut_19[4] , \nLeftOut_19[3] , 
        \nLeftOut_19[2] , \nLeftOut_19[1] , \nLeftOut_19[0] }), .outright({
        \nRightOut_19[8] , \nRightOut_19[7] , \nRightOut_19[6] , 
        \nRightOut_19[5] , \nRightOut_19[4] , \nRightOut_19[3] , 
        \nRightOut_19[2] , \nRightOut_19[1] , \nRightOut_19[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s2_SCAN1 node_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_17[8] , \nLeftOut_17[7] , 
        \nLeftOut_17[6] , \nLeftOut_17[5] , \nLeftOut_17[4] , \nLeftOut_17[3] , 
        \nLeftOut_17[2] , \nLeftOut_17[1] , \nLeftOut_17[0] }), .inright({
        \nLeftOut_19[8] , \nLeftOut_19[7] , \nLeftOut_19[6] , \nLeftOut_19[5] , 
        \nLeftOut_19[4] , \nLeftOut_19[3] , \nLeftOut_19[2] , \nLeftOut_19[1] , 
        \nLeftOut_19[0] }), .outleft({\nLeftOut_25[8] , \nLeftOut_25[7] , 
        \nLeftOut_25[6] , \nLeftOut_25[5] , \nLeftOut_25[4] , \nLeftOut_25[3] , 
        \nLeftOut_25[2] , \nLeftOut_25[1] , \nLeftOut_25[0] }), .outright({
        \nRightOut_25[8] , \nRightOut_25[7] , \nRightOut_25[6] , 
        \nRightOut_25[5] , \nRightOut_25[4] , \nRightOut_25[3] , 
        \nRightOut_25[2] , \nRightOut_25[1] , \nRightOut_25[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_14[8] , \nLeftOut_14[7] , 
        \nLeftOut_14[6] , \nLeftOut_14[5] , \nLeftOut_14[4] , \nLeftOut_14[3] , 
        \nLeftOut_14[2] , \nLeftOut_14[1] , \nLeftOut_14[0] }), .inright({
        \nLeftOut_15[8] , \nLeftOut_15[7] , \nLeftOut_15[6] , \nLeftOut_15[5] , 
        \nLeftOut_15[4] , \nLeftOut_15[3] , \nLeftOut_15[2] , \nLeftOut_15[1] , 
        \nLeftOut_15[0] }), .outleft({\nLeftOut_22[8] , \nLeftOut_22[7] , 
        \nLeftOut_22[6] , \nLeftOut_22[5] , \nLeftOut_22[4] , \nLeftOut_22[3] , 
        \nLeftOut_22[2] , \nLeftOut_22[1] , \nLeftOut_22[0] }), .outright({
        \nRightOut_22[8] , \nRightOut_22[7] , \nRightOut_22[6] , 
        \nRightOut_22[5] , \nRightOut_22[4] , \nRightOut_22[3] , 
        \nRightOut_22[2] , \nRightOut_22[1] , \nRightOut_22[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s7_SCAN1 node_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_27[8] , \nRightOut_27[7] , 
        \nRightOut_27[6] , \nRightOut_27[5] , \nRightOut_27[4] , 
        \nRightOut_27[3] , \nRightOut_27[2] , \nRightOut_27[1] , 
        \nRightOut_27[0] }), .inright({\nRightOut_31[8] , \nRightOut_31[7] , 
        \nRightOut_31[6] , \nRightOut_31[5] , \nRightOut_31[4] , 
        \nRightOut_31[3] , \nRightOut_31[2] , \nRightOut_31[1] , 
        \nRightOut_31[0] }), .outleft({\nLeftOut_39[8] , \nLeftOut_39[7] , 
        \nLeftOut_39[6] , \nLeftOut_39[5] , \nLeftOut_39[4] , \nLeftOut_39[3] , 
        \nLeftOut_39[2] , \nLeftOut_39[1] , \nLeftOut_39[0] }), .outright({
        \nRightOut_39[8] , \nRightOut_39[7] , \nRightOut_39[6] , 
        \nRightOut_39[5] , \nRightOut_39[4] , \nRightOut_39[3] , 
        \nRightOut_39[2] , \nRightOut_39[1] , \nRightOut_39[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_8[8] , \nLeftOut_8[7] , 
        \nLeftOut_8[6] , \nLeftOut_8[5] , \nLeftOut_8[4] , \nLeftOut_8[3] , 
        \nLeftOut_8[2] , \nLeftOut_8[1] , \nLeftOut_8[0] }), .inright({
        \nLeftOut_9[8] , \nLeftOut_9[7] , \nLeftOut_9[6] , \nLeftOut_9[5] , 
        \nLeftOut_9[4] , \nLeftOut_9[3] , \nLeftOut_9[2] , \nLeftOut_9[1] , 
        \nLeftOut_9[0] }), .outleft({\nLeftOut_16[8] , \nLeftOut_16[7] , 
        \nLeftOut_16[6] , \nLeftOut_16[5] , \nLeftOut_16[4] , \nLeftOut_16[3] , 
        \nLeftOut_16[2] , \nLeftOut_16[1] , \nLeftOut_16[0] }), .outright({
        \nRightOut_16[8] , \nRightOut_16[7] , \nRightOut_16[6] , 
        \nRightOut_16[5] , \nRightOut_16[4] , \nRightOut_16[3] , 
        \nRightOut_16[2] , \nRightOut_16[1] , \nRightOut_16[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_8[8] , \nRightOut_8[7] , 
        \nRightOut_8[6] , \nRightOut_8[5] , \nRightOut_8[4] , \nRightOut_8[3] , 
        \nRightOut_8[2] , \nRightOut_8[1] , \nRightOut_8[0] }), .inright({
        \nRightOut_9[8] , \nRightOut_9[7] , \nRightOut_9[6] , \nRightOut_9[5] , 
        \nRightOut_9[4] , \nRightOut_9[3] , \nRightOut_9[2] , \nRightOut_9[1] , 
        \nRightOut_9[0] }), .outleft({\nLeftOut_17[8] , \nLeftOut_17[7] , 
        \nLeftOut_17[6] , \nLeftOut_17[5] , \nLeftOut_17[4] , \nLeftOut_17[3] , 
        \nLeftOut_17[2] , \nLeftOut_17[1] , \nLeftOut_17[0] }), .outright({
        \nRightOut_17[8] , \nRightOut_17[7] , \nRightOut_17[6] , 
        \nRightOut_17[5] , \nRightOut_17[4] , \nRightOut_17[3] , 
        \nRightOut_17[2] , \nRightOut_17[1] , \nRightOut_17[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_14[8] , \nRightOut_14[7] , 
        \nRightOut_14[6] , \nRightOut_14[5] , \nRightOut_14[4] , 
        \nRightOut_14[3] , \nRightOut_14[2] , \nRightOut_14[1] , 
        \nRightOut_14[0] }), .inright({\nRightOut_15[8] , \nRightOut_15[7] , 
        \nRightOut_15[6] , \nRightOut_15[5] , \nRightOut_15[4] , 
        \nRightOut_15[3] , \nRightOut_15[2] , \nRightOut_15[1] , 
        \nRightOut_15[0] }), .outleft({\nLeftOut_23[8] , \nLeftOut_23[7] , 
        \nLeftOut_23[6] , \nLeftOut_23[5] , \nLeftOut_23[4] , \nLeftOut_23[3] , 
        \nLeftOut_23[2] , \nLeftOut_23[1] , \nLeftOut_23[0] }), .outright({
        \nRightOut_23[8] , \nRightOut_23[7] , \nRightOut_23[6] , 
        \nRightOut_23[5] , \nRightOut_23[4] , \nRightOut_23[3] , 
        \nRightOut_23[2] , \nRightOut_23[1] , \nRightOut_23[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_20[8] , \nRightOut_20[7] , 
        \nRightOut_20[6] , \nRightOut_20[5] , \nRightOut_20[4] , 
        \nRightOut_20[3] , \nRightOut_20[2] , \nRightOut_20[1] , 
        \nRightOut_20[0] }), .inright({\nRightOut_22[8] , \nRightOut_22[7] , 
        \nRightOut_22[6] , \nRightOut_22[5] , \nRightOut_22[4] , 
        \nRightOut_22[3] , \nRightOut_22[2] , \nRightOut_22[1] , 
        \nRightOut_22[0] }), .outleft({\nLeftOut_30[8] , \nLeftOut_30[7] , 
        \nLeftOut_30[6] , \nLeftOut_30[5] , \nLeftOut_30[4] , \nLeftOut_30[3] , 
        \nLeftOut_30[2] , \nLeftOut_30[1] , \nLeftOut_30[0] }), .outright({
        \nRightOut_30[8] , \nRightOut_30[7] , \nRightOut_30[6] , 
        \nRightOut_30[5] , \nRightOut_30[4] , \nRightOut_30[3] , 
        \nRightOut_30[2] , \nRightOut_30[1] , \nRightOut_30[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink13[7] , \ScanLink13[6] , \ScanLink13[5] , 
        \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , \ScanLink13[1] , 
        \ScanLink13[0] }), .ScanOut({\ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_34[8] , \nRightOut_34[7] , \nRightOut_34[6] , 
        \nRightOut_34[5] , \nRightOut_34[4] , \nRightOut_34[3] , 
        \nRightOut_34[2] , \nRightOut_34[1] , \nRightOut_34[0] }), .inright({
        \nRightOut_35[8] , \nRightOut_35[7] , \nRightOut_35[6] , 
        \nRightOut_35[5] , \nRightOut_35[4] , \nRightOut_35[3] , 
        \nRightOut_35[2] , \nRightOut_35[1] , \nRightOut_35[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s6_SCAN1 node_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_26[8] , \nRightOut_26[7] , 
        \nRightOut_26[6] , \nRightOut_26[5] , \nRightOut_26[4] , 
        \nRightOut_26[3] , \nRightOut_26[2] , \nRightOut_26[1] , 
        \nRightOut_26[0] }), .inright({\nRightOut_30[8] , \nRightOut_30[7] , 
        \nRightOut_30[6] , \nRightOut_30[5] , \nRightOut_30[4] , 
        \nRightOut_30[3] , \nRightOut_30[2] , \nRightOut_30[1] , 
        \nRightOut_30[0] }), .outleft({\nLeftOut_38[8] , \nLeftOut_38[7] , 
        \nLeftOut_38[6] , \nLeftOut_38[5] , \nLeftOut_38[4] , \nLeftOut_38[3] , 
        \nLeftOut_38[2] , \nLeftOut_38[1] , \nLeftOut_38[0] }), .outright({
        \nRightOut_38[8] , \nRightOut_38[7] , \nRightOut_38[6] , 
        \nRightOut_38[5] , \nRightOut_38[4] , \nRightOut_38[3] , 
        \nRightOut_38[2] , \nRightOut_38[1] , \nRightOut_38[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink12[7] , \ScanLink12[6] , \ScanLink12[5] , 
        \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , \ScanLink12[1] , 
        \ScanLink12[0] }), .ScanOut({\ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_32[8] , \nRightOut_32[7] , \nRightOut_32[6] , 
        \nRightOut_32[5] , \nRightOut_32[4] , \nRightOut_32[3] , 
        \nRightOut_32[2] , \nRightOut_32[1] , \nRightOut_32[0] }), .inright({
        \nRightOut_33[8] , \nRightOut_33[7] , \nRightOut_33[6] , 
        \nRightOut_33[5] , \nRightOut_33[4] , \nRightOut_33[3] , 
        \nRightOut_33[2] , \nRightOut_33[1] , \nRightOut_33[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s6_SCAN1 node_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_21[8] , \nRightOut_21[7] , 
        \nRightOut_21[6] , \nRightOut_21[5] , \nRightOut_21[4] , 
        \nRightOut_21[3] , \nRightOut_21[2] , \nRightOut_21[1] , 
        \nRightOut_21[0] }), .inright({\nRightOut_23[8] , \nRightOut_23[7] , 
        \nRightOut_23[6] , \nRightOut_23[5] , \nRightOut_23[4] , 
        \nRightOut_23[3] , \nRightOut_23[2] , \nRightOut_23[1] , 
        \nRightOut_23[0] }), .outleft({\nLeftOut_31[8] , \nLeftOut_31[7] , 
        \nLeftOut_31[6] , \nLeftOut_31[5] , \nLeftOut_31[4] , \nLeftOut_31[3] , 
        \nLeftOut_31[2] , \nLeftOut_31[1] , \nLeftOut_31[0] }), .outright({
        \nRightOut_31[8] , \nRightOut_31[7] , \nRightOut_31[6] , 
        \nRightOut_31[5] , \nRightOut_31[4] , \nRightOut_31[3] , 
        \nRightOut_31[2] , \nRightOut_31[1] , \nRightOut_31[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink5[7] , \ScanLink5[6] , \ScanLink5[5] , 
        \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , \ScanLink5[1] , 
        \ScanLink5[0] }), .ScanOut({\ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_5[8] , \nLeftOut_5[7] , \nLeftOut_5[6] , \nLeftOut_5[5] , 
        \nLeftOut_5[4] , \nLeftOut_5[3] , \nLeftOut_5[2] , \nLeftOut_5[1] , 
        \nLeftOut_5[0] }), .inright({\nRightOut_5[8] , \nRightOut_5[7] , 
        \nRightOut_5[6] , \nRightOut_5[5] , \nRightOut_5[4] , \nRightOut_5[3] , 
        \nRightOut_5[2] , \nRightOut_5[1] , \nRightOut_5[0] }), .outleft({
        \nLeftOut_5[8] , \nLeftOut_5[7] , \nLeftOut_5[6] , \nLeftOut_5[5] , 
        \nLeftOut_5[4] , \nLeftOut_5[3] , \nLeftOut_5[2] , \nLeftOut_5[1] , 
        \nLeftOut_5[0] }), .outright({\nRightOut_5[8] , \nRightOut_5[7] , 
        \nRightOut_5[6] , \nRightOut_5[5] , \nRightOut_5[4] , \nRightOut_5[3] , 
        \nRightOut_5[2] , \nRightOut_5[1] , \nRightOut_5[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink7[7] , \ScanLink7[6] , \ScanLink7[5] , 
        \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , \ScanLink7[1] , 
        \ScanLink7[0] }), .ScanOut({\ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_7[8] , \nLeftOut_7[7] , \nLeftOut_7[6] , \nLeftOut_7[5] , 
        \nLeftOut_7[4] , \nLeftOut_7[3] , \nLeftOut_7[2] , \nLeftOut_7[1] , 
        \nLeftOut_7[0] }), .inright({\nRightOut_7[8] , \nRightOut_7[7] , 
        \nRightOut_7[6] , \nRightOut_7[5] , \nRightOut_7[4] , \nRightOut_7[3] , 
        \nRightOut_7[2] , \nRightOut_7[1] , \nRightOut_7[0] }), .outleft({
        \nLeftOut_7[8] , \nLeftOut_7[7] , \nLeftOut_7[6] , \nLeftOut_7[5] , 
        \nLeftOut_7[4] , \nLeftOut_7[3] , \nLeftOut_7[2] , \nLeftOut_7[1] , 
        \nLeftOut_7[0] }), .outright({\nRightOut_7[8] , \nRightOut_7[7] , 
        \nRightOut_7[6] , \nRightOut_7[5] , \nRightOut_7[4] , \nRightOut_7[3] , 
        \nRightOut_7[2] , \nRightOut_7[1] , \nRightOut_7[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_3[8] , \nLeftOut_3[7] , 
        \nLeftOut_3[6] , \nLeftOut_3[5] , \nLeftOut_3[4] , \nLeftOut_3[3] , 
        \nLeftOut_3[2] , \nLeftOut_3[1] , \nLeftOut_3[0] }), .inright({
        \nRightOut_3[8] , \nRightOut_3[7] , \nRightOut_3[6] , \nRightOut_3[5] , 
        \nRightOut_3[4] , \nRightOut_3[3] , \nRightOut_3[2] , \nRightOut_3[1] , 
        \nRightOut_3[0] }), .outleft({\nLeftOut_11[8] , \nLeftOut_11[7] , 
        \nLeftOut_11[6] , \nLeftOut_11[5] , \nLeftOut_11[4] , \nLeftOut_11[3] , 
        \nLeftOut_11[2] , \nLeftOut_11[1] , \nLeftOut_11[0] }), .outright({
        \nRightOut_11[8] , \nRightOut_11[7] , \nRightOut_11[6] , 
        \nRightOut_11[5] , \nRightOut_11[4] , \nRightOut_11[3] , 
        \nRightOut_11[2] , \nRightOut_11[1] , \nRightOut_11[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_24[8] , \nRightOut_24[7] , 
        \nRightOut_24[6] , \nRightOut_24[5] , \nRightOut_24[4] , 
        \nRightOut_24[3] , \nRightOut_24[2] , \nRightOut_24[1] , 
        \nRightOut_24[0] }), .inright({\nRightOut_28[8] , \nRightOut_28[7] , 
        \nRightOut_28[6] , \nRightOut_28[5] , \nRightOut_28[4] , 
        \nRightOut_28[3] , \nRightOut_28[2] , \nRightOut_28[1] , 
        \nRightOut_28[0] }), .outleft({\nLeftOut_36[8] , \nLeftOut_36[7] , 
        \nLeftOut_36[6] , \nLeftOut_36[5] , \nLeftOut_36[4] , \nLeftOut_36[3] , 
        \nLeftOut_36[2] , \nLeftOut_36[1] , \nLeftOut_36[0] }), .outright({
        \nRightOut_36[8] , \nRightOut_36[7] , \nRightOut_36[6] , 
        \nRightOut_36[5] , \nRightOut_36[4] , \nRightOut_36[3] , 
        \nRightOut_36[2] , \nRightOut_36[1] , \nRightOut_36[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_5[8] , \nLeftOut_5[7] , 
        \nLeftOut_5[6] , \nLeftOut_5[5] , \nLeftOut_5[4] , \nLeftOut_5[3] , 
        \nLeftOut_5[2] , \nLeftOut_5[1] , \nLeftOut_5[0] }), .inright({
        \nRightOut_5[8] , \nRightOut_5[7] , \nRightOut_5[6] , \nRightOut_5[5] , 
        \nRightOut_5[4] , \nRightOut_5[3] , \nRightOut_5[2] , \nRightOut_5[1] , 
        \nRightOut_5[0] }), .outleft({\nLeftOut_13[8] , \nLeftOut_13[7] , 
        \nLeftOut_13[6] , \nLeftOut_13[5] , \nLeftOut_13[4] , \nLeftOut_13[3] , 
        \nLeftOut_13[2] , \nLeftOut_13[1] , \nLeftOut_13[0] }), .outright({
        \nRightOut_13[8] , \nRightOut_13[7] , \nRightOut_13[6] , 
        \nRightOut_13[5] , \nRightOut_13[4] , \nRightOut_13[3] , 
        \nRightOut_13[2] , \nRightOut_13[1] , \nRightOut_13[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_10[8] , \nLeftOut_10[7] , 
        \nLeftOut_10[6] , \nLeftOut_10[5] , \nLeftOut_10[4] , \nLeftOut_10[3] , 
        \nLeftOut_10[2] , \nLeftOut_10[1] , \nLeftOut_10[0] }), .inright({
        \nLeftOut_11[8] , \nLeftOut_11[7] , \nLeftOut_11[6] , \nLeftOut_11[5] , 
        \nLeftOut_11[4] , \nLeftOut_11[3] , \nLeftOut_11[2] , \nLeftOut_11[1] , 
        \nLeftOut_11[0] }), .outleft({\nLeftOut_18[8] , \nLeftOut_18[7] , 
        \nLeftOut_18[6] , \nLeftOut_18[5] , \nLeftOut_18[4] , \nLeftOut_18[3] , 
        \nLeftOut_18[2] , \nLeftOut_18[1] , \nLeftOut_18[0] }), .outright({
        \nRightOut_18[8] , \nRightOut_18[7] , \nRightOut_18[6] , 
        \nRightOut_18[5] , \nRightOut_18[4] , \nRightOut_18[3] , 
        \nRightOut_18[2] , \nRightOut_18[1] , \nRightOut_18[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink11[7] , \ScanLink11[6] , \ScanLink11[5] , 
        \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , \ScanLink11[1] , 
        \ScanLink11[0] }), .ScanOut({\ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_38[8] , \nLeftOut_38[7] , \nLeftOut_38[6] , \nLeftOut_38[5] , 
        \nLeftOut_38[4] , \nLeftOut_38[3] , \nLeftOut_38[2] , \nLeftOut_38[1] , 
        \nLeftOut_38[0] }), .inright({\nLeftOut_39[8] , \nLeftOut_39[7] , 
        \nLeftOut_39[6] , \nLeftOut_39[5] , \nLeftOut_39[4] , \nLeftOut_39[3] , 
        \nLeftOut_39[2] , \nLeftOut_39[1] , \nLeftOut_39[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_16[8] , \nLeftOut_16[7] , 
        \nLeftOut_16[6] , \nLeftOut_16[5] , \nLeftOut_16[4] , \nLeftOut_16[3] , 
        \nLeftOut_16[2] , \nLeftOut_16[1] , \nLeftOut_16[0] }), .inright({
        \nLeftOut_18[8] , \nLeftOut_18[7] , \nLeftOut_18[6] , \nLeftOut_18[5] , 
        \nLeftOut_18[4] , \nLeftOut_18[3] , \nLeftOut_18[2] , \nLeftOut_18[1] , 
        \nLeftOut_18[0] }), .outleft({\nLeftOut_24[8] , \nLeftOut_24[7] , 
        \nLeftOut_24[6] , \nLeftOut_24[5] , \nLeftOut_24[4] , \nLeftOut_24[3] , 
        \nLeftOut_24[2] , \nLeftOut_24[1] , \nLeftOut_24[0] }), .outright({
        \nRightOut_24[8] , \nRightOut_24[7] , \nRightOut_24[6] , 
        \nRightOut_24[5] , \nRightOut_24[4] , \nRightOut_24[3] , 
        \nRightOut_24[2] , \nRightOut_24[1] , \nRightOut_24[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink9[7] , \ScanLink9[6] , \ScanLink9[5] , 
        \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , \ScanLink9[1] , 
        \ScanLink9[0] }), .ScanOut({\ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_34[8] , \nLeftOut_34[7] , \nLeftOut_34[6] , \nLeftOut_34[5] , 
        \nLeftOut_34[4] , \nLeftOut_34[3] , \nLeftOut_34[2] , \nLeftOut_34[1] , 
        \nLeftOut_34[0] }), .inright({\nLeftOut_35[8] , \nLeftOut_35[7] , 
        \nLeftOut_35[6] , \nLeftOut_35[5] , \nLeftOut_35[4] , \nLeftOut_35[3] , 
        \nLeftOut_35[2] , \nLeftOut_35[1] , \nLeftOut_35[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s2_SCAN1 node_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_26[8] , \nLeftOut_26[7] , 
        \nLeftOut_26[6] , \nLeftOut_26[5] , \nLeftOut_26[4] , \nLeftOut_26[3] , 
        \nLeftOut_26[2] , \nLeftOut_26[1] , \nLeftOut_26[0] }), .inright({
        \nLeftOut_30[8] , \nLeftOut_30[7] , \nLeftOut_30[6] , \nLeftOut_30[5] , 
        \nLeftOut_30[4] , \nLeftOut_30[3] , \nLeftOut_30[2] , \nLeftOut_30[1] , 
        \nLeftOut_30[0] }), .outleft({\nLeftOut_34[8] , \nLeftOut_34[7] , 
        \nLeftOut_34[6] , \nLeftOut_34[5] , \nLeftOut_34[4] , \nLeftOut_34[3] , 
        \nLeftOut_34[2] , \nLeftOut_34[1] , \nLeftOut_34[0] }), .outright({
        \nRightOut_34[8] , \nRightOut_34[7] , \nRightOut_34[6] , 
        \nRightOut_34[5] , \nRightOut_34[4] , \nRightOut_34[3] , 
        \nRightOut_34[2] , \nRightOut_34[1] , \nRightOut_34[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_9 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .ScanIn({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_1[8] , \nLeftOut_1[7] , \nLeftOut_1[6] , \nLeftOut_1[5] , 
        \nLeftOut_1[4] , \nLeftOut_1[3] , \nLeftOut_1[2] , \nLeftOut_1[1] , 
        \nLeftOut_1[0] }), .inright({\nRightOut_1[8] , \nRightOut_1[7] , 
        \nRightOut_1[6] , \nRightOut_1[5] , \nRightOut_1[4] , \nRightOut_1[3] , 
        \nRightOut_1[2] , \nRightOut_1[1] , \nRightOut_1[0] }), .outleft({
        \nLeftOut_9[8] , \nLeftOut_9[7] , \nLeftOut_9[6] , \nLeftOut_9[5] , 
        \nLeftOut_9[4] , \nLeftOut_9[3] , \nLeftOut_9[2] , \nLeftOut_9[1] , 
        \nLeftOut_9[0] }), .outright({\nRightOut_9[8] , \nRightOut_9[7] , 
        \nRightOut_9[6] , \nRightOut_9[5] , \nRightOut_9[4] , \nRightOut_9[3] , 
        \nRightOut_9[2] , \nRightOut_9[1] , \nRightOut_9[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_16[8] , \nRightOut_16[7] , 
        \nRightOut_16[6] , \nRightOut_16[5] , \nRightOut_16[4] , 
        \nRightOut_16[3] , \nRightOut_16[2] , \nRightOut_16[1] , 
        \nRightOut_16[0] }), .inright({\nRightOut_18[8] , \nRightOut_18[7] , 
        \nRightOut_18[6] , \nRightOut_18[5] , \nRightOut_18[4] , 
        \nRightOut_18[3] , \nRightOut_18[2] , \nRightOut_18[1] , 
        \nRightOut_18[0] }), .outleft({\nLeftOut_26[8] , \nLeftOut_26[7] , 
        \nLeftOut_26[6] , \nLeftOut_26[5] , \nLeftOut_26[4] , \nLeftOut_26[3] , 
        \nLeftOut_26[2] , \nLeftOut_26[1] , \nLeftOut_26[0] }), .outright({
        \nRightOut_26[8] , \nRightOut_26[7] , \nRightOut_26[6] , 
        \nRightOut_26[5] , \nRightOut_26[4] , \nRightOut_26[3] , 
        \nRightOut_26[2] , \nRightOut_26[1] , \nRightOut_26[0] }) );
    FFT_Control_SIZE8_IDWIDTH1_SCAN1 node_Control ( .Clk(Clk), .Reset(Reset), 
        .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink16[7] , \ScanLink16[6] , \ScanLink16[5] , 
        \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , \ScanLink16[1] , 
        \ScanLink16[0] }), .ScanOut({\ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(\ScanEnable[0] ), 
        .ScanId(1'b1), .Id(1'b0), .Enable(\nEnable[0] ) );
    FFT_Node_SIZE8_IDWIDTH1_s4_SCAN1 node_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_12[8] , \nRightOut_12[7] , 
        \nRightOut_12[6] , \nRightOut_12[5] , \nRightOut_12[4] , 
        \nRightOut_12[3] , \nRightOut_12[2] , \nRightOut_12[1] , 
        \nRightOut_12[0] }), .inright({\nRightOut_13[8] , \nRightOut_13[7] , 
        \nRightOut_13[6] , \nRightOut_13[5] , \nRightOut_13[4] , 
        \nRightOut_13[3] , \nRightOut_13[2] , \nRightOut_13[1] , 
        \nRightOut_13[0] }), .outleft({\nLeftOut_21[8] , \nLeftOut_21[7] , 
        \nLeftOut_21[6] , \nLeftOut_21[5] , \nLeftOut_21[4] , \nLeftOut_21[3] , 
        \nLeftOut_21[2] , \nLeftOut_21[1] , \nLeftOut_21[0] }), .outright({
        \nRightOut_21[8] , \nRightOut_21[7] , \nRightOut_21[6] , 
        \nRightOut_21[5] , \nRightOut_21[4] , \nRightOut_21[3] , 
        \nRightOut_21[2] , \nRightOut_21[1] , \nRightOut_21[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink1[7] , \ScanLink1[6] , \ScanLink1[5] , 
        \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , \ScanLink1[1] , 
        \ScanLink1[0] }), .ScanOut({\ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_1[8] , \nLeftOut_1[7] , \nLeftOut_1[6] , \nLeftOut_1[5] , 
        \nLeftOut_1[4] , \nLeftOut_1[3] , \nLeftOut_1[2] , \nLeftOut_1[1] , 
        \nLeftOut_1[0] }), .inright({\nRightOut_1[8] , \nRightOut_1[7] , 
        \nRightOut_1[6] , \nRightOut_1[5] , \nRightOut_1[4] , \nRightOut_1[3] , 
        \nRightOut_1[2] , \nRightOut_1[1] , \nRightOut_1[0] }), .outleft({
        \nLeftOut_1[8] , \nLeftOut_1[7] , \nLeftOut_1[6] , \nLeftOut_1[5] , 
        \nLeftOut_1[4] , \nLeftOut_1[3] , \nLeftOut_1[2] , \nLeftOut_1[1] , 
        \nLeftOut_1[0] }), .outright({\nRightOut_1[8] , \nRightOut_1[7] , 
        \nRightOut_1[6] , \nRightOut_1[5] , \nRightOut_1[4] , \nRightOut_1[3] , 
        \nRightOut_1[2] , \nRightOut_1[1] , \nRightOut_1[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_8 ( .Clk(Clk), .Reset(Reset), .RD(RD
        ), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .ScanIn({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ScanEnable(1'b0), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_0[8] , \nLeftOut_0[7] , \nLeftOut_0[6] , \nLeftOut_0[5] , 
        \nLeftOut_0[4] , \nLeftOut_0[3] , \nLeftOut_0[2] , \nLeftOut_0[1] , 
        \nLeftOut_0[0] }), .inright({\nRightOut_0[8] , \nRightOut_0[7] , 
        \nRightOut_0[6] , \nRightOut_0[5] , \nRightOut_0[4] , \nRightOut_0[3] , 
        \nRightOut_0[2] , \nRightOut_0[1] , \nRightOut_0[0] }), .outleft({
        \nLeftOut_8[8] , \nLeftOut_8[7] , \nLeftOut_8[6] , \nLeftOut_8[5] , 
        \nLeftOut_8[4] , \nLeftOut_8[3] , \nLeftOut_8[2] , \nLeftOut_8[1] , 
        \nLeftOut_8[0] }), .outright({\nRightOut_8[8] , \nRightOut_8[7] , 
        \nRightOut_8[6] , \nRightOut_8[5] , \nRightOut_8[4] , \nRightOut_8[3] , 
        \nRightOut_8[2] , \nRightOut_8[1] , \nRightOut_8[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_6[8] , \nLeftOut_6[7] , 
        \nLeftOut_6[6] , \nLeftOut_6[5] , \nLeftOut_6[4] , \nLeftOut_6[3] , 
        \nLeftOut_6[2] , \nLeftOut_6[1] , \nLeftOut_6[0] }), .inright({
        \nRightOut_6[8] , \nRightOut_6[7] , \nRightOut_6[6] , \nRightOut_6[5] , 
        \nRightOut_6[4] , \nRightOut_6[3] , \nRightOut_6[2] , \nRightOut_6[1] , 
        \nRightOut_6[0] }), .outleft({\nLeftOut_14[8] , \nLeftOut_14[7] , 
        \nLeftOut_14[6] , \nLeftOut_14[5] , \nLeftOut_14[4] , \nLeftOut_14[3] , 
        \nLeftOut_14[2] , \nLeftOut_14[1] , \nLeftOut_14[0] }), .outright({
        \nRightOut_14[8] , \nRightOut_14[7] , \nRightOut_14[6] , 
        \nRightOut_14[5] , \nRightOut_14[4] , \nRightOut_14[3] , 
        \nRightOut_14[2] , \nRightOut_14[1] , \nRightOut_14[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s1_SCAN1 node_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_25[8] , \nLeftOut_25[7] , 
        \nLeftOut_25[6] , \nLeftOut_25[5] , \nLeftOut_25[4] , \nLeftOut_25[3] , 
        \nLeftOut_25[2] , \nLeftOut_25[1] , \nLeftOut_25[0] }), .inright({
        \nLeftOut_29[8] , \nLeftOut_29[7] , \nLeftOut_29[6] , \nLeftOut_29[5] , 
        \nLeftOut_29[4] , \nLeftOut_29[3] , \nLeftOut_29[2] , \nLeftOut_29[1] , 
        \nLeftOut_29[0] }), .outleft({\nLeftOut_33[8] , \nLeftOut_33[7] , 
        \nLeftOut_33[6] , \nLeftOut_33[5] , \nLeftOut_33[4] , \nLeftOut_33[3] , 
        \nLeftOut_33[2] , \nLeftOut_33[1] , \nLeftOut_33[0] }), .outright({
        \nRightOut_33[8] , \nRightOut_33[7] , \nRightOut_33[6] , 
        \nRightOut_33[5] , \nRightOut_33[4] , \nRightOut_33[3] , 
        \nRightOut_33[2] , \nRightOut_33[1] , \nRightOut_33[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_12[8] , \nLeftOut_12[7] , 
        \nLeftOut_12[6] , \nLeftOut_12[5] , \nLeftOut_12[4] , \nLeftOut_12[3] , 
        \nLeftOut_12[2] , \nLeftOut_12[1] , \nLeftOut_12[0] }), .inright({
        \nLeftOut_13[8] , \nLeftOut_13[7] , \nLeftOut_13[6] , \nLeftOut_13[5] , 
        \nLeftOut_13[4] , \nLeftOut_13[3] , \nLeftOut_13[2] , \nLeftOut_13[1] , 
        \nLeftOut_13[0] }), .outleft({\nLeftOut_20[8] , \nLeftOut_20[7] , 
        \nLeftOut_20[6] , \nLeftOut_20[5] , \nLeftOut_20[4] , \nLeftOut_20[3] , 
        \nLeftOut_20[2] , \nLeftOut_20[1] , \nLeftOut_20[0] }), .outright({
        \nRightOut_20[8] , \nRightOut_20[7] , \nRightOut_20[6] , 
        \nRightOut_20[5] , \nRightOut_20[4] , \nRightOut_20[3] , 
        \nRightOut_20[2] , \nRightOut_20[1] , \nRightOut_20[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_20[8] , \nLeftOut_20[7] , 
        \nLeftOut_20[6] , \nLeftOut_20[5] , \nLeftOut_20[4] , \nLeftOut_20[3] , 
        \nLeftOut_20[2] , \nLeftOut_20[1] , \nLeftOut_20[0] }), .inright({
        \nLeftOut_22[8] , \nLeftOut_22[7] , \nLeftOut_22[6] , \nLeftOut_22[5] , 
        \nLeftOut_22[4] , \nLeftOut_22[3] , \nLeftOut_22[2] , \nLeftOut_22[1] , 
        \nLeftOut_22[0] }), .outleft({\nLeftOut_28[8] , \nLeftOut_28[7] , 
        \nLeftOut_28[6] , \nLeftOut_28[5] , \nLeftOut_28[4] , \nLeftOut_28[3] , 
        \nLeftOut_28[2] , \nLeftOut_28[1] , \nLeftOut_28[0] }), .outright({
        \nRightOut_28[8] , \nRightOut_28[7] , \nRightOut_28[6] , 
        \nRightOut_28[5] , \nRightOut_28[4] , \nRightOut_28[3] , 
        \nRightOut_28[2] , \nRightOut_28[1] , \nRightOut_28[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink14[7] , \ScanLink14[6] , \ScanLink14[5] , 
        \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , \ScanLink14[1] , 
        \ScanLink14[0] }), .ScanOut({\ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_36[8] , \nRightOut_36[7] , \nRightOut_36[6] , 
        \nRightOut_36[5] , \nRightOut_36[4] , \nRightOut_36[3] , 
        \nRightOut_36[2] , \nRightOut_36[1] , \nRightOut_36[0] }), .inright({
        \nRightOut_37[8] , \nRightOut_37[7] , \nRightOut_37[6] , 
        \nRightOut_37[5] , \nRightOut_37[4] , \nRightOut_37[3] , 
        \nRightOut_37[2] , \nRightOut_37[1] , \nRightOut_37[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_7[8] , \nLeftOut_7[7] , 
        \nLeftOut_7[6] , \nLeftOut_7[5] , \nLeftOut_7[4] , \nLeftOut_7[3] , 
        \nLeftOut_7[2] , \nLeftOut_7[1] , \nLeftOut_7[0] }), .inright({
        \nRightOut_7[8] , \nRightOut_7[7] , \nRightOut_7[6] , \nRightOut_7[5] , 
        \nRightOut_7[4] , \nRightOut_7[3] , \nRightOut_7[2] , \nRightOut_7[1] , 
        \nRightOut_7[0] }), .outleft({\nLeftOut_15[8] , \nLeftOut_15[7] , 
        \nLeftOut_15[6] , \nLeftOut_15[5] , \nLeftOut_15[4] , \nLeftOut_15[3] , 
        \nLeftOut_15[2] , \nLeftOut_15[1] , \nLeftOut_15[0] }), .outright({
        \nRightOut_15[8] , \nRightOut_15[7] , \nRightOut_15[6] , 
        \nRightOut_15[5] , \nRightOut_15[4] , \nRightOut_15[3] , 
        \nRightOut_15[2] , \nRightOut_15[1] , \nRightOut_15[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s2_SCAN1 node_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_21[8] , \nLeftOut_21[7] , 
        \nLeftOut_21[6] , \nLeftOut_21[5] , \nLeftOut_21[4] , \nLeftOut_21[3] , 
        \nLeftOut_21[2] , \nLeftOut_21[1] , \nLeftOut_21[0] }), .inright({
        \nLeftOut_23[8] , \nLeftOut_23[7] , \nLeftOut_23[6] , \nLeftOut_23[5] , 
        \nLeftOut_23[4] , \nLeftOut_23[3] , \nLeftOut_23[2] , \nLeftOut_23[1] , 
        \nLeftOut_23[0] }), .outleft({\nLeftOut_29[8] , \nLeftOut_29[7] , 
        \nLeftOut_29[6] , \nLeftOut_29[5] , \nLeftOut_29[4] , \nLeftOut_29[3] , 
        \nLeftOut_29[2] , \nLeftOut_29[1] , \nLeftOut_29[0] }), .outright({
        \nRightOut_29[8] , \nRightOut_29[7] , \nRightOut_29[6] , 
        \nRightOut_29[5] , \nRightOut_29[4] , \nRightOut_29[3] , 
        \nRightOut_29[2] , \nRightOut_29[1] , \nRightOut_29[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink15[7] , \ScanLink15[6] , \ScanLink15[5] , 
        \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , \ScanLink15[1] , 
        \ScanLink15[0] }), .ScanOut({\ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(\ScanEnable[0] ), 
        .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nRightOut_38[8] , \nRightOut_38[7] , \nRightOut_38[6] , 
        \nRightOut_38[5] , \nRightOut_38[4] , \nRightOut_38[3] , 
        \nRightOut_38[2] , \nRightOut_38[1] , \nRightOut_38[0] }), .inright({
        \nRightOut_39[8] , \nRightOut_39[7] , \nRightOut_39[6] , 
        \nRightOut_39[5] , \nRightOut_39[4] , \nRightOut_39[3] , 
        \nRightOut_39[2] , \nRightOut_39[1] , \nRightOut_39[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_24[8] , \nLeftOut_24[7] , 
        \nLeftOut_24[6] , \nLeftOut_24[5] , \nLeftOut_24[4] , \nLeftOut_24[3] , 
        \nLeftOut_24[2] , \nLeftOut_24[1] , \nLeftOut_24[0] }), .inright({
        \nLeftOut_28[8] , \nLeftOut_28[7] , \nLeftOut_28[6] , \nLeftOut_28[5] , 
        \nLeftOut_28[4] , \nLeftOut_28[3] , \nLeftOut_28[2] , \nLeftOut_28[1] , 
        \nLeftOut_28[0] }), .outleft({\nLeftOut_32[8] , \nLeftOut_32[7] , 
        \nLeftOut_32[6] , \nLeftOut_32[5] , \nLeftOut_32[4] , \nLeftOut_32[3] , 
        \nLeftOut_32[2] , \nLeftOut_32[1] , \nLeftOut_32[0] }), .outright({
        \nRightOut_32[8] , \nRightOut_32[7] , \nRightOut_32[6] , 
        \nRightOut_32[5] , \nRightOut_32[4] , \nRightOut_32[3] , 
        \nRightOut_32[2] , \nRightOut_32[1] , \nRightOut_32[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink6[7] , \ScanLink6[6] , \ScanLink6[5] , 
        \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , \ScanLink6[1] , 
        \ScanLink6[0] }), .ScanOut({\ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_6[8] , \nLeftOut_6[7] , \nLeftOut_6[6] , \nLeftOut_6[5] , 
        \nLeftOut_6[4] , \nLeftOut_6[3] , \nLeftOut_6[2] , \nLeftOut_6[1] , 
        \nLeftOut_6[0] }), .inright({\nRightOut_6[8] , \nRightOut_6[7] , 
        \nRightOut_6[6] , \nRightOut_6[5] , \nRightOut_6[4] , \nRightOut_6[3] , 
        \nRightOut_6[2] , \nRightOut_6[1] , \nRightOut_6[0] }), .outleft({
        \nLeftOut_6[8] , \nLeftOut_6[7] , \nLeftOut_6[6] , \nLeftOut_6[5] , 
        \nLeftOut_6[4] , \nLeftOut_6[3] , \nLeftOut_6[2] , \nLeftOut_6[1] , 
        \nLeftOut_6[0] }), .outright({\nRightOut_6[8] , \nRightOut_6[7] , 
        \nRightOut_6[6] , \nRightOut_6[5] , \nRightOut_6[4] , \nRightOut_6[3] , 
        \nRightOut_6[2] , \nRightOut_6[1] , \nRightOut_6[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s0_SCAN1 node_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_4[8] , \nLeftOut_4[7] , 
        \nLeftOut_4[6] , \nLeftOut_4[5] , \nLeftOut_4[4] , \nLeftOut_4[3] , 
        \nLeftOut_4[2] , \nLeftOut_4[1] , \nLeftOut_4[0] }), .inright({
        \nRightOut_4[8] , \nRightOut_4[7] , \nRightOut_4[6] , \nRightOut_4[5] , 
        \nRightOut_4[4] , \nRightOut_4[3] , \nRightOut_4[2] , \nRightOut_4[1] , 
        \nRightOut_4[0] }), .outleft({\nLeftOut_12[8] , \nLeftOut_12[7] , 
        \nLeftOut_12[6] , \nLeftOut_12[5] , \nLeftOut_12[4] , \nLeftOut_12[3] , 
        \nLeftOut_12[2] , \nLeftOut_12[1] , \nLeftOut_12[0] }), .outright({
        \nRightOut_12[8] , \nRightOut_12[7] , \nRightOut_12[6] , 
        \nRightOut_12[5] , \nRightOut_12[4] , \nRightOut_12[3] , 
        \nRightOut_12[2] , \nRightOut_12[1] , \nRightOut_12[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s6_SCAN1 node_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nRightOut_17[8] , \nRightOut_17[7] , 
        \nRightOut_17[6] , \nRightOut_17[5] , \nRightOut_17[4] , 
        \nRightOut_17[3] , \nRightOut_17[2] , \nRightOut_17[1] , 
        \nRightOut_17[0] }), .inright({\nRightOut_19[8] , \nRightOut_19[7] , 
        \nRightOut_19[6] , \nRightOut_19[5] , \nRightOut_19[4] , 
        \nRightOut_19[3] , \nRightOut_19[2] , \nRightOut_19[1] , 
        \nRightOut_19[0] }), .outleft({\nLeftOut_27[8] , \nLeftOut_27[7] , 
        \nLeftOut_27[6] , \nLeftOut_27[5] , \nLeftOut_27[4] , \nLeftOut_27[3] , 
        \nLeftOut_27[2] , \nLeftOut_27[1] , \nLeftOut_27[0] }), .outright({
        \nRightOut_27[8] , \nRightOut_27[7] , \nRightOut_27[6] , 
        \nRightOut_27[5] , \nRightOut_27[4] , \nRightOut_27[3] , 
        \nRightOut_27[2] , \nRightOut_27[1] , \nRightOut_27[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s3_SCAN1 node_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .ScanEnable(1'b0), .Idl(1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(
        \nEnable[0] ), .inleft({\nLeftOut_27[8] , \nLeftOut_27[7] , 
        \nLeftOut_27[6] , \nLeftOut_27[5] , \nLeftOut_27[4] , \nLeftOut_27[3] , 
        \nLeftOut_27[2] , \nLeftOut_27[1] , \nLeftOut_27[0] }), .inright({
        \nLeftOut_31[8] , \nLeftOut_31[7] , \nLeftOut_31[6] , \nLeftOut_31[5] , 
        \nLeftOut_31[4] , \nLeftOut_31[3] , \nLeftOut_31[2] , \nLeftOut_31[1] , 
        \nLeftOut_31[0] }), .outleft({\nLeftOut_35[8] , \nLeftOut_35[7] , 
        \nLeftOut_35[6] , \nLeftOut_35[5] , \nLeftOut_35[4] , \nLeftOut_35[3] , 
        \nLeftOut_35[2] , \nLeftOut_35[1] , \nLeftOut_35[0] }), .outright({
        \nRightOut_35[8] , \nRightOut_35[7] , \nRightOut_35[6] , 
        \nRightOut_35[5] , \nRightOut_35[4] , \nRightOut_35[3] , 
        \nRightOut_35[2] , \nRightOut_35[1] , \nRightOut_35[0] }) );
    FFT_Node_SIZE8_IDWIDTH1_s17_SCAN1 node_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\ScanLink8[7] , \ScanLink8[6] , \ScanLink8[5] , 
        \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , \ScanLink8[1] , 
        \ScanLink8[0] }), .ScanOut({\ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(\ScanEnable[0] ), .Idl(
        1'b0), .Idr(1'b0), .Ids(1'b0), .Enable(\nEnable[0] ), .inleft({
        \nLeftOut_32[8] , \nLeftOut_32[7] , \nLeftOut_32[6] , \nLeftOut_32[5] , 
        \nLeftOut_32[4] , \nLeftOut_32[3] , \nLeftOut_32[2] , \nLeftOut_32[1] , 
        \nLeftOut_32[0] }), .inright({\nLeftOut_33[8] , \nLeftOut_33[7] , 
        \nLeftOut_33[6] , \nLeftOut_33[5] , \nLeftOut_33[4] , \nLeftOut_33[3] , 
        \nLeftOut_33[2] , \nLeftOut_33[1] , \nLeftOut_33[0] }) );
endmodule

