
module EdgeAux_DW01_add_16_0 ( A, B, CI, SUM, CO );
input  [15:0] A;
input  [15:0] B;
output [15:0] SUM;
input  CI;
output CO;
    wire \carry[15] , \carry[13] , \carry[9] , \carry[4] , \carry[6] , 
        \carry[2] , \carry[14] , \carry[11] , \carry[10] , \carry[12] , 
        \carry[8] , \carry[7] , \carry[3] , \carry[5] , \carry[1] , n1;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(
        \carry[9] ) );
    VMW_FADD U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(
        \carry[8] ) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(
        \carry[10] ) );
    VMW_FADD U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
    VMW_FADD U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
    VMW_FADD U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]) );
    VMW_FADD U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
    VMW_FADD U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
endmodule


module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [9:0] Eid;
input  [9:0] WeightAddr;
input  [15:0] InEdge;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire \Weight[11] , \Weight[6] , \Weight[15] , \Weight[2] , \Weight[0] , 
        \Weight[9] , \Weight[13] , \Weight[4] , \Weight[12] , \Weight[5] , 
        \Weight[1] , \Weight[8] , \Weight[14] , \Weight[3] , \Weight[10] , 
        \Weight[7] , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101, n102, n103, n104, n105, n106;
    VMW_PULLDOWN U15 ( .Z(n106) );
    VMW_AO22 U16 ( .A(\Weight[9] ), .B(n76), .C(WeightData[9]), .D(n77), .Z(
        n96) );
    VMW_AO22 U17 ( .A(\Weight[8] ), .B(n76), .C(WeightData[8]), .D(n77), .Z(
        n97) );
    VMW_AO22 U18 ( .A(\Weight[7] ), .B(n76), .C(WeightData[7]), .D(n77), .Z(
        n98) );
    VMW_AO22 U19 ( .A(\Weight[6] ), .B(n76), .C(WeightData[6]), .D(n77), .Z(
        n99) );
    VMW_AO22 U20 ( .A(\Weight[5] ), .B(n76), .C(WeightData[5]), .D(n77), .Z(
        n100) );
    VMW_AO22 U21 ( .A(\Weight[4] ), .B(n76), .C(WeightData[4]), .D(n77), .Z(
        n101) );
    VMW_AO22 U22 ( .A(\Weight[3] ), .B(n76), .C(WeightData[3]), .D(n77), .Z(
        n102) );
    VMW_AO22 U23 ( .A(\Weight[2] ), .B(n76), .C(WeightData[2]), .D(n77), .Z(
        n103) );
    VMW_AO22 U24 ( .A(\Weight[1] ), .B(n76), .C(WeightData[1]), .D(n77), .Z(
        n104) );
    VMW_AO22 U25 ( .A(\Weight[15] ), .B(n76), .C(WeightData[15]), .D(n77), .Z(
        n90) );
    VMW_AO22 U26 ( .A(\Weight[14] ), .B(n76), .C(WeightData[14]), .D(n77), .Z(
        n91) );
    VMW_AO22 U27 ( .A(\Weight[13] ), .B(n76), .C(WeightData[13]), .D(n77), .Z(
        n92) );
    VMW_AO22 U28 ( .A(\Weight[12] ), .B(n76), .C(WeightData[12]), .D(n77), .Z(
        n93) );
    VMW_AO22 U29 ( .A(\Weight[11] ), .B(n76), .C(WeightData[11]), .D(n77), .Z(
        n94) );
    VMW_AO22 U30 ( .A(\Weight[10] ), .B(n76), .C(WeightData[10]), .D(n77), .Z(
        n95) );
    VMW_AO22 U31 ( .A(\Weight[0] ), .B(n76), .C(WeightData[0]), .D(n77), .Z(
        n105) );
    VMW_AND5 U32 ( .A(n79), .B(n80), .C(n81), .D(n82), .E(n83), .Z(n78) );
    VMW_AND3 U33 ( .A(n85), .B(n86), .C(n87), .Z(n84) );
    VMW_AND4 U34 ( .A(n88), .B(n89), .C(n84), .D(n78), .Z(n77) );
    VMW_XNOR2 U35 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n80) );
    VMW_XNOR2 U36 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n79) );
    VMW_XNOR2 U37 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n81) );
    VMW_XNOR2 U38 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n83) );
    VMW_XNOR2 U39 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n82) );
    VMW_XNOR2 U40 ( .A(WeightAddr[9]), .B(Eid[9]), .Z(n86) );
    VMW_XNOR2 U41 ( .A(WeightAddr[6]), .B(Eid[6]), .Z(n85) );
    VMW_XNOR2 U42 ( .A(WeightAddr[7]), .B(Eid[7]), .Z(n87) );
    VMW_XNOR2 U43 ( .A(WeightAddr[8]), .B(Eid[8]), .Z(n89) );
    VMW_XNOR2 U44 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n88) );
    VMW_INV U45 ( .A(n77), .Z(n76) );
    VMW_FD \Weight_reg[15]  ( .D(n90), .CP(Clk), .Q(\Weight[15] ) );
    VMW_FD \Weight_reg[14]  ( .D(n91), .CP(Clk), .Q(\Weight[14] ) );
    VMW_FD \Weight_reg[13]  ( .D(n92), .CP(Clk), .Q(\Weight[13] ) );
    VMW_FD \Weight_reg[12]  ( .D(n93), .CP(Clk), .Q(\Weight[12] ) );
    VMW_FD \Weight_reg[11]  ( .D(n94), .CP(Clk), .Q(\Weight[11] ) );
    VMW_FD \Weight_reg[10]  ( .D(n95), .CP(Clk), .Q(\Weight[10] ) );
    VMW_FD \Weight_reg[9]  ( .D(n96), .CP(Clk), .Q(\Weight[9] ) );
    VMW_FD \Weight_reg[8]  ( .D(n97), .CP(Clk), .Q(\Weight[8] ) );
    VMW_FD \Weight_reg[7]  ( .D(n98), .CP(Clk), .Q(\Weight[7] ) );
    VMW_FD \Weight_reg[6]  ( .D(n99), .CP(Clk), .Q(\Weight[6] ) );
    VMW_FD \Weight_reg[5]  ( .D(n100), .CP(Clk), .Q(\Weight[5] ) );
    VMW_FD \Weight_reg[4]  ( .D(n101), .CP(Clk), .Q(\Weight[4] ) );
    VMW_FD \Weight_reg[3]  ( .D(n102), .CP(Clk), .Q(\Weight[3] ) );
    VMW_FD \Weight_reg[2]  ( .D(n103), .CP(Clk), .Q(\Weight[2] ) );
    VMW_FD \Weight_reg[1]  ( .D(n104), .CP(Clk), .Q(\Weight[1] ) );
    VMW_FD \Weight_reg[0]  ( .D(n105), .CP(Clk), .Q(\Weight[0] ) );
    EdgeAux_DW01_add_16_0 add_92 ( .A({\Weight[15] , \Weight[14] , 
        \Weight[13] , \Weight[12] , \Weight[11] , \Weight[10] , \Weight[9] , 
        \Weight[8] , \Weight[7] , \Weight[6] , \Weight[5] , \Weight[4] , 
        \Weight[3] , \Weight[2] , \Weight[1] , \Weight[0] }), .B(InEdge), .CI(
        n106), .SUM(OutEdge) );
endmodule


module NodeAux_INDEGREE1_SOURCE1_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , n267, n268, n269, n270, 
        n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n282) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(InEdges[15]), .D(n268), .Z(
        \OutEdge96[15] ) );
    VMW_AO22 U48 ( .A(OutEdge[14]), .B(n267), .C(InEdges[14]), .D(n268), .Z(
        \OutEdge96[14] ) );
    VMW_AO22 U49 ( .A(OutEdge[13]), .B(n267), .C(InEdges[13]), .D(n268), .Z(
        \OutEdge96[13] ) );
    VMW_AO22 U50 ( .A(OutEdge[12]), .B(n267), .C(InEdges[12]), .D(n268), .Z(
        \OutEdge96[12] ) );
    VMW_AO22 U51 ( .A(OutEdge[11]), .B(n267), .C(InEdges[11]), .D(n268), .Z(
        \OutEdge96[11] ) );
    VMW_AO22 U52 ( .A(OutEdge[10]), .B(n267), .C(InEdges[10]), .D(n268), .Z(
        \OutEdge96[10] ) );
    VMW_AO22 U53 ( .A(OutEdge[9]), .B(n267), .C(InEdges[9]), .D(n268), .Z(
        \OutEdge96[9] ) );
    VMW_AO22 U54 ( .A(OutEdge[8]), .B(n267), .C(InEdges[8]), .D(n268), .Z(
        \OutEdge96[8] ) );
    VMW_AO22 U55 ( .A(OutEdge[7]), .B(n267), .C(InEdges[7]), .D(n268), .Z(
        \OutEdge96[7] ) );
    VMW_AO22 U56 ( .A(OutEdge[6]), .B(n267), .C(InEdges[6]), .D(n268), .Z(
        \OutEdge96[6] ) );
    VMW_AO22 U57 ( .A(OutEdge[5]), .B(n267), .C(InEdges[5]), .D(n268), .Z(
        \OutEdge96[5] ) );
    VMW_AO22 U58 ( .A(OutEdge[4]), .B(n267), .C(InEdges[4]), .D(n268), .Z(
        \OutEdge96[4] ) );
    VMW_AO22 U59 ( .A(OutEdge[3]), .B(n267), .C(InEdges[3]), .D(n268), .Z(
        \OutEdge96[3] ) );
    VMW_AO22 U60 ( .A(OutEdge[2]), .B(n267), .C(InEdges[2]), .D(n268), .Z(
        \OutEdge96[2] ) );
    VMW_AO22 U61 ( .A(OutEdge[1]), .B(n267), .C(InEdges[1]), .D(n268), .Z(
        \OutEdge96[1] ) );
    VMW_AO22 U62 ( .A(OutEdge[0]), .B(n267), .C(InEdges[0]), .D(n268), .Z(
        \OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(Start), .B(\path[1] ), .C(n267), .Z(n281) );
    VMW_AO21 U64 ( .A(\path[2] ), .B(Start), .C(n267), .Z(n280) );
    VMW_AO21 U65 ( .A(Start), .B(\path[0] ), .C(n267), .Z(n279) );
    VMW_NOR2 U66 ( .A(n269), .B(Start), .Z(n268) );
    VMW_NOR2 U67 ( .A(Start), .B(n82), .Z(n267) );
    VMW_AND4 U68 ( .A(n271), .B(n272), .C(n273), .D(n274), .Z(n270) );
    VMW_AND4 U69 ( .A(n275), .B(n276), .C(n277), .D(n270), .Z(n278) );
    VMW_XNOR2 U70 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n274) );
    VMW_XNOR2 U71 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n273) );
    VMW_XNOR2 U72 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n272) );
    VMW_XNOR2 U73 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n271) );
    VMW_XNOR2 U74 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n276) );
    VMW_XNOR2 U75 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n275) );
    VMW_XNOR2 U76 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n277) );
    VMW_INV U77 ( .A(n82), .Z(n269) );
    VMW_BUFIZ U78 ( .A(\path[1] ), .E(n278), .Z(\PathData[1] ) );
    VMW_BUFIZ U79 ( .A(\path[0] ), .E(n278), .Z(\PathData[0] ) );
    VMW_BUFIZ U80 ( .A(\path[2] ), .E(n278), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n279), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n280), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n281), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE1_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n282), .TC(n282), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE1_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , n82, \OutEdge96[11] , \OutEdge96[5] , 
        \OutEdge96[15] , \OutEdge96[8] , \OutEdge96[1] , \OutEdge96[3] , 
        \OutEdge96[7] , \OutEdge96[13] , \OutEdge96[6] , \OutEdge96[12] , 
        \OutEdge96[2] , \OutEdge96[9] , \OutEdge96[14] , \OutEdge96[0] , 
        \OutEdge96[10] , \OutEdge96[4] , \path[1] , n267, n268, n269, n270, 
        n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
        n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
        n295, n296, n297;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U46 ( .Z(n297) );
    VMW_AO22 U47 ( .A(OutEdge[15]), .B(n267), .C(n268), .D(InEdges[15]), .Z(
        \OutEdge96[15] ) );
    VMW_OR2 U48 ( .A(n269), .B(Start), .Z(\OutEdge96[14] ) );
    VMW_OR2 U49 ( .A(n270), .B(Start), .Z(\OutEdge96[13] ) );
    VMW_OR2 U50 ( .A(n271), .B(Start), .Z(\OutEdge96[12] ) );
    VMW_OR2 U51 ( .A(n272), .B(Start), .Z(\OutEdge96[11] ) );
    VMW_OR2 U52 ( .A(n273), .B(Start), .Z(\OutEdge96[10] ) );
    VMW_OR2 U53 ( .A(n274), .B(Start), .Z(\OutEdge96[9] ) );
    VMW_OR2 U54 ( .A(n275), .B(Start), .Z(\OutEdge96[8] ) );
    VMW_OR2 U55 ( .A(n276), .B(Start), .Z(\OutEdge96[7] ) );
    VMW_OR2 U56 ( .A(n277), .B(Start), .Z(\OutEdge96[6] ) );
    VMW_OR2 U57 ( .A(n278), .B(Start), .Z(\OutEdge96[5] ) );
    VMW_OR2 U58 ( .A(n279), .B(Start), .Z(\OutEdge96[4] ) );
    VMW_OR2 U59 ( .A(n280), .B(Start), .Z(\OutEdge96[3] ) );
    VMW_OR2 U60 ( .A(n281), .B(Start), .Z(\OutEdge96[2] ) );
    VMW_OR2 U61 ( .A(n282), .B(Start), .Z(\OutEdge96[1] ) );
    VMW_OR2 U62 ( .A(n283), .B(Start), .Z(\OutEdge96[0] ) );
    VMW_AO21 U63 ( .A(\path[1] ), .B(Start), .C(n267), .Z(n296) );
    VMW_AO21 U64 ( .A(Start), .B(\path[2] ), .C(n267), .Z(n295) );
    VMW_AO21 U65 ( .A(\path[0] ), .B(Start), .C(n267), .Z(n294) );
    VMW_INV U66 ( .A(n82), .Z(n284) );
    VMW_NOR2 U67 ( .A(Start), .B(n82), .Z(n267) );
    VMW_AND4 U68 ( .A(n286), .B(n287), .C(n288), .D(n289), .Z(n285) );
    VMW_NOR2 U69 ( .A(Start), .B(n284), .Z(n268) );
    VMW_AND4 U70 ( .A(n290), .B(n291), .C(n292), .D(n285), .Z(n293) );
    VMW_XNOR2 U71 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n289) );
    VMW_XNOR2 U72 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n288) );
    VMW_XNOR2 U73 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n287) );
    VMW_XNOR2 U74 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n286) );
    VMW_XNOR2 U75 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n291) );
    VMW_XNOR2 U76 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n290) );
    VMW_XNOR2 U77 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n292) );
    VMW_AO22 U78 ( .A(InEdges[9]), .B(n82), .C(OutEdge[9]), .D(n284), .Z(n274)
         );
    VMW_AO22 U79 ( .A(InEdges[8]), .B(n82), .C(OutEdge[8]), .D(n284), .Z(n275)
         );
    VMW_AO22 U80 ( .A(InEdges[7]), .B(n82), .C(OutEdge[7]), .D(n284), .Z(n276)
         );
    VMW_AO22 U81 ( .A(InEdges[6]), .B(n82), .C(OutEdge[6]), .D(n284), .Z(n277)
         );
    VMW_AO22 U82 ( .A(InEdges[5]), .B(n82), .C(OutEdge[5]), .D(n284), .Z(n278)
         );
    VMW_AO22 U83 ( .A(InEdges[4]), .B(n82), .C(OutEdge[4]), .D(n284), .Z(n279)
         );
    VMW_AO22 U84 ( .A(InEdges[3]), .B(n82), .C(OutEdge[3]), .D(n284), .Z(n280)
         );
    VMW_AO22 U85 ( .A(InEdges[2]), .B(n82), .C(OutEdge[2]), .D(n284), .Z(n281)
         );
    VMW_AO22 U86 ( .A(InEdges[1]), .B(n82), .C(OutEdge[1]), .D(n284), .Z(n282)
         );
    VMW_AO22 U87 ( .A(InEdges[14]), .B(n82), .C(OutEdge[14]), .D(n284), .Z(
        n269) );
    VMW_AO22 U88 ( .A(InEdges[13]), .B(n82), .C(OutEdge[13]), .D(n284), .Z(
        n270) );
    VMW_AO22 U89 ( .A(InEdges[12]), .B(n82), .C(OutEdge[12]), .D(n284), .Z(
        n271) );
    VMW_AO22 U90 ( .A(InEdges[11]), .B(n82), .C(OutEdge[11]), .D(n284), .Z(
        n272) );
    VMW_AO22 U91 ( .A(InEdges[10]), .B(n82), .C(OutEdge[10]), .D(n284), .Z(
        n273) );
    VMW_AO22 U92 ( .A(InEdges[0]), .B(n82), .C(OutEdge[0]), .D(n284), .Z(n283)
         );
    VMW_BUFIZ U93 ( .A(\path[1] ), .E(n293), .Z(\PathData[1] ) );
    VMW_BUFIZ U94 ( .A(\path[0] ), .E(n293), .Z(\PathData[0] ) );
    VMW_BUFIZ U95 ( .A(\path[2] ), .E(n293), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n294), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n295), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n296), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge96[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge96[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge96[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge96[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge96[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge96[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge96[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge96[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge96[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge96[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge96[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge96[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge96[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge96[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge96[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge96[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE1_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges), 
        .LEQ(n297), .TC(n297), .GE_GT(n82) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n85) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n85), .D(n82), .Z(n86) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n86), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n93) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n93), .D(n90), .Z(n94) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n94), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n96), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n111), .C(n107), .D(n102), .Z(n110) );
    VMW_NAND2 U30 ( .A(n111), .B(A[13]), .Z(n112) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n112), .D(n110), .Z(n113) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n114), .C(n113), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n114) );
    VMW_INV U48 ( .A(B[13]), .Z(n111) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp180[1] , \temp180[8] , \OutEdge106[5] , \temp180[5] , 
        \OutEdge106[8] , \OutEdge106[1] , \path[2] , \path[0] , 
        \OutEdge106[3] , \temp180[7] , \OutEdge106[7] , \temp180[3] , 
        \OutEdge106[13] , \temp180[12] , \temp180[10] , \OutEdge106[11] , 
        \OutEdge106[15] , \temp180[14] , n84, \OutEdge106[14] , \temp180[15] , 
        \temp180[11] , \OutEdge106[10] , \OutEdge106[12] , \temp180[13] , 
        \OutEdge106[6] , \temp180[2] , \path[1] , n92, \OutEdge106[2] , 
        \temp180[6] , \temp180[4] , \OutEdge106[9] , \OutEdge106[0] , 
        \temp180[0] , \temp180[9] , \OutEdge106[4] , n367, n368, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
        n395, n396, n397, n398, n399, n400, n401;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U55 ( .Z(n400) );
    VMW_PULLDOWN U56 ( .Z(n401) );
    VMW_NOR2 U57 ( .A(Start), .B(n367), .Z(\OutEdge106[15] ) );
    VMW_NAND2 U58 ( .A(n368), .B(n369), .Z(\OutEdge106[14] ) );
    VMW_NAND2 U59 ( .A(n370), .B(n369), .Z(\OutEdge106[13] ) );
    VMW_NAND2 U60 ( .A(n371), .B(n369), .Z(\OutEdge106[12] ) );
    VMW_NAND2 U61 ( .A(n372), .B(n369), .Z(\OutEdge106[11] ) );
    VMW_NAND2 U62 ( .A(n373), .B(n369), .Z(\OutEdge106[10] ) );
    VMW_NAND2 U63 ( .A(n374), .B(n369), .Z(\OutEdge106[9] ) );
    VMW_NAND2 U64 ( .A(n375), .B(n369), .Z(\OutEdge106[8] ) );
    VMW_NAND2 U65 ( .A(n376), .B(n369), .Z(\OutEdge106[7] ) );
    VMW_NAND2 U66 ( .A(n377), .B(n369), .Z(\OutEdge106[6] ) );
    VMW_NAND2 U67 ( .A(n378), .B(n369), .Z(\OutEdge106[5] ) );
    VMW_NAND2 U68 ( .A(n379), .B(n369), .Z(\OutEdge106[4] ) );
    VMW_NAND2 U69 ( .A(n380), .B(n369), .Z(\OutEdge106[3] ) );
    VMW_NAND2 U70 ( .A(n381), .B(n369), .Z(\OutEdge106[2] ) );
    VMW_NAND2 U71 ( .A(n382), .B(n369), .Z(\OutEdge106[1] ) );
    VMW_NAND2 U72 ( .A(n383), .B(n369), .Z(\OutEdge106[0] ) );
    VMW_AO21 U73 ( .A(Start), .B(\path[1] ), .C(n384), .Z(n399) );
    VMW_AO21 U74 ( .A(\path[2] ), .B(Start), .C(n384), .Z(n398) );
    VMW_OR2 U75 ( .A(n386), .B(n92), .Z(n385) );
    VMW_AO22 U76 ( .A(OutEdge[15]), .B(n386), .C(InEdges[15]), .D(n84), .Z(
        \temp180[15] ) );
    VMW_OAI22 U77 ( .A(\path[0] ), .B(n369), .C(n385), .D(Start), .Z(n387) );
    VMW_MUX2I U78 ( .A(\temp180[15] ), .B(InEdges[31]), .S(n92), .Z(n367) );
    VMW_AND4 U79 ( .A(n389), .B(n390), .C(n391), .D(n392), .Z(n388) );
    VMW_NOR3 U80 ( .A(Start), .B(n84), .C(n92), .Z(n384) );
    VMW_AND4 U81 ( .A(n393), .B(n394), .C(n395), .D(n388), .Z(n396) );
    VMW_XNOR2 U82 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n392) );
    VMW_XNOR2 U83 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n391) );
    VMW_XNOR2 U84 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n390) );
    VMW_XNOR2 U85 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n389) );
    VMW_XNOR2 U86 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n394) );
    VMW_XNOR2 U87 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n393) );
    VMW_XNOR2 U88 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n395) );
    VMW_AO22 U89 ( .A(OutEdge[9]), .B(n386), .C(InEdges[9]), .D(n84), .Z(
        \temp180[9] ) );
    VMW_AO22 U90 ( .A(OutEdge[8]), .B(n386), .C(InEdges[8]), .D(n84), .Z(
        \temp180[8] ) );
    VMW_AO22 U91 ( .A(OutEdge[7]), .B(n386), .C(InEdges[7]), .D(n84), .Z(
        \temp180[7] ) );
    VMW_AO22 U92 ( .A(OutEdge[6]), .B(n386), .C(InEdges[6]), .D(n84), .Z(
        \temp180[6] ) );
    VMW_AO22 U93 ( .A(OutEdge[5]), .B(n386), .C(InEdges[5]), .D(n84), .Z(
        \temp180[5] ) );
    VMW_AO22 U94 ( .A(OutEdge[4]), .B(n386), .C(InEdges[4]), .D(n84), .Z(
        \temp180[4] ) );
    VMW_AO22 U95 ( .A(OutEdge[3]), .B(n386), .C(InEdges[3]), .D(n84), .Z(
        \temp180[3] ) );
    VMW_AO22 U96 ( .A(OutEdge[2]), .B(n386), .C(InEdges[2]), .D(n84), .Z(
        \temp180[2] ) );
    VMW_AO22 U97 ( .A(OutEdge[1]), .B(n386), .C(InEdges[1]), .D(n84), .Z(
        \temp180[1] ) );
    VMW_AO22 U98 ( .A(OutEdge[14]), .B(n386), .C(InEdges[14]), .D(n84), .Z(
        \temp180[14] ) );
    VMW_AO22 U99 ( .A(OutEdge[13]), .B(n386), .C(InEdges[13]), .D(n84), .Z(
        \temp180[13] ) );
    VMW_AO22 U100 ( .A(OutEdge[12]), .B(n386), .C(InEdges[12]), .D(n84), .Z(
        \temp180[12] ) );
    VMW_AO22 U101 ( .A(OutEdge[11]), .B(n386), .C(InEdges[11]), .D(n84), .Z(
        \temp180[11] ) );
    VMW_AO22 U102 ( .A(OutEdge[10]), .B(n386), .C(InEdges[10]), .D(n84), .Z(
        \temp180[10] ) );
    VMW_AO22 U103 ( .A(OutEdge[0]), .B(n386), .C(InEdges[0]), .D(n84), .Z(
        \temp180[0] ) );
    VMW_MUX2I U104 ( .A(\temp180[9] ), .B(InEdges[25]), .S(n92), .Z(n374) );
    VMW_MUX2I U105 ( .A(\temp180[8] ), .B(InEdges[24]), .S(n92), .Z(n375) );
    VMW_MUX2I U106 ( .A(\temp180[7] ), .B(InEdges[23]), .S(n92), .Z(n376) );
    VMW_MUX2I U107 ( .A(\temp180[6] ), .B(InEdges[22]), .S(n92), .Z(n377) );
    VMW_MUX2I U108 ( .A(\temp180[5] ), .B(InEdges[21]), .S(n92), .Z(n378) );
    VMW_MUX2I U109 ( .A(\temp180[4] ), .B(InEdges[20]), .S(n92), .Z(n379) );
    VMW_MUX2I U110 ( .A(\temp180[3] ), .B(InEdges[19]), .S(n92), .Z(n380) );
    VMW_MUX2I U111 ( .A(\temp180[2] ), .B(InEdges[18]), .S(n92), .Z(n381) );
    VMW_MUX2I U112 ( .A(\temp180[1] ), .B(InEdges[17]), .S(n92), .Z(n382) );
    VMW_MUX2I U113 ( .A(\temp180[14] ), .B(InEdges[30]), .S(n92), .Z(n368) );
    VMW_MUX2I U114 ( .A(\temp180[13] ), .B(InEdges[29]), .S(n92), .Z(n370) );
    VMW_MUX2I U115 ( .A(\temp180[12] ), .B(InEdges[28]), .S(n92), .Z(n371) );
    VMW_MUX2I U116 ( .A(\temp180[11] ), .B(InEdges[27]), .S(n92), .Z(n372) );
    VMW_MUX2I U117 ( .A(\temp180[10] ), .B(InEdges[26]), .S(n92), .Z(n373) );
    VMW_MUX2I U118 ( .A(\temp180[0] ), .B(InEdges[16]), .S(n92), .Z(n383) );
    VMW_INV U119 ( .A(n84), .Z(n386) );
    VMW_INV U120 ( .A(Start), .Z(n369) );
    VMW_INV U121 ( .A(n387), .Z(n397) );
    VMW_BUFIZ U122 ( .A(\path[1] ), .E(n396), .Z(\PathData[1] ) );
    VMW_BUFIZ U123 ( .A(\path[0] ), .E(n396), .Z(\PathData[0] ) );
    VMW_BUFIZ U124 ( .A(\path[2] ), .E(n396), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n397), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n398), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n399), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge106[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge106[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge106[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge106[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge106[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge106[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge106[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge106[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge106[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge106[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge106[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge106[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge106[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge106[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge106[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge106[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n401), .TC(n401), .GE_GT(n84) );
    NodeAux_INDEGREE2_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp180[15] , 
        \temp180[14] , \temp180[13] , \temp180[12] , \temp180[11] , 
        \temp180[10] , \temp180[9] , \temp180[8] , \temp180[7] , \temp180[6] , 
        \temp180[5] , \temp180[4] , \temp180[3] , \temp180[2] , \temp180[1] , 
        \temp180[0] }), .B(InEdges[31:16]), .LEQ(n400), .TC(n400), .GE_GT(n92)
         );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, 
        n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, 
        n108, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n87), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n95), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n96) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n88), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n104), .B(B[12]), .Z(n103) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n96), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n104), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n103), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n104) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n95) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n87) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
        n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n119), .B(B[2]), .Z(n118) );
    VMW_AO22 U5 ( .A(n121), .B(B[0]), .C(n122), .D(B[1]), .Z(n120) );
    VMW_OR2 U6 ( .A(B[2]), .B(n119), .Z(n123) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n122), .C(n123), .D(n120), .Z(n124) );
    VMW_NAND2 U8 ( .A(n126), .B(B[4]), .Z(n125) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n128), .C(n124), .D(n118), .Z(n127) );
    VMW_OR2 U10 ( .A(B[4]), .B(n126), .Z(n129) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n131), .C(n129), .D(n127), .Z(n130) );
    VMW_NAND2 U12 ( .A(n133), .B(B[6]), .Z(n132) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n135), .C(n130), .D(n125), .Z(n134) );
    VMW_OR2 U14 ( .A(B[6]), .B(n133), .Z(n136) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n138), .C(n136), .D(n134), .Z(n137) );
    VMW_NAND2 U16 ( .A(n140), .B(B[8]), .Z(n139) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n142), .C(n137), .D(n132), .Z(n141) );
    VMW_OR2 U18 ( .A(B[8]), .B(n140), .Z(n143) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n145), .C(n143), .D(n141), .Z(n144) );
    VMW_NAND2 U20 ( .A(n147), .B(B[10]), .Z(n146) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n149), .C(n144), .D(n139), .Z(n148) );
    VMW_NAND2 U22 ( .A(n149), .B(A[9]), .Z(n150) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n147), .C(n150), .D(n148), .Z(n151) );
    VMW_NAND2 U24 ( .A(n153), .B(B[12]), .Z(n152) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n155), .C(n151), .D(n146), .Z(n154) );
    VMW_NAND2 U26 ( .A(n155), .B(A[11]), .Z(n156) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n153), .C(n156), .D(n154), .Z(n157) );
    VMW_NAND2 U28 ( .A(n159), .B(B[14]), .Z(n158) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n161), .C(n157), .D(n152), .Z(n160) );
    VMW_NAND2 U30 ( .A(n161), .B(A[13]), .Z(n162) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n159), .C(n162), .D(n160), .Z(n163) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n164), .C(n163), .D(n158), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n153) );
    VMW_INV U34 ( .A(B[7]), .Z(n142) );
    VMW_INV U35 ( .A(A[7]), .Z(n145) );
    VMW_INV U36 ( .A(A[3]), .Z(n131) );
    VMW_INV U37 ( .A(B[3]), .Z(n128) );
    VMW_INV U38 ( .A(A[10]), .Z(n147) );
    VMW_INV U39 ( .A(B[9]), .Z(n149) );
    VMW_INV U40 ( .A(A[4]), .Z(n126) );
    VMW_INV U41 ( .A(A[8]), .Z(n140) );
    VMW_INV U42 ( .A(A[14]), .Z(n159) );
    VMW_INV U43 ( .A(B[11]), .Z(n155) );
    VMW_INV U44 ( .A(A[5]), .Z(n138) );
    VMW_INV U45 ( .A(B[5]), .Z(n135) );
    VMW_INV U46 ( .A(A[1]), .Z(n122) );
    VMW_INV U47 ( .A(B[15]), .Z(n164) );
    VMW_INV U48 ( .A(B[13]), .Z(n161) );
    VMW_INV U49 ( .A(A[6]), .Z(n133) );
    VMW_INV U50 ( .A(A[2]), .Z(n119) );
    VMW_INV U51 ( .A(A[0]), .Z(n121) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp284[0] , \OutEdge116[6] , \temp284[9] , \temp284[11] , 
        \temp190[2] , \OutEdge116[2] , \temp284[4] , \temp190[6] , 
        \temp284[15] , \path[2] , \OutEdge116[9] , \path[0] , \temp190[4] , 
        \OutEdge116[0] , \temp284[6] , \temp284[13] , \temp190[0] , 
        \temp284[2] , \OutEdge116[4] , \temp190[9] , \temp190[10] , 
        \OutEdge116[11] , \OutEdge116[15] , \temp190[14] , \OutEdge116[13] , 
        \temp190[12] , n94, \OutEdge116[12] , \temp190[13] , n86, 
        \OutEdge116[14] , \temp190[15] , \temp190[11] , \OutEdge116[10] , 
        \temp284[12] , \temp190[1] , \temp284[3] , \OutEdge116[5] , 
        \temp190[8] , \path[1] , \OutEdge116[8] , \temp190[5] , 
        \OutEdge116[1] , \temp284[7] , n102, \OutEdge116[3] , \temp284[5] , 
        \temp190[7] , \temp284[14] , \temp284[1] , \OutEdge116[7] , 
        \temp284[8] , \temp284[10] , \temp190[3] , n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U64 ( .Z(n504) );
    VMW_PULLDOWN U65 ( .Z(n506) );
    VMW_PULLDOWN U66 ( .Z(n505) );
    VMW_AND2 U67 ( .A(n467), .B(n468), .Z(\OutEdge116[15] ) );
    VMW_OR2 U68 ( .A(n469), .B(Start), .Z(\OutEdge116[14] ) );
    VMW_OR2 U69 ( .A(n470), .B(Start), .Z(\OutEdge116[13] ) );
    VMW_OR2 U70 ( .A(n471), .B(Start), .Z(\OutEdge116[12] ) );
    VMW_OR2 U71 ( .A(n472), .B(Start), .Z(\OutEdge116[11] ) );
    VMW_OR2 U72 ( .A(n473), .B(Start), .Z(\OutEdge116[10] ) );
    VMW_OR2 U73 ( .A(n474), .B(Start), .Z(\OutEdge116[9] ) );
    VMW_OR2 U74 ( .A(n475), .B(Start), .Z(\OutEdge116[8] ) );
    VMW_OR2 U75 ( .A(n476), .B(Start), .Z(\OutEdge116[7] ) );
    VMW_OR2 U76 ( .A(n477), .B(Start), .Z(\OutEdge116[6] ) );
    VMW_OR2 U77 ( .A(n478), .B(Start), .Z(\OutEdge116[5] ) );
    VMW_OR2 U78 ( .A(n479), .B(Start), .Z(\OutEdge116[4] ) );
    VMW_OR2 U79 ( .A(n480), .B(Start), .Z(\OutEdge116[3] ) );
    VMW_OR2 U80 ( .A(n481), .B(Start), .Z(\OutEdge116[2] ) );
    VMW_OR2 U81 ( .A(n482), .B(Start), .Z(\OutEdge116[1] ) );
    VMW_OR2 U82 ( .A(n483), .B(Start), .Z(\OutEdge116[0] ) );
    VMW_OR2 U83 ( .A(n484), .B(n485), .Z(n503) );
    VMW_AO22 U84 ( .A(\path[2] ), .B(Start), .C(n486), .D(n485), .Z(n502) );
    VMW_AO22 U85 ( .A(\temp190[15] ), .B(n487), .C(InEdges[31]), .D(n94), .Z(
        \temp284[15] ) );
    VMW_AND3 U86 ( .A(n467), .B(n488), .C(n487), .Z(n485) );
    VMW_INV U87 ( .A(Start), .Z(n467) );
    VMW_AO22 U88 ( .A(n490), .B(n467), .C(n491), .D(Start), .Z(n489) );
    VMW_AO22 U89 ( .A(\temp284[15] ), .B(n486), .C(InEdges[47]), .D(n102), .Z(
        n468) );
    VMW_AND4 U90 ( .A(n493), .B(n494), .C(n495), .D(n496), .Z(n492) );
    VMW_INV U91 ( .A(n102), .Z(n486) );
    VMW_AND4 U92 ( .A(n497), .B(n498), .C(n499), .D(n492), .Z(n500) );
    VMW_XNOR2 U93 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n496) );
    VMW_XNOR2 U94 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n495) );
    VMW_XNOR2 U95 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n494) );
    VMW_XNOR2 U96 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n493) );
    VMW_XNOR2 U97 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n498) );
    VMW_XNOR2 U98 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n497) );
    VMW_XNOR2 U99 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n499) );
    VMW_AO22 U100 ( .A(InEdges[9]), .B(n86), .C(OutEdge[9]), .D(n488), .Z(
        \temp190[9] ) );
    VMW_AO22 U101 ( .A(\temp190[9] ), .B(n487), .C(InEdges[25]), .D(n94), .Z(
        \temp284[9] ) );
    VMW_AO22 U102 ( .A(InEdges[8]), .B(n86), .C(OutEdge[8]), .D(n488), .Z(
        \temp190[8] ) );
    VMW_AO22 U103 ( .A(\temp190[8] ), .B(n487), .C(InEdges[24]), .D(n94), .Z(
        \temp284[8] ) );
    VMW_AO22 U104 ( .A(InEdges[7]), .B(n86), .C(OutEdge[7]), .D(n488), .Z(
        \temp190[7] ) );
    VMW_AO22 U105 ( .A(\temp190[7] ), .B(n487), .C(InEdges[23]), .D(n94), .Z(
        \temp284[7] ) );
    VMW_AO22 U106 ( .A(InEdges[6]), .B(n86), .C(OutEdge[6]), .D(n488), .Z(
        \temp190[6] ) );
    VMW_AO22 U107 ( .A(\temp190[6] ), .B(n487), .C(InEdges[22]), .D(n94), .Z(
        \temp284[6] ) );
    VMW_AO22 U108 ( .A(InEdges[5]), .B(n86), .C(OutEdge[5]), .D(n488), .Z(
        \temp190[5] ) );
    VMW_AO22 U109 ( .A(\temp190[5] ), .B(n487), .C(InEdges[21]), .D(n94), .Z(
        \temp284[5] ) );
    VMW_AO22 U110 ( .A(InEdges[4]), .B(n86), .C(OutEdge[4]), .D(n488), .Z(
        \temp190[4] ) );
    VMW_AO22 U111 ( .A(\temp190[4] ), .B(n487), .C(InEdges[20]), .D(n94), .Z(
        \temp284[4] ) );
    VMW_AO22 U112 ( .A(InEdges[3]), .B(n86), .C(OutEdge[3]), .D(n488), .Z(
        \temp190[3] ) );
    VMW_AO22 U113 ( .A(\temp190[3] ), .B(n487), .C(InEdges[19]), .D(n94), .Z(
        \temp284[3] ) );
    VMW_AO22 U114 ( .A(InEdges[2]), .B(n86), .C(OutEdge[2]), .D(n488), .Z(
        \temp190[2] ) );
    VMW_AO22 U115 ( .A(\temp190[2] ), .B(n487), .C(InEdges[18]), .D(n94), .Z(
        \temp284[2] ) );
    VMW_AO22 U116 ( .A(InEdges[1]), .B(n86), .C(OutEdge[1]), .D(n488), .Z(
        \temp190[1] ) );
    VMW_AO22 U117 ( .A(\temp190[1] ), .B(n487), .C(InEdges[17]), .D(n94), .Z(
        \temp284[1] ) );
    VMW_AO22 U118 ( .A(InEdges[15]), .B(n86), .C(OutEdge[15]), .D(n488), .Z(
        \temp190[15] ) );
    VMW_AO22 U119 ( .A(InEdges[14]), .B(n86), .C(OutEdge[14]), .D(n488), .Z(
        \temp190[14] ) );
    VMW_AO22 U120 ( .A(\temp190[14] ), .B(n487), .C(InEdges[30]), .D(n94), .Z(
        \temp284[14] ) );
    VMW_AO22 U121 ( .A(InEdges[13]), .B(n86), .C(OutEdge[13]), .D(n488), .Z(
        \temp190[13] ) );
    VMW_AO22 U122 ( .A(\temp190[13] ), .B(n487), .C(InEdges[29]), .D(n94), .Z(
        \temp284[13] ) );
    VMW_AO22 U123 ( .A(InEdges[12]), .B(n86), .C(OutEdge[12]), .D(n488), .Z(
        \temp190[12] ) );
    VMW_AO22 U124 ( .A(\temp190[12] ), .B(n487), .C(InEdges[28]), .D(n94), .Z(
        \temp284[12] ) );
    VMW_AO22 U125 ( .A(InEdges[11]), .B(n86), .C(OutEdge[11]), .D(n488), .Z(
        \temp190[11] ) );
    VMW_AO22 U126 ( .A(\temp190[11] ), .B(n487), .C(InEdges[27]), .D(n94), .Z(
        \temp284[11] ) );
    VMW_AO22 U127 ( .A(InEdges[10]), .B(n86), .C(OutEdge[10]), .D(n488), .Z(
        \temp190[10] ) );
    VMW_AO22 U128 ( .A(\temp190[10] ), .B(n487), .C(InEdges[26]), .D(n94), .Z(
        \temp284[10] ) );
    VMW_AO22 U129 ( .A(InEdges[0]), .B(n86), .C(OutEdge[0]), .D(n488), .Z(
        \temp190[0] ) );
    VMW_AO22 U130 ( .A(\temp190[0] ), .B(n487), .C(InEdges[16]), .D(n94), .Z(
        \temp284[0] ) );
    VMW_AO22 U131 ( .A(\path[1] ), .B(Start), .C(n102), .D(n467), .Z(n484) );
    VMW_AO21 U132 ( .A(n487), .B(n86), .C(n102), .Z(n490) );
    VMW_AO22 U133 ( .A(\temp284[9] ), .B(n486), .C(InEdges[41]), .D(n102), .Z(
        n474) );
    VMW_AO22 U134 ( .A(\temp284[8] ), .B(n486), .C(InEdges[40]), .D(n102), .Z(
        n475) );
    VMW_AO22 U135 ( .A(\temp284[7] ), .B(n486), .C(InEdges[39]), .D(n102), .Z(
        n476) );
    VMW_AO22 U136 ( .A(\temp284[6] ), .B(n486), .C(InEdges[38]), .D(n102), .Z(
        n477) );
    VMW_AO22 U137 ( .A(\temp284[5] ), .B(n486), .C(InEdges[37]), .D(n102), .Z(
        n478) );
    VMW_AO22 U138 ( .A(\temp284[4] ), .B(n486), .C(InEdges[36]), .D(n102), .Z(
        n479) );
    VMW_AO22 U139 ( .A(\temp284[3] ), .B(n486), .C(InEdges[35]), .D(n102), .Z(
        n480) );
    VMW_AO22 U140 ( .A(\temp284[2] ), .B(n486), .C(InEdges[34]), .D(n102), .Z(
        n481) );
    VMW_AO22 U141 ( .A(\temp284[1] ), .B(n486), .C(InEdges[33]), .D(n102), .Z(
        n482) );
    VMW_AO22 U142 ( .A(\temp284[14] ), .B(n486), .C(InEdges[46]), .D(n102), 
        .Z(n469) );
    VMW_AO22 U143 ( .A(\temp284[13] ), .B(n486), .C(InEdges[45]), .D(n102), 
        .Z(n470) );
    VMW_AO22 U144 ( .A(\temp284[12] ), .B(n486), .C(InEdges[44]), .D(n102), 
        .Z(n471) );
    VMW_AO22 U145 ( .A(\temp284[11] ), .B(n486), .C(InEdges[43]), .D(n102), 
        .Z(n472) );
    VMW_AO22 U146 ( .A(\temp284[10] ), .B(n486), .C(InEdges[42]), .D(n102), 
        .Z(n473) );
    VMW_AO22 U147 ( .A(\temp284[0] ), .B(n486), .C(InEdges[32]), .D(n102), .Z(
        n483) );
    VMW_INV U148 ( .A(n86), .Z(n488) );
    VMW_INV U149 ( .A(n94), .Z(n487) );
    VMW_INV U150 ( .A(n489), .Z(n501) );
    VMW_INV U151 ( .A(\path[0] ), .Z(n491) );
    VMW_BUFIZ U152 ( .A(\path[1] ), .E(n500), .Z(\PathData[1] ) );
    VMW_BUFIZ U153 ( .A(\path[0] ), .E(n500), .Z(\PathData[0] ) );
    VMW_BUFIZ U154 ( .A(\path[2] ), .E(n500), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n501), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n502), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n503), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge116[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge116[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge116[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge116[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge116[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge116[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge116[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge116[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge116[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge116[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge116[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge116[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge116[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge116[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge116[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge116[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp190[15] , 
        \temp190[14] , \temp190[13] , \temp190[12] , \temp190[11] , 
        \temp190[10] , \temp190[9] , \temp190[8] , \temp190[7] , \temp190[6] , 
        \temp190[5] , \temp190[4] , \temp190[3] , \temp190[2] , \temp190[1] , 
        \temp190[0] }), .B(InEdges[31:16]), .LEQ(n506), .TC(n506), .GE_GT(n94)
         );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_1 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n505), .TC(n505), .GE_GT(n86) );
    NodeAux_INDEGREE3_SOURCE0_DW01_cmp2_16_0 lte_55_2 ( .A({\temp284[15] , 
        \temp284[14] , \temp284[13] , \temp284[12] , \temp284[11] , 
        \temp284[10] , \temp284[9] , \temp284[8] , \temp284[7] , \temp284[6] , 
        \temp284[5] , \temp284[4] , \temp284[3] , \temp284[2] , \temp284[1] , 
        \temp284[0] }), .B(InEdges[47:32]), .LEQ(n504), .TC(n504), .GE_GT(n102
        ) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, 
        n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, 
        n108, n109, n110, n111, n113, n114, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n89), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n90) );
    VMW_OR2 U18 ( .A(B[8]), .B(n89), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n90), .Z(n93) );
    VMW_NAND2 U20 ( .A(n97), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n98) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n97), .C(n100), .D(n98), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n106), .C(n101), .D(n95), .Z(n105) );
    VMW_NAND2 U26 ( .A(n106), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n105), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n113), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n113), .B(A[13]), .Z(n114) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n114), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n97) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n89) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n106) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n113) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n127), .B(B[4]), .Z(n126) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n129), .C(n125), .D(n119), .Z(n128) );
    VMW_OR2 U10 ( .A(B[4]), .B(n127), .Z(n130) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n132), .C(n130), .D(n128), .Z(n131) );
    VMW_NAND2 U12 ( .A(n134), .B(B[6]), .Z(n133) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n136), .C(n131), .D(n126), .Z(n135) );
    VMW_OR2 U14 ( .A(B[6]), .B(n134), .Z(n137) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n139), .C(n137), .D(n135), .Z(n138) );
    VMW_NAND2 U16 ( .A(n141), .B(B[8]), .Z(n140) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n143), .C(n138), .D(n133), .Z(n142) );
    VMW_OR2 U18 ( .A(B[8]), .B(n141), .Z(n144) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n146), .C(n144), .D(n142), .Z(n145) );
    VMW_NAND2 U20 ( .A(n148), .B(B[10]), .Z(n147) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n150), .C(n145), .D(n140), .Z(n149) );
    VMW_NAND2 U22 ( .A(n150), .B(A[9]), .Z(n151) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n148), .C(n151), .D(n149), .Z(n152) );
    VMW_NAND2 U24 ( .A(n154), .B(B[12]), .Z(n153) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n156), .C(n152), .D(n147), .Z(n155) );
    VMW_NAND2 U26 ( .A(n156), .B(A[11]), .Z(n157) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n154), .C(n157), .D(n155), .Z(n158) );
    VMW_NAND2 U28 ( .A(n160), .B(B[14]), .Z(n159) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n162), .C(n158), .D(n153), .Z(n161) );
    VMW_NAND2 U30 ( .A(n162), .B(A[13]), .Z(n163) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n160), .C(n163), .D(n161), .Z(n164) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n165), .C(n164), .D(n159), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n154) );
    VMW_INV U34 ( .A(B[7]), .Z(n143) );
    VMW_INV U35 ( .A(A[7]), .Z(n146) );
    VMW_INV U36 ( .A(A[3]), .Z(n132) );
    VMW_INV U37 ( .A(B[3]), .Z(n129) );
    VMW_INV U38 ( .A(A[10]), .Z(n148) );
    VMW_INV U39 ( .A(B[9]), .Z(n150) );
    VMW_INV U40 ( .A(A[4]), .Z(n127) );
    VMW_INV U41 ( .A(A[8]), .Z(n141) );
    VMW_INV U42 ( .A(A[14]), .Z(n160) );
    VMW_INV U43 ( .A(B[11]), .Z(n156) );
    VMW_INV U44 ( .A(A[5]), .Z(n139) );
    VMW_INV U45 ( .A(B[5]), .Z(n136) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n165) );
    VMW_INV U48 ( .A(B[13]), .Z(n162) );
    VMW_INV U49 ( .A(A[6]), .Z(n134) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
        n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
        n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
        n213, n214;
    VMW_OAI21 U3 ( .A(B[15]), .B(n166), .C(n167), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n169), .B(B[2]), .Z(n168) );
    VMW_AO22 U5 ( .A(n171), .B(B[0]), .C(n172), .D(B[1]), .Z(n170) );
    VMW_OR2 U6 ( .A(B[2]), .B(n169), .Z(n173) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n172), .C(n173), .D(n170), .Z(n174) );
    VMW_NAND2 U8 ( .A(n176), .B(B[4]), .Z(n175) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n178), .C(n174), .D(n168), .Z(n177) );
    VMW_OR2 U10 ( .A(B[4]), .B(n176), .Z(n179) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n181), .C(n179), .D(n177), .Z(n180) );
    VMW_NAND2 U12 ( .A(n183), .B(B[6]), .Z(n182) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n185), .C(n180), .D(n175), .Z(n184) );
    VMW_OR2 U14 ( .A(B[6]), .B(n183), .Z(n186) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n188), .C(n186), .D(n184), .Z(n187) );
    VMW_NAND2 U16 ( .A(n190), .B(B[8]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n192), .C(n187), .D(n182), .Z(n191) );
    VMW_OR2 U18 ( .A(B[8]), .B(n190), .Z(n193) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n195), .C(n193), .D(n191), .Z(n194) );
    VMW_NAND2 U20 ( .A(n197), .B(B[10]), .Z(n196) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n199), .C(n194), .D(n189), .Z(n198) );
    VMW_NAND2 U22 ( .A(n199), .B(A[9]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n197), .C(n200), .D(n198), .Z(n201) );
    VMW_NAND2 U24 ( .A(n203), .B(B[12]), .Z(n202) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n205), .C(n201), .D(n196), .Z(n204) );
    VMW_NAND2 U26 ( .A(n205), .B(A[11]), .Z(n206) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n203), .C(n206), .D(n204), .Z(n207) );
    VMW_NAND2 U28 ( .A(n209), .B(B[14]), .Z(n208) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n211), .C(n207), .D(n202), .Z(n210) );
    VMW_NAND2 U30 ( .A(n211), .B(A[13]), .Z(n212) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n209), .C(n212), .D(n210), .Z(n213) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n214), .C(n213), .D(n208), .Z(n167) );
    VMW_INV U33 ( .A(A[12]), .Z(n203) );
    VMW_INV U34 ( .A(B[7]), .Z(n192) );
    VMW_INV U35 ( .A(A[7]), .Z(n195) );
    VMW_INV U36 ( .A(A[3]), .Z(n181) );
    VMW_INV U37 ( .A(B[3]), .Z(n178) );
    VMW_INV U38 ( .A(A[10]), .Z(n197) );
    VMW_INV U39 ( .A(B[9]), .Z(n199) );
    VMW_INV U40 ( .A(A[4]), .Z(n176) );
    VMW_INV U41 ( .A(A[8]), .Z(n190) );
    VMW_INV U42 ( .A(A[14]), .Z(n209) );
    VMW_INV U43 ( .A(B[11]), .Z(n205) );
    VMW_INV U44 ( .A(A[5]), .Z(n188) );
    VMW_INV U45 ( .A(B[5]), .Z(n185) );
    VMW_INV U46 ( .A(A[1]), .Z(n172) );
    VMW_INV U47 ( .A(B[15]), .Z(n214) );
    VMW_INV U48 ( .A(B[13]), .Z(n211) );
    VMW_INV U49 ( .A(A[6]), .Z(n183) );
    VMW_INV U50 ( .A(A[2]), .Z(n169) );
    VMW_INV U51 ( .A(A[0]), .Z(n171) );
    VMW_INV U52 ( .A(A[15]), .Z(n166) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp200[0] , \temp384[15] , \OutEdge126[12] , \temp200[15] , 
        \temp200[9] , \temp384[6] , \temp294[3] , n112, \temp294[13] , 
        \temp384[11] , \temp200[4] , \temp294[7] , \temp384[2] , \path[2] , 
        \temp200[11] , \temp200[13] , \path[0] , \temp294[5] , \temp384[0] , 
        \temp384[13] , \temp200[6] , \temp384[9] , \OutEdge126[14] , 
        \temp294[11] , \temp384[4] , \temp294[1] , \OutEdge126[10] , 
        \temp294[15] , \temp200[2] , \temp294[8] , \OutEdge126[8] , 
        \OutEdge126[1] , \OutEdge126[5] , n96, \OutEdge126[7] , 
        \OutEdge126[3] , \OutEdge126[2] , \OutEdge126[6] , \OutEdge126[4] , 
        n104, \OutEdge126[9] , n88, \OutEdge126[0] , \temp384[5] , 
        \temp294[0] , \OutEdge126[11] , \temp294[14] , \temp200[3] , 
        \temp294[9] , \path[1] , \temp200[12] , \temp294[4] , \temp384[1] , 
        \temp384[12] , \temp384[8] , \temp200[7] , \OutEdge126[15] , 
        \temp294[10] , \temp294[12] , \temp384[10] , \temp200[5] , 
        \temp294[6] , \temp384[3] , \temp200[10] , \temp200[1] , \temp384[14] , 
        \OutEdge126[13] , \temp200[14] , \temp384[7] , \temp200[8] , 
        \temp294[2] , n567, n568, n569, n570, n571, n572, n573, n574, n575, 
        n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
        n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
        n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U73 ( .Z(n607) );
    VMW_PULLDOWN U74 ( .Z(n608) );
    VMW_PULLDOWN U75 ( .Z(n609) );
    VMW_PULLDOWN U76 ( .Z(n610) );
    VMW_NOR2 U77 ( .A(Start), .B(n567), .Z(\OutEdge126[15] ) );
    VMW_NAND2 U78 ( .A(n568), .B(n569), .Z(\OutEdge126[14] ) );
    VMW_NAND2 U79 ( .A(n570), .B(n569), .Z(\OutEdge126[13] ) );
    VMW_NAND2 U80 ( .A(n571), .B(n569), .Z(\OutEdge126[12] ) );
    VMW_NAND2 U81 ( .A(n572), .B(n569), .Z(\OutEdge126[11] ) );
    VMW_NAND2 U82 ( .A(n573), .B(n569), .Z(\OutEdge126[10] ) );
    VMW_NAND2 U83 ( .A(n574), .B(n569), .Z(\OutEdge126[9] ) );
    VMW_NAND2 U84 ( .A(n575), .B(n569), .Z(\OutEdge126[8] ) );
    VMW_NAND2 U85 ( .A(n576), .B(n569), .Z(\OutEdge126[7] ) );
    VMW_NAND2 U86 ( .A(n577), .B(n569), .Z(\OutEdge126[6] ) );
    VMW_NAND2 U87 ( .A(n578), .B(n569), .Z(\OutEdge126[5] ) );
    VMW_NAND2 U88 ( .A(n579), .B(n569), .Z(\OutEdge126[4] ) );
    VMW_NAND2 U89 ( .A(n580), .B(n569), .Z(\OutEdge126[3] ) );
    VMW_NAND2 U90 ( .A(n581), .B(n569), .Z(\OutEdge126[2] ) );
    VMW_NAND2 U91 ( .A(n582), .B(n569), .Z(\OutEdge126[1] ) );
    VMW_NAND2 U92 ( .A(n583), .B(n569), .Z(\OutEdge126[0] ) );
    VMW_OAI211 U93 ( .A(n96), .B(n88), .C(n585), .D(n586), .Z(n584) );
    VMW_NAND2 U94 ( .A(n585), .B(n588), .Z(n587) );
    VMW_AO22 U95 ( .A(\temp294[15] ), .B(n586), .C(InEdges[47]), .D(n104), .Z(
        \temp384[15] ) );
    VMW_INV U96 ( .A(n88), .Z(n589) );
    VMW_OAI22 U97 ( .A(n591), .B(Start), .C(\path[2] ), .D(n569), .Z(n590) );
    VMW_OAI22 U98 ( .A(n584), .B(Start), .C(\path[1] ), .D(n569), .Z(n592) );
    VMW_OAI22 U99 ( .A(n587), .B(Start), .C(\path[0] ), .D(n569), .Z(n593) );
    VMW_MUX2I U100 ( .A(\temp384[15] ), .B(InEdges[63]), .S(n112), .Z(n567) );
    VMW_AND4 U101 ( .A(n595), .B(n596), .C(n597), .D(n598), .Z(n594) );
    VMW_INV U102 ( .A(Start), .Z(n569) );
    VMW_INV U103 ( .A(n96), .Z(n599) );
    VMW_OAI21 U104 ( .A(n96), .B(n589), .C(n586), .Z(n588) );
    VMW_AND4 U105 ( .A(n600), .B(n601), .C(n602), .D(n594), .Z(n603) );
    VMW_XNOR2 U106 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n598) );
    VMW_XNOR2 U107 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n597) );
    VMW_XNOR2 U108 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n596) );
    VMW_XNOR2 U109 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n595) );
    VMW_XNOR2 U110 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n601) );
    VMW_XNOR2 U111 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n600) );
    VMW_XNOR2 U112 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n602) );
    VMW_AO22 U113 ( .A(InEdges[9]), .B(n88), .C(OutEdge[9]), .D(n589), .Z(
        \temp200[9] ) );
    VMW_AO22 U114 ( .A(InEdges[25]), .B(n96), .C(\temp200[9] ), .D(n599), .Z(
        \temp294[9] ) );
    VMW_AO22 U115 ( .A(\temp294[9] ), .B(n586), .C(InEdges[41]), .D(n104), .Z(
        \temp384[9] ) );
    VMW_AO22 U116 ( .A(InEdges[8]), .B(n88), .C(OutEdge[8]), .D(n589), .Z(
        \temp200[8] ) );
    VMW_AO22 U117 ( .A(InEdges[24]), .B(n96), .C(\temp200[8] ), .D(n599), .Z(
        \temp294[8] ) );
    VMW_AO22 U118 ( .A(\temp294[8] ), .B(n586), .C(InEdges[40]), .D(n104), .Z(
        \temp384[8] ) );
    VMW_AO22 U119 ( .A(InEdges[7]), .B(n88), .C(OutEdge[7]), .D(n589), .Z(
        \temp200[7] ) );
    VMW_AO22 U120 ( .A(InEdges[23]), .B(n96), .C(\temp200[7] ), .D(n599), .Z(
        \temp294[7] ) );
    VMW_AO22 U121 ( .A(\temp294[7] ), .B(n586), .C(InEdges[39]), .D(n104), .Z(
        \temp384[7] ) );
    VMW_AO22 U122 ( .A(InEdges[6]), .B(n88), .C(OutEdge[6]), .D(n589), .Z(
        \temp200[6] ) );
    VMW_AO22 U123 ( .A(InEdges[22]), .B(n96), .C(\temp200[6] ), .D(n599), .Z(
        \temp294[6] ) );
    VMW_AO22 U124 ( .A(\temp294[6] ), .B(n586), .C(InEdges[38]), .D(n104), .Z(
        \temp384[6] ) );
    VMW_AO22 U125 ( .A(InEdges[5]), .B(n88), .C(OutEdge[5]), .D(n589), .Z(
        \temp200[5] ) );
    VMW_AO22 U126 ( .A(InEdges[21]), .B(n96), .C(\temp200[5] ), .D(n599), .Z(
        \temp294[5] ) );
    VMW_AO22 U127 ( .A(\temp294[5] ), .B(n586), .C(InEdges[37]), .D(n104), .Z(
        \temp384[5] ) );
    VMW_AO22 U128 ( .A(InEdges[4]), .B(n88), .C(OutEdge[4]), .D(n589), .Z(
        \temp200[4] ) );
    VMW_AO22 U129 ( .A(InEdges[20]), .B(n96), .C(\temp200[4] ), .D(n599), .Z(
        \temp294[4] ) );
    VMW_AO22 U130 ( .A(\temp294[4] ), .B(n586), .C(InEdges[36]), .D(n104), .Z(
        \temp384[4] ) );
    VMW_AO22 U131 ( .A(InEdges[3]), .B(n88), .C(OutEdge[3]), .D(n589), .Z(
        \temp200[3] ) );
    VMW_AO22 U132 ( .A(InEdges[19]), .B(n96), .C(\temp200[3] ), .D(n599), .Z(
        \temp294[3] ) );
    VMW_AO22 U133 ( .A(\temp294[3] ), .B(n586), .C(InEdges[35]), .D(n104), .Z(
        \temp384[3] ) );
    VMW_AO22 U134 ( .A(InEdges[2]), .B(n88), .C(OutEdge[2]), .D(n589), .Z(
        \temp200[2] ) );
    VMW_AO22 U135 ( .A(InEdges[18]), .B(n96), .C(\temp200[2] ), .D(n599), .Z(
        \temp294[2] ) );
    VMW_AO22 U136 ( .A(\temp294[2] ), .B(n586), .C(InEdges[34]), .D(n104), .Z(
        \temp384[2] ) );
    VMW_AO22 U137 ( .A(InEdges[1]), .B(n88), .C(OutEdge[1]), .D(n589), .Z(
        \temp200[1] ) );
    VMW_AO22 U138 ( .A(InEdges[17]), .B(n96), .C(\temp200[1] ), .D(n599), .Z(
        \temp294[1] ) );
    VMW_AO22 U139 ( .A(\temp294[1] ), .B(n586), .C(InEdges[33]), .D(n104), .Z(
        \temp384[1] ) );
    VMW_AO22 U140 ( .A(InEdges[15]), .B(n88), .C(OutEdge[15]), .D(n589), .Z(
        \temp200[15] ) );
    VMW_AO22 U141 ( .A(InEdges[31]), .B(n96), .C(\temp200[15] ), .D(n599), .Z(
        \temp294[15] ) );
    VMW_AO22 U142 ( .A(InEdges[14]), .B(n88), .C(OutEdge[14]), .D(n589), .Z(
        \temp200[14] ) );
    VMW_AO22 U143 ( .A(InEdges[30]), .B(n96), .C(\temp200[14] ), .D(n599), .Z(
        \temp294[14] ) );
    VMW_AO22 U144 ( .A(\temp294[14] ), .B(n586), .C(InEdges[46]), .D(n104), 
        .Z(\temp384[14] ) );
    VMW_AO22 U145 ( .A(InEdges[13]), .B(n88), .C(OutEdge[13]), .D(n589), .Z(
        \temp200[13] ) );
    VMW_AO22 U146 ( .A(InEdges[29]), .B(n96), .C(\temp200[13] ), .D(n599), .Z(
        \temp294[13] ) );
    VMW_AO22 U147 ( .A(\temp294[13] ), .B(n586), .C(InEdges[45]), .D(n104), 
        .Z(\temp384[13] ) );
    VMW_AO22 U148 ( .A(InEdges[12]), .B(n88), .C(OutEdge[12]), .D(n589), .Z(
        \temp200[12] ) );
    VMW_AO22 U149 ( .A(InEdges[28]), .B(n96), .C(\temp200[12] ), .D(n599), .Z(
        \temp294[12] ) );
    VMW_AO22 U150 ( .A(\temp294[12] ), .B(n586), .C(InEdges[44]), .D(n104), 
        .Z(\temp384[12] ) );
    VMW_AO22 U151 ( .A(InEdges[11]), .B(n88), .C(OutEdge[11]), .D(n589), .Z(
        \temp200[11] ) );
    VMW_AO22 U152 ( .A(InEdges[27]), .B(n96), .C(\temp200[11] ), .D(n599), .Z(
        \temp294[11] ) );
    VMW_AO22 U153 ( .A(\temp294[11] ), .B(n586), .C(InEdges[43]), .D(n104), 
        .Z(\temp384[11] ) );
    VMW_AO22 U154 ( .A(InEdges[10]), .B(n88), .C(OutEdge[10]), .D(n589), .Z(
        \temp200[10] ) );
    VMW_AO22 U155 ( .A(InEdges[26]), .B(n96), .C(\temp200[10] ), .D(n599), .Z(
        \temp294[10] ) );
    VMW_AO22 U156 ( .A(\temp294[10] ), .B(n586), .C(InEdges[42]), .D(n104), 
        .Z(\temp384[10] ) );
    VMW_AO22 U157 ( .A(InEdges[0]), .B(n88), .C(OutEdge[0]), .D(n589), .Z(
        \temp200[0] ) );
    VMW_AO22 U158 ( .A(InEdges[16]), .B(n96), .C(\temp200[0] ), .D(n599), .Z(
        \temp294[0] ) );
    VMW_AO22 U159 ( .A(\temp294[0] ), .B(n586), .C(InEdges[32]), .D(n104), .Z(
        \temp384[0] ) );
    VMW_AND4 U160 ( .A(n599), .B(n586), .C(n589), .D(n585), .Z(n591) );
    VMW_MUX2I U161 ( .A(\temp384[9] ), .B(InEdges[57]), .S(n112), .Z(n574) );
    VMW_MUX2I U162 ( .A(\temp384[8] ), .B(InEdges[56]), .S(n112), .Z(n575) );
    VMW_MUX2I U163 ( .A(\temp384[7] ), .B(InEdges[55]), .S(n112), .Z(n576) );
    VMW_MUX2I U164 ( .A(\temp384[6] ), .B(InEdges[54]), .S(n112), .Z(n577) );
    VMW_MUX2I U165 ( .A(\temp384[5] ), .B(InEdges[53]), .S(n112), .Z(n578) );
    VMW_MUX2I U166 ( .A(\temp384[4] ), .B(InEdges[52]), .S(n112), .Z(n579) );
    VMW_MUX2I U167 ( .A(\temp384[3] ), .B(InEdges[51]), .S(n112), .Z(n580) );
    VMW_MUX2I U168 ( .A(\temp384[2] ), .B(InEdges[50]), .S(n112), .Z(n581) );
    VMW_MUX2I U169 ( .A(\temp384[1] ), .B(InEdges[49]), .S(n112), .Z(n582) );
    VMW_MUX2I U170 ( .A(\temp384[14] ), .B(InEdges[62]), .S(n112), .Z(n568) );
    VMW_MUX2I U171 ( .A(\temp384[13] ), .B(InEdges[61]), .S(n112), .Z(n570) );
    VMW_MUX2I U172 ( .A(\temp384[12] ), .B(InEdges[60]), .S(n112), .Z(n571) );
    VMW_MUX2I U173 ( .A(\temp384[11] ), .B(InEdges[59]), .S(n112), .Z(n572) );
    VMW_MUX2I U174 ( .A(\temp384[10] ), .B(InEdges[58]), .S(n112), .Z(n573) );
    VMW_MUX2I U175 ( .A(\temp384[0] ), .B(InEdges[48]), .S(n112), .Z(n583) );
    VMW_INV U176 ( .A(n104), .Z(n586) );
    VMW_INV U177 ( .A(n112), .Z(n585) );
    VMW_INV U178 ( .A(n590), .Z(n605) );
    VMW_INV U179 ( .A(n592), .Z(n606) );
    VMW_INV U180 ( .A(n593), .Z(n604) );
    VMW_BUFIZ U181 ( .A(\path[1] ), .E(n603), .Z(\PathData[1] ) );
    VMW_BUFIZ U182 ( .A(\path[0] ), .E(n603), .Z(\PathData[0] ) );
    VMW_BUFIZ U183 ( .A(\path[2] ), .E(n603), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n604), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n605), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n606), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge126[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge126[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge126[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge126[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge126[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge126[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge126[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge126[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge126[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge126[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge126[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge126[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge126[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge126[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge126[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge126[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n610), .TC(n610), .GE_GT(n88) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_2 lte_55_1 ( .A({\temp200[15] , 
        \temp200[14] , \temp200[13] , \temp200[12] , \temp200[11] , 
        \temp200[10] , \temp200[9] , \temp200[8] , \temp200[7] , \temp200[6] , 
        \temp200[5] , \temp200[4] , \temp200[3] , \temp200[2] , \temp200[1] , 
        \temp200[0] }), .B(InEdges[31:16]), .LEQ(n609), .TC(n609), .GE_GT(n96)
         );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp294[15] , 
        \temp294[14] , \temp294[13] , \temp294[12] , \temp294[11] , 
        \temp294[10] , \temp294[9] , \temp294[8] , \temp294[7] , \temp294[6] , 
        \temp294[5] , \temp294[4] , \temp294[3] , \temp294[2] , \temp294[1] , 
        \temp294[0] }), .B(InEdges[47:32]), .LEQ(n608), .TC(n608), .GE_GT(n104
        ) );
    NodeAux_INDEGREE4_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp384[15] , 
        \temp384[14] , \temp384[13] , \temp384[12] , \temp384[11] , 
        \temp384[10] , \temp384[9] , \temp384[8] , \temp384[7] , \temp384[6] , 
        \temp384[5] , \temp384[4] , \temp384[3] , \temp384[2] , \temp384[1] , 
        \temp384[0] }), .B(InEdges[63:48]), .LEQ(n607), .TC(n607), .GE_GT(n112
        ) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, 
        n93, n94, n95, n96, n97, n99, n100, n101, n102, n103, n104, n105, n107, 
        n108, n109, n110, n111, n112, n113, n115, n116;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n91), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n92) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n92), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n99), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n99), .B(A[9]), .Z(n100) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n100), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n107) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n107), .D(n104), .Z(n108) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n108), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n115) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n116), .C(n115), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n91) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n99) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n116) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n123), .B(B[0]), .C(n124), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n124), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n135), .B(B[6]), .Z(n134) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n137), .C(n132), .D(n127), .Z(n136) );
    VMW_OR2 U14 ( .A(B[6]), .B(n135), .Z(n138) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n140), .C(n138), .D(n136), .Z(n139) );
    VMW_NAND2 U16 ( .A(n142), .B(B[8]), .Z(n141) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n144), .C(n139), .D(n134), .Z(n143) );
    VMW_OR2 U18 ( .A(B[8]), .B(n142), .Z(n145) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n147), .C(n145), .D(n143), .Z(n146) );
    VMW_NAND2 U20 ( .A(n149), .B(B[10]), .Z(n148) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n151), .C(n146), .D(n141), .Z(n150) );
    VMW_NAND2 U22 ( .A(n151), .B(A[9]), .Z(n152) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n149), .C(n152), .D(n150), .Z(n153) );
    VMW_NAND2 U24 ( .A(n155), .B(B[12]), .Z(n154) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n157), .C(n153), .D(n148), .Z(n156) );
    VMW_NAND2 U26 ( .A(n157), .B(A[11]), .Z(n158) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n155), .C(n158), .D(n156), .Z(n159) );
    VMW_NAND2 U28 ( .A(n161), .B(B[14]), .Z(n160) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n163), .C(n159), .D(n154), .Z(n162) );
    VMW_NAND2 U30 ( .A(n163), .B(A[13]), .Z(n164) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n161), .C(n164), .D(n162), .Z(n165) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n166), .C(n165), .D(n160), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n155) );
    VMW_INV U34 ( .A(B[7]), .Z(n144) );
    VMW_INV U35 ( .A(A[7]), .Z(n147) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n149) );
    VMW_INV U39 ( .A(B[9]), .Z(n151) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n142) );
    VMW_INV U42 ( .A(A[14]), .Z(n161) );
    VMW_INV U43 ( .A(B[11]), .Z(n157) );
    VMW_INV U44 ( .A(A[5]), .Z(n140) );
    VMW_INV U45 ( .A(B[5]), .Z(n137) );
    VMW_INV U46 ( .A(A[1]), .Z(n124) );
    VMW_INV U47 ( .A(B[15]), .Z(n166) );
    VMW_INV U48 ( .A(B[13]), .Z(n163) );
    VMW_INV U49 ( .A(A[6]), .Z(n135) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n123) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
        n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
        n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
        n214, n215;
    VMW_OAI21 U3 ( .A(B[15]), .B(n167), .C(n168), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n170), .B(B[2]), .Z(n169) );
    VMW_AO22 U5 ( .A(n172), .B(B[0]), .C(n173), .D(B[1]), .Z(n171) );
    VMW_OR2 U6 ( .A(B[2]), .B(n170), .Z(n174) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n173), .C(n174), .D(n171), .Z(n175) );
    VMW_NAND2 U8 ( .A(n177), .B(B[4]), .Z(n176) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n179), .C(n175), .D(n169), .Z(n178) );
    VMW_OR2 U10 ( .A(B[4]), .B(n177), .Z(n180) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n182), .C(n180), .D(n178), .Z(n181) );
    VMW_NAND2 U12 ( .A(n184), .B(B[6]), .Z(n183) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n186), .C(n181), .D(n176), .Z(n185) );
    VMW_OR2 U14 ( .A(B[6]), .B(n184), .Z(n187) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n189), .C(n187), .D(n185), .Z(n188) );
    VMW_NAND2 U16 ( .A(n191), .B(B[8]), .Z(n190) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n193), .C(n188), .D(n183), .Z(n192) );
    VMW_OR2 U18 ( .A(B[8]), .B(n191), .Z(n194) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n196), .C(n194), .D(n192), .Z(n195) );
    VMW_NAND2 U20 ( .A(n198), .B(B[10]), .Z(n197) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n200), .C(n195), .D(n190), .Z(n199) );
    VMW_NAND2 U22 ( .A(n200), .B(A[9]), .Z(n201) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n198), .C(n201), .D(n199), .Z(n202) );
    VMW_NAND2 U24 ( .A(n204), .B(B[12]), .Z(n203) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n206), .C(n202), .D(n197), .Z(n205) );
    VMW_NAND2 U26 ( .A(n206), .B(A[11]), .Z(n207) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n204), .C(n207), .D(n205), .Z(n208) );
    VMW_NAND2 U28 ( .A(n210), .B(B[14]), .Z(n209) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n212), .C(n208), .D(n203), .Z(n211) );
    VMW_NAND2 U30 ( .A(n212), .B(A[13]), .Z(n213) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n210), .C(n213), .D(n211), .Z(n214) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n215), .C(n214), .D(n209), .Z(n168) );
    VMW_INV U33 ( .A(A[12]), .Z(n204) );
    VMW_INV U34 ( .A(B[7]), .Z(n193) );
    VMW_INV U35 ( .A(A[7]), .Z(n196) );
    VMW_INV U36 ( .A(A[3]), .Z(n182) );
    VMW_INV U37 ( .A(B[3]), .Z(n179) );
    VMW_INV U38 ( .A(A[10]), .Z(n198) );
    VMW_INV U39 ( .A(B[9]), .Z(n200) );
    VMW_INV U40 ( .A(A[4]), .Z(n177) );
    VMW_INV U41 ( .A(A[8]), .Z(n191) );
    VMW_INV U42 ( .A(A[14]), .Z(n210) );
    VMW_INV U43 ( .A(B[11]), .Z(n206) );
    VMW_INV U44 ( .A(A[5]), .Z(n189) );
    VMW_INV U45 ( .A(B[5]), .Z(n186) );
    VMW_INV U46 ( .A(A[1]), .Z(n173) );
    VMW_INV U47 ( .A(B[15]), .Z(n215) );
    VMW_INV U48 ( .A(B[13]), .Z(n212) );
    VMW_INV U49 ( .A(A[6]), .Z(n184) );
    VMW_INV U50 ( .A(A[2]), .Z(n170) );
    VMW_INV U51 ( .A(A[0]), .Z(n172) );
    VMW_INV U52 ( .A(A[15]), .Z(n167) );
endmodule


module NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264;
    VMW_OAI21 U3 ( .A(B[15]), .B(n216), .C(n217), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n219), .B(B[2]), .Z(n218) );
    VMW_AO22 U5 ( .A(n221), .B(B[0]), .C(n222), .D(B[1]), .Z(n220) );
    VMW_OR2 U6 ( .A(B[2]), .B(n219), .Z(n223) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n222), .C(n223), .D(n220), .Z(n224) );
    VMW_NAND2 U8 ( .A(n226), .B(B[4]), .Z(n225) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n228), .C(n224), .D(n218), .Z(n227) );
    VMW_OR2 U10 ( .A(B[4]), .B(n226), .Z(n229) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n231), .C(n229), .D(n227), .Z(n230) );
    VMW_NAND2 U12 ( .A(n233), .B(B[6]), .Z(n232) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n235), .C(n230), .D(n225), .Z(n234) );
    VMW_OR2 U14 ( .A(B[6]), .B(n233), .Z(n236) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n238), .C(n236), .D(n234), .Z(n237) );
    VMW_NAND2 U16 ( .A(n240), .B(B[8]), .Z(n239) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n242), .C(n237), .D(n232), .Z(n241) );
    VMW_OR2 U18 ( .A(B[8]), .B(n240), .Z(n243) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n245), .C(n243), .D(n241), .Z(n244) );
    VMW_NAND2 U20 ( .A(n247), .B(B[10]), .Z(n246) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n249), .C(n244), .D(n239), .Z(n248) );
    VMW_NAND2 U22 ( .A(n249), .B(A[9]), .Z(n250) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n247), .C(n250), .D(n248), .Z(n251) );
    VMW_NAND2 U24 ( .A(n253), .B(B[12]), .Z(n252) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n255), .C(n251), .D(n246), .Z(n254) );
    VMW_NAND2 U26 ( .A(n255), .B(A[11]), .Z(n256) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n253), .C(n256), .D(n254), .Z(n257) );
    VMW_NAND2 U28 ( .A(n259), .B(B[14]), .Z(n258) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n261), .C(n257), .D(n252), .Z(n260) );
    VMW_NAND2 U30 ( .A(n261), .B(A[13]), .Z(n262) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n259), .C(n262), .D(n260), .Z(n263) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n264), .C(n263), .D(n258), .Z(n217) );
    VMW_INV U33 ( .A(A[12]), .Z(n253) );
    VMW_INV U34 ( .A(B[7]), .Z(n242) );
    VMW_INV U35 ( .A(A[7]), .Z(n245) );
    VMW_INV U36 ( .A(A[3]), .Z(n231) );
    VMW_INV U37 ( .A(B[3]), .Z(n228) );
    VMW_INV U38 ( .A(A[10]), .Z(n247) );
    VMW_INV U39 ( .A(B[9]), .Z(n249) );
    VMW_INV U40 ( .A(A[4]), .Z(n226) );
    VMW_INV U41 ( .A(A[8]), .Z(n240) );
    VMW_INV U42 ( .A(A[14]), .Z(n259) );
    VMW_INV U43 ( .A(B[11]), .Z(n255) );
    VMW_INV U44 ( .A(A[5]), .Z(n238) );
    VMW_INV U45 ( .A(B[5]), .Z(n235) );
    VMW_INV U46 ( .A(A[1]), .Z(n222) );
    VMW_INV U47 ( .A(B[15]), .Z(n264) );
    VMW_INV U48 ( .A(B[13]), .Z(n261) );
    VMW_INV U49 ( .A(A[6]), .Z(n233) );
    VMW_INV U50 ( .A(A[2]), .Z(n219) );
    VMW_INV U51 ( .A(A[0]), .Z(n221) );
    VMW_INV U52 ( .A(A[15]), .Z(n216) );
endmodule


module NodeAux_INDEGREE5_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp210[13] , \temp484[4] , \temp394[5] , \temp304[13] , 
        \temp210[3] , \temp394[13] , \OutEdge136[14] , \temp394[1] , 
        \temp484[0] , \OutEdge136[10] , \path[2] , \temp394[8] , \temp210[7] , 
        \temp484[9] , \temp394[15] , \path[0] , \temp210[5] , \OutEdge136[12] , 
        \temp210[15] , \temp304[15] , \temp394[3] , \temp484[2] , \temp210[1] , 
        n90, \temp394[11] , \temp484[6] , \temp394[7] , \temp210[8] , 
        \temp304[11] , \temp210[11] , n98, n114, \OutEdge136[2] , \temp304[4] , 
        \OutEdge136[6] , \temp304[9] , \temp304[0] , \temp484[13] , n106, 
        \temp304[2] , \temp484[11] , \OutEdge136[4] , \temp484[15] , 
        \temp304[6] , \OutEdge136[9] , \OutEdge136[0] , \temp484[14] , 
        \OutEdge136[8] , \temp304[7] , \OutEdge136[1] , \temp304[3] , 
        \temp484[10] , \OutEdge136[5] , \OutEdge136[7] , \temp304[8] , 
        \temp304[1] , \temp484[12] , \OutEdge136[3] , \temp304[5] , 
        \temp394[10] , \temp210[0] , \temp484[7] , \temp210[9] , \temp304[10] , 
        \temp394[6] , \temp210[10] , \temp210[4] , \path[1] , \temp394[14] , 
        \OutEdge136[13] , \temp210[14] , \temp394[2] , n122, \temp304[14] , 
        \temp484[3] , \temp394[0] , \temp484[1] , \OutEdge136[11] , 
        \temp210[6] , \temp394[9] , \temp484[8] , \temp210[12] , \temp484[5] , 
        \temp304[12] , \temp394[4] , \OutEdge136[15] , \temp394[12] , 
        \temp210[2] , n667, n668, n669, n670, n671, n672, n673, n674, n675, 
        n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
        n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
        n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
        n712, n713;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U82 ( .Z(n712) );
    VMW_PULLDOWN U83 ( .Z(n709) );
    VMW_PULLDOWN U84 ( .Z(n711) );
    VMW_PULLDOWN U85 ( .Z(n710) );
    VMW_PULLDOWN U86 ( .Z(n713) );
    VMW_AO21 U87 ( .A(\temp484[15] ), .B(n667), .C(n668), .Z(\OutEdge136[15] )
         );
    VMW_NAND2 U88 ( .A(n669), .B(n670), .Z(\OutEdge136[14] ) );
    VMW_NAND2 U89 ( .A(n671), .B(n670), .Z(\OutEdge136[13] ) );
    VMW_NAND2 U90 ( .A(n672), .B(n670), .Z(\OutEdge136[12] ) );
    VMW_NAND2 U91 ( .A(n673), .B(n670), .Z(\OutEdge136[11] ) );
    VMW_NAND2 U92 ( .A(n674), .B(n670), .Z(\OutEdge136[10] ) );
    VMW_NAND2 U93 ( .A(n675), .B(n670), .Z(\OutEdge136[9] ) );
    VMW_NAND2 U94 ( .A(n676), .B(n670), .Z(\OutEdge136[8] ) );
    VMW_NAND2 U95 ( .A(n677), .B(n670), .Z(\OutEdge136[7] ) );
    VMW_NAND2 U96 ( .A(n678), .B(n670), .Z(\OutEdge136[6] ) );
    VMW_NAND2 U97 ( .A(n679), .B(n670), .Z(\OutEdge136[5] ) );
    VMW_NAND2 U98 ( .A(n680), .B(n670), .Z(\OutEdge136[4] ) );
    VMW_NAND2 U99 ( .A(n681), .B(n670), .Z(\OutEdge136[3] ) );
    VMW_NAND2 U100 ( .A(n682), .B(n670), .Z(\OutEdge136[2] ) );
    VMW_NAND2 U101 ( .A(n683), .B(n670), .Z(\OutEdge136[1] ) );
    VMW_NAND2 U102 ( .A(n684), .B(n670), .Z(\OutEdge136[0] ) );
    VMW_AO22 U103 ( .A(\path[1] ), .B(Start), .C(n667), .D(n685), .Z(n708) );
    VMW_OAI21 U104 ( .A(n670), .B(n686), .C(n687), .Z(n706) );
    VMW_OR2 U105 ( .A(n122), .B(n689), .Z(n688) );
    VMW_AO22 U106 ( .A(InEdges[63]), .B(n114), .C(\temp394[15] ), .D(n690), 
        .Z(\temp484[15] ) );
    VMW_INV U107 ( .A(Start), .Z(n670) );
    VMW_OR2 U108 ( .A(Start), .B(n122), .Z(n691) );
    VMW_OAI22 U109 ( .A(\path[2] ), .B(n670), .C(n688), .D(Start), .Z(n692) );
    VMW_AND4 U110 ( .A(n694), .B(n695), .C(n696), .D(n697), .Z(n693) );
    VMW_INV U111 ( .A(n114), .Z(n690) );
    VMW_INV U112 ( .A(n106), .Z(n698) );
    VMW_NOR4 U113 ( .A(n98), .B(n106), .C(n90), .D(n114), .Z(n689) );
    VMW_OAI211 U114 ( .A(n90), .B(n98), .C(n698), .D(n690), .Z(n685) );
    VMW_OAI21 U115 ( .A(n98), .B(n700), .C(n698), .Z(n699) );
    VMW_AO21 U116 ( .A(n690), .B(n699), .C(n691), .Z(n687) );
    VMW_AND4 U117 ( .A(n701), .B(n702), .C(n703), .D(n693), .Z(n705) );
    VMW_AND3 U118 ( .A(n122), .B(n670), .C(InEdges[79]), .Z(n668) );
    VMW_XNOR2 U119 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n697) );
    VMW_XNOR2 U120 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n696) );
    VMW_XNOR2 U121 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n695) );
    VMW_XNOR2 U122 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n694) );
    VMW_XNOR2 U123 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n702) );
    VMW_XNOR2 U124 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n701) );
    VMW_XNOR2 U125 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n703) );
    VMW_AO22 U126 ( .A(OutEdge[9]), .B(n700), .C(InEdges[9]), .D(n90), .Z(
        \temp210[9] ) );
    VMW_AO22 U127 ( .A(\temp210[9] ), .B(n704), .C(InEdges[25]), .D(n98), .Z(
        \temp304[9] ) );
    VMW_AO22 U128 ( .A(\temp304[9] ), .B(n698), .C(InEdges[41]), .D(n106), .Z(
        \temp394[9] ) );
    VMW_AO22 U129 ( .A(\temp394[9] ), .B(n690), .C(InEdges[57]), .D(n114), .Z(
        \temp484[9] ) );
    VMW_AO22 U130 ( .A(OutEdge[8]), .B(n700), .C(InEdges[8]), .D(n90), .Z(
        \temp210[8] ) );
    VMW_AO22 U131 ( .A(\temp210[8] ), .B(n704), .C(InEdges[24]), .D(n98), .Z(
        \temp304[8] ) );
    VMW_AO22 U132 ( .A(\temp304[8] ), .B(n698), .C(InEdges[40]), .D(n106), .Z(
        \temp394[8] ) );
    VMW_AO22 U133 ( .A(\temp394[8] ), .B(n690), .C(InEdges[56]), .D(n114), .Z(
        \temp484[8] ) );
    VMW_AO22 U134 ( .A(OutEdge[7]), .B(n700), .C(InEdges[7]), .D(n90), .Z(
        \temp210[7] ) );
    VMW_AO22 U135 ( .A(\temp210[7] ), .B(n704), .C(InEdges[23]), .D(n98), .Z(
        \temp304[7] ) );
    VMW_AO22 U136 ( .A(\temp304[7] ), .B(n698), .C(InEdges[39]), .D(n106), .Z(
        \temp394[7] ) );
    VMW_AO22 U137 ( .A(\temp394[7] ), .B(n690), .C(InEdges[55]), .D(n114), .Z(
        \temp484[7] ) );
    VMW_AO22 U138 ( .A(OutEdge[6]), .B(n700), .C(InEdges[6]), .D(n90), .Z(
        \temp210[6] ) );
    VMW_AO22 U139 ( .A(\temp210[6] ), .B(n704), .C(InEdges[22]), .D(n98), .Z(
        \temp304[6] ) );
    VMW_AO22 U140 ( .A(\temp304[6] ), .B(n698), .C(InEdges[38]), .D(n106), .Z(
        \temp394[6] ) );
    VMW_AO22 U141 ( .A(\temp394[6] ), .B(n690), .C(InEdges[54]), .D(n114), .Z(
        \temp484[6] ) );
    VMW_AO22 U142 ( .A(OutEdge[5]), .B(n700), .C(InEdges[5]), .D(n90), .Z(
        \temp210[5] ) );
    VMW_AO22 U143 ( .A(\temp210[5] ), .B(n704), .C(InEdges[21]), .D(n98), .Z(
        \temp304[5] ) );
    VMW_AO22 U144 ( .A(\temp304[5] ), .B(n698), .C(InEdges[37]), .D(n106), .Z(
        \temp394[5] ) );
    VMW_AO22 U145 ( .A(\temp394[5] ), .B(n690), .C(InEdges[53]), .D(n114), .Z(
        \temp484[5] ) );
    VMW_AO22 U146 ( .A(OutEdge[4]), .B(n700), .C(InEdges[4]), .D(n90), .Z(
        \temp210[4] ) );
    VMW_AO22 U147 ( .A(\temp210[4] ), .B(n704), .C(InEdges[20]), .D(n98), .Z(
        \temp304[4] ) );
    VMW_AO22 U148 ( .A(\temp304[4] ), .B(n698), .C(InEdges[36]), .D(n106), .Z(
        \temp394[4] ) );
    VMW_AO22 U149 ( .A(\temp394[4] ), .B(n690), .C(InEdges[52]), .D(n114), .Z(
        \temp484[4] ) );
    VMW_AO22 U150 ( .A(OutEdge[3]), .B(n700), .C(InEdges[3]), .D(n90), .Z(
        \temp210[3] ) );
    VMW_AO22 U151 ( .A(\temp210[3] ), .B(n704), .C(InEdges[19]), .D(n98), .Z(
        \temp304[3] ) );
    VMW_AO22 U152 ( .A(\temp304[3] ), .B(n698), .C(InEdges[35]), .D(n106), .Z(
        \temp394[3] ) );
    VMW_AO22 U153 ( .A(\temp394[3] ), .B(n690), .C(InEdges[51]), .D(n114), .Z(
        \temp484[3] ) );
    VMW_AO22 U154 ( .A(OutEdge[2]), .B(n700), .C(InEdges[2]), .D(n90), .Z(
        \temp210[2] ) );
    VMW_AO22 U155 ( .A(\temp210[2] ), .B(n704), .C(InEdges[18]), .D(n98), .Z(
        \temp304[2] ) );
    VMW_AO22 U156 ( .A(\temp304[2] ), .B(n698), .C(InEdges[34]), .D(n106), .Z(
        \temp394[2] ) );
    VMW_AO22 U157 ( .A(\temp394[2] ), .B(n690), .C(InEdges[50]), .D(n114), .Z(
        \temp484[2] ) );
    VMW_AO22 U158 ( .A(OutEdge[1]), .B(n700), .C(InEdges[1]), .D(n90), .Z(
        \temp210[1] ) );
    VMW_AO22 U159 ( .A(\temp210[1] ), .B(n704), .C(InEdges[17]), .D(n98), .Z(
        \temp304[1] ) );
    VMW_AO22 U160 ( .A(\temp304[1] ), .B(n698), .C(InEdges[33]), .D(n106), .Z(
        \temp394[1] ) );
    VMW_AO22 U161 ( .A(\temp394[1] ), .B(n690), .C(InEdges[49]), .D(n114), .Z(
        \temp484[1] ) );
    VMW_AO22 U162 ( .A(OutEdge[15]), .B(n700), .C(InEdges[15]), .D(n90), .Z(
        \temp210[15] ) );
    VMW_AO22 U163 ( .A(\temp210[15] ), .B(n704), .C(InEdges[31]), .D(n98), .Z(
        \temp304[15] ) );
    VMW_AO22 U164 ( .A(\temp304[15] ), .B(n698), .C(InEdges[47]), .D(n106), 
        .Z(\temp394[15] ) );
    VMW_AO22 U165 ( .A(OutEdge[14]), .B(n700), .C(InEdges[14]), .D(n90), .Z(
        \temp210[14] ) );
    VMW_AO22 U166 ( .A(\temp210[14] ), .B(n704), .C(InEdges[30]), .D(n98), .Z(
        \temp304[14] ) );
    VMW_AO22 U167 ( .A(\temp304[14] ), .B(n698), .C(InEdges[46]), .D(n106), 
        .Z(\temp394[14] ) );
    VMW_AO22 U168 ( .A(\temp394[14] ), .B(n690), .C(InEdges[62]), .D(n114), 
        .Z(\temp484[14] ) );
    VMW_AO22 U169 ( .A(OutEdge[13]), .B(n700), .C(InEdges[13]), .D(n90), .Z(
        \temp210[13] ) );
    VMW_AO22 U170 ( .A(\temp210[13] ), .B(n704), .C(InEdges[29]), .D(n98), .Z(
        \temp304[13] ) );
    VMW_AO22 U171 ( .A(\temp304[13] ), .B(n698), .C(InEdges[45]), .D(n106), 
        .Z(\temp394[13] ) );
    VMW_AO22 U172 ( .A(\temp394[13] ), .B(n690), .C(InEdges[61]), .D(n114), 
        .Z(\temp484[13] ) );
    VMW_AO22 U173 ( .A(OutEdge[12]), .B(n700), .C(InEdges[12]), .D(n90), .Z(
        \temp210[12] ) );
    VMW_AO22 U174 ( .A(\temp210[12] ), .B(n704), .C(InEdges[28]), .D(n98), .Z(
        \temp304[12] ) );
    VMW_AO22 U175 ( .A(\temp304[12] ), .B(n698), .C(InEdges[44]), .D(n106), 
        .Z(\temp394[12] ) );
    VMW_AO22 U176 ( .A(\temp394[12] ), .B(n690), .C(InEdges[60]), .D(n114), 
        .Z(\temp484[12] ) );
    VMW_AO22 U177 ( .A(OutEdge[11]), .B(n700), .C(InEdges[11]), .D(n90), .Z(
        \temp210[11] ) );
    VMW_AO22 U178 ( .A(\temp210[11] ), .B(n704), .C(InEdges[27]), .D(n98), .Z(
        \temp304[11] ) );
    VMW_AO22 U179 ( .A(\temp304[11] ), .B(n698), .C(InEdges[43]), .D(n106), 
        .Z(\temp394[11] ) );
    VMW_AO22 U180 ( .A(\temp394[11] ), .B(n690), .C(InEdges[59]), .D(n114), 
        .Z(\temp484[11] ) );
    VMW_AO22 U181 ( .A(OutEdge[10]), .B(n700), .C(InEdges[10]), .D(n90), .Z(
        \temp210[10] ) );
    VMW_AO22 U182 ( .A(\temp210[10] ), .B(n704), .C(InEdges[26]), .D(n98), .Z(
        \temp304[10] ) );
    VMW_AO22 U183 ( .A(\temp304[10] ), .B(n698), .C(InEdges[42]), .D(n106), 
        .Z(\temp394[10] ) );
    VMW_AO22 U184 ( .A(\temp394[10] ), .B(n690), .C(InEdges[58]), .D(n114), 
        .Z(\temp484[10] ) );
    VMW_AO22 U185 ( .A(OutEdge[0]), .B(n700), .C(InEdges[0]), .D(n90), .Z(
        \temp210[0] ) );
    VMW_AO22 U186 ( .A(\temp210[0] ), .B(n704), .C(InEdges[16]), .D(n98), .Z(
        \temp304[0] ) );
    VMW_AO22 U187 ( .A(\temp304[0] ), .B(n698), .C(InEdges[32]), .D(n106), .Z(
        \temp394[0] ) );
    VMW_AO22 U188 ( .A(\temp394[0] ), .B(n690), .C(InEdges[48]), .D(n114), .Z(
        \temp484[0] ) );
    VMW_MUX2I U189 ( .A(\temp484[9] ), .B(InEdges[73]), .S(n122), .Z(n675) );
    VMW_MUX2I U190 ( .A(\temp484[8] ), .B(InEdges[72]), .S(n122), .Z(n676) );
    VMW_MUX2I U191 ( .A(\temp484[7] ), .B(InEdges[71]), .S(n122), .Z(n677) );
    VMW_MUX2I U192 ( .A(\temp484[6] ), .B(InEdges[70]), .S(n122), .Z(n678) );
    VMW_MUX2I U193 ( .A(\temp484[5] ), .B(InEdges[69]), .S(n122), .Z(n679) );
    VMW_MUX2I U194 ( .A(\temp484[4] ), .B(InEdges[68]), .S(n122), .Z(n680) );
    VMW_MUX2I U195 ( .A(\temp484[3] ), .B(InEdges[67]), .S(n122), .Z(n681) );
    VMW_MUX2I U196 ( .A(\temp484[2] ), .B(InEdges[66]), .S(n122), .Z(n682) );
    VMW_MUX2I U197 ( .A(\temp484[1] ), .B(InEdges[65]), .S(n122), .Z(n683) );
    VMW_MUX2I U198 ( .A(\temp484[14] ), .B(InEdges[78]), .S(n122), .Z(n669) );
    VMW_MUX2I U199 ( .A(\temp484[13] ), .B(InEdges[77]), .S(n122), .Z(n671) );
    VMW_MUX2I U200 ( .A(\temp484[12] ), .B(InEdges[76]), .S(n122), .Z(n672) );
    VMW_MUX2I U201 ( .A(\temp484[11] ), .B(InEdges[75]), .S(n122), .Z(n673) );
    VMW_MUX2I U202 ( .A(\temp484[10] ), .B(InEdges[74]), .S(n122), .Z(n674) );
    VMW_MUX2I U203 ( .A(\temp484[0] ), .B(InEdges[64]), .S(n122), .Z(n684) );
    VMW_INV U204 ( .A(n90), .Z(n700) );
    VMW_INV U205 ( .A(n98), .Z(n704) );
    VMW_INV U206 ( .A(n691), .Z(n667) );
    VMW_INV U207 ( .A(n692), .Z(n707) );
    VMW_INV U208 ( .A(\path[0] ), .Z(n686) );
    VMW_BUFIZ U209 ( .A(\path[1] ), .E(n705), .Z(\PathData[1] ) );
    VMW_BUFIZ U210 ( .A(\path[0] ), .E(n705), .Z(\PathData[0] ) );
    VMW_BUFIZ U211 ( .A(\path[2] ), .E(n705), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n706), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n707), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n708), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge136[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge136[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge136[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge136[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge136[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge136[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge136[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge136[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge136[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge136[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge136[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge136[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge136[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge136[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge136[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge136[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_4 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n713), .TC(n713), .GE_GT(n90) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp484[15] , 
        \temp484[14] , \temp484[13] , \temp484[12] , \temp484[11] , 
        \temp484[10] , \temp484[9] , \temp484[8] , \temp484[7] , \temp484[6] , 
        \temp484[5] , \temp484[4] , \temp484[3] , \temp484[2] , \temp484[1] , 
        \temp484[0] }), .B(InEdges[79:64]), .LEQ(n712), .TC(n712), .GE_GT(n122
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_2 lte_55_2 ( .A({\temp304[15] , 
        \temp304[14] , \temp304[13] , \temp304[12] , \temp304[11] , 
        \temp304[10] , \temp304[9] , \temp304[8] , \temp304[7] , \temp304[6] , 
        \temp304[5] , \temp304[4] , \temp304[3] , \temp304[2] , \temp304[1] , 
        \temp304[0] }), .B(InEdges[47:32]), .LEQ(n711), .TC(n711), .GE_GT(n106
        ) );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_1 lte_55_1 ( .A({\temp210[15] , 
        \temp210[14] , \temp210[13] , \temp210[12] , \temp210[11] , 
        \temp210[10] , \temp210[9] , \temp210[8] , \temp210[7] , \temp210[6] , 
        \temp210[5] , \temp210[4] , \temp210[3] , \temp210[2] , \temp210[1] , 
        \temp210[0] }), .B(InEdges[31:16]), .LEQ(n710), .TC(n710), .GE_GT(n98)
         );
    NodeAux_INDEGREE5_SOURCE0_DW01_cmp2_16_0 lte_55_3 ( .A({\temp394[15] , 
        \temp394[14] , \temp394[13] , \temp394[12] , \temp394[11] , 
        \temp394[10] , \temp394[9] , \temp394[8] , \temp394[7] , \temp394[6] , 
        \temp394[5] , \temp394[4] , \temp394[3] , \temp394[2] , \temp394[1] , 
        \temp394[0] }), .B(InEdges[63:48]), .LEQ(n709), .TC(n709), .GE_GT(n114
        ) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, 
        n107, n109, n110, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n94), .C(n91), .D(n89), .Z(n93) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n93), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n101) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n102) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n101), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n110), .B(B[14]), .Z(n109) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n109), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n94) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n110) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, 
        n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n166, n167;
    VMW_OAI21 U3 ( .A(B[15]), .B(n117), .C(n118), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n125) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n125), .D(n121), .Z(n126) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n126), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n134), .C(n131), .D(n129), .Z(n133) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n133), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n143), .B(B[8]), .Z(n142) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n145), .C(n140), .D(n135), .Z(n144) );
    VMW_OR2 U18 ( .A(B[8]), .B(n143), .Z(n146) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n148), .C(n146), .D(n144), .Z(n147) );
    VMW_NAND2 U20 ( .A(n150), .B(B[10]), .Z(n149) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n152), .C(n147), .D(n142), .Z(n151) );
    VMW_NAND2 U22 ( .A(n152), .B(A[9]), .Z(n153) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U24 ( .A(n156), .B(B[12]), .Z(n155) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_NAND2 U26 ( .A(n158), .B(A[11]), .Z(n159) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_NAND2 U28 ( .A(n162), .B(B[14]), .Z(n161) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_NAND2 U30 ( .A(n164), .B(A[13]), .Z(n165) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n162), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n167), .C(n166), .D(n161), .Z(n118) );
    VMW_INV U33 ( .A(A[12]), .Z(n156) );
    VMW_INV U34 ( .A(B[7]), .Z(n145) );
    VMW_INV U35 ( .A(A[7]), .Z(n148) );
    VMW_INV U36 ( .A(A[3]), .Z(n134) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n150) );
    VMW_INV U39 ( .A(B[9]), .Z(n152) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n143) );
    VMW_INV U42 ( .A(A[14]), .Z(n162) );
    VMW_INV U43 ( .A(B[11]), .Z(n158) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n167) );
    VMW_INV U48 ( .A(B[13]), .Z(n164) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n117) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216;
    VMW_OAI21 U3 ( .A(B[15]), .B(n168), .C(n169), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n171), .B(B[2]), .Z(n170) );
    VMW_AO22 U5 ( .A(n173), .B(B[0]), .C(n174), .D(B[1]), .Z(n172) );
    VMW_OR2 U6 ( .A(B[2]), .B(n171), .Z(n175) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n174), .C(n175), .D(n172), .Z(n176) );
    VMW_NAND2 U8 ( .A(n178), .B(B[4]), .Z(n177) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n180), .C(n176), .D(n170), .Z(n179) );
    VMW_OR2 U10 ( .A(B[4]), .B(n178), .Z(n181) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n183), .C(n181), .D(n179), .Z(n182) );
    VMW_NAND2 U12 ( .A(n185), .B(B[6]), .Z(n184) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n187), .C(n182), .D(n177), .Z(n186) );
    VMW_OR2 U14 ( .A(B[6]), .B(n185), .Z(n188) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n190), .C(n188), .D(n186), .Z(n189) );
    VMW_NAND2 U16 ( .A(n192), .B(B[8]), .Z(n191) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n194), .C(n189), .D(n184), .Z(n193) );
    VMW_OR2 U18 ( .A(B[8]), .B(n192), .Z(n195) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n197), .C(n195), .D(n193), .Z(n196) );
    VMW_NAND2 U20 ( .A(n199), .B(B[10]), .Z(n198) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n201), .C(n196), .D(n191), .Z(n200) );
    VMW_NAND2 U22 ( .A(n201), .B(A[9]), .Z(n202) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n199), .C(n202), .D(n200), .Z(n203) );
    VMW_NAND2 U24 ( .A(n205), .B(B[12]), .Z(n204) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n207), .C(n203), .D(n198), .Z(n206) );
    VMW_NAND2 U26 ( .A(n207), .B(A[11]), .Z(n208) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n205), .C(n208), .D(n206), .Z(n209) );
    VMW_NAND2 U28 ( .A(n211), .B(B[14]), .Z(n210) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n213), .C(n209), .D(n204), .Z(n212) );
    VMW_NAND2 U30 ( .A(n213), .B(A[13]), .Z(n214) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n211), .C(n214), .D(n212), .Z(n215) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n216), .C(n215), .D(n210), .Z(n169) );
    VMW_INV U33 ( .A(A[12]), .Z(n205) );
    VMW_INV U34 ( .A(B[7]), .Z(n194) );
    VMW_INV U35 ( .A(A[7]), .Z(n197) );
    VMW_INV U36 ( .A(A[3]), .Z(n183) );
    VMW_INV U37 ( .A(B[3]), .Z(n180) );
    VMW_INV U38 ( .A(A[10]), .Z(n199) );
    VMW_INV U39 ( .A(B[9]), .Z(n201) );
    VMW_INV U40 ( .A(A[4]), .Z(n178) );
    VMW_INV U41 ( .A(A[8]), .Z(n192) );
    VMW_INV U42 ( .A(A[14]), .Z(n211) );
    VMW_INV U43 ( .A(B[11]), .Z(n207) );
    VMW_INV U44 ( .A(A[5]), .Z(n190) );
    VMW_INV U45 ( .A(B[5]), .Z(n187) );
    VMW_INV U46 ( .A(A[1]), .Z(n174) );
    VMW_INV U47 ( .A(B[15]), .Z(n216) );
    VMW_INV U48 ( .A(B[13]), .Z(n213) );
    VMW_INV U49 ( .A(A[6]), .Z(n185) );
    VMW_INV U50 ( .A(A[2]), .Z(n171) );
    VMW_INV U51 ( .A(A[0]), .Z(n173) );
    VMW_INV U52 ( .A(A[15]), .Z(n168) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265;
    VMW_OAI21 U3 ( .A(B[15]), .B(n217), .C(n218), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n220), .B(B[2]), .Z(n219) );
    VMW_AO22 U5 ( .A(n222), .B(B[0]), .C(n223), .D(B[1]), .Z(n221) );
    VMW_OR2 U6 ( .A(B[2]), .B(n220), .Z(n224) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n223), .C(n224), .D(n221), .Z(n225) );
    VMW_NAND2 U8 ( .A(n227), .B(B[4]), .Z(n226) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n229), .C(n225), .D(n219), .Z(n228) );
    VMW_OR2 U10 ( .A(B[4]), .B(n227), .Z(n230) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n232), .C(n230), .D(n228), .Z(n231) );
    VMW_NAND2 U12 ( .A(n234), .B(B[6]), .Z(n233) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n236), .C(n231), .D(n226), .Z(n235) );
    VMW_OR2 U14 ( .A(B[6]), .B(n234), .Z(n237) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n239), .C(n237), .D(n235), .Z(n238) );
    VMW_NAND2 U16 ( .A(n241), .B(B[8]), .Z(n240) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n243), .C(n238), .D(n233), .Z(n242) );
    VMW_OR2 U18 ( .A(B[8]), .B(n241), .Z(n244) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n246), .C(n244), .D(n242), .Z(n245) );
    VMW_NAND2 U20 ( .A(n248), .B(B[10]), .Z(n247) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n250), .C(n245), .D(n240), .Z(n249) );
    VMW_NAND2 U22 ( .A(n250), .B(A[9]), .Z(n251) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n248), .C(n251), .D(n249), .Z(n252) );
    VMW_NAND2 U24 ( .A(n254), .B(B[12]), .Z(n253) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n256), .C(n252), .D(n247), .Z(n255) );
    VMW_NAND2 U26 ( .A(n256), .B(A[11]), .Z(n257) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n254), .C(n257), .D(n255), .Z(n258) );
    VMW_NAND2 U28 ( .A(n260), .B(B[14]), .Z(n259) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n262), .C(n258), .D(n253), .Z(n261) );
    VMW_NAND2 U30 ( .A(n262), .B(A[13]), .Z(n263) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n260), .C(n263), .D(n261), .Z(n264) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n265), .C(n264), .D(n259), .Z(n218) );
    VMW_INV U33 ( .A(A[12]), .Z(n254) );
    VMW_INV U34 ( .A(B[7]), .Z(n243) );
    VMW_INV U35 ( .A(A[7]), .Z(n246) );
    VMW_INV U36 ( .A(A[3]), .Z(n232) );
    VMW_INV U37 ( .A(B[3]), .Z(n229) );
    VMW_INV U38 ( .A(A[10]), .Z(n248) );
    VMW_INV U39 ( .A(B[9]), .Z(n250) );
    VMW_INV U40 ( .A(A[4]), .Z(n227) );
    VMW_INV U41 ( .A(A[8]), .Z(n241) );
    VMW_INV U42 ( .A(A[14]), .Z(n260) );
    VMW_INV U43 ( .A(B[11]), .Z(n256) );
    VMW_INV U44 ( .A(A[5]), .Z(n239) );
    VMW_INV U45 ( .A(B[5]), .Z(n236) );
    VMW_INV U46 ( .A(A[1]), .Z(n223) );
    VMW_INV U47 ( .A(B[15]), .Z(n265) );
    VMW_INV U48 ( .A(B[13]), .Z(n262) );
    VMW_INV U49 ( .A(A[6]), .Z(n234) );
    VMW_INV U50 ( .A(A[2]), .Z(n220) );
    VMW_INV U51 ( .A(A[0]), .Z(n222) );
    VMW_INV U52 ( .A(A[15]), .Z(n217) );
endmodule


module NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314;
    VMW_OAI21 U3 ( .A(B[15]), .B(n266), .C(n267), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n269), .B(B[2]), .Z(n268) );
    VMW_AO22 U5 ( .A(n271), .B(B[0]), .C(n272), .D(B[1]), .Z(n270) );
    VMW_OR2 U6 ( .A(B[2]), .B(n269), .Z(n273) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n272), .C(n273), .D(n270), .Z(n274) );
    VMW_NAND2 U8 ( .A(n276), .B(B[4]), .Z(n275) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n278), .C(n274), .D(n268), .Z(n277) );
    VMW_OR2 U10 ( .A(B[4]), .B(n276), .Z(n279) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n281), .C(n279), .D(n277), .Z(n280) );
    VMW_NAND2 U12 ( .A(n283), .B(B[6]), .Z(n282) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n285), .C(n280), .D(n275), .Z(n284) );
    VMW_OR2 U14 ( .A(B[6]), .B(n283), .Z(n286) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n288), .C(n286), .D(n284), .Z(n287) );
    VMW_NAND2 U16 ( .A(n290), .B(B[8]), .Z(n289) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n292), .C(n287), .D(n282), .Z(n291) );
    VMW_OR2 U18 ( .A(B[8]), .B(n290), .Z(n293) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n295), .C(n293), .D(n291), .Z(n294) );
    VMW_NAND2 U20 ( .A(n297), .B(B[10]), .Z(n296) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n299), .C(n294), .D(n289), .Z(n298) );
    VMW_NAND2 U22 ( .A(n299), .B(A[9]), .Z(n300) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n297), .C(n300), .D(n298), .Z(n301) );
    VMW_NAND2 U24 ( .A(n303), .B(B[12]), .Z(n302) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n305), .C(n301), .D(n296), .Z(n304) );
    VMW_NAND2 U26 ( .A(n305), .B(A[11]), .Z(n306) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n303), .C(n306), .D(n304), .Z(n307) );
    VMW_NAND2 U28 ( .A(n309), .B(B[14]), .Z(n308) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n311), .C(n307), .D(n302), .Z(n310) );
    VMW_NAND2 U30 ( .A(n311), .B(A[13]), .Z(n312) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n309), .C(n312), .D(n310), .Z(n313) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n314), .C(n313), .D(n308), .Z(n267) );
    VMW_INV U33 ( .A(A[12]), .Z(n303) );
    VMW_INV U34 ( .A(B[7]), .Z(n292) );
    VMW_INV U35 ( .A(A[7]), .Z(n295) );
    VMW_INV U36 ( .A(A[3]), .Z(n281) );
    VMW_INV U37 ( .A(B[3]), .Z(n278) );
    VMW_INV U38 ( .A(A[10]), .Z(n297) );
    VMW_INV U39 ( .A(B[9]), .Z(n299) );
    VMW_INV U40 ( .A(A[4]), .Z(n276) );
    VMW_INV U41 ( .A(A[8]), .Z(n290) );
    VMW_INV U42 ( .A(A[14]), .Z(n309) );
    VMW_INV U43 ( .A(B[11]), .Z(n305) );
    VMW_INV U44 ( .A(A[5]), .Z(n288) );
    VMW_INV U45 ( .A(B[5]), .Z(n285) );
    VMW_INV U46 ( .A(A[1]), .Z(n272) );
    VMW_INV U47 ( .A(B[15]), .Z(n314) );
    VMW_INV U48 ( .A(B[13]), .Z(n311) );
    VMW_INV U49 ( .A(A[6]), .Z(n283) );
    VMW_INV U50 ( .A(A[2]), .Z(n269) );
    VMW_INV U51 ( .A(A[0]), .Z(n271) );
    VMW_INV U52 ( .A(A[15]), .Z(n266) );
endmodule


module NodeAux_INDEGREE6_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \temp494[7] , \temp584[2] , n100, \OutEdge146[7] , \temp314[15] , 
        \OutEdge146[12] , \temp314[11] , \OutEdge146[3] , \temp494[3] , 
        \temp584[6] , \path[2] , \path[0] , \temp314[13] , \temp494[1] , 
        \OutEdge146[1] , \temp584[4] , \OutEdge146[8] , \temp494[8] , n132, 
        \OutEdge146[10] , \temp584[0] , \OutEdge146[5] , \temp494[5] , 
        \OutEdge146[14] , \temp584[9] , \temp220[10] , \temp220[4] , 
        \temp314[7] , \temp494[11] , \temp404[6] , \temp584[13] , 
        \temp404[11] , \temp404[2] , \temp220[0] , \temp314[3] , \temp494[15] , 
        \temp220[14] , \temp404[15] , \temp220[9] , \temp404[9] , \temp314[8] , 
        \temp220[2] , \temp404[0] , \temp314[1] , \temp584[15] , n108, 
        \temp404[13] , \temp584[11] , \temp220[12] , \temp220[6] , 
        \temp314[5] , \temp404[4] , \temp494[13] , \temp404[12] , 
        \temp584[10] , \temp220[7] , \temp314[4] , n124, \temp494[12] , 
        \temp220[13] , \temp404[5] , \temp404[8] , \temp314[9] , \temp404[1] , 
        \temp220[3] , \temp314[0] , \temp584[14] , \temp404[3] , \temp220[15] , 
        \temp220[1] , \temp314[2] , \temp494[14] , \temp220[8] , \temp404[14] , 
        n116, \temp220[5] , \temp314[6] , \temp494[10] , \temp220[11] , 
        \temp404[7] , \temp584[12] , \temp404[10] , \temp584[1] , 
        \OutEdge146[4] , \temp494[4] , \OutEdge146[15] , \temp584[8] , 
        \path[1] , \temp494[0] , \OutEdge146[0] , \temp314[12] , n92, 
        \temp584[5] , \OutEdge146[9] , \temp494[9] , \OutEdge146[11] , 
        \OutEdge146[13] , \temp494[2] , \OutEdge146[2] , \temp314[10] , 
        \temp584[7] , \temp584[3] , \temp314[14] , \temp494[6] , 
        \OutEdge146[6] , n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
        n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
        n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
        n812, n813, n814, n815, n816;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U91 ( .Z(n815) );
    VMW_PULLDOWN U92 ( .Z(n814) );
    VMW_PULLDOWN U93 ( .Z(n813) );
    VMW_PULLDOWN U94 ( .Z(n812) );
    VMW_PULLDOWN U95 ( .Z(n816) );
    VMW_PULLDOWN U96 ( .Z(n811) );
    VMW_NOR2 U97 ( .A(Start), .B(n767), .Z(\OutEdge146[15] ) );
    VMW_NAND2 U98 ( .A(n768), .B(n769), .Z(\OutEdge146[14] ) );
    VMW_NAND2 U99 ( .A(n770), .B(n769), .Z(\OutEdge146[13] ) );
    VMW_NAND2 U100 ( .A(n771), .B(n769), .Z(\OutEdge146[12] ) );
    VMW_NAND2 U101 ( .A(n772), .B(n769), .Z(\OutEdge146[11] ) );
    VMW_NAND2 U102 ( .A(n773), .B(n769), .Z(\OutEdge146[10] ) );
    VMW_NAND2 U103 ( .A(n774), .B(n769), .Z(\OutEdge146[9] ) );
    VMW_NAND2 U104 ( .A(n775), .B(n769), .Z(\OutEdge146[8] ) );
    VMW_NAND2 U105 ( .A(n776), .B(n769), .Z(\OutEdge146[7] ) );
    VMW_NAND2 U106 ( .A(n777), .B(n769), .Z(\OutEdge146[6] ) );
    VMW_NAND2 U107 ( .A(n778), .B(n769), .Z(\OutEdge146[5] ) );
    VMW_NAND2 U108 ( .A(n779), .B(n769), .Z(\OutEdge146[4] ) );
    VMW_NAND2 U109 ( .A(n780), .B(n769), .Z(\OutEdge146[3] ) );
    VMW_NAND2 U110 ( .A(n781), .B(n769), .Z(\OutEdge146[2] ) );
    VMW_NAND2 U111 ( .A(n782), .B(n769), .Z(\OutEdge146[1] ) );
    VMW_NAND2 U112 ( .A(n783), .B(n769), .Z(\OutEdge146[0] ) );
    VMW_AND4 U113 ( .A(n785), .B(n786), .C(n787), .D(n788), .Z(n784) );
    VMW_OR3 U114 ( .A(n784), .B(n124), .C(n132), .Z(n789) );
    VMW_OR2 U115 ( .A(n132), .B(n791), .Z(n790) );
    VMW_AO22 U116 ( .A(\temp494[15] ), .B(n792), .C(InEdges[79]), .D(n124), 
        .Z(\temp584[15] ) );
    VMW_OAI22 U117 ( .A(\path[2] ), .B(n769), .C(n789), .D(Start), .Z(n793) );
    VMW_OAI22 U118 ( .A(\path[1] ), .B(n769), .C(n795), .D(Start), .Z(n794) );
    VMW_OAI22 U119 ( .A(\path[0] ), .B(n769), .C(n790), .D(Start), .Z(n796) );
    VMW_MUX2I U120 ( .A(\temp584[15] ), .B(InEdges[95]), .S(n132), .Z(n767) );
    VMW_AND4 U121 ( .A(n798), .B(n799), .C(n800), .D(n801), .Z(n797) );
    VMW_INV U122 ( .A(Start), .Z(n769) );
    VMW_INV U123 ( .A(n116), .Z(n786) );
    VMW_AOI211 U124 ( .A(n785), .B(n787), .C(n108), .D(n116), .Z(n802) );
    VMW_OAI21 U125 ( .A(n100), .B(n785), .C(n788), .Z(n803) );
    VMW_AOI21 U126 ( .A(n786), .B(n803), .C(n124), .Z(n791) );
    VMW_AND4 U127 ( .A(n804), .B(n805), .C(n806), .D(n797), .Z(n807) );
    VMW_XNOR2 U128 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n801) );
    VMW_XNOR2 U129 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n800) );
    VMW_XNOR2 U130 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n799) );
    VMW_XNOR2 U131 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n798) );
    VMW_XNOR2 U132 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n805) );
    VMW_XNOR2 U133 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n804) );
    VMW_XNOR2 U134 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n806) );
    VMW_AO22 U135 ( .A(OutEdge[9]), .B(n785), .C(InEdges[9]), .D(n92), .Z(
        \temp220[9] ) );
    VMW_AO22 U136 ( .A(\temp220[9] ), .B(n787), .C(InEdges[25]), .D(n100), .Z(
        \temp314[9] ) );
    VMW_AO22 U137 ( .A(\temp314[9] ), .B(n788), .C(InEdges[41]), .D(n108), .Z(
        \temp404[9] ) );
    VMW_AO22 U138 ( .A(\temp404[9] ), .B(n786), .C(InEdges[57]), .D(n116), .Z(
        \temp494[9] ) );
    VMW_AO22 U139 ( .A(\temp494[9] ), .B(n792), .C(InEdges[73]), .D(n124), .Z(
        \temp584[9] ) );
    VMW_AO22 U140 ( .A(OutEdge[8]), .B(n785), .C(InEdges[8]), .D(n92), .Z(
        \temp220[8] ) );
    VMW_AO22 U141 ( .A(\temp220[8] ), .B(n787), .C(InEdges[24]), .D(n100), .Z(
        \temp314[8] ) );
    VMW_AO22 U142 ( .A(\temp314[8] ), .B(n788), .C(InEdges[40]), .D(n108), .Z(
        \temp404[8] ) );
    VMW_AO22 U143 ( .A(\temp404[8] ), .B(n786), .C(InEdges[56]), .D(n116), .Z(
        \temp494[8] ) );
    VMW_AO22 U144 ( .A(\temp494[8] ), .B(n792), .C(InEdges[72]), .D(n124), .Z(
        \temp584[8] ) );
    VMW_AO22 U145 ( .A(OutEdge[7]), .B(n785), .C(InEdges[7]), .D(n92), .Z(
        \temp220[7] ) );
    VMW_AO22 U146 ( .A(\temp220[7] ), .B(n787), .C(InEdges[23]), .D(n100), .Z(
        \temp314[7] ) );
    VMW_AO22 U147 ( .A(\temp314[7] ), .B(n788), .C(InEdges[39]), .D(n108), .Z(
        \temp404[7] ) );
    VMW_AO22 U148 ( .A(\temp404[7] ), .B(n786), .C(InEdges[55]), .D(n116), .Z(
        \temp494[7] ) );
    VMW_AO22 U149 ( .A(\temp494[7] ), .B(n792), .C(InEdges[71]), .D(n124), .Z(
        \temp584[7] ) );
    VMW_AO22 U150 ( .A(OutEdge[6]), .B(n785), .C(InEdges[6]), .D(n92), .Z(
        \temp220[6] ) );
    VMW_AO22 U151 ( .A(\temp220[6] ), .B(n787), .C(InEdges[22]), .D(n100), .Z(
        \temp314[6] ) );
    VMW_AO22 U152 ( .A(\temp314[6] ), .B(n788), .C(InEdges[38]), .D(n108), .Z(
        \temp404[6] ) );
    VMW_AO22 U153 ( .A(\temp404[6] ), .B(n786), .C(InEdges[54]), .D(n116), .Z(
        \temp494[6] ) );
    VMW_AO22 U154 ( .A(\temp494[6] ), .B(n792), .C(InEdges[70]), .D(n124), .Z(
        \temp584[6] ) );
    VMW_AO22 U155 ( .A(OutEdge[5]), .B(n785), .C(InEdges[5]), .D(n92), .Z(
        \temp220[5] ) );
    VMW_AO22 U156 ( .A(\temp220[5] ), .B(n787), .C(InEdges[21]), .D(n100), .Z(
        \temp314[5] ) );
    VMW_AO22 U157 ( .A(\temp314[5] ), .B(n788), .C(InEdges[37]), .D(n108), .Z(
        \temp404[5] ) );
    VMW_AO22 U158 ( .A(\temp404[5] ), .B(n786), .C(InEdges[53]), .D(n116), .Z(
        \temp494[5] ) );
    VMW_AO22 U159 ( .A(\temp494[5] ), .B(n792), .C(InEdges[69]), .D(n124), .Z(
        \temp584[5] ) );
    VMW_AO22 U160 ( .A(OutEdge[4]), .B(n785), .C(InEdges[4]), .D(n92), .Z(
        \temp220[4] ) );
    VMW_AO22 U161 ( .A(\temp220[4] ), .B(n787), .C(InEdges[20]), .D(n100), .Z(
        \temp314[4] ) );
    VMW_AO22 U162 ( .A(\temp314[4] ), .B(n788), .C(InEdges[36]), .D(n108), .Z(
        \temp404[4] ) );
    VMW_AO22 U163 ( .A(\temp404[4] ), .B(n786), .C(InEdges[52]), .D(n116), .Z(
        \temp494[4] ) );
    VMW_AO22 U164 ( .A(\temp494[4] ), .B(n792), .C(InEdges[68]), .D(n124), .Z(
        \temp584[4] ) );
    VMW_AO22 U165 ( .A(OutEdge[3]), .B(n785), .C(InEdges[3]), .D(n92), .Z(
        \temp220[3] ) );
    VMW_AO22 U166 ( .A(\temp220[3] ), .B(n787), .C(InEdges[19]), .D(n100), .Z(
        \temp314[3] ) );
    VMW_AO22 U167 ( .A(\temp314[3] ), .B(n788), .C(InEdges[35]), .D(n108), .Z(
        \temp404[3] ) );
    VMW_AO22 U168 ( .A(\temp404[3] ), .B(n786), .C(InEdges[51]), .D(n116), .Z(
        \temp494[3] ) );
    VMW_AO22 U169 ( .A(\temp494[3] ), .B(n792), .C(InEdges[67]), .D(n124), .Z(
        \temp584[3] ) );
    VMW_AO22 U170 ( .A(OutEdge[2]), .B(n785), .C(InEdges[2]), .D(n92), .Z(
        \temp220[2] ) );
    VMW_AO22 U171 ( .A(\temp220[2] ), .B(n787), .C(InEdges[18]), .D(n100), .Z(
        \temp314[2] ) );
    VMW_AO22 U172 ( .A(\temp314[2] ), .B(n788), .C(InEdges[34]), .D(n108), .Z(
        \temp404[2] ) );
    VMW_AO22 U173 ( .A(\temp404[2] ), .B(n786), .C(InEdges[50]), .D(n116), .Z(
        \temp494[2] ) );
    VMW_AO22 U174 ( .A(\temp494[2] ), .B(n792), .C(InEdges[66]), .D(n124), .Z(
        \temp584[2] ) );
    VMW_AO22 U175 ( .A(OutEdge[1]), .B(n785), .C(InEdges[1]), .D(n92), .Z(
        \temp220[1] ) );
    VMW_AO22 U176 ( .A(\temp220[1] ), .B(n787), .C(InEdges[17]), .D(n100), .Z(
        \temp314[1] ) );
    VMW_AO22 U177 ( .A(\temp314[1] ), .B(n788), .C(InEdges[33]), .D(n108), .Z(
        \temp404[1] ) );
    VMW_AO22 U178 ( .A(\temp404[1] ), .B(n786), .C(InEdges[49]), .D(n116), .Z(
        \temp494[1] ) );
    VMW_AO22 U179 ( .A(\temp494[1] ), .B(n792), .C(InEdges[65]), .D(n124), .Z(
        \temp584[1] ) );
    VMW_AO22 U180 ( .A(OutEdge[15]), .B(n785), .C(InEdges[15]), .D(n92), .Z(
        \temp220[15] ) );
    VMW_AO22 U181 ( .A(\temp220[15] ), .B(n787), .C(InEdges[31]), .D(n100), 
        .Z(\temp314[15] ) );
    VMW_AO22 U182 ( .A(\temp314[15] ), .B(n788), .C(InEdges[47]), .D(n108), 
        .Z(\temp404[15] ) );
    VMW_AO22 U183 ( .A(\temp404[15] ), .B(n786), .C(InEdges[63]), .D(n116), 
        .Z(\temp494[15] ) );
    VMW_AO22 U184 ( .A(OutEdge[14]), .B(n785), .C(InEdges[14]), .D(n92), .Z(
        \temp220[14] ) );
    VMW_AO22 U185 ( .A(\temp220[14] ), .B(n787), .C(InEdges[30]), .D(n100), 
        .Z(\temp314[14] ) );
    VMW_AO22 U186 ( .A(\temp314[14] ), .B(n788), .C(InEdges[46]), .D(n108), 
        .Z(\temp404[14] ) );
    VMW_AO22 U187 ( .A(\temp404[14] ), .B(n786), .C(InEdges[62]), .D(n116), 
        .Z(\temp494[14] ) );
    VMW_AO22 U188 ( .A(\temp494[14] ), .B(n792), .C(InEdges[78]), .D(n124), 
        .Z(\temp584[14] ) );
    VMW_AO22 U189 ( .A(OutEdge[13]), .B(n785), .C(InEdges[13]), .D(n92), .Z(
        \temp220[13] ) );
    VMW_AO22 U190 ( .A(\temp220[13] ), .B(n787), .C(InEdges[29]), .D(n100), 
        .Z(\temp314[13] ) );
    VMW_AO22 U191 ( .A(\temp314[13] ), .B(n788), .C(InEdges[45]), .D(n108), 
        .Z(\temp404[13] ) );
    VMW_AO22 U192 ( .A(\temp404[13] ), .B(n786), .C(InEdges[61]), .D(n116), 
        .Z(\temp494[13] ) );
    VMW_AO22 U193 ( .A(\temp494[13] ), .B(n792), .C(InEdges[77]), .D(n124), 
        .Z(\temp584[13] ) );
    VMW_AO22 U194 ( .A(OutEdge[12]), .B(n785), .C(InEdges[12]), .D(n92), .Z(
        \temp220[12] ) );
    VMW_AO22 U195 ( .A(\temp220[12] ), .B(n787), .C(InEdges[28]), .D(n100), 
        .Z(\temp314[12] ) );
    VMW_AO22 U196 ( .A(\temp314[12] ), .B(n788), .C(InEdges[44]), .D(n108), 
        .Z(\temp404[12] ) );
    VMW_AO22 U197 ( .A(\temp404[12] ), .B(n786), .C(InEdges[60]), .D(n116), 
        .Z(\temp494[12] ) );
    VMW_AO22 U198 ( .A(\temp494[12] ), .B(n792), .C(InEdges[76]), .D(n124), 
        .Z(\temp584[12] ) );
    VMW_AO22 U199 ( .A(OutEdge[11]), .B(n785), .C(InEdges[11]), .D(n92), .Z(
        \temp220[11] ) );
    VMW_AO22 U200 ( .A(\temp220[11] ), .B(n787), .C(InEdges[27]), .D(n100), 
        .Z(\temp314[11] ) );
    VMW_AO22 U201 ( .A(\temp314[11] ), .B(n788), .C(InEdges[43]), .D(n108), 
        .Z(\temp404[11] ) );
    VMW_AO22 U202 ( .A(\temp404[11] ), .B(n786), .C(InEdges[59]), .D(n116), 
        .Z(\temp494[11] ) );
    VMW_AO22 U203 ( .A(\temp494[11] ), .B(n792), .C(InEdges[75]), .D(n124), 
        .Z(\temp584[11] ) );
    VMW_AO22 U204 ( .A(OutEdge[10]), .B(n785), .C(InEdges[10]), .D(n92), .Z(
        \temp220[10] ) );
    VMW_AO22 U205 ( .A(\temp220[10] ), .B(n787), .C(InEdges[26]), .D(n100), 
        .Z(\temp314[10] ) );
    VMW_AO22 U206 ( .A(\temp314[10] ), .B(n788), .C(InEdges[42]), .D(n108), 
        .Z(\temp404[10] ) );
    VMW_AO22 U207 ( .A(\temp404[10] ), .B(n786), .C(InEdges[58]), .D(n116), 
        .Z(\temp494[10] ) );
    VMW_AO22 U208 ( .A(\temp494[10] ), .B(n792), .C(InEdges[74]), .D(n124), 
        .Z(\temp584[10] ) );
    VMW_AO22 U209 ( .A(OutEdge[0]), .B(n785), .C(InEdges[0]), .D(n92), .Z(
        \temp220[0] ) );
    VMW_AO22 U210 ( .A(\temp220[0] ), .B(n787), .C(InEdges[16]), .D(n100), .Z(
        \temp314[0] ) );
    VMW_AO22 U211 ( .A(\temp314[0] ), .B(n788), .C(InEdges[32]), .D(n108), .Z(
        \temp404[0] ) );
    VMW_AO22 U212 ( .A(\temp404[0] ), .B(n786), .C(InEdges[48]), .D(n116), .Z(
        \temp494[0] ) );
    VMW_AO22 U213 ( .A(\temp494[0] ), .B(n792), .C(InEdges[64]), .D(n124), .Z(
        \temp584[0] ) );
    VMW_NOR3 U214 ( .A(n132), .B(n124), .C(n802), .Z(n795) );
    VMW_MUX2I U215 ( .A(\temp584[9] ), .B(InEdges[89]), .S(n132), .Z(n774) );
    VMW_MUX2I U216 ( .A(\temp584[8] ), .B(InEdges[88]), .S(n132), .Z(n775) );
    VMW_MUX2I U217 ( .A(\temp584[7] ), .B(InEdges[87]), .S(n132), .Z(n776) );
    VMW_MUX2I U218 ( .A(\temp584[6] ), .B(InEdges[86]), .S(n132), .Z(n777) );
    VMW_MUX2I U219 ( .A(\temp584[5] ), .B(InEdges[85]), .S(n132), .Z(n778) );
    VMW_MUX2I U220 ( .A(\temp584[4] ), .B(InEdges[84]), .S(n132), .Z(n779) );
    VMW_MUX2I U221 ( .A(\temp584[3] ), .B(InEdges[83]), .S(n132), .Z(n780) );
    VMW_MUX2I U222 ( .A(\temp584[2] ), .B(InEdges[82]), .S(n132), .Z(n781) );
    VMW_MUX2I U223 ( .A(\temp584[1] ), .B(InEdges[81]), .S(n132), .Z(n782) );
    VMW_MUX2I U224 ( .A(\temp584[14] ), .B(InEdges[94]), .S(n132), .Z(n768) );
    VMW_MUX2I U225 ( .A(\temp584[13] ), .B(InEdges[93]), .S(n132), .Z(n770) );
    VMW_MUX2I U226 ( .A(\temp584[12] ), .B(InEdges[92]), .S(n132), .Z(n771) );
    VMW_MUX2I U227 ( .A(\temp584[11] ), .B(InEdges[91]), .S(n132), .Z(n772) );
    VMW_MUX2I U228 ( .A(\temp584[10] ), .B(InEdges[90]), .S(n132), .Z(n773) );
    VMW_MUX2I U229 ( .A(\temp584[0] ), .B(InEdges[80]), .S(n132), .Z(n783) );
    VMW_INV U230 ( .A(n100), .Z(n787) );
    VMW_INV U231 ( .A(n92), .Z(n785) );
    VMW_INV U232 ( .A(n108), .Z(n788) );
    VMW_INV U233 ( .A(n124), .Z(n792) );
    VMW_INV U234 ( .A(n793), .Z(n809) );
    VMW_INV U235 ( .A(n794), .Z(n810) );
    VMW_INV U236 ( .A(n796), .Z(n808) );
    VMW_BUFIZ U237 ( .A(\path[1] ), .E(n807), .Z(\PathData[1] ) );
    VMW_BUFIZ U238 ( .A(\path[0] ), .E(n807), .Z(\PathData[0] ) );
    VMW_BUFIZ U239 ( .A(\path[2] ), .E(n807), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n808), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n809), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n810), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge146[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge146[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge146[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge146[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge146[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge146[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge146[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge146[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge146[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge146[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge146[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge146[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge146[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge146[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge146[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge146[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_5 lte_55_1 ( .A({\temp220[15] , 
        \temp220[14] , \temp220[13] , \temp220[12] , \temp220[11] , 
        \temp220[10] , \temp220[9] , \temp220[8] , \temp220[7] , \temp220[6] , 
        \temp220[5] , \temp220[4] , \temp220[3] , \temp220[2] , \temp220[1] , 
        \temp220[0] }), .B(InEdges[31:16]), .LEQ(n816), .TC(n816), .GE_GT(n100
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_4 lte_55_5 ( .A({\temp584[15] , 
        \temp584[14] , \temp584[13] , \temp584[12] , \temp584[11] , 
        \temp584[10] , \temp584[9] , \temp584[8] , \temp584[7] , \temp584[6] , 
        \temp584[5] , \temp584[4] , \temp584[3] , \temp584[2] , \temp584[1] , 
        \temp584[0] }), .B(InEdges[95:80]), .LEQ(n815), .TC(n815), .GE_GT(n132
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_3 lte_55_4 ( .A({\temp494[15] , 
        \temp494[14] , \temp494[13] , \temp494[12] , \temp494[11] , 
        \temp494[10] , \temp494[9] , \temp494[8] , \temp494[7] , \temp494[6] , 
        \temp494[5] , \temp494[4] , \temp494[3] , \temp494[2] , \temp494[1] , 
        \temp494[0] }), .B(InEdges[79:64]), .LEQ(n814), .TC(n814), .GE_GT(n124
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_2 lte_55_3 ( .A({\temp404[15] , 
        \temp404[14] , \temp404[13] , \temp404[12] , \temp404[11] , 
        \temp404[10] , \temp404[9] , \temp404[8] , \temp404[7] , \temp404[6] , 
        \temp404[5] , \temp404[4] , \temp404[3] , \temp404[2] , \temp404[1] , 
        \temp404[0] }), .B(InEdges[63:48]), .LEQ(n813), .TC(n813), .GE_GT(n116
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp314[15] , 
        \temp314[14] , \temp314[13] , \temp314[12] , \temp314[11] , 
        \temp314[10] , \temp314[9] , \temp314[8] , \temp314[7] , \temp314[6] , 
        \temp314[5] , \temp314[4] , \temp314[3] , \temp314[2] , \temp314[1] , 
        \temp314[0] }), .B(InEdges[47:32]), .LEQ(n812), .TC(n812), .GE_GT(n108
        ) );
    NodeAux_INDEGREE6_SOURCE0_DW01_cmp2_16_0 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n811), .TC(n811), .GE_GT(n92) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63;
    VMW_OAI21 U3 ( .A(B[15]), .B(n15), .C(n16), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n18), .B(B[2]), .Z(n17) );
    VMW_AO22 U5 ( .A(n20), .B(B[0]), .C(n21), .D(B[1]), .Z(n19) );
    VMW_OR2 U6 ( .A(B[2]), .B(n18), .Z(n22) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n21), .C(n22), .D(n19), .Z(n23) );
    VMW_NAND2 U8 ( .A(n25), .B(B[4]), .Z(n24) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n27), .C(n23), .D(n17), .Z(n26) );
    VMW_OR2 U10 ( .A(B[4]), .B(n25), .Z(n28) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n30), .C(n28), .D(n26), .Z(n29) );
    VMW_NAND2 U12 ( .A(n32), .B(B[6]), .Z(n31) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n34), .C(n29), .D(n24), .Z(n33) );
    VMW_OR2 U14 ( .A(B[6]), .B(n32), .Z(n35) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n37), .C(n35), .D(n33), .Z(n36) );
    VMW_NAND2 U16 ( .A(n39), .B(B[8]), .Z(n38) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n41), .C(n36), .D(n31), .Z(n40) );
    VMW_OR2 U18 ( .A(B[8]), .B(n39), .Z(n42) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n44), .C(n42), .D(n40), .Z(n43) );
    VMW_NAND2 U20 ( .A(n46), .B(B[10]), .Z(n45) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n48), .C(n43), .D(n38), .Z(n47) );
    VMW_NAND2 U22 ( .A(n48), .B(A[9]), .Z(n49) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n46), .C(n49), .D(n47), .Z(n50) );
    VMW_NAND2 U24 ( .A(n52), .B(B[12]), .Z(n51) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n54), .C(n50), .D(n45), .Z(n53) );
    VMW_NAND2 U26 ( .A(n54), .B(A[11]), .Z(n55) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n52), .C(n55), .D(n53), .Z(n56) );
    VMW_NAND2 U28 ( .A(n58), .B(B[14]), .Z(n57) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n60), .C(n56), .D(n51), .Z(n59) );
    VMW_NAND2 U30 ( .A(n60), .B(A[13]), .Z(n61) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n58), .C(n61), .D(n59), .Z(n62) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n63), .C(n62), .D(n57), .Z(n16) );
    VMW_INV U33 ( .A(A[12]), .Z(n52) );
    VMW_INV U34 ( .A(B[7]), .Z(n41) );
    VMW_INV U35 ( .A(A[7]), .Z(n44) );
    VMW_INV U36 ( .A(A[3]), .Z(n30) );
    VMW_INV U37 ( .A(B[3]), .Z(n27) );
    VMW_INV U38 ( .A(A[10]), .Z(n46) );
    VMW_INV U39 ( .A(B[9]), .Z(n48) );
    VMW_INV U40 ( .A(A[4]), .Z(n25) );
    VMW_INV U41 ( .A(A[8]), .Z(n39) );
    VMW_INV U42 ( .A(A[14]), .Z(n58) );
    VMW_INV U43 ( .A(B[11]), .Z(n54) );
    VMW_INV U44 ( .A(A[5]), .Z(n37) );
    VMW_INV U45 ( .A(B[5]), .Z(n34) );
    VMW_INV U46 ( .A(A[1]), .Z(n21) );
    VMW_INV U47 ( .A(B[15]), .Z(n63) );
    VMW_INV U48 ( .A(B[13]), .Z(n60) );
    VMW_INV U49 ( .A(A[6]), .Z(n32) );
    VMW_INV U50 ( .A(A[2]), .Z(n18) );
    VMW_INV U51 ( .A(A[0]), .Z(n20) );
    VMW_INV U52 ( .A(A[15]), .Z(n15) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, 
        n107, n108, n109, n111, n112, n113, n114, n115;
    VMW_OAI21 U3 ( .A(B[15]), .B(n64), .C(n65), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n67), .B(B[2]), .Z(n66) );
    VMW_AO22 U5 ( .A(n69), .B(B[0]), .C(n70), .D(B[1]), .Z(n68) );
    VMW_OR2 U6 ( .A(B[2]), .B(n67), .Z(n71) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n70), .C(n71), .D(n68), .Z(n72) );
    VMW_NAND2 U8 ( .A(n74), .B(B[4]), .Z(n73) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n76), .C(n72), .D(n66), .Z(n75) );
    VMW_OR2 U10 ( .A(B[4]), .B(n74), .Z(n77) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n79), .C(n77), .D(n75), .Z(n78) );
    VMW_NAND2 U12 ( .A(n81), .B(B[6]), .Z(n80) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n83), .C(n78), .D(n73), .Z(n82) );
    VMW_OR2 U14 ( .A(B[6]), .B(n81), .Z(n84) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n86), .C(n84), .D(n82), .Z(n85) );
    VMW_NAND2 U16 ( .A(n88), .B(B[8]), .Z(n87) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n90), .C(n85), .D(n80), .Z(n89) );
    VMW_OR2 U18 ( .A(B[8]), .B(n88), .Z(n91) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n93), .C(n91), .D(n89), .Z(n92) );
    VMW_NAND2 U20 ( .A(n96), .B(B[10]), .Z(n95) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n98), .C(n92), .D(n87), .Z(n97) );
    VMW_NAND2 U22 ( .A(n98), .B(A[9]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n96), .C(n99), .D(n97), .Z(n100) );
    VMW_NAND2 U24 ( .A(n103), .B(B[12]), .Z(n101) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_NAND2 U26 ( .A(n105), .B(A[11]), .Z(n106) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n103), .C(n106), .D(n104), .Z(n107) );
    VMW_NAND2 U28 ( .A(n109), .B(B[14]), .Z(n108) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n112), .C(n107), .D(n101), .Z(n111) );
    VMW_NAND2 U30 ( .A(n112), .B(A[13]), .Z(n113) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n109), .C(n113), .D(n111), .Z(n114) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n115), .C(n114), .D(n108), .Z(n65) );
    VMW_INV U33 ( .A(A[12]), .Z(n103) );
    VMW_INV U34 ( .A(B[7]), .Z(n90) );
    VMW_INV U35 ( .A(A[7]), .Z(n93) );
    VMW_INV U36 ( .A(A[3]), .Z(n79) );
    VMW_INV U37 ( .A(B[3]), .Z(n76) );
    VMW_INV U38 ( .A(A[10]), .Z(n96) );
    VMW_INV U39 ( .A(B[9]), .Z(n98) );
    VMW_INV U40 ( .A(A[4]), .Z(n74) );
    VMW_INV U41 ( .A(A[8]), .Z(n88) );
    VMW_INV U42 ( .A(A[14]), .Z(n109) );
    VMW_INV U43 ( .A(B[11]), .Z(n105) );
    VMW_INV U44 ( .A(A[5]), .Z(n86) );
    VMW_INV U45 ( .A(B[5]), .Z(n83) );
    VMW_INV U46 ( .A(A[1]), .Z(n70) );
    VMW_INV U47 ( .A(B[15]), .Z(n115) );
    VMW_INV U48 ( .A(B[13]), .Z(n112) );
    VMW_INV U49 ( .A(A[6]), .Z(n81) );
    VMW_INV U50 ( .A(A[2]), .Z(n67) );
    VMW_INV U51 ( .A(A[0]), .Z(n69) );
    VMW_INV U52 ( .A(A[15]), .Z(n64) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n117, n119, n120, n121, n122, n123, n124, n125, n127, n128, 
        n129, n130, n131, n132, n133, n135, n136, n137, n138, n139, n140, n141, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168;
    VMW_OAI21 U3 ( .A(B[15]), .B(n116), .C(n117), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n120), .B(B[2]), .Z(n119) );
    VMW_AO22 U5 ( .A(n122), .B(B[0]), .C(n123), .D(B[1]), .Z(n121) );
    VMW_OR2 U6 ( .A(B[2]), .B(n120), .Z(n124) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n123), .C(n124), .D(n121), .Z(n125) );
    VMW_NAND2 U8 ( .A(n128), .B(B[4]), .Z(n127) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n130), .C(n125), .D(n119), .Z(n129) );
    VMW_OR2 U10 ( .A(B[4]), .B(n128), .Z(n131) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n133), .C(n131), .D(n129), .Z(n132) );
    VMW_NAND2 U12 ( .A(n136), .B(B[6]), .Z(n135) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n138), .C(n132), .D(n127), .Z(n137) );
    VMW_OR2 U14 ( .A(B[6]), .B(n136), .Z(n139) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n141), .C(n139), .D(n137), .Z(n140) );
    VMW_NAND2 U16 ( .A(n144), .B(B[8]), .Z(n143) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n146), .C(n140), .D(n135), .Z(n145) );
    VMW_OR2 U18 ( .A(B[8]), .B(n144), .Z(n147) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n149), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U20 ( .A(n151), .B(B[10]), .Z(n150) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n153), .C(n148), .D(n143), .Z(n152) );
    VMW_NAND2 U22 ( .A(n153), .B(A[9]), .Z(n154) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U24 ( .A(n157), .B(B[12]), .Z(n156) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_NAND2 U26 ( .A(n159), .B(A[11]), .Z(n160) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_NAND2 U28 ( .A(n163), .B(B[14]), .Z(n162) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_NAND2 U30 ( .A(n165), .B(A[13]), .Z(n166) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n163), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n168), .C(n167), .D(n162), .Z(n117) );
    VMW_INV U33 ( .A(A[12]), .Z(n157) );
    VMW_INV U34 ( .A(B[7]), .Z(n146) );
    VMW_INV U35 ( .A(A[7]), .Z(n149) );
    VMW_INV U36 ( .A(A[3]), .Z(n133) );
    VMW_INV U37 ( .A(B[3]), .Z(n130) );
    VMW_INV U38 ( .A(A[10]), .Z(n151) );
    VMW_INV U39 ( .A(B[9]), .Z(n153) );
    VMW_INV U40 ( .A(A[4]), .Z(n128) );
    VMW_INV U41 ( .A(A[8]), .Z(n144) );
    VMW_INV U42 ( .A(A[14]), .Z(n163) );
    VMW_INV U43 ( .A(B[11]), .Z(n159) );
    VMW_INV U44 ( .A(A[5]), .Z(n141) );
    VMW_INV U45 ( .A(B[5]), .Z(n138) );
    VMW_INV U46 ( .A(A[1]), .Z(n123) );
    VMW_INV U47 ( .A(B[15]), .Z(n168) );
    VMW_INV U48 ( .A(B[13]), .Z(n165) );
    VMW_INV U49 ( .A(A[6]), .Z(n136) );
    VMW_INV U50 ( .A(A[2]), .Z(n120) );
    VMW_INV U51 ( .A(A[0]), .Z(n122) );
    VMW_INV U52 ( .A(A[15]), .Z(n116) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
        n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
        n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
        n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
        n216, n217;
    VMW_OAI21 U3 ( .A(B[15]), .B(n169), .C(n170), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n172), .B(B[2]), .Z(n171) );
    VMW_AO22 U5 ( .A(n174), .B(B[0]), .C(n175), .D(B[1]), .Z(n173) );
    VMW_OR2 U6 ( .A(B[2]), .B(n172), .Z(n176) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n175), .C(n176), .D(n173), .Z(n177) );
    VMW_NAND2 U8 ( .A(n179), .B(B[4]), .Z(n178) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n181), .C(n177), .D(n171), .Z(n180) );
    VMW_OR2 U10 ( .A(B[4]), .B(n179), .Z(n182) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n184), .C(n182), .D(n180), .Z(n183) );
    VMW_NAND2 U12 ( .A(n186), .B(B[6]), .Z(n185) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n188), .C(n183), .D(n178), .Z(n187) );
    VMW_OR2 U14 ( .A(B[6]), .B(n186), .Z(n189) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n191), .C(n189), .D(n187), .Z(n190) );
    VMW_NAND2 U16 ( .A(n193), .B(B[8]), .Z(n192) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n195), .C(n190), .D(n185), .Z(n194) );
    VMW_OR2 U18 ( .A(B[8]), .B(n193), .Z(n196) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n198), .C(n196), .D(n194), .Z(n197) );
    VMW_NAND2 U20 ( .A(n200), .B(B[10]), .Z(n199) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n202), .C(n197), .D(n192), .Z(n201) );
    VMW_NAND2 U22 ( .A(n202), .B(A[9]), .Z(n203) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n200), .C(n203), .D(n201), .Z(n204) );
    VMW_NAND2 U24 ( .A(n206), .B(B[12]), .Z(n205) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n208), .C(n204), .D(n199), .Z(n207) );
    VMW_NAND2 U26 ( .A(n208), .B(A[11]), .Z(n209) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n206), .C(n209), .D(n207), .Z(n210) );
    VMW_NAND2 U28 ( .A(n212), .B(B[14]), .Z(n211) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n214), .C(n210), .D(n205), .Z(n213) );
    VMW_NAND2 U30 ( .A(n214), .B(A[13]), .Z(n215) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n212), .C(n215), .D(n213), .Z(n216) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n217), .C(n216), .D(n211), .Z(n170) );
    VMW_INV U33 ( .A(A[12]), .Z(n206) );
    VMW_INV U34 ( .A(B[7]), .Z(n195) );
    VMW_INV U35 ( .A(A[7]), .Z(n198) );
    VMW_INV U36 ( .A(A[3]), .Z(n184) );
    VMW_INV U37 ( .A(B[3]), .Z(n181) );
    VMW_INV U38 ( .A(A[10]), .Z(n200) );
    VMW_INV U39 ( .A(B[9]), .Z(n202) );
    VMW_INV U40 ( .A(A[4]), .Z(n179) );
    VMW_INV U41 ( .A(A[8]), .Z(n193) );
    VMW_INV U42 ( .A(A[14]), .Z(n212) );
    VMW_INV U43 ( .A(B[11]), .Z(n208) );
    VMW_INV U44 ( .A(A[5]), .Z(n191) );
    VMW_INV U45 ( .A(B[5]), .Z(n188) );
    VMW_INV U46 ( .A(A[1]), .Z(n175) );
    VMW_INV U47 ( .A(B[15]), .Z(n217) );
    VMW_INV U48 ( .A(B[13]), .Z(n214) );
    VMW_INV U49 ( .A(A[6]), .Z(n186) );
    VMW_INV U50 ( .A(A[2]), .Z(n172) );
    VMW_INV U51 ( .A(A[0]), .Z(n174) );
    VMW_INV U52 ( .A(A[15]), .Z(n169) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266;
    VMW_OAI21 U3 ( .A(B[15]), .B(n218), .C(n219), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n221), .B(B[2]), .Z(n220) );
    VMW_AO22 U5 ( .A(n223), .B(B[0]), .C(n224), .D(B[1]), .Z(n222) );
    VMW_OR2 U6 ( .A(B[2]), .B(n221), .Z(n225) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n224), .C(n225), .D(n222), .Z(n226) );
    VMW_NAND2 U8 ( .A(n228), .B(B[4]), .Z(n227) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n230), .C(n226), .D(n220), .Z(n229) );
    VMW_OR2 U10 ( .A(B[4]), .B(n228), .Z(n231) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n233), .C(n231), .D(n229), .Z(n232) );
    VMW_NAND2 U12 ( .A(n235), .B(B[6]), .Z(n234) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n237), .C(n232), .D(n227), .Z(n236) );
    VMW_OR2 U14 ( .A(B[6]), .B(n235), .Z(n238) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n240), .C(n238), .D(n236), .Z(n239) );
    VMW_NAND2 U16 ( .A(n242), .B(B[8]), .Z(n241) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n244), .C(n239), .D(n234), .Z(n243) );
    VMW_OR2 U18 ( .A(B[8]), .B(n242), .Z(n245) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n247), .C(n245), .D(n243), .Z(n246) );
    VMW_NAND2 U20 ( .A(n249), .B(B[10]), .Z(n248) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n251), .C(n246), .D(n241), .Z(n250) );
    VMW_NAND2 U22 ( .A(n251), .B(A[9]), .Z(n252) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n249), .C(n252), .D(n250), .Z(n253) );
    VMW_NAND2 U24 ( .A(n255), .B(B[12]), .Z(n254) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n257), .C(n253), .D(n248), .Z(n256) );
    VMW_NAND2 U26 ( .A(n257), .B(A[11]), .Z(n258) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n255), .C(n258), .D(n256), .Z(n259) );
    VMW_NAND2 U28 ( .A(n261), .B(B[14]), .Z(n260) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n263), .C(n259), .D(n254), .Z(n262) );
    VMW_NAND2 U30 ( .A(n263), .B(A[13]), .Z(n264) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n261), .C(n264), .D(n262), .Z(n265) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n266), .C(n265), .D(n260), .Z(n219) );
    VMW_INV U33 ( .A(A[12]), .Z(n255) );
    VMW_INV U34 ( .A(B[7]), .Z(n244) );
    VMW_INV U35 ( .A(A[7]), .Z(n247) );
    VMW_INV U36 ( .A(A[3]), .Z(n233) );
    VMW_INV U37 ( .A(B[3]), .Z(n230) );
    VMW_INV U38 ( .A(A[10]), .Z(n249) );
    VMW_INV U39 ( .A(B[9]), .Z(n251) );
    VMW_INV U40 ( .A(A[4]), .Z(n228) );
    VMW_INV U41 ( .A(A[8]), .Z(n242) );
    VMW_INV U42 ( .A(A[14]), .Z(n261) );
    VMW_INV U43 ( .A(B[11]), .Z(n257) );
    VMW_INV U44 ( .A(A[5]), .Z(n240) );
    VMW_INV U45 ( .A(B[5]), .Z(n237) );
    VMW_INV U46 ( .A(A[1]), .Z(n224) );
    VMW_INV U47 ( .A(B[15]), .Z(n266) );
    VMW_INV U48 ( .A(B[13]), .Z(n263) );
    VMW_INV U49 ( .A(A[6]), .Z(n235) );
    VMW_INV U50 ( .A(A[2]), .Z(n221) );
    VMW_INV U51 ( .A(A[0]), .Z(n223) );
    VMW_INV U52 ( .A(A[15]), .Z(n218) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315;
    VMW_OAI21 U3 ( .A(B[15]), .B(n267), .C(n268), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n270), .B(B[2]), .Z(n269) );
    VMW_AO22 U5 ( .A(n272), .B(B[0]), .C(n273), .D(B[1]), .Z(n271) );
    VMW_OR2 U6 ( .A(B[2]), .B(n270), .Z(n274) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n273), .C(n274), .D(n271), .Z(n275) );
    VMW_NAND2 U8 ( .A(n277), .B(B[4]), .Z(n276) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n279), .C(n275), .D(n269), .Z(n278) );
    VMW_OR2 U10 ( .A(B[4]), .B(n277), .Z(n280) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n282), .C(n280), .D(n278), .Z(n281) );
    VMW_NAND2 U12 ( .A(n284), .B(B[6]), .Z(n283) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n286), .C(n281), .D(n276), .Z(n285) );
    VMW_OR2 U14 ( .A(B[6]), .B(n284), .Z(n287) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n289), .C(n287), .D(n285), .Z(n288) );
    VMW_NAND2 U16 ( .A(n291), .B(B[8]), .Z(n290) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n293), .C(n288), .D(n283), .Z(n292) );
    VMW_OR2 U18 ( .A(B[8]), .B(n291), .Z(n294) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n296), .C(n294), .D(n292), .Z(n295) );
    VMW_NAND2 U20 ( .A(n298), .B(B[10]), .Z(n297) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n300), .C(n295), .D(n290), .Z(n299) );
    VMW_NAND2 U22 ( .A(n300), .B(A[9]), .Z(n301) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n298), .C(n301), .D(n299), .Z(n302) );
    VMW_NAND2 U24 ( .A(n304), .B(B[12]), .Z(n303) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n306), .C(n302), .D(n297), .Z(n305) );
    VMW_NAND2 U26 ( .A(n306), .B(A[11]), .Z(n307) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n304), .C(n307), .D(n305), .Z(n308) );
    VMW_NAND2 U28 ( .A(n310), .B(B[14]), .Z(n309) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n312), .C(n308), .D(n303), .Z(n311) );
    VMW_NAND2 U30 ( .A(n312), .B(A[13]), .Z(n313) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n310), .C(n313), .D(n311), .Z(n314) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n315), .C(n314), .D(n309), .Z(n268) );
    VMW_INV U33 ( .A(A[12]), .Z(n304) );
    VMW_INV U34 ( .A(B[7]), .Z(n293) );
    VMW_INV U35 ( .A(A[7]), .Z(n296) );
    VMW_INV U36 ( .A(A[3]), .Z(n282) );
    VMW_INV U37 ( .A(B[3]), .Z(n279) );
    VMW_INV U38 ( .A(A[10]), .Z(n298) );
    VMW_INV U39 ( .A(B[9]), .Z(n300) );
    VMW_INV U40 ( .A(A[4]), .Z(n277) );
    VMW_INV U41 ( .A(A[8]), .Z(n291) );
    VMW_INV U42 ( .A(A[14]), .Z(n310) );
    VMW_INV U43 ( .A(B[11]), .Z(n306) );
    VMW_INV U44 ( .A(A[5]), .Z(n289) );
    VMW_INV U45 ( .A(B[5]), .Z(n286) );
    VMW_INV U46 ( .A(A[1]), .Z(n273) );
    VMW_INV U47 ( .A(B[15]), .Z(n315) );
    VMW_INV U48 ( .A(B[13]), .Z(n312) );
    VMW_INV U49 ( .A(A[6]), .Z(n284) );
    VMW_INV U50 ( .A(A[2]), .Z(n270) );
    VMW_INV U51 ( .A(A[0]), .Z(n272) );
    VMW_INV U52 ( .A(A[15]), .Z(n267) );
endmodule


module NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 ( A, B, LEQ, TC, LT_LE, GE_GT
     );
input  [15:0] A;
input  [15:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
        n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
        n363, n364;
    VMW_OAI21 U3 ( .A(B[15]), .B(n316), .C(n317), .Z(GE_GT) );
    VMW_NAND2 U4 ( .A(n319), .B(B[2]), .Z(n318) );
    VMW_AO22 U5 ( .A(n321), .B(B[0]), .C(n322), .D(B[1]), .Z(n320) );
    VMW_OR2 U6 ( .A(B[2]), .B(n319), .Z(n323) );
    VMW_OAI211 U7 ( .A(B[1]), .B(n322), .C(n323), .D(n320), .Z(n324) );
    VMW_NAND2 U8 ( .A(n326), .B(B[4]), .Z(n325) );
    VMW_OAI211 U9 ( .A(A[3]), .B(n328), .C(n324), .D(n318), .Z(n327) );
    VMW_OR2 U10 ( .A(B[4]), .B(n326), .Z(n329) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n331), .C(n329), .D(n327), .Z(n330) );
    VMW_NAND2 U12 ( .A(n333), .B(B[6]), .Z(n332) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n335), .C(n330), .D(n325), .Z(n334) );
    VMW_OR2 U14 ( .A(B[6]), .B(n333), .Z(n336) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n338), .C(n336), .D(n334), .Z(n337) );
    VMW_NAND2 U16 ( .A(n340), .B(B[8]), .Z(n339) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n342), .C(n337), .D(n332), .Z(n341) );
    VMW_OR2 U18 ( .A(B[8]), .B(n340), .Z(n343) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n345), .C(n343), .D(n341), .Z(n344) );
    VMW_NAND2 U20 ( .A(n347), .B(B[10]), .Z(n346) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n349), .C(n344), .D(n339), .Z(n348) );
    VMW_NAND2 U22 ( .A(n349), .B(A[9]), .Z(n350) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n347), .C(n350), .D(n348), .Z(n351) );
    VMW_NAND2 U24 ( .A(n353), .B(B[12]), .Z(n352) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n355), .C(n351), .D(n346), .Z(n354) );
    VMW_NAND2 U26 ( .A(n355), .B(A[11]), .Z(n356) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n353), .C(n356), .D(n354), .Z(n357) );
    VMW_NAND2 U28 ( .A(n359), .B(B[14]), .Z(n358) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n361), .C(n357), .D(n352), .Z(n360) );
    VMW_NAND2 U30 ( .A(n361), .B(A[13]), .Z(n362) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n359), .C(n362), .D(n360), .Z(n363) );
    VMW_OAI211 U32 ( .A(A[15]), .B(n364), .C(n363), .D(n358), .Z(n317) );
    VMW_INV U33 ( .A(A[12]), .Z(n353) );
    VMW_INV U34 ( .A(B[7]), .Z(n342) );
    VMW_INV U35 ( .A(A[7]), .Z(n345) );
    VMW_INV U36 ( .A(A[3]), .Z(n331) );
    VMW_INV U37 ( .A(B[3]), .Z(n328) );
    VMW_INV U38 ( .A(A[10]), .Z(n347) );
    VMW_INV U39 ( .A(B[9]), .Z(n349) );
    VMW_INV U40 ( .A(A[4]), .Z(n326) );
    VMW_INV U41 ( .A(A[8]), .Z(n340) );
    VMW_INV U42 ( .A(A[14]), .Z(n359) );
    VMW_INV U43 ( .A(B[11]), .Z(n355) );
    VMW_INV U44 ( .A(A[5]), .Z(n338) );
    VMW_INV U45 ( .A(B[5]), .Z(n335) );
    VMW_INV U46 ( .A(A[1]), .Z(n322) );
    VMW_INV U47 ( .A(B[15]), .Z(n364) );
    VMW_INV U48 ( .A(B[13]), .Z(n361) );
    VMW_INV U49 ( .A(A[6]), .Z(n333) );
    VMW_INV U50 ( .A(A[2]), .Z(n319) );
    VMW_INV U51 ( .A(A[0]), .Z(n321) );
    VMW_INV U52 ( .A(A[15]), .Z(n316) );
endmodule


module NodeAux_INDEGREE7_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [6:0] Nid;
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \OutEdge156[4] , \temp324[9] , \temp594[1] , \temp324[0] , 
        \temp594[8] , \OutEdge156[10] , \OutEdge156[0] , \temp594[5] , 
        \temp684[12] , \OutEdge156[14] , \path[2] , \OutEdge156[9] , 
        \temp324[4] , \path[0] , \temp324[6] , \temp684[10] , \temp594[7] , 
        \OutEdge156[2] , \OutEdge156[12] , \temp324[2] , \OutEdge156[6] , 
        \temp594[3] , \temp684[14] , \temp504[15] , \temp684[8] , \temp504[9] , 
        \temp414[5] , \temp230[7] , \temp504[0] , \temp594[15] , \temp684[1] , 
        \temp414[13] , \temp414[8] , \temp504[11] , \temp684[5] , 
        \temp594[11] , \temp324[12] , \temp230[3] , \temp504[4] , \temp414[1] , 
        \temp230[12] , \temp230[1] , \temp504[6] , \temp414[3] , \temp230[10] , 
        n126, \temp594[13] , \temp684[7] , \temp324[10] , \temp504[13] , 
        \temp230[8] , \temp414[11] , \temp324[14] , \temp684[3] , 
        \temp230[14] , \temp414[7] , \temp230[5] , \temp504[2] , \temp414[15] , 
        n134, \temp324[15] , n118, \temp684[2] , \temp414[6] , \temp230[15] , 
        n94, \temp504[3] , \temp230[4] , \temp414[14] , \temp230[0] , 
        \temp504[7] , \temp230[11] , \temp414[2] , \temp684[6] , \temp594[12] , 
        \temp324[11] , \temp504[12] , \temp230[9] , \temp414[10] , 
        \temp414[9] , \temp414[12] , \temp504[10] , \temp684[4] , 
        \temp594[10] , \temp324[13] , \temp230[2] , \temp504[5] , 
        \temp230[13] , \temp414[0] , \temp504[14] , \temp684[9] , \temp504[8] , 
        \temp414[4] , \temp230[6] , \temp504[1] , \temp684[0] , \temp594[14] , 
        \OutEdge156[13] , \temp324[3] , \OutEdge156[7] , \temp594[2] , 
        \temp684[15] , \temp324[7] , \path[1] , \temp684[11] , \temp594[6] , 
        \OutEdge156[3] , n102, \temp594[4] , \OutEdge156[1] , \temp684[13] , 
        \OutEdge156[15] , \temp324[5] , \OutEdge156[8] , \OutEdge156[5] , n142, 
        \temp324[8] , \temp594[0] , \OutEdge156[11] , \temp594[9] , 
        \temp324[1] , n110, n867, n868, n869, n870, n871, n872, n873, n874, 
        n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, 
        n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, 
        n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, 
        n911, n912, n913, n914, n915, n916, n917, n918, n919;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_PULLDOWN U100 ( .Z(n915) );
    VMW_PULLDOWN U101 ( .Z(n919) );
    VMW_PULLDOWN U102 ( .Z(n917) );
    VMW_PULLDOWN U103 ( .Z(n918) );
    VMW_PULLDOWN U104 ( .Z(n914) );
    VMW_PULLDOWN U105 ( .Z(n913) );
    VMW_PULLDOWN U106 ( .Z(n916) );
    VMW_NOR2 U107 ( .A(Start), .B(n867), .Z(\OutEdge156[15] ) );
    VMW_NAND2 U108 ( .A(n868), .B(n869), .Z(\OutEdge156[14] ) );
    VMW_NAND2 U109 ( .A(n870), .B(n869), .Z(\OutEdge156[13] ) );
    VMW_NAND2 U110 ( .A(n871), .B(n869), .Z(\OutEdge156[12] ) );
    VMW_NAND2 U111 ( .A(n872), .B(n869), .Z(\OutEdge156[11] ) );
    VMW_NAND2 U112 ( .A(n873), .B(n869), .Z(\OutEdge156[10] ) );
    VMW_NAND2 U113 ( .A(n874), .B(n869), .Z(\OutEdge156[9] ) );
    VMW_NAND2 U114 ( .A(n875), .B(n869), .Z(\OutEdge156[8] ) );
    VMW_NAND2 U115 ( .A(n876), .B(n869), .Z(\OutEdge156[7] ) );
    VMW_NAND2 U116 ( .A(n877), .B(n869), .Z(\OutEdge156[6] ) );
    VMW_NAND2 U117 ( .A(n878), .B(n869), .Z(\OutEdge156[5] ) );
    VMW_NAND2 U118 ( .A(n879), .B(n869), .Z(\OutEdge156[4] ) );
    VMW_NAND2 U119 ( .A(n880), .B(n869), .Z(\OutEdge156[3] ) );
    VMW_NAND2 U120 ( .A(n881), .B(n869), .Z(\OutEdge156[2] ) );
    VMW_NAND2 U121 ( .A(n882), .B(n869), .Z(\OutEdge156[1] ) );
    VMW_NAND2 U122 ( .A(n883), .B(n869), .Z(\OutEdge156[0] ) );
    VMW_AND4 U123 ( .A(n885), .B(n886), .C(n887), .D(n888), .Z(n884) );
    VMW_OR4 U124 ( .A(n142), .B(n126), .C(n134), .D(n884), .Z(n889) );
    VMW_NOR3 U125 ( .A(n134), .B(n126), .C(n891), .Z(n890) );
    VMW_OR2 U126 ( .A(n890), .B(n142), .Z(n892) );
    VMW_AO22 U127 ( .A(InEdges[95]), .B(n134), .C(\temp594[15] ), .D(n893), 
        .Z(\temp684[15] ) );
    VMW_OAI22 U128 ( .A(n889), .B(Start), .C(\path[2] ), .D(n869), .Z(n894) );
    VMW_OAI22 U129 ( .A(n892), .B(Start), .C(\path[1] ), .D(n869), .Z(n895) );
    VMW_OAI22 U130 ( .A(n897), .B(Start), .C(\path[0] ), .D(n869), .Z(n896) );
    VMW_MUX2I U131 ( .A(\temp684[15] ), .B(InEdges[111]), .S(n142), .Z(n867)
         );
    VMW_AND4 U132 ( .A(n899), .B(n900), .C(n901), .D(n902), .Z(n898) );
    VMW_INV U133 ( .A(Start), .Z(n869) );
    VMW_INV U134 ( .A(n118), .Z(n886) );
    VMW_INV U135 ( .A(n134), .Z(n893) );
    VMW_AOI211 U136 ( .A(n885), .B(n887), .C(n110), .D(n118), .Z(n891) );
    VMW_OAI21 U137 ( .A(n102), .B(n885), .C(n888), .Z(n903) );
    VMW_AO21 U138 ( .A(n886), .B(n903), .C(n126), .Z(n904) );
    VMW_AND4 U139 ( .A(n905), .B(n906), .C(n907), .D(n898), .Z(n909) );
    VMW_XNOR2 U140 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n902) );
    VMW_XNOR2 U141 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n901) );
    VMW_XNOR2 U142 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n900) );
    VMW_XNOR2 U143 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n899) );
    VMW_XNOR2 U144 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n906) );
    VMW_XNOR2 U145 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n905) );
    VMW_XNOR2 U146 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n907) );
    VMW_AO22 U147 ( .A(InEdges[9]), .B(n94), .C(OutEdge[9]), .D(n885), .Z(
        \temp230[9] ) );
    VMW_AO22 U148 ( .A(InEdges[25]), .B(n102), .C(\temp230[9] ), .D(n887), .Z(
        \temp324[9] ) );
    VMW_AO22 U149 ( .A(\temp324[9] ), .B(n888), .C(InEdges[41]), .D(n110), .Z(
        \temp414[9] ) );
    VMW_AO22 U150 ( .A(InEdges[57]), .B(n118), .C(\temp414[9] ), .D(n886), .Z(
        \temp504[9] ) );
    VMW_AO22 U151 ( .A(\temp504[9] ), .B(n908), .C(InEdges[73]), .D(n126), .Z(
        \temp594[9] ) );
    VMW_AO22 U152 ( .A(InEdges[89]), .B(n134), .C(\temp594[9] ), .D(n893), .Z(
        \temp684[9] ) );
    VMW_AO22 U153 ( .A(InEdges[8]), .B(n94), .C(OutEdge[8]), .D(n885), .Z(
        \temp230[8] ) );
    VMW_AO22 U154 ( .A(InEdges[24]), .B(n102), .C(\temp230[8] ), .D(n887), .Z(
        \temp324[8] ) );
    VMW_AO22 U155 ( .A(\temp324[8] ), .B(n888), .C(InEdges[40]), .D(n110), .Z(
        \temp414[8] ) );
    VMW_AO22 U156 ( .A(InEdges[56]), .B(n118), .C(\temp414[8] ), .D(n886), .Z(
        \temp504[8] ) );
    VMW_AO22 U157 ( .A(\temp504[8] ), .B(n908), .C(InEdges[72]), .D(n126), .Z(
        \temp594[8] ) );
    VMW_AO22 U158 ( .A(InEdges[88]), .B(n134), .C(\temp594[8] ), .D(n893), .Z(
        \temp684[8] ) );
    VMW_AO22 U159 ( .A(InEdges[7]), .B(n94), .C(OutEdge[7]), .D(n885), .Z(
        \temp230[7] ) );
    VMW_AO22 U160 ( .A(InEdges[23]), .B(n102), .C(\temp230[7] ), .D(n887), .Z(
        \temp324[7] ) );
    VMW_AO22 U161 ( .A(\temp324[7] ), .B(n888), .C(InEdges[39]), .D(n110), .Z(
        \temp414[7] ) );
    VMW_AO22 U162 ( .A(InEdges[55]), .B(n118), .C(\temp414[7] ), .D(n886), .Z(
        \temp504[7] ) );
    VMW_AO22 U163 ( .A(\temp504[7] ), .B(n908), .C(InEdges[71]), .D(n126), .Z(
        \temp594[7] ) );
    VMW_AO22 U164 ( .A(InEdges[87]), .B(n134), .C(\temp594[7] ), .D(n893), .Z(
        \temp684[7] ) );
    VMW_AO22 U165 ( .A(InEdges[6]), .B(n94), .C(OutEdge[6]), .D(n885), .Z(
        \temp230[6] ) );
    VMW_AO22 U166 ( .A(InEdges[22]), .B(n102), .C(\temp230[6] ), .D(n887), .Z(
        \temp324[6] ) );
    VMW_AO22 U167 ( .A(\temp324[6] ), .B(n888), .C(InEdges[38]), .D(n110), .Z(
        \temp414[6] ) );
    VMW_AO22 U168 ( .A(InEdges[54]), .B(n118), .C(\temp414[6] ), .D(n886), .Z(
        \temp504[6] ) );
    VMW_AO22 U169 ( .A(\temp504[6] ), .B(n908), .C(InEdges[70]), .D(n126), .Z(
        \temp594[6] ) );
    VMW_AO22 U170 ( .A(InEdges[86]), .B(n134), .C(\temp594[6] ), .D(n893), .Z(
        \temp684[6] ) );
    VMW_AO22 U171 ( .A(InEdges[5]), .B(n94), .C(OutEdge[5]), .D(n885), .Z(
        \temp230[5] ) );
    VMW_AO22 U172 ( .A(InEdges[21]), .B(n102), .C(\temp230[5] ), .D(n887), .Z(
        \temp324[5] ) );
    VMW_AO22 U173 ( .A(\temp324[5] ), .B(n888), .C(InEdges[37]), .D(n110), .Z(
        \temp414[5] ) );
    VMW_AO22 U174 ( .A(InEdges[53]), .B(n118), .C(\temp414[5] ), .D(n886), .Z(
        \temp504[5] ) );
    VMW_AO22 U175 ( .A(\temp504[5] ), .B(n908), .C(InEdges[69]), .D(n126), .Z(
        \temp594[5] ) );
    VMW_AO22 U176 ( .A(InEdges[85]), .B(n134), .C(\temp594[5] ), .D(n893), .Z(
        \temp684[5] ) );
    VMW_AO22 U177 ( .A(InEdges[4]), .B(n94), .C(OutEdge[4]), .D(n885), .Z(
        \temp230[4] ) );
    VMW_AO22 U178 ( .A(InEdges[20]), .B(n102), .C(\temp230[4] ), .D(n887), .Z(
        \temp324[4] ) );
    VMW_AO22 U179 ( .A(\temp324[4] ), .B(n888), .C(InEdges[36]), .D(n110), .Z(
        \temp414[4] ) );
    VMW_AO22 U180 ( .A(InEdges[52]), .B(n118), .C(\temp414[4] ), .D(n886), .Z(
        \temp504[4] ) );
    VMW_AO22 U181 ( .A(\temp504[4] ), .B(n908), .C(InEdges[68]), .D(n126), .Z(
        \temp594[4] ) );
    VMW_AO22 U182 ( .A(InEdges[84]), .B(n134), .C(\temp594[4] ), .D(n893), .Z(
        \temp684[4] ) );
    VMW_AO22 U183 ( .A(InEdges[3]), .B(n94), .C(OutEdge[3]), .D(n885), .Z(
        \temp230[3] ) );
    VMW_AO22 U184 ( .A(InEdges[19]), .B(n102), .C(\temp230[3] ), .D(n887), .Z(
        \temp324[3] ) );
    VMW_AO22 U185 ( .A(\temp324[3] ), .B(n888), .C(InEdges[35]), .D(n110), .Z(
        \temp414[3] ) );
    VMW_AO22 U186 ( .A(InEdges[51]), .B(n118), .C(\temp414[3] ), .D(n886), .Z(
        \temp504[3] ) );
    VMW_AO22 U187 ( .A(\temp504[3] ), .B(n908), .C(InEdges[67]), .D(n126), .Z(
        \temp594[3] ) );
    VMW_AO22 U188 ( .A(InEdges[83]), .B(n134), .C(\temp594[3] ), .D(n893), .Z(
        \temp684[3] ) );
    VMW_AO22 U189 ( .A(InEdges[2]), .B(n94), .C(OutEdge[2]), .D(n885), .Z(
        \temp230[2] ) );
    VMW_AO22 U190 ( .A(InEdges[18]), .B(n102), .C(\temp230[2] ), .D(n887), .Z(
        \temp324[2] ) );
    VMW_AO22 U191 ( .A(\temp324[2] ), .B(n888), .C(InEdges[34]), .D(n110), .Z(
        \temp414[2] ) );
    VMW_AO22 U192 ( .A(InEdges[50]), .B(n118), .C(\temp414[2] ), .D(n886), .Z(
        \temp504[2] ) );
    VMW_AO22 U193 ( .A(\temp504[2] ), .B(n908), .C(InEdges[66]), .D(n126), .Z(
        \temp594[2] ) );
    VMW_AO22 U194 ( .A(InEdges[82]), .B(n134), .C(\temp594[2] ), .D(n893), .Z(
        \temp684[2] ) );
    VMW_AO22 U195 ( .A(InEdges[1]), .B(n94), .C(OutEdge[1]), .D(n885), .Z(
        \temp230[1] ) );
    VMW_AO22 U196 ( .A(InEdges[17]), .B(n102), .C(\temp230[1] ), .D(n887), .Z(
        \temp324[1] ) );
    VMW_AO22 U197 ( .A(\temp324[1] ), .B(n888), .C(InEdges[33]), .D(n110), .Z(
        \temp414[1] ) );
    VMW_AO22 U198 ( .A(InEdges[49]), .B(n118), .C(\temp414[1] ), .D(n886), .Z(
        \temp504[1] ) );
    VMW_AO22 U199 ( .A(\temp504[1] ), .B(n908), .C(InEdges[65]), .D(n126), .Z(
        \temp594[1] ) );
    VMW_AO22 U200 ( .A(InEdges[81]), .B(n134), .C(\temp594[1] ), .D(n893), .Z(
        \temp684[1] ) );
    VMW_AO22 U201 ( .A(InEdges[15]), .B(n94), .C(OutEdge[15]), .D(n885), .Z(
        \temp230[15] ) );
    VMW_AO22 U202 ( .A(InEdges[31]), .B(n102), .C(\temp230[15] ), .D(n887), 
        .Z(\temp324[15] ) );
    VMW_AO22 U203 ( .A(\temp324[15] ), .B(n888), .C(InEdges[47]), .D(n110), 
        .Z(\temp414[15] ) );
    VMW_AO22 U204 ( .A(InEdges[63]), .B(n118), .C(\temp414[15] ), .D(n886), 
        .Z(\temp504[15] ) );
    VMW_AO22 U205 ( .A(\temp504[15] ), .B(n908), .C(InEdges[79]), .D(n126), 
        .Z(\temp594[15] ) );
    VMW_AO22 U206 ( .A(InEdges[14]), .B(n94), .C(OutEdge[14]), .D(n885), .Z(
        \temp230[14] ) );
    VMW_AO22 U207 ( .A(InEdges[30]), .B(n102), .C(\temp230[14] ), .D(n887), 
        .Z(\temp324[14] ) );
    VMW_AO22 U208 ( .A(\temp324[14] ), .B(n888), .C(InEdges[46]), .D(n110), 
        .Z(\temp414[14] ) );
    VMW_AO22 U209 ( .A(InEdges[62]), .B(n118), .C(\temp414[14] ), .D(n886), 
        .Z(\temp504[14] ) );
    VMW_AO22 U210 ( .A(\temp504[14] ), .B(n908), .C(InEdges[78]), .D(n126), 
        .Z(\temp594[14] ) );
    VMW_AO22 U211 ( .A(InEdges[94]), .B(n134), .C(\temp594[14] ), .D(n893), 
        .Z(\temp684[14] ) );
    VMW_AO22 U212 ( .A(InEdges[13]), .B(n94), .C(OutEdge[13]), .D(n885), .Z(
        \temp230[13] ) );
    VMW_AO22 U213 ( .A(InEdges[29]), .B(n102), .C(\temp230[13] ), .D(n887), 
        .Z(\temp324[13] ) );
    VMW_AO22 U214 ( .A(\temp324[13] ), .B(n888), .C(InEdges[45]), .D(n110), 
        .Z(\temp414[13] ) );
    VMW_AO22 U215 ( .A(InEdges[61]), .B(n118), .C(\temp414[13] ), .D(n886), 
        .Z(\temp504[13] ) );
    VMW_AO22 U216 ( .A(\temp504[13] ), .B(n908), .C(InEdges[77]), .D(n126), 
        .Z(\temp594[13] ) );
    VMW_AO22 U217 ( .A(InEdges[93]), .B(n134), .C(\temp594[13] ), .D(n893), 
        .Z(\temp684[13] ) );
    VMW_AO22 U218 ( .A(InEdges[12]), .B(n94), .C(OutEdge[12]), .D(n885), .Z(
        \temp230[12] ) );
    VMW_AO22 U219 ( .A(InEdges[28]), .B(n102), .C(\temp230[12] ), .D(n887), 
        .Z(\temp324[12] ) );
    VMW_AO22 U220 ( .A(\temp324[12] ), .B(n888), .C(InEdges[44]), .D(n110), 
        .Z(\temp414[12] ) );
    VMW_AO22 U221 ( .A(InEdges[60]), .B(n118), .C(\temp414[12] ), .D(n886), 
        .Z(\temp504[12] ) );
    VMW_AO22 U222 ( .A(\temp504[12] ), .B(n908), .C(InEdges[76]), .D(n126), 
        .Z(\temp594[12] ) );
    VMW_AO22 U223 ( .A(InEdges[92]), .B(n134), .C(\temp594[12] ), .D(n893), 
        .Z(\temp684[12] ) );
    VMW_AO22 U224 ( .A(InEdges[11]), .B(n94), .C(OutEdge[11]), .D(n885), .Z(
        \temp230[11] ) );
    VMW_AO22 U225 ( .A(InEdges[27]), .B(n102), .C(\temp230[11] ), .D(n887), 
        .Z(\temp324[11] ) );
    VMW_AO22 U226 ( .A(\temp324[11] ), .B(n888), .C(InEdges[43]), .D(n110), 
        .Z(\temp414[11] ) );
    VMW_AO22 U227 ( .A(InEdges[59]), .B(n118), .C(\temp414[11] ), .D(n886), 
        .Z(\temp504[11] ) );
    VMW_AO22 U228 ( .A(\temp504[11] ), .B(n908), .C(InEdges[75]), .D(n126), 
        .Z(\temp594[11] ) );
    VMW_AO22 U229 ( .A(InEdges[91]), .B(n134), .C(\temp594[11] ), .D(n893), 
        .Z(\temp684[11] ) );
    VMW_AO22 U230 ( .A(InEdges[10]), .B(n94), .C(OutEdge[10]), .D(n885), .Z(
        \temp230[10] ) );
    VMW_AO22 U231 ( .A(InEdges[26]), .B(n102), .C(\temp230[10] ), .D(n887), 
        .Z(\temp324[10] ) );
    VMW_AO22 U232 ( .A(\temp324[10] ), .B(n888), .C(InEdges[42]), .D(n110), 
        .Z(\temp414[10] ) );
    VMW_AO22 U233 ( .A(InEdges[58]), .B(n118), .C(\temp414[10] ), .D(n886), 
        .Z(\temp504[10] ) );
    VMW_AO22 U234 ( .A(\temp504[10] ), .B(n908), .C(InEdges[74]), .D(n126), 
        .Z(\temp594[10] ) );
    VMW_AO22 U235 ( .A(InEdges[90]), .B(n134), .C(\temp594[10] ), .D(n893), 
        .Z(\temp684[10] ) );
    VMW_AO22 U236 ( .A(InEdges[0]), .B(n94), .C(OutEdge[0]), .D(n885), .Z(
        \temp230[0] ) );
    VMW_AO22 U237 ( .A(InEdges[16]), .B(n102), .C(\temp230[0] ), .D(n887), .Z(
        \temp324[0] ) );
    VMW_AO22 U238 ( .A(\temp324[0] ), .B(n888), .C(InEdges[32]), .D(n110), .Z(
        \temp414[0] ) );
    VMW_AO22 U239 ( .A(InEdges[48]), .B(n118), .C(\temp414[0] ), .D(n886), .Z(
        \temp504[0] ) );
    VMW_AO22 U240 ( .A(\temp504[0] ), .B(n908), .C(InEdges[64]), .D(n126), .Z(
        \temp594[0] ) );
    VMW_AO22 U241 ( .A(InEdges[80]), .B(n134), .C(\temp594[0] ), .D(n893), .Z(
        \temp684[0] ) );
    VMW_AOI21 U242 ( .A(n893), .B(n904), .C(n142), .Z(n897) );
    VMW_MUX2I U243 ( .A(\temp684[9] ), .B(InEdges[105]), .S(n142), .Z(n874) );
    VMW_MUX2I U244 ( .A(\temp684[8] ), .B(InEdges[104]), .S(n142), .Z(n875) );
    VMW_MUX2I U245 ( .A(\temp684[7] ), .B(InEdges[103]), .S(n142), .Z(n876) );
    VMW_MUX2I U246 ( .A(\temp684[6] ), .B(InEdges[102]), .S(n142), .Z(n877) );
    VMW_MUX2I U247 ( .A(\temp684[5] ), .B(InEdges[101]), .S(n142), .Z(n878) );
    VMW_MUX2I U248 ( .A(\temp684[4] ), .B(InEdges[100]), .S(n142), .Z(n879) );
    VMW_MUX2I U249 ( .A(\temp684[3] ), .B(InEdges[99]), .S(n142), .Z(n880) );
    VMW_MUX2I U250 ( .A(\temp684[2] ), .B(InEdges[98]), .S(n142), .Z(n881) );
    VMW_MUX2I U251 ( .A(\temp684[1] ), .B(InEdges[97]), .S(n142), .Z(n882) );
    VMW_MUX2I U252 ( .A(\temp684[14] ), .B(InEdges[110]), .S(n142), .Z(n868)
         );
    VMW_MUX2I U253 ( .A(\temp684[13] ), .B(InEdges[109]), .S(n142), .Z(n870)
         );
    VMW_MUX2I U254 ( .A(\temp684[12] ), .B(InEdges[108]), .S(n142), .Z(n871)
         );
    VMW_MUX2I U255 ( .A(\temp684[11] ), .B(InEdges[107]), .S(n142), .Z(n872)
         );
    VMW_MUX2I U256 ( .A(\temp684[10] ), .B(InEdges[106]), .S(n142), .Z(n873)
         );
    VMW_MUX2I U257 ( .A(\temp684[0] ), .B(InEdges[96]), .S(n142), .Z(n883) );
    VMW_INV U258 ( .A(n102), .Z(n887) );
    VMW_INV U259 ( .A(n94), .Z(n885) );
    VMW_INV U260 ( .A(n110), .Z(n888) );
    VMW_INV U261 ( .A(n126), .Z(n908) );
    VMW_INV U262 ( .A(n894), .Z(n911) );
    VMW_INV U263 ( .A(n895), .Z(n912) );
    VMW_INV U264 ( .A(n896), .Z(n910) );
    VMW_BUFIZ U265 ( .A(\path[1] ), .E(n909), .Z(\PathData[1] ) );
    VMW_BUFIZ U266 ( .A(\path[0] ), .E(n909), .Z(\PathData[0] ) );
    VMW_BUFIZ U267 ( .A(\path[2] ), .E(n909), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n910), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n911), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n912), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[15]  ( .D(\OutEdge156[15] ), .CP(Clk), .Q(OutEdge[15])
         );
    VMW_FD \OutEdge_reg[14]  ( .D(\OutEdge156[14] ), .CP(Clk), .Q(OutEdge[14])
         );
    VMW_FD \OutEdge_reg[13]  ( .D(\OutEdge156[13] ), .CP(Clk), .Q(OutEdge[13])
         );
    VMW_FD \OutEdge_reg[12]  ( .D(\OutEdge156[12] ), .CP(Clk), .Q(OutEdge[12])
         );
    VMW_FD \OutEdge_reg[11]  ( .D(\OutEdge156[11] ), .CP(Clk), .Q(OutEdge[11])
         );
    VMW_FD \OutEdge_reg[10]  ( .D(\OutEdge156[10] ), .CP(Clk), .Q(OutEdge[10])
         );
    VMW_FD \OutEdge_reg[9]  ( .D(\OutEdge156[9] ), .CP(Clk), .Q(OutEdge[9]) );
    VMW_FD \OutEdge_reg[8]  ( .D(\OutEdge156[8] ), .CP(Clk), .Q(OutEdge[8]) );
    VMW_FD \OutEdge_reg[7]  ( .D(\OutEdge156[7] ), .CP(Clk), .Q(OutEdge[7]) );
    VMW_FD \OutEdge_reg[6]  ( .D(\OutEdge156[6] ), .CP(Clk), .Q(OutEdge[6]) );
    VMW_FD \OutEdge_reg[5]  ( .D(\OutEdge156[5] ), .CP(Clk), .Q(OutEdge[5]) );
    VMW_FD \OutEdge_reg[4]  ( .D(\OutEdge156[4] ), .CP(Clk), .Q(OutEdge[4]) );
    VMW_FD \OutEdge_reg[3]  ( .D(\OutEdge156[3] ), .CP(Clk), .Q(OutEdge[3]) );
    VMW_FD \OutEdge_reg[2]  ( .D(\OutEdge156[2] ), .CP(Clk), .Q(OutEdge[2]) );
    VMW_FD \OutEdge_reg[1]  ( .D(\OutEdge156[1] ), .CP(Clk), .Q(OutEdge[1]) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge156[0] ), .CP(Clk), .Q(OutEdge[0]) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_6 lte_55_5 ( .A({\temp594[15] , 
        \temp594[14] , \temp594[13] , \temp594[12] , \temp594[11] , 
        \temp594[10] , \temp594[9] , \temp594[8] , \temp594[7] , \temp594[6] , 
        \temp594[5] , \temp594[4] , \temp594[3] , \temp594[2] , \temp594[1] , 
        \temp594[0] }), .B(InEdges[95:80]), .LEQ(n919), .TC(n919), .GE_GT(n134
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_5 lte_55_3 ( .A({\temp414[15] , 
        \temp414[14] , \temp414[13] , \temp414[12] , \temp414[11] , 
        \temp414[10] , \temp414[9] , \temp414[8] , \temp414[7] , \temp414[6] , 
        \temp414[5] , \temp414[4] , \temp414[3] , \temp414[2] , \temp414[1] , 
        \temp414[0] }), .B(InEdges[63:48]), .LEQ(n918), .TC(n918), .GE_GT(n118
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_4 lte_55_4 ( .A({\temp504[15] , 
        \temp504[14] , \temp504[13] , \temp504[12] , \temp504[11] , 
        \temp504[10] , \temp504[9] , \temp504[8] , \temp504[7] , \temp504[6] , 
        \temp504[5] , \temp504[4] , \temp504[3] , \temp504[2] , \temp504[1] , 
        \temp504[0] }), .B(InEdges[79:64]), .LEQ(n917), .TC(n917), .GE_GT(n126
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_3 lte_55 ( .A(OutEdge), .B(InEdges
        [15:0]), .LEQ(n916), .TC(n916), .GE_GT(n94) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_2 lte_55_6 ( .A({\temp684[15] , 
        \temp684[14] , \temp684[13] , \temp684[12] , \temp684[11] , 
        \temp684[10] , \temp684[9] , \temp684[8] , \temp684[7] , \temp684[6] , 
        \temp684[5] , \temp684[4] , \temp684[3] , \temp684[2] , \temp684[1] , 
        \temp684[0] }), .B(InEdges[111:96]), .LEQ(n915), .TC(n915), .GE_GT(
        n142) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_1 lte_55_2 ( .A({\temp324[15] , 
        \temp324[14] , \temp324[13] , \temp324[12] , \temp324[11] , 
        \temp324[10] , \temp324[9] , \temp324[8] , \temp324[7] , \temp324[6] , 
        \temp324[5] , \temp324[4] , \temp324[3] , \temp324[2] , \temp324[1] , 
        \temp324[0] }), .B(InEdges[47:32]), .LEQ(n914), .TC(n914), .GE_GT(n110
        ) );
    NodeAux_INDEGREE7_SOURCE0_DW01_cmp2_16_0 lte_55_1 ( .A({\temp230[15] , 
        \temp230[14] , \temp230[13] , \temp230[12] , \temp230[11] , 
        \temp230[10] , \temp230[9] , \temp230[8] , \temp230[7] , \temp230[6] , 
        \temp230[5] , \temp230[4] , \temp230[3] , \temp230[2] , \temp230[1] , 
        \temp230[0] }), .B(InEdges[31:16]), .LEQ(n913), .TC(n913), .GE_GT(n102
        ) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
input  [9:0] WeightAddr;
input  [9:0] Eid;
output [2:0] PathData;
input  [15:0] WeightData;
input  [6:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[15:0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE1 n_1_1 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE0 n_1_0 ( .Nid(Nid), .InEdges(InEdges[15:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges[63:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE5_SOURCE0 n_5_0 ( .Nid(Nid), .InEdges(InEdges[79:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[31:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE0 n_6_0 ( .Nid(Nid), .InEdges(InEdges[95:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE7_SOURCE0 n_7_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[47:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID16_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID17_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID18_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID19_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID64 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID65 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID66 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID67 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID68 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID69 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID20_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID70 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID71 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID72 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID73 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID21_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID74 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID75 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID22_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID76 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID77 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID78 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID23_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID79 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID24_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID80 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID81 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID82 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID83 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID84 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID85 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID86 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID25_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID87 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID88 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID26_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID89 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID90 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID91 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID92 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID27_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID93 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID94 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID95 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID96 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID97 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID98 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID28_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID99 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID29_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID30_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID31_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID32_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID33_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID34_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID35_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID36_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID37_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID38_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID39_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID40_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID41_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID42_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID43_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID44_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID45_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID46_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID47_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID48_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID49_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID50_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID51_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID52_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID53_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID54_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID55_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID56_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID57_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID224 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID225 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID226 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID58_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID227 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID228 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID229 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID230 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID231 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID232 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID59_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID233 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID234 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID235 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID236 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID237 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID238 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID60_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID239 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID240 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID241 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID242 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID243 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID61_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID244 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID62_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID245 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID246 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID247 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID248 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID249 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID250 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID63_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID251 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID252 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID253 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID254 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID255 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID256 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID64_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID257 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID258 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID259 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID260 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID261 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID65_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID262 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID263 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID264 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID66_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID265 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID266 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID267 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID268 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID269 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID67_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID270 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID271 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID272 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID68_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID273 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID274 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID275 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID276 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID277 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID278 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID279 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID69_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID280 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID281 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID70_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID282 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID283 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID284 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID285 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID71_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID286 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID287 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID288 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID289 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID290 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID291 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID292 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID72_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID293 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID294 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID295 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID73_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID296 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID297 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID298 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID299 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID300 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID301 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID74_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID302 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID75_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID303 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID304 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID305 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID306 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID307 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID308 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID76_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID309 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID77_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID310 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID311 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID312 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID313 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID314 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID315 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID316 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID78_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID317 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID318 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID319 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID79_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID320 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID321 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID322 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID80_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID323 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID324 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID81_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID325 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID326 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID82_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID327 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID83_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID328 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID329 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID330 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID331 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID332 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID333 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID334 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID84_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID335 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID336 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID337 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID338 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID339 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID85_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID340 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID86_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID341 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID342 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID343 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID344 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID87_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID345 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID346 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID347 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID348 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID349 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID350 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID88_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID351 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID352 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID353 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID354 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID355 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID89_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID356 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID357 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID358 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID359 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID360 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID90_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID361 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID362 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID363 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID364 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID365 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID91_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID366 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID367 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID368 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID369 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID370 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID92_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID371 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID372 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID373 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID374 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID375 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID376 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID377 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID93_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID378 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID379 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID380 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID94_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID381 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID95_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID382 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID383 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID384 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID385 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID96_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID386 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID387 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID388 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID97_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID389 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID390 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID391 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID392 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID98_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID393 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID394 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID395 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID396 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID397 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID398 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID99_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID399 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID400 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID401 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID100_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID402 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID403 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID404 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID405 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID101_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID406 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID407 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID408 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID409 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID102_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID410 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID411 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID412 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID413 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID414 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID415 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID416 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID103_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID417 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID104_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID418 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID419 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID420 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID421 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID105_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID422 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID423 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID424 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID425 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID426 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID427 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID106_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID428 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID429 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID430 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID431 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID107_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID432 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID433 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID434 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID435 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID436 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID437 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID438 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID108_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID439 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID440 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID441 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID442 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID443 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID109_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID444 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID110_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID445 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID446 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID111_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID447 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID448 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID449 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID450 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID451 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID112_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID452 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID453 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID454 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID455 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID456 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID457 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID458 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID113_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [111:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID459 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID460 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID461 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID462 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID463 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID464 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID465 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID114_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [15:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID466 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID115_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID467 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID468 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID116_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID469 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID470 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID471 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID472 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID473 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID474 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID117_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID475 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID476 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID477 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID118_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID478 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID479 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID480 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID119_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [95:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID481 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID482 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID483 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID484 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID485 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID486 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID120_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID487 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID488 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID489 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID490 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID491 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID121_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID492 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID493 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID494 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID122_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID495 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID496 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID123_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [47:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID497 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID498 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID499 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID124_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID500 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID501 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID502 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID503 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID125_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [31:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID504 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID505 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID126_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [63:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID506 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID507 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID508 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID509 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID127_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [79:0] InEdges;
output [15:0] OutEdge;
input  [6:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID510 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID511 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID512 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID513 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID514 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [15:0] InEdge;
input  [9:0] WeightAddr;
output [15:0] OutEdge;
input  [15:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [9:0] WeightAddr;
input  [15:0] WeightData;
input  [6:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire [15:0] In0;
    wire [15:0] Out0;
    wire [47:0] In1;
    wire [15:0] Out1;
    wire [47:0] In2;
    wire [15:0] Out2;
    wire [47:0] In3;
    wire [15:0] Out3;
    wire [31:0] In4;
    wire [15:0] Out4;
    wire [111:0] In5;
    wire [15:0] Out5;
    wire [111:0] In6;
    wire [15:0] Out6;
    wire [63:0] In7;
    wire [15:0] Out7;
    wire [95:0] In8;
    wire [15:0] Out8;
    wire [15:0] In9;
    wire [15:0] Out9;
    wire [63:0] In10;
    wire [15:0] Out10;
    wire [15:0] In11;
    wire [15:0] Out11;
    wire [31:0] In12;
    wire [15:0] Out12;
    wire [95:0] In13;
    wire [15:0] Out13;
    wire [31:0] In14;
    wire [15:0] Out14;
    wire [31:0] In15;
    wire [15:0] Out15;
    wire [15:0] In16;
    wire [15:0] Out16;
    wire [95:0] In17;
    wire [15:0] Out17;
    wire [47:0] In18;
    wire [15:0] Out18;
    wire [95:0] In19;
    wire [15:0] Out19;
    wire [63:0] In20;
    wire [15:0] Out20;
    wire [31:0] In21;
    wire [15:0] Out21;
    wire [47:0] In22;
    wire [15:0] Out22;
    wire [15:0] In23;
    wire [15:0] Out23;
    wire [111:0] In24;
    wire [15:0] Out24;
    wire [31:0] In25;
    wire [15:0] Out25;
    wire [63:0] In26;
    wire [15:0] Out26;
    wire [95:0] In27;
    wire [15:0] Out27;
    wire [95:0] In28;
    wire [15:0] Out28;
    wire [31:0] In29;
    wire [15:0] Out29;
    wire [95:0] In30;
    wire [15:0] Out30;
    wire [95:0] In31;
    wire [15:0] Out31;
    wire [111:0] In32;
    wire [15:0] Out32;
    wire [47:0] In33;
    wire [15:0] Out33;
    wire [79:0] In34;
    wire [15:0] Out34;
    wire [111:0] In35;
    wire [15:0] Out35;
    wire [63:0] In36;
    wire [15:0] Out36;
    wire [31:0] In37;
    wire [15:0] Out37;
    wire [79:0] In38;
    wire [15:0] Out38;
    wire [79:0] In39;
    wire [15:0] Out39;
    wire [15:0] In40;
    wire [15:0] Out40;
    wire [15:0] In41;
    wire [15:0] Out41;
    wire [111:0] In42;
    wire [15:0] Out42;
    wire [63:0] In43;
    wire [15:0] Out43;
    wire [79:0] In44;
    wire [15:0] Out44;
    wire [31:0] In45;
    wire [15:0] Out45;
    wire [95:0] In46;
    wire [15:0] Out46;
    wire [111:0] In47;
    wire [15:0] Out47;
    wire [31:0] In48;
    wire [15:0] Out48;
    wire [31:0] In49;
    wire [15:0] Out49;
    wire [95:0] In50;
    wire [15:0] Out50;
    wire [15:0] In51;
    wire [15:0] Out51;
    wire [63:0] In52;
    wire [15:0] Out52;
    wire [79:0] In53;
    wire [15:0] Out53;
    wire [79:0] In54;
    wire [15:0] Out54;
    wire [79:0] In55;
    wire [15:0] Out55;
    wire [31:0] In56;
    wire [15:0] Out56;
    wire [79:0] In57;
    wire [15:0] Out57;
    wire [95:0] In58;
    wire [15:0] Out58;
    wire [95:0] In59;
    wire [15:0] Out59;
    wire [79:0] In60;
    wire [15:0] Out60;
    wire [15:0] In61;
    wire [15:0] Out61;
    wire [95:0] In62;
    wire [15:0] Out62;
    wire [95:0] In63;
    wire [15:0] Out63;
    wire [79:0] In64;
    wire [15:0] Out64;
    wire [47:0] In65;
    wire [15:0] Out65;
    wire [79:0] In66;
    wire [15:0] Out66;
    wire [47:0] In67;
    wire [15:0] Out67;
    wire [111:0] In68;
    wire [15:0] Out68;
    wire [31:0] In69;
    wire [15:0] Out69;
    wire [63:0] In70;
    wire [15:0] Out70;
    wire [111:0] In71;
    wire [15:0] Out71;
    wire [47:0] In72;
    wire [15:0] Out72;
    wire [95:0] In73;
    wire [15:0] Out73;
    wire [15:0] In74;
    wire [15:0] Out74;
    wire [95:0] In75;
    wire [15:0] Out75;
    wire [15:0] In76;
    wire [15:0] Out76;
    wire [111:0] In77;
    wire [15:0] Out77;
    wire [47:0] In78;
    wire [15:0] Out78;
    wire [47:0] In79;
    wire [15:0] Out79;
    wire [31:0] In80;
    wire [15:0] Out80;
    wire [31:0] In81;
    wire [15:0] Out81;
    wire [15:0] In82;
    wire [15:0] Out82;
    wire [111:0] In83;
    wire [15:0] Out83;
    wire [79:0] In84;
    wire [15:0] Out84;
    wire [15:0] In85;
    wire [15:0] Out85;
    wire [63:0] In86;
    wire [15:0] Out86;
    wire [95:0] In87;
    wire [15:0] Out87;
    wire [79:0] In88;
    wire [15:0] Out88;
    wire [79:0] In89;
    wire [15:0] Out89;
    wire [79:0] In90;
    wire [15:0] Out90;
    wire [79:0] In91;
    wire [15:0] Out91;
    wire [111:0] In92;
    wire [15:0] Out92;
    wire [47:0] In93;
    wire [15:0] Out93;
    wire [15:0] In94;
    wire [15:0] Out94;
    wire [63:0] In95;
    wire [15:0] Out95;
    wire [47:0] In96;
    wire [15:0] Out96;
    wire [63:0] In97;
    wire [15:0] Out97;
    wire [95:0] In98;
    wire [15:0] Out98;
    wire [47:0] In99;
    wire [15:0] Out99;
    wire [63:0] In100;
    wire [15:0] Out100;
    wire [63:0] In101;
    wire [15:0] Out101;
    wire [111:0] In102;
    wire [15:0] Out102;
    wire [15:0] In103;
    wire [15:0] Out103;
    wire [63:0] In104;
    wire [15:0] Out104;
    wire [95:0] In105;
    wire [15:0] Out105;
    wire [63:0] In106;
    wire [15:0] Out106;
    wire [111:0] In107;
    wire [15:0] Out107;
    wire [79:0] In108;
    wire [15:0] Out108;
    wire [15:0] In109;
    wire [15:0] Out109;
    wire [31:0] In110;
    wire [15:0] Out110;
    wire [79:0] In111;
    wire [15:0] Out111;
    wire [111:0] In112;
    wire [15:0] Out112;
    wire [111:0] In113;
    wire [15:0] Out113;
    wire [15:0] In114;
    wire [15:0] Out114;
    wire [31:0] In115;
    wire [15:0] Out115;
    wire [95:0] In116;
    wire [15:0] Out116;
    wire [47:0] In117;
    wire [15:0] Out117;
    wire [47:0] In118;
    wire [15:0] Out118;
    wire [95:0] In119;
    wire [15:0] Out119;
    wire [79:0] In120;
    wire [15:0] Out120;
    wire [47:0] In121;
    wire [15:0] Out121;
    wire [31:0] In122;
    wire [15:0] Out122;
    wire [47:0] In123;
    wire [15:0] Out123;
    wire [63:0] In124;
    wire [15:0] Out124;
    wire [31:0] In125;
    wire [15:0] Out125;
    wire [63:0] In126;
    wire [15:0] Out126;
    wire [79:0] In127;
    wire [15:0] Out127;

    Node_NID0_INDEGREE1 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out103), .OutEdge(In0[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE3 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out55), .OutEdge(In1[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out122), .OutEdge(In1[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out32), .OutEdge(In1[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE3 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out94), .OutEdge(In2[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out76), .OutEdge(In2[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out51), .OutEdge(In2[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE3 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out23), .OutEdge(In3[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out70), .OutEdge(In3[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out80), .OutEdge(In3[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE2 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out33), .OutEdge(In4[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out44), .OutEdge(In4[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE7 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out54), .OutEdge(In5[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out70), .OutEdge(In5[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out124), .OutEdge(In5[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out15), .OutEdge(In5[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out78), .OutEdge(In5[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out76), .OutEdge(In5[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out75), .OutEdge(In5[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE7 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out28), .OutEdge(In6[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out83), .OutEdge(In6[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out8), .OutEdge(In6[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out97), .OutEdge(In6[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out5), .OutEdge(In6[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out85), .OutEdge(In6[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out47), .OutEdge(In6[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE4 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out19), .OutEdge(In7[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out69), .OutEdge(In7[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out39), .OutEdge(In7[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out22), .OutEdge(In7[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE6 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out120), .OutEdge(In8[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out23), .OutEdge(In8[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out32), .OutEdge(In8[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out89), .OutEdge(In8[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out55), .OutEdge(In8[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out21), .OutEdge(In8[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE1 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out87), .OutEdge(In9[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE4 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out2), .OutEdge(In10[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out13), .OutEdge(In10[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out107), .OutEdge(In10[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out18), .OutEdge(In10[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE1 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out7), .OutEdge(In11[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE2 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out125), .OutEdge(In12[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out54), .OutEdge(In12[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE6 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out107), .OutEdge(In13[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out63), .OutEdge(In13[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out94), .OutEdge(In13[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out65), .OutEdge(In13[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out116), .OutEdge(In13[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out122), .OutEdge(In13[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE2 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out16), .OutEdge(In14[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out2), .OutEdge(In14[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE2 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out66), .OutEdge(In15[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out33), .OutEdge(In15[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID16_INDEGREE1 n16 ( .InEdges(In16), .OutEdge(Out16),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out120), .OutEdge(In16[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID17_INDEGREE6 n17 ( .InEdges(In17), .OutEdge(Out17),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out127), .OutEdge(In17[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out119), .OutEdge(In17[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out32), .OutEdge(In17[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out117), .OutEdge(In17[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out50), .OutEdge(In17[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out86), .OutEdge(In17[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID18_INDEGREE3 n18 ( .InEdges(In18), .OutEdge(Out18),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out93), .OutEdge(In18[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out96), .OutEdge(In18[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out3), .OutEdge(In18[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID19_INDEGREE6 n19 ( .InEdges(In19), .OutEdge(Out19),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID64 e64 ( .InEdge(Out9), .OutEdge(In19[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID65 e65 ( .InEdge(Out59), .OutEdge(In19[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID66 e66 ( .InEdge(Out98), .OutEdge(In19[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID67 e67 ( .InEdge(Out30), .OutEdge(In19[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID68 e68 ( .InEdge(Out92), .OutEdge(In19[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID69 e69 ( .InEdge(Out11), .OutEdge(In19[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID20_INDEGREE4 n20 ( .InEdges(In20), .OutEdge(Out20),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID70 e70 ( .InEdge(Out40), .OutEdge(In20[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID71 e71 ( .InEdge(Out59), .OutEdge(In20[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID72 e72 ( .InEdge(Out113), .OutEdge(In20[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID73 e73 ( .InEdge(Out24), .OutEdge(In20[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID21_INDEGREE2 n21 ( .InEdges(In21), .OutEdge(Out21),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID74 e74 ( .InEdge(Out25), .OutEdge(In21[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID75 e75 ( .InEdge(Out72), .OutEdge(In21[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID22_INDEGREE3 n22 ( .InEdges(In22), .OutEdge(Out22),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID76 e76 ( .InEdge(Out35), .OutEdge(In22[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID77 e77 ( .InEdge(Out37), .OutEdge(In22[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID78 e78 ( .InEdge(Out63), .OutEdge(In22[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID23_INDEGREE1 n23 ( .InEdges(In23), .OutEdge(Out23),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID79 e79 ( .InEdge(Out68), .OutEdge(In23[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID24_INDEGREE7 n24 ( .InEdges(In24), .OutEdge(Out24),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID80 e80 ( .InEdge(Out50), .OutEdge(In24[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID81 e81 ( .InEdge(Out93), .OutEdge(In24[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID82 e82 ( .InEdge(Out107), .OutEdge(In24[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID83 e83 ( .InEdge(Out103), .OutEdge(In24[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID84 e84 ( .InEdge(Out94), .OutEdge(In24[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID85 e85 ( .InEdge(Out65), .OutEdge(In24[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID86 e86 ( .InEdge(Out61), .OutEdge(In24[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID25_INDEGREE2 n25 ( .InEdges(In25), .OutEdge(Out25),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID87 e87 ( .InEdge(Out93), .OutEdge(In25[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID88 e88 ( .InEdge(Out115), .OutEdge(In25[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID26_INDEGREE4 n26 ( .InEdges(In26), .OutEdge(Out26),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID89 e89 ( .InEdge(Out123), .OutEdge(In26[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID90 e90 ( .InEdge(Out69), .OutEdge(In26[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID91 e91 ( .InEdge(Out70), .OutEdge(In26[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID92 e92 ( .InEdge(Out52), .OutEdge(In26[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID27_INDEGREE6 n27 ( .InEdges(In27), .OutEdge(Out27),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID93 e93 ( .InEdge(Out78), .OutEdge(In27[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID94 e94 ( .InEdge(Out125), .OutEdge(In27[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID95 e95 ( .InEdge(Out96), .OutEdge(In27[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID96 e96 ( .InEdge(Out50), .OutEdge(In27[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID97 e97 ( .InEdge(Out68), .OutEdge(In27[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID98 e98 ( .InEdge(Out6), .OutEdge(In27[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID28_INDEGREE6 n28 ( .InEdges(In28), .OutEdge(Out28),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID99 e99 ( .InEdge(Out3), .OutEdge(In28[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID100 e100 ( .InEdge(Out69), .OutEdge(In28[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID101 e101 ( .InEdge(Out60), .OutEdge(In28[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID102 e102 ( .InEdge(Out109), .OutEdge(In28[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID103 e103 ( .InEdge(Out122), .OutEdge(In28[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID104 e104 ( .InEdge(Out35), .OutEdge(In28[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID29_INDEGREE2 n29 ( .InEdges(In29), .OutEdge(Out29),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID105 e105 ( .InEdge(Out120), .OutEdge(In29[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID106 e106 ( .InEdge(Out75), .OutEdge(In29[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID30_INDEGREE6 n30 ( .InEdges(In30), .OutEdge(Out30),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID107 e107 ( .InEdge(Out76), .OutEdge(In30[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID108 e108 ( .InEdge(Out78), .OutEdge(In30[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID109 e109 ( .InEdge(Out45), .OutEdge(In30[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID110 e110 ( .InEdge(Out35), .OutEdge(In30[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID111 e111 ( .InEdge(Out80), .OutEdge(In30[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID112 e112 ( .InEdge(Out70), .OutEdge(In30[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID31_INDEGREE6 n31 ( .InEdges(In31), .OutEdge(Out31),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID113 e113 ( .InEdge(Out33), .OutEdge(In31[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID114 e114 ( .InEdge(Out87), .OutEdge(In31[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID115 e115 ( .InEdge(Out4), .OutEdge(In31[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID116 e116 ( .InEdge(Out88), .OutEdge(In31[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID117 e117 ( .InEdge(Out103), .OutEdge(In31[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID118 e118 ( .InEdge(Out100), .OutEdge(In31[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID32_INDEGREE7 n32 ( .InEdges(In32), .OutEdge(Out32),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID119 e119 ( .InEdge(Out101), .OutEdge(In32[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID120 e120 ( .InEdge(Out119), .OutEdge(In32[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID121 e121 ( .InEdge(Out55), .OutEdge(In32[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID122 e122 ( .InEdge(Out16), .OutEdge(In32[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID123 e123 ( .InEdge(Out121), .OutEdge(In32[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID124 e124 ( .InEdge(Out35), .OutEdge(In32[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID125 e125 ( .InEdge(Out85), .OutEdge(In32[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID33_INDEGREE3 n33 ( .InEdges(In33), .OutEdge(Out33),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID126 e126 ( .InEdge(Out60), .OutEdge(In33[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID127 e127 ( .InEdge(Out103), .OutEdge(In33[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID128 e128 ( .InEdge(Out7), .OutEdge(In33[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID34_INDEGREE5 n34 ( .InEdges(In34), .OutEdge(Out34),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID129 e129 ( .InEdge(Out114), .OutEdge(In34[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID130 e130 ( .InEdge(Out58), .OutEdge(In34[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID131 e131 ( .InEdge(Out99), .OutEdge(In34[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID132 e132 ( .InEdge(Out35), .OutEdge(In34[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID133 e133 ( .InEdge(Out42), .OutEdge(In34[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID35_INDEGREE7 n35 ( .InEdges(In35), .OutEdge(Out35),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID134 e134 ( .InEdge(Out15), .OutEdge(In35[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID135 e135 ( .InEdge(Out25), .OutEdge(In35[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID136 e136 ( .InEdge(Out116), .OutEdge(In35[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID137 e137 ( .InEdge(Out105), .OutEdge(In35[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID138 e138 ( .InEdge(Out22), .OutEdge(In35[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID139 e139 ( .InEdge(Out111), .OutEdge(In35[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID140 e140 ( .InEdge(Out34), .OutEdge(In35[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID36_INDEGREE4 n36 ( .InEdges(In36), .OutEdge(Out36),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID141 e141 ( .InEdge(Out113), .OutEdge(In36[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID142 e142 ( .InEdge(Out22), .OutEdge(In36[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID143 e143 ( .InEdge(Out106), .OutEdge(In36[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID144 e144 ( .InEdge(Out61), .OutEdge(In36[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID37_INDEGREE2 n37 ( .InEdges(In37), .OutEdge(Out37),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID145 e145 ( .InEdge(Out121), .OutEdge(In37[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID146 e146 ( .InEdge(Out117), .OutEdge(In37[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID38_INDEGREE5 n38 ( .InEdges(In38), .OutEdge(Out38),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID147 e147 ( .InEdge(Out1), .OutEdge(In38[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID148 e148 ( .InEdge(Out78), .OutEdge(In38[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID149 e149 ( .InEdge(Out74), .OutEdge(In38[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID150 e150 ( .InEdge(Out109), .OutEdge(In38[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID151 e151 ( .InEdge(Out0), .OutEdge(In38[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID39_INDEGREE5 n39 ( .InEdges(In39), .OutEdge(Out39),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID152 e152 ( .InEdge(Out101), .OutEdge(In39[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID153 e153 ( .InEdge(Out8), .OutEdge(In39[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID154 e154 ( .InEdge(Out66), .OutEdge(In39[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID155 e155 ( .InEdge(Out10), .OutEdge(In39[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID156 e156 ( .InEdge(Out37), .OutEdge(In39[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID40_INDEGREE1 n40 ( .InEdges(In40), .OutEdge(Out40),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID157 e157 ( .InEdge(Out79), .OutEdge(In40[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID41_INDEGREE1 n41 ( .InEdges(In41), .OutEdge(Out41),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID158 e158 ( .InEdge(Out78), .OutEdge(In41[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID42_INDEGREE7 n42 ( .InEdges(In42), .OutEdge(Out42),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID159 e159 ( .InEdge(Out66), .OutEdge(In42[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID160 e160 ( .InEdge(Out122), .OutEdge(In42[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID161 e161 ( .InEdge(Out104), .OutEdge(In42[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID162 e162 ( .InEdge(Out19), .OutEdge(In42[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID163 e163 ( .InEdge(Out102), .OutEdge(In42[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID164 e164 ( .InEdge(Out12), .OutEdge(In42[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID165 e165 ( .InEdge(Out13), .OutEdge(In42[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID43_INDEGREE4 n43 ( .InEdges(In43), .OutEdge(Out43),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID166 e166 ( .InEdge(Out44), .OutEdge(In43[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID167 e167 ( .InEdge(Out124), .OutEdge(In43[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID168 e168 ( .InEdge(Out67), .OutEdge(In43[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID169 e169 ( .InEdge(Out78), .OutEdge(In43[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID44_INDEGREE5 n44 ( .InEdges(In44), .OutEdge(Out44),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID170 e170 ( .InEdge(Out33), .OutEdge(In44[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID171 e171 ( .InEdge(Out112), .OutEdge(In44[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID172 e172 ( .InEdge(Out90), .OutEdge(In44[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID173 e173 ( .InEdge(Out45), .OutEdge(In44[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID174 e174 ( .InEdge(Out23), .OutEdge(In44[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID45_INDEGREE2 n45 ( .InEdges(In45), .OutEdge(Out45),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID175 e175 ( .InEdge(Out14), .OutEdge(In45[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID176 e176 ( .InEdge(Out58), .OutEdge(In45[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID46_INDEGREE6 n46 ( .InEdges(In46), .OutEdge(Out46),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID177 e177 ( .InEdge(Out84), .OutEdge(In46[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID178 e178 ( .InEdge(Out108), .OutEdge(In46[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID179 e179 ( .InEdge(Out54), .OutEdge(In46[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID180 e180 ( .InEdge(Out72), .OutEdge(In46[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID181 e181 ( .InEdge(Out34), .OutEdge(In46[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID182 e182 ( .InEdge(Out95), .OutEdge(In46[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID47_INDEGREE7 n47 ( .InEdges(In47), .OutEdge(Out47),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID183 e183 ( .InEdge(Out20), .OutEdge(In47[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID184 e184 ( .InEdge(Out62), .OutEdge(In47[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID185 e185 ( .InEdge(Out82), .OutEdge(In47[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID186 e186 ( .InEdge(Out89), .OutEdge(In47[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID187 e187 ( .InEdge(Out33), .OutEdge(In47[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID188 e188 ( .InEdge(Out65), .OutEdge(In47[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID189 e189 ( .InEdge(Out80), .OutEdge(In47[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID48_INDEGREE2 n48 ( .InEdges(In48), .OutEdge(Out48),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID190 e190 ( .InEdge(Out116), .OutEdge(In48[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID191 e191 ( .InEdge(Out40), .OutEdge(In48[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID49_INDEGREE2 n49 ( .InEdges(In49), .OutEdge(Out49),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID192 e192 ( .InEdge(Out18), .OutEdge(In49[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID193 e193 ( .InEdge(Out114), .OutEdge(In49[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID50_INDEGREE6 n50 ( .InEdges(In50), .OutEdge(Out50),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID194 e194 ( .InEdge(Out119), .OutEdge(In50[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID195 e195 ( .InEdge(Out71), .OutEdge(In50[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID196 e196 ( .InEdge(Out40), .OutEdge(In50[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID197 e197 ( .InEdge(Out126), .OutEdge(In50[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID198 e198 ( .InEdge(Out108), .OutEdge(In50[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID199 e199 ( .InEdge(Out56), .OutEdge(In50[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID51_INDEGREE1 n51 ( .InEdges(In51), .OutEdge(Out51),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID200 e200 ( .InEdge(Out45), .OutEdge(In51[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID52_INDEGREE4 n52 ( .InEdges(In52), .OutEdge(Out52),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID201 e201 ( .InEdge(Out110), .OutEdge(In52[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID202 e202 ( .InEdge(Out93), .OutEdge(In52[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID203 e203 ( .InEdge(Out67), .OutEdge(In52[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID204 e204 ( .InEdge(Out55), .OutEdge(In52[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID53_INDEGREE5 n53 ( .InEdges(In53), .OutEdge(Out53),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID205 e205 ( .InEdge(Out113), .OutEdge(In53[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID206 e206 ( .InEdge(Out20), .OutEdge(In53[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID207 e207 ( .InEdge(Out46), .OutEdge(In53[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID208 e208 ( .InEdge(Out80), .OutEdge(In53[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID209 e209 ( .InEdge(Out4), .OutEdge(In53[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID54_INDEGREE5 n54 ( .InEdges(In54), .OutEdge(Out54),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID210 e210 ( .InEdge(Out83), .OutEdge(In54[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID211 e211 ( .InEdge(Out17), .OutEdge(In54[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID212 e212 ( .InEdge(Out55), .OutEdge(In54[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID213 e213 ( .InEdge(Out4), .OutEdge(In54[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID214 e214 ( .InEdge(Out123), .OutEdge(In54[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID55_INDEGREE5 n55 ( .InEdges(In55), .OutEdge(Out55),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID215 e215 ( .InEdge(Out46), .OutEdge(In55[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID216 e216 ( .InEdge(Out42), .OutEdge(In55[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID217 e217 ( .InEdge(Out32), .OutEdge(In55[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID218 e218 ( .InEdge(Out115), .OutEdge(In55[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID219 e219 ( .InEdge(Out98), .OutEdge(In55[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID56_INDEGREE2 n56 ( .InEdges(In56), .OutEdge(Out56),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID220 e220 ( .InEdge(Out60), .OutEdge(In56[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID221 e221 ( .InEdge(Out124), .OutEdge(In56[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID57_INDEGREE5 n57 ( .InEdges(In57), .OutEdge(Out57),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID222 e222 ( .InEdge(Out106), .OutEdge(In57[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID223 e223 ( .InEdge(Out63), .OutEdge(In57[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID224 e224 ( .InEdge(Out109), .OutEdge(In57[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID225 e225 ( .InEdge(Out24), .OutEdge(In57[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID226 e226 ( .InEdge(Out64), .OutEdge(In57[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID58_INDEGREE6 n58 ( .InEdges(In58), .OutEdge(Out58),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID227 e227 ( .InEdge(Out86), .OutEdge(In58[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID228 e228 ( .InEdge(Out37), .OutEdge(In58[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID229 e229 ( .InEdge(Out79), .OutEdge(In58[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID230 e230 ( .InEdge(Out112), .OutEdge(In58[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID231 e231 ( .InEdge(Out46), .OutEdge(In58[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID232 e232 ( .InEdge(Out76), .OutEdge(In58[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID59_INDEGREE6 n59 ( .InEdges(In59), .OutEdge(Out59),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID233 e233 ( .InEdge(Out31), .OutEdge(In59[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID234 e234 ( .InEdge(Out22), .OutEdge(In59[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID235 e235 ( .InEdge(Out70), .OutEdge(In59[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID236 e236 ( .InEdge(Out120), .OutEdge(In59[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID237 e237 ( .InEdge(Out39), .OutEdge(In59[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID238 e238 ( .InEdge(Out49), .OutEdge(In59[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID60_INDEGREE5 n60 ( .InEdges(In60), .OutEdge(Out60),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID239 e239 ( .InEdge(Out59), .OutEdge(In60[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID240 e240 ( .InEdge(Out118), .OutEdge(In60[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID241 e241 ( .InEdge(Out3), .OutEdge(In60[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID242 e242 ( .InEdge(Out98), .OutEdge(In60[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID243 e243 ( .InEdge(Out77), .OutEdge(In60[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID61_INDEGREE1 n61 ( .InEdges(In61), .OutEdge(Out61),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID244 e244 ( .InEdge(Out110), .OutEdge(In61[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID62_INDEGREE6 n62 ( .InEdges(In62), .OutEdge(Out62),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID245 e245 ( .InEdge(Out7), .OutEdge(In62[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID246 e246 ( .InEdge(Out38), .OutEdge(In62[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID247 e247 ( .InEdge(Out88), .OutEdge(In62[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID248 e248 ( .InEdge(Out33), .OutEdge(In62[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID249 e249 ( .InEdge(Out41), .OutEdge(In62[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID250 e250 ( .InEdge(Out28), .OutEdge(In62[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID63_INDEGREE6 n63 ( .InEdges(In63), .OutEdge(Out63),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID251 e251 ( .InEdge(Out93), .OutEdge(In63[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID252 e252 ( .InEdge(Out49), .OutEdge(In63[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID253 e253 ( .InEdge(Out33), .OutEdge(In63[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID254 e254 ( .InEdge(Out72), .OutEdge(In63[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID255 e255 ( .InEdge(Out48), .OutEdge(In63[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID256 e256 ( .InEdge(Out69), .OutEdge(In63[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID64_INDEGREE5 n64 ( .InEdges(In64), .OutEdge(Out64),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID257 e257 ( .InEdge(Out90), .OutEdge(In64[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID258 e258 ( .InEdge(Out13), .OutEdge(In64[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID259 e259 ( .InEdge(Out82), .OutEdge(In64[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID260 e260 ( .InEdge(Out83), .OutEdge(In64[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID261 e261 ( .InEdge(Out68), .OutEdge(In64[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID65_INDEGREE3 n65 ( .InEdges(In65), .OutEdge(Out65),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID262 e262 ( .InEdge(Out124), .OutEdge(In65[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID263 e263 ( .InEdge(Out119), .OutEdge(In65[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID264 e264 ( .InEdge(Out26), .OutEdge(In65[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID66_INDEGREE5 n66 ( .InEdges(In66), .OutEdge(Out66),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID265 e265 ( .InEdge(Out70), .OutEdge(In66[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID266 e266 ( .InEdge(Out68), .OutEdge(In66[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID267 e267 ( .InEdge(Out116), .OutEdge(In66[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID268 e268 ( .InEdge(Out114), .OutEdge(In66[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID269 e269 ( .InEdge(Out111), .OutEdge(In66[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID67_INDEGREE3 n67 ( .InEdges(In67), .OutEdge(Out67),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID270 e270 ( .InEdge(Out29), .OutEdge(In67[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID271 e271 ( .InEdge(Out56), .OutEdge(In67[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID272 e272 ( .InEdge(Out90), .OutEdge(In67[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID68_INDEGREE7 n68 ( .InEdges(In68), .OutEdge(Out68),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID273 e273 ( .InEdge(Out33), .OutEdge(In68[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID274 e274 ( .InEdge(Out82), .OutEdge(In68[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID275 e275 ( .InEdge(Out77), .OutEdge(In68[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID276 e276 ( .InEdge(Out14), .OutEdge(In68[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID277 e277 ( .InEdge(Out48), .OutEdge(In68[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID278 e278 ( .InEdge(Out64), .OutEdge(In68[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID279 e279 ( .InEdge(Out103), .OutEdge(In68[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID69_INDEGREE2 n69 ( .InEdges(In69), .OutEdge(Out69),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID280 e280 ( .InEdge(Out21), .OutEdge(In69[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID281 e281 ( .InEdge(Out31), .OutEdge(In69[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID70_INDEGREE4 n70 ( .InEdges(In70), .OutEdge(Out70),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID282 e282 ( .InEdge(Out126), .OutEdge(In70[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID283 e283 ( .InEdge(Out107), .OutEdge(In70[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID284 e284 ( .InEdge(Out63), .OutEdge(In70[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID285 e285 ( .InEdge(Out6), .OutEdge(In70[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID71_INDEGREE7 n71 ( .InEdges(In71), .OutEdge(Out71),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID286 e286 ( .InEdge(Out98), .OutEdge(In71[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID287 e287 ( .InEdge(Out94), .OutEdge(In71[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID288 e288 ( .InEdge(Out74), .OutEdge(In71[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID289 e289 ( .InEdge(Out6), .OutEdge(In71[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID290 e290 ( .InEdge(Out112), .OutEdge(In71[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID291 e291 ( .InEdge(Out124), .OutEdge(In71[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID292 e292 ( .InEdge(Out31), .OutEdge(In71[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID72_INDEGREE3 n72 ( .InEdges(In72), .OutEdge(Out72),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID293 e293 ( .InEdge(Out47), .OutEdge(In72[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID294 e294 ( .InEdge(Out49), .OutEdge(In72[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID295 e295 ( .InEdge(Out100), .OutEdge(In72[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID73_INDEGREE6 n73 ( .InEdges(In73), .OutEdge(Out73),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID296 e296 ( .InEdge(Out33), .OutEdge(In73[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID297 e297 ( .InEdge(Out7), .OutEdge(In73[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID298 e298 ( .InEdge(Out16), .OutEdge(In73[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID299 e299 ( .InEdge(Out23), .OutEdge(In73[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID300 e300 ( .InEdge(Out64), .OutEdge(In73[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID301 e301 ( .InEdge(Out86), .OutEdge(In73[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID74_INDEGREE1 n74 ( .InEdges(In74), .OutEdge(Out74),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID302 e302 ( .InEdge(Out55), .OutEdge(In74[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID75_INDEGREE6 n75 ( .InEdges(In75), .OutEdge(Out75),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID303 e303 ( .InEdge(Out90), .OutEdge(In75[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID304 e304 ( .InEdge(Out18), .OutEdge(In75[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID305 e305 ( .InEdge(Out14), .OutEdge(In75[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID306 e306 ( .InEdge(Out2), .OutEdge(In75[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID307 e307 ( .InEdge(Out76), .OutEdge(In75[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID308 e308 ( .InEdge(Out74), .OutEdge(In75[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID76_INDEGREE1 n76 ( .InEdges(In76), .OutEdge(Out76),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID309 e309 ( .InEdge(Out9), .OutEdge(In76[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID77_INDEGREE7 n77 ( .InEdges(In77), .OutEdge(Out77),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID310 e310 ( .InEdge(Out118), .OutEdge(In77[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID311 e311 ( .InEdge(Out104), .OutEdge(In77[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID312 e312 ( .InEdge(Out92), .OutEdge(In77[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID313 e313 ( .InEdge(Out2), .OutEdge(In77[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID314 e314 ( .InEdge(Out4), .OutEdge(In77[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID315 e315 ( .InEdge(Out58), .OutEdge(In77[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID316 e316 ( .InEdge(Out73), .OutEdge(In77[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID78_INDEGREE3 n78 ( .InEdges(In78), .OutEdge(Out78),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID317 e317 ( .InEdge(Out46), .OutEdge(In78[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID318 e318 ( .InEdge(Out34), .OutEdge(In78[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID319 e319 ( .InEdge(Out127), .OutEdge(In78[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID79_INDEGREE3 n79 ( .InEdges(In79), .OutEdge(Out79),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID320 e320 ( .InEdge(Out69), .OutEdge(In79[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID321 e321 ( .InEdge(Out78), .OutEdge(In79[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID322 e322 ( .InEdge(Out105), .OutEdge(In79[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID80_INDEGREE2 n80 ( .InEdges(In80), .OutEdge(Out80),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID323 e323 ( .InEdge(Out99), .OutEdge(In80[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID324 e324 ( .InEdge(Out42), .OutEdge(In80[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID81_INDEGREE2 n81 ( .InEdges(In81), .OutEdge(Out81),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID325 e325 ( .InEdge(Out99), .OutEdge(In81[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID326 e326 ( .InEdge(Out10), .OutEdge(In81[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID82_INDEGREE1 n82 ( .InEdges(In82), .OutEdge(Out82),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID327 e327 ( .InEdge(Out26), .OutEdge(In82[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID83_INDEGREE7 n83 ( .InEdges(In83), .OutEdge(Out83),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID328 e328 ( .InEdge(Out42), .OutEdge(In83[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID329 e329 ( .InEdge(Out20), .OutEdge(In83[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID330 e330 ( .InEdge(Out59), .OutEdge(In83[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID331 e331 ( .InEdge(Out99), .OutEdge(In83[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID332 e332 ( .InEdge(Out95), .OutEdge(In83[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID333 e333 ( .InEdge(Out54), .OutEdge(In83[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID334 e334 ( .InEdge(Out43), .OutEdge(In83[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID84_INDEGREE5 n84 ( .InEdges(In84), .OutEdge(Out84),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID335 e335 ( .InEdge(Out4), .OutEdge(In84[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID336 e336 ( .InEdge(Out45), .OutEdge(In84[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID337 e337 ( .InEdge(Out57), .OutEdge(In84[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID338 e338 ( .InEdge(Out93), .OutEdge(In84[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID339 e339 ( .InEdge(Out59), .OutEdge(In84[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID85_INDEGREE1 n85 ( .InEdges(In85), .OutEdge(Out85),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID340 e340 ( .InEdge(Out0), .OutEdge(In85[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID86_INDEGREE4 n86 ( .InEdges(In86), .OutEdge(Out86),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID341 e341 ( .InEdge(Out16), .OutEdge(In86[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID342 e342 ( .InEdge(Out0), .OutEdge(In86[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID343 e343 ( .InEdge(Out89), .OutEdge(In86[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID344 e344 ( .InEdge(Out31), .OutEdge(In86[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID87_INDEGREE6 n87 ( .InEdges(In87), .OutEdge(Out87),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID345 e345 ( .InEdge(Out119), .OutEdge(In87[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID346 e346 ( .InEdge(Out91), .OutEdge(In87[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID347 e347 ( .InEdge(Out68), .OutEdge(In87[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID348 e348 ( .InEdge(Out86), .OutEdge(In87[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID349 e349 ( .InEdge(Out53), .OutEdge(In87[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID350 e350 ( .InEdge(Out85), .OutEdge(In87[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID88_INDEGREE5 n88 ( .InEdges(In88), .OutEdge(Out88),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID351 e351 ( .InEdge(Out91), .OutEdge(In88[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID352 e352 ( .InEdge(Out38), .OutEdge(In88[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID353 e353 ( .InEdge(Out89), .OutEdge(In88[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID354 e354 ( .InEdge(Out118), .OutEdge(In88[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID355 e355 ( .InEdge(Out96), .OutEdge(In88[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID89_INDEGREE5 n89 ( .InEdges(In89), .OutEdge(Out89),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID356 e356 ( .InEdge(Out83), .OutEdge(In89[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID357 e357 ( .InEdge(Out78), .OutEdge(In89[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID358 e358 ( .InEdge(Out17), .OutEdge(In89[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID359 e359 ( .InEdge(Out126), .OutEdge(In89[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID360 e360 ( .InEdge(Out101), .OutEdge(In89[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID90_INDEGREE5 n90 ( .InEdges(In90), .OutEdge(Out90),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID361 e361 ( .InEdge(Out79), .OutEdge(In90[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID362 e362 ( .InEdge(Out30), .OutEdge(In90[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID363 e363 ( .InEdge(Out33), .OutEdge(In90[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID364 e364 ( .InEdge(Out48), .OutEdge(In90[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID365 e365 ( .InEdge(Out107), .OutEdge(In90[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID91_INDEGREE5 n91 ( .InEdges(In91), .OutEdge(Out91),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID366 e366 ( .InEdge(Out92), .OutEdge(In91[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID367 e367 ( .InEdge(Out69), .OutEdge(In91[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID368 e368 ( .InEdge(Out20), .OutEdge(In91[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID369 e369 ( .InEdge(Out35), .OutEdge(In91[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID370 e370 ( .InEdge(Out34), .OutEdge(In91[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID92_INDEGREE7 n92 ( .InEdges(In92), .OutEdge(Out92),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID371 e371 ( .InEdge(Out81), .OutEdge(In92[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID372 e372 ( .InEdge(Out51), .OutEdge(In92[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID373 e373 ( .InEdge(Out121), .OutEdge(In92[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID374 e374 ( .InEdge(Out58), .OutEdge(In92[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID375 e375 ( .InEdge(Out67), .OutEdge(In92[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID376 e376 ( .InEdge(Out24), .OutEdge(In92[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID377 e377 ( .InEdge(Out17), .OutEdge(In92[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID93_INDEGREE3 n93 ( .InEdges(In93), .OutEdge(Out93),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID378 e378 ( .InEdge(Out116), .OutEdge(In93[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID379 e379 ( .InEdge(Out31), .OutEdge(In93[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID380 e380 ( .InEdge(Out109), .OutEdge(In93[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID94_INDEGREE1 n94 ( .InEdges(In94), .OutEdge(Out94),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID381 e381 ( .InEdge(Out99), .OutEdge(In94[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID95_INDEGREE4 n95 ( .InEdges(In95), .OutEdge(Out95),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID382 e382 ( .InEdge(Out122), .OutEdge(In95[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID383 e383 ( .InEdge(Out24), .OutEdge(In95[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID384 e384 ( .InEdge(Out60), .OutEdge(In95[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID385 e385 ( .InEdge(Out107), .OutEdge(In95[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID96_INDEGREE3 n96 ( .InEdges(In96), .OutEdge(Out96),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID386 e386 ( .InEdge(Out61), .OutEdge(In96[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID387 e387 ( .InEdge(Out105), .OutEdge(In96[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID388 e388 ( .InEdge(Out69), .OutEdge(In96[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID97_INDEGREE4 n97 ( .InEdges(In97), .OutEdge(Out97),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID389 e389 ( .InEdge(Out109), .OutEdge(In97[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID390 e390 ( .InEdge(Out43), .OutEdge(In97[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID391 e391 ( .InEdge(Out37), .OutEdge(In97[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID392 e392 ( .InEdge(Out27), .OutEdge(In97[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID98_INDEGREE6 n98 ( .InEdges(In98), .OutEdge(Out98),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID393 e393 ( .InEdge(Out33), .OutEdge(In98[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID394 e394 ( .InEdge(Out26), .OutEdge(In98[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID395 e395 ( .InEdge(Out89), .OutEdge(In98[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID396 e396 ( .InEdge(Out5), .OutEdge(In98[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID397 e397 ( .InEdge(Out74), .OutEdge(In98[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID398 e398 ( .InEdge(Out22), .OutEdge(In98[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID99_INDEGREE3 n99 ( .InEdges(In99), .OutEdge(Out99),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID399 e399 ( .InEdge(Out111), .OutEdge(In99[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID400 e400 ( .InEdge(Out98), .OutEdge(In99[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID401 e401 ( .InEdge(Out77), .OutEdge(In99[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID100_INDEGREE4 n100 ( .InEdges(In100), .OutEdge(Out100),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID402 e402 ( .InEdge(Out72), .OutEdge(In100[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID403 e403 ( .InEdge(Out8), .OutEdge(In100[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID404 e404 ( .InEdge(Out5), .OutEdge(In100[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID405 e405 ( .InEdge(Out61), .OutEdge(In100[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID101_INDEGREE4 n101 ( .InEdges(In101), .OutEdge(Out101),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID406 e406 ( .InEdge(Out13), .OutEdge(In101[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID407 e407 ( .InEdge(Out95), .OutEdge(In101[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID408 e408 ( .InEdge(Out94), .OutEdge(In101[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID409 e409 ( .InEdge(Out44), .OutEdge(In101[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID102_INDEGREE7 n102 ( .InEdges(In102), .OutEdge(Out102),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID410 e410 ( .InEdge(Out91), .OutEdge(In102[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID411 e411 ( .InEdge(Out99), .OutEdge(In102[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID412 e412 ( .InEdge(Out92), .OutEdge(In102[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID413 e413 ( .InEdge(Out60), .OutEdge(In102[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID414 e414 ( .InEdge(Out45), .OutEdge(In102[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID415 e415 ( .InEdge(Out107), .OutEdge(In102[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID416 e416 ( .InEdge(Out50), .OutEdge(In102[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID103_INDEGREE1 n103 ( .InEdges(In103), .OutEdge(Out103),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID417 e417 ( .InEdge(Out33), .OutEdge(In103[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID104_INDEGREE4 n104 ( .InEdges(In104), .OutEdge(Out104),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID418 e418 ( .InEdge(Out5), .OutEdge(In104[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID419 e419 ( .InEdge(Out21), .OutEdge(In104[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID420 e420 ( .InEdge(Out78), .OutEdge(In104[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID421 e421 ( .InEdge(Out29), .OutEdge(In104[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID105_INDEGREE6 n105 ( .InEdges(In105), .OutEdge(Out105),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID422 e422 ( .InEdge(Out80), .OutEdge(In105[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID423 e423 ( .InEdge(Out40), .OutEdge(In105[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID424 e424 ( .InEdge(Out118), .OutEdge(In105[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID425 e425 ( .InEdge(Out107), .OutEdge(In105[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID426 e426 ( .InEdge(Out8), .OutEdge(In105[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID427 e427 ( .InEdge(Out19), .OutEdge(In105[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID106_INDEGREE4 n106 ( .InEdges(In106), .OutEdge(Out106),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID428 e428 ( .InEdge(Out54), .OutEdge(In106[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID429 e429 ( .InEdge(Out95), .OutEdge(In106[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID430 e430 ( .InEdge(Out58), .OutEdge(In106[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID431 e431 ( .InEdge(Out73), .OutEdge(In106[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID107_INDEGREE7 n107 ( .InEdges(In107), .OutEdge(Out107),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID432 e432 ( .InEdge(Out125), .OutEdge(In107[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID433 e433 ( .InEdge(Out91), .OutEdge(In107[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID434 e434 ( .InEdge(Out100), .OutEdge(In107[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID435 e435 ( .InEdge(Out121), .OutEdge(In107[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID436 e436 ( .InEdge(Out81), .OutEdge(In107[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID437 e437 ( .InEdge(Out93), .OutEdge(In107[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID438 e438 ( .InEdge(Out74), .OutEdge(In107[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID108_INDEGREE5 n108 ( .InEdges(In108), .OutEdge(Out108),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID439 e439 ( .InEdge(Out99), .OutEdge(In108[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID440 e440 ( .InEdge(Out96), .OutEdge(In108[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID441 e441 ( .InEdge(Out103), .OutEdge(In108[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID442 e442 ( .InEdge(Out62), .OutEdge(In108[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID443 e443 ( .InEdge(Out67), .OutEdge(In108[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID109_INDEGREE1 n109 ( .InEdges(In109), .OutEdge(Out109),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID444 e444 ( .InEdge(Out35), .OutEdge(In109[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID110_INDEGREE2 n110 ( .InEdges(In110), .OutEdge(Out110),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID445 e445 ( .InEdge(Out101), .OutEdge(In110[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID446 e446 ( .InEdge(Out99), .OutEdge(In110[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID111_INDEGREE5 n111 ( .InEdges(In111), .OutEdge(Out111),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID447 e447 ( .InEdge(Out31), .OutEdge(In111[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID448 e448 ( .InEdge(Out16), .OutEdge(In111[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID449 e449 ( .InEdge(Out57), .OutEdge(In111[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID450 e450 ( .InEdge(Out38), .OutEdge(In111[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID451 e451 ( .InEdge(Out32), .OutEdge(In111[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID112_INDEGREE7 n112 ( .InEdges(In112), .OutEdge(Out112),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID452 e452 ( .InEdge(Out113), .OutEdge(In112[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID453 e453 ( .InEdge(Out104), .OutEdge(In112[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID454 e454 ( .InEdge(Out95), .OutEdge(In112[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID455 e455 ( .InEdge(Out24), .OutEdge(In112[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID456 e456 ( .InEdge(Out33), .OutEdge(In112[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID457 e457 ( .InEdge(Out126), .OutEdge(In112[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID458 e458 ( .InEdge(Out34), .OutEdge(In112[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID113_INDEGREE7 n113 ( .InEdges(In113), .OutEdge(Out113),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID459 e459 ( .InEdge(Out88), .OutEdge(In113[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID460 e460 ( .InEdge(Out123), .OutEdge(In113[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID461 e461 ( .InEdge(Out29), .OutEdge(In113[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID462 e462 ( .InEdge(Out12), .OutEdge(In113[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID463 e463 ( .InEdge(Out93), .OutEdge(In113[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID464 e464 ( .InEdge(Out52), .OutEdge(In113[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID465 e465 ( .InEdge(Out57), .OutEdge(In113[111:96]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID114_INDEGREE1 n114 ( .InEdges(In114), .OutEdge(Out114),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID466 e466 ( .InEdge(Out72), .OutEdge(In114[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID115_INDEGREE2 n115 ( .InEdges(In115), .OutEdge(Out115),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID467 e467 ( .InEdge(Out108), .OutEdge(In115[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID468 e468 ( .InEdge(Out98), .OutEdge(In115[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID116_INDEGREE6 n116 ( .InEdges(In116), .OutEdge(Out116),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID469 e469 ( .InEdge(Out72), .OutEdge(In116[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID470 e470 ( .InEdge(Out53), .OutEdge(In116[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID471 e471 ( .InEdge(Out45), .OutEdge(In116[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID472 e472 ( .InEdge(Out11), .OutEdge(In116[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID473 e473 ( .InEdge(Out118), .OutEdge(In116[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID474 e474 ( .InEdge(Out50), .OutEdge(In116[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID117_INDEGREE3 n117 ( .InEdges(In117), .OutEdge(Out117),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID475 e475 ( .InEdge(Out80), .OutEdge(In117[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID476 e476 ( .InEdge(Out7), .OutEdge(In117[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID477 e477 ( .InEdge(Out98), .OutEdge(In117[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID118_INDEGREE3 n118 ( .InEdges(In118), .OutEdge(Out118),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID478 e478 ( .InEdge(Out80), .OutEdge(In118[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID479 e479 ( .InEdge(Out42), .OutEdge(In118[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID480 e480 ( .InEdge(Out55), .OutEdge(In118[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID119_INDEGREE6 n119 ( .InEdges(In119), .OutEdge(Out119),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID481 e481 ( .InEdge(Out43), .OutEdge(In119[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID482 e482 ( .InEdge(Out103), .OutEdge(In119[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID483 e483 ( .InEdge(Out61), .OutEdge(In119[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID484 e484 ( .InEdge(Out62), .OutEdge(In119[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID485 e485 ( .InEdge(Out121), .OutEdge(In119[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID486 e486 ( .InEdge(Out8), .OutEdge(In119[95:80]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID120_INDEGREE5 n120 ( .InEdges(In120), .OutEdge(Out120),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID487 e487 ( .InEdge(Out3), .OutEdge(In120[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID488 e488 ( .InEdge(Out88), .OutEdge(In120[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID489 e489 ( .InEdge(Out67), .OutEdge(In120[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID490 e490 ( .InEdge(Out16), .OutEdge(In120[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID491 e491 ( .InEdge(Out84), .OutEdge(In120[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID121_INDEGREE3 n121 ( .InEdges(In121), .OutEdge(Out121),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID492 e492 ( .InEdge(Out55), .OutEdge(In121[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID493 e493 ( .InEdge(Out109), .OutEdge(In121[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID494 e494 ( .InEdge(Out76), .OutEdge(In121[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID122_INDEGREE2 n122 ( .InEdges(In122), .OutEdge(Out122),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID495 e495 ( .InEdge(Out16), .OutEdge(In122[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID496 e496 ( .InEdge(Out105), .OutEdge(In122[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID123_INDEGREE3 n123 ( .InEdges(In123), .OutEdge(Out123),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID497 e497 ( .InEdge(Out44), .OutEdge(In123[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID498 e498 ( .InEdge(Out21), .OutEdge(In123[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID499 e499 ( .InEdge(Out70), .OutEdge(In123[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID124_INDEGREE4 n124 ( .InEdges(In124), .OutEdge(Out124),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID500 e500 ( .InEdge(Out81), .OutEdge(In124[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID501 e501 ( .InEdge(Out15), .OutEdge(In124[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID502 e502 ( .InEdge(Out10), .OutEdge(In124[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID503 e503 ( .InEdge(Out90), .OutEdge(In124[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID125_INDEGREE2 n125 ( .InEdges(In125), .OutEdge(Out125),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID504 e504 ( .InEdge(Out91), .OutEdge(In125[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID505 e505 ( .InEdge(Out49), .OutEdge(In125[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID126_INDEGREE4 n126 ( .InEdges(In126), .OutEdge(Out126),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID506 e506 ( .InEdge(Out25), .OutEdge(In126[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID507 e507 ( .InEdge(Out1), .OutEdge(In126[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID508 e508 ( .InEdge(Out31), .OutEdge(In126[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID509 e509 ( .InEdge(Out114), .OutEdge(In126[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID127_INDEGREE5 n127 ( .InEdges(In127), .OutEdge(Out127),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID510 e510 ( .InEdge(Out1), .OutEdge(In127[15:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID511 e511 ( .InEdge(Out49), .OutEdge(In127[31:16]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID512 e512 ( .InEdge(Out11), .OutEdge(In127[47:32]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID513 e513 ( .InEdge(Out51), .OutEdge(In127[63:48]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID514 e514 ( .InEdge(Out94), .OutEdge(In127[79:64]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
