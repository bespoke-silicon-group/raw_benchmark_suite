
module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n185, n182, \ScanOut[1]1 , 
        n184, \ScanOut[0]1 , n183, \ScanOut[6]1 , \ScanOut[3]1 , n176, 
        \ScanOut[2]1 , n181, n186, n178, n179, n177, n180;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO22 U28 ( .A(ScanIn[1]), .B(n176), .C(\ScanOut[1]1 ), .D(n177), .Z(
        n185) );
    VMW_AO22 U33 ( .A(ScanIn[6]), .B(n176), .C(\ScanOut[6]1 ), .D(n177), .Z(
        n180) );
    VMW_AO22 U34 ( .A(ScanIn[7]), .B(n176), .C(\ScanOut[7] ), .D(n177), .Z(
        n179) );
    VMW_NOR2 U35 ( .A(ScanEnable), .B(Reset), .Z(n177) );
    VMW_AO22 U27 ( .A(ScanIn[0]), .B(n176), .C(\ScanOut[0]1 ), .D(n177), .Z(
        n186) );
    VMW_FD \Out_reg[5]  ( .D(n181), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U29 ( .A(ScanIn[2]), .B(n176), .C(\ScanOut[2]1 ), .D(n177), .Z(
        n184) );
    VMW_FD \Out_reg[7]  ( .D(n179), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n183), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_FD \Out_reg[1]  ( .D(n185), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_AO22 U32 ( .A(ScanIn[5]), .B(n176), .C(\ScanOut[5]1 ), .D(n177), .Z(
        n181) );
    VMW_AO22 U30 ( .A(ScanIn[3]), .B(n176), .C(\ScanOut[3]1 ), .D(n177), .Z(
        n183) );
    VMW_FD \Out_reg[6]  ( .D(n180), .CP(Clk), .Q(\ScanOut[6]1 ) );
    VMW_AO22 U31 ( .A(ScanIn[4]), .B(n176), .C(\ScanOut[4]1 ), .D(n177), .Z(
        n182) );
    VMW_NOR2 U36 ( .A(n178), .B(Reset), .Z(n176) );
    VMW_INV U37 ( .A(ScanEnable), .Z(n178) );
    VMW_FD \Out_reg[2]  ( .D(n184), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_FD \Out_reg[4]  ( .D(n182), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n186), .CP(Clk), .Q(\ScanOut[0]1 ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n1, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n1), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_AND2 U1 ( .A(A[0]), .B(B[0]), .Z(\carry[1] ) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .CO(\carry[2] ) );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .CO(\carry[7] ), .S(
        SUM[6]) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .CO(\carry[3] ), .S(
        SUM[2]) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .CO(\carry[4] ), .S(
        SUM[3]) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .CO(\carry[5] ), .S(
        SUM[4]) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .CO(\carry[6] ), .S(
        SUM[5]) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 ( A, B, CI, 
    SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n3, \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n3) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_FADD U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(
        \carry[7] ) );
    VMW_FADD U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(
        \carry[4] ) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(
        \carry[6] ) );
endmodule


module Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Enable, NorthIn, SouthIn, 
    EastIn, WestIn, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] SouthIn;
input  [7:0] ScanIn;
output [7:0] Out;
output [7:0] ScanOut;
input  [7:0] NorthIn;
input  [7:0] WestIn;
input  [7:0] EastIn;
input  Clk, Reset, RD, WR, ScanEnable, Enable;
    wire \ScanOut[7] , \ScanOut[5]1 , \ScanOut[4]1 , n222, n217, n225, n219, 
        n210, \ScanOut[6]1 , n224, \a184[4] , \n161[4] , \ScanOut[1]1 , n218, 
        \n158[4] , \ScanOut[0]1 , n211, n216, \n158[2] , n223, \n161[2] , 
        \n158[6] , \a184[6] , \n161[6] , \ScanOut[3]1 , \n158[7] , n214, 
        \n161[7] , \a184[7] , n206, n221, \n158[3] , \ScanOut[2]1 , \a184[3] , 
        \n161[3] , \n161[1] , \n158[8] , n226, \a184[8] , \n161[8] , \n158[1] , 
        n213, \a184[5] , n208, \n161[5] , \n158[5] , n209, n212, n215, n207, 
        n220;
    wire UNCONNECTED_1 , UNCONNECTED_2 ;
    assign ScanOut[7] = \ScanOut[7] ;
    assign ScanOut[6] = \ScanOut[6]1 ;
    assign ScanOut[5] = \ScanOut[5]1 ;
    assign ScanOut[4] = \ScanOut[4]1 ;
    assign ScanOut[3] = \ScanOut[3]1 ;
    assign ScanOut[2] = \ScanOut[2]1 ;
    assign ScanOut[1] = \ScanOut[1]1 ;
    assign ScanOut[0] = \ScanOut[0]1 ;
    assign Out[7] = \ScanOut[7] ;
    assign Out[6] = \ScanOut[6]1 ;
    assign Out[5] = \ScanOut[5]1 ;
    assign Out[4] = \ScanOut[4]1 ;
    assign Out[3] = \ScanOut[3]1 ;
    assign Out[2] = \ScanOut[2]1 ;
    assign Out[1] = \ScanOut[1]1 ;
    assign Out[0] = \ScanOut[0]1 ;
    VMW_AO21 U33 ( .A(\ScanOut[0]1 ), .B(n206), .C(n207), .Z(n223) );
    VMW_AO21 U34 ( .A(\ScanOut[1]1 ), .B(n206), .C(n208), .Z(n222) );
    VMW_NOR2 U41 ( .A(n214), .B(Reset), .Z(n213) );
    VMW_AO22 U46 ( .A(ScanIn[3]), .B(n213), .C(\a184[6] ), .D(n215), .Z(n210)
         );
    VMW_AO21 U35 ( .A(\ScanOut[2]1 ), .B(n206), .C(n209), .Z(n221) );
    VMW_AO22 U48 ( .A(ScanIn[1]), .B(n213), .C(\a184[4] ), .D(n215), .Z(n208)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_1 add_98 ( .A({
        \n158[1] , \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , 
        \n158[7] , \n158[8] }), .B(WestIn), .CI(n225), .SUM({\a184[8] , 
        \a184[7] , \a184[6] , \a184[5] , \a184[4] , \a184[3] , UNCONNECTED_1, 
        UNCONNECTED_2}) );
    VMW_PULLDOWN U32 ( .Z(n224) );
    VMW_AO22 U40 ( .A(\ScanOut[7] ), .B(n206), .C(ScanIn[7]), .D(n213), .Z(
        n216) );
    VMW_FD \Out_reg[5]  ( .D(n218), .CP(Clk), .Q(\ScanOut[5]1 ) );
    VMW_AO22 U47 ( .A(ScanIn[2]), .B(n213), .C(\a184[5] ), .D(n215), .Z(n209)
         );
    VMW_AO22 U49 ( .A(ScanIn[0]), .B(n213), .C(\a184[3] ), .D(n215), .Z(n207)
         );
    VMW_FD \Out_reg[1]  ( .D(n222), .CP(Clk), .Q(\ScanOut[1]1 ) );
    VMW_FD \Out_reg[7]  ( .D(n216), .CP(Clk), .Q(\ScanOut[7] ) );
    VMW_FD \Out_reg[3]  ( .D(n220), .CP(Clk), .Q(\ScanOut[3]1 ) );
    VMW_PULLDOWN U30 ( .Z(n225) );
    VMW_AO22 U39 ( .A(\ScanOut[6]1 ), .B(n206), .C(ScanIn[6]), .D(n213), .Z(
        n217) );
    VMW_FD \Out_reg[6]  ( .D(n217), .CP(Clk), .Q(\ScanOut[6]1 ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_0 add_98_2 ( .A(
        NorthIn), .B(SouthIn), .CI(n224), .SUM({\n161[1] , \n161[2] , 
        \n161[3] , \n161[4] , \n161[5] , \n161[6] , \n161[7] , \n161[8] }) );
    VMW_PULLDOWN U31 ( .Z(n226) );
    VMW_AO21 U36 ( .A(\ScanOut[3]1 ), .B(n206), .C(n210), .Z(n220) );
    VMW_AO21 U37 ( .A(\ScanOut[4]1 ), .B(n206), .C(n211), .Z(n219) );
    VMW_NOR3 U42 ( .A(ScanEnable), .B(Reset), .C(Enable), .Z(n206) );
    VMW_AO22 U45 ( .A(ScanIn[4]), .B(n213), .C(\a184[7] ), .D(n215), .Z(n211)
         );
    VMW_FD \Out_reg[2]  ( .D(n221), .CP(Clk), .Q(\ScanOut[2]1 ) );
    VMW_INV U50 ( .A(ScanEnable), .Z(n214) );
    VMW_FD \Out_reg[4]  ( .D(n219), .CP(Clk), .Q(\ScanOut[4]1 ) );
    VMW_FD \Out_reg[0]  ( .D(n223), .CP(Clk), .Q(\ScanOut[0]1 ) );
    VMW_AO21 U38 ( .A(\ScanOut[5]1 ), .B(n206), .C(n212), .Z(n218) );
    VMW_NOR3 U43 ( .A(Reset), .B(ScanEnable), .C(n206), .Z(n215) );
    VMW_AO22 U44 ( .A(ScanIn[5]), .B(n213), .C(\a184[8] ), .D(n215), .Z(n212)
         );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1_DW01_add_8_2 add_98_1 ( .A({
        \n161[1] , \n161[2] , \n161[3] , \n161[4] , \n161[5] , \n161[6] , 
        \n161[7] , \n161[8] }), .B(EastIn), .CI(n226), .SUM({\n158[1] , 
        \n158[2] , \n158[3] , \n158[4] , \n158[5] , \n158[6] , \n158[7] , 
        \n158[8] }) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 ( A, SUM );
input  [6:0] A;
output [6:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[2]), .C(n6), .Z(SUM[2]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n9), .Z(SUM[1]) );
    VMW_INV U6 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO22 U14 ( .A(A[5]), .B(n13), .C(n12), .D(n10), .Z(SUM[5]) );
    VMW_AO21 U7 ( .A(n8), .B(A[4]), .C(n10), .Z(SUM[4]) );
    VMW_AND2 U8 ( .A(n10), .B(n12), .Z(n11) );
    VMW_XOR2 U13 ( .A(A[6]), .B(n11), .Z(SUM[6]) );
    VMW_OR2 U9 ( .A(A[0]), .B(A[1]), .Z(n5) );
    VMW_NOR2 U12 ( .A(n8), .B(A[4]), .Z(n10) );
    VMW_INV U15 ( .A(A[5]), .Z(n12) );
    VMW_INV U17 ( .A(A[3]), .Z(n7) );
    VMW_NOR2 U10 ( .A(n5), .B(A[2]), .Z(n6) );
    VMW_NAND2 U11 ( .A(n6), .B(n7), .Z(n8) );
    VMW_OAI21 U4 ( .A(n6), .B(n7), .C(n8), .Z(SUM[3]) );
    VMW_INV U18 ( .A(n5), .Z(n9) );
    VMW_INV U16 ( .A(n10), .Z(n13) );
endmodule


module Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [7:0] ScanIn;
output [7:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n379, \count[2] , n387, n362, n406, n395, \count[6] , n370, n389, 
        n408, n377, n392, \count[4] , n380, n401, n365, \count[0] , n393, n376, 
        \ScanReg[2] , n409, \count260[3] , n388, n364, n400, n381, 
        \ScanReg[6] , n386, n407, \ScanReg[4] , n363, \count260[5] , n378, 
        \count260[1] , \ScanReg[0] , n371, n394, \count260[0] , \ScanReg[1] , 
        \ScanReg[7] , n405, n384, \ScanReg[5] , \count260[4] , n396, n373, 
        n368, n374, \count260[6] , n383, n391, n410, n402, n366, n390, n398, 
        \count260[2] , \ScanReg[3] , n411, n375, \count[1] , n399, n367, n382, 
        n403, n385, \count[5] , n404, n369, \count[3] , n372, n397;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_PULLDOWN U54 ( .Z(n372) );
    VMW_PULLDOWN U73 ( .Z(n399) );
    VMW_INV U113 ( .A(n370), .Z(ScanEnable) );
    VMW_BUFIZ U134 ( .A(n393), .E(n377), .Z(\arr[3] ) );
    VMW_PULLDOWN U68 ( .Z(n391) );
    VMW_AND2 U96 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_AO22 U108 ( .A(\count[0] ), .B(n366), .C(\ScanReg[0] ), .D(n365), .Z(
        n373) );
    VMW_BUFIZ U141 ( .A(n400), .E(n377), .Z(\arr[18] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n405), .CP(Clk), .Q(\count[6] ) );
    VMW_PULLDOWN U61 ( .Z(n382) );
    VMW_AO22 U84 ( .A(ScanOut[4]), .B(n363), .C(\count260[4] ), .D(n364), .Z(
        n407) );
    VMW_FD \count_reg[2]  ( .D(n409), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_PULLDOWN U66 ( .Z(n389) );
    VMW_XNOR2 U101 ( .A(Addr[0]), .B(ScanId), .Z(n371) );
    VMW_AO22 U106 ( .A(\count[2] ), .B(n366), .C(\ScanReg[2] ), .D(n365), .Z(
        n388) );
    VMW_BUFIZ U121 ( .A(n380), .E(n377), .Z(\arr[14] ) );
    VMW_BUFIZ U126 ( .A(n385), .E(n377), .Z(\arr[31] ) );
    VMW_PULLDOWN U74 ( .Z(n400) );
    VMW_AO22 U83 ( .A(ScanOut[3]), .B(n363), .C(\count260[3] ), .D(n364), .Z(
        n408) );
    VMW_FD \count_reg[0]  ( .D(n411), .CP(Clk), .Q(\count[0] ) );
    VMW_NOR2 U91 ( .A(n367), .B(n368), .Z(n364) );
    VMW_AND2 U98 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_BUFIZ U128 ( .A(n387), .E(n377), .Z(\arr[28] ) );
    VMW_FD \count_reg[4]  ( .D(n407), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U114 ( .A(n372), .E(n377), .Z(\arr[19] ) );
    VMW_BUFIZ U133 ( .A(n392), .E(n377), .Z(\arr[20] ) );
    VMW_AND2 U99 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_PULLDOWN U55 ( .Z(n374) );
    VMW_PULLDOWN U67 ( .Z(n390) );
    VMW_AO22 U82 ( .A(ScanOut[2]), .B(n363), .C(\count260[2] ), .D(n364), .Z(
        n409) );
    VMW_AO22 U107 ( .A(\count[1] ), .B(n366), .C(\ScanReg[1] ), .D(n365), .Z(
        n403) );
    VMW_BUFIZ U120 ( .A(n379), .E(n377), .Z(\arr[27] ) );
    VMW_PULLDOWN U69 ( .Z(n392) );
    VMW_PULLDOWN U75 ( .Z(n401) );
    VMW_BUFIZ U115 ( .A(n373), .E(n377), .Z(\arr[0] ) );
    VMW_BUFIZ U132 ( .A(n391), .E(n377), .Z(\arr[29] ) );
    VMW_OAI21 U90 ( .A(n368), .B(Enable), .C(n369), .Z(n367) );
    VMW_OR4 U109 ( .A(\count[3] ), .B(\count[4] ), .C(\count[5] ), .D(
        \count[6] ), .Z(n362) );
    VMW_BUFIZ U129 ( .A(n388), .E(n377), .Z(\arr[2] ) );
    VMW_PULLDOWN U72 ( .Z(n398) );
    VMW_AND2 U97 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U140 ( .A(n399), .E(n377), .Z(\arr[15] ) );
    VMW_INV U112 ( .A(Reset), .Z(n369) );
    VMW_BUFIZ U135 ( .A(n394), .E(n377), .Z(\arr[24] ) );
    VMW_PULLDOWN U60 ( .Z(n381) );
    VMW_AO22 U85 ( .A(ScanOut[5]), .B(n363), .C(\count260[5] ), .D(n364), .Z(
        n406) );
    VMW_OAI21 U100 ( .A(WR), .B(RD), .C(n371), .Z(n370) );
    VMW_BUFIZ U127 ( .A(n386), .E(n377), .Z(\arr[21] ) );
    VMW_PULLDOWN U56 ( .Z(n375) );
    VMW_PULLDOWN U57 ( .Z(n376) );
    VMW_BUFIZ U137 ( .A(n396), .E(n377), .Z(\arr[7] ) );
    VMW_PULLDOWN U58 ( .Z(n379) );
    VMW_PULLDOWN U59 ( .Z(n380) );
    VMW_PULLDOWN U62 ( .Z(n383) );
    VMW_PULLDOWN U70 ( .Z(n394) );
    VMW_AND2 U79 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U95 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AND2 U110 ( .A(n366), .B(WR), .Z(n368) );
    VMW_BUFIZ U119 ( .A(n378), .E(n377), .Z(\arr[4] ) );
    VMW_BUFIZ U142 ( .A(n401), .E(n377), .Z(\arr[22] ) );
    VMW_AND2 U87 ( .A(\ScanReg[7] ), .B(n365), .Z(n396) );
    VMW_BUFIZ U125 ( .A(n384), .E(n377), .Z(\arr[6] ) );
    VMW_PULLDOWN U65 ( .Z(n387) );
    VMW_AO22 U102 ( .A(\count[6] ), .B(n366), .C(\ScanReg[6] ), .D(n365), .Z(
        n384) );
    VMW_AO22 U105 ( .A(\count[3] ), .B(n366), .C(\ScanReg[3] ), .D(n365), .Z(
        n393) );
    VMW_AO22 U80 ( .A(ScanOut[0]), .B(n363), .C(\count260[0] ), .D(n364), .Z(
        n411) );
    VMW_BUFIZ U122 ( .A(n381), .E(n377), .Z(\arr[25] ) );
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 sub_189 ( .A({
        \count[6] , \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[6] , \count260[5] , \count260[4] , 
        \count260[3] , \count260[2] , \count260[1] , \count260[0] }) );
    VMW_BUFIZ U139 ( .A(n398), .E(n377), .Z(\arr[26] ) );
    VMW_PULLDOWN U77 ( .Z(n404) );
    VMW_XOR2 U89 ( .A(Addr[0]), .B(Id), .Z(n365) );
    VMW_NOR2 U92 ( .A(n367), .B(n365), .Z(n363) );
    VMW_BUFIZ U145 ( .A(n404), .E(n377), .Z(\arr[8] ) );
    VMW_BUFIZ U117 ( .A(n375), .E(n377), .Z(\arr[10] ) );
    VMW_BUFIZ U130 ( .A(n389), .E(n377), .Z(\arr[13] ) );
    VMW_BUFIZ U138 ( .A(n397), .E(n377), .Z(\arr[5] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n406), .CP(Clk), .Q(\count[5] ) );
    VMW_PULLDOWN U64 ( .Z(n386) );
    VMW_AO22 U81 ( .A(ScanOut[1]), .B(n363), .C(\count260[1] ), .D(n364), .Z(
        n410) );
    VMW_AO22 U104 ( .A(\count[4] ), .B(n366), .C(\ScanReg[4] ), .D(n365), .Z(
        n378) );
    VMW_PULLDOWN U76 ( .Z(n402) );
    VMW_BUFIZ U116 ( .A(n374), .E(n377), .Z(\arr[23] ) );
    VMW_BUFIZ U123 ( .A(n382), .E(n377), .Z(\arr[16] ) );
    VMW_AO21 U88 ( .A(RD), .B(ScanEnable), .C(n366), .Z(n377) );
    VMW_AND2 U93 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_BUFIZ U131 ( .A(n390), .E(n377), .Z(\arr[30] ) );
    VMW_FD \count_reg[1]  ( .D(n410), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_BUFIZ U143 ( .A(n402), .E(n377), .Z(\arr[11] ) );
    VMW_BUFIZ U144 ( .A(n403), .E(n377), .Z(\arr[1] ) );
    VMW_FD \count_reg[3]  ( .D(n408), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n395), .E(n377), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_PULLDOWN U63 ( .Z(n385) );
    VMW_PULLDOWN U71 ( .Z(n395) );
    VMW_INV U111 ( .A(n365), .Z(n366) );
    VMW_BUFIZ U124 ( .A(n383), .E(n377), .Z(\arr[12] ) );
    VMW_OR4 U78 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n362), 
        .Z(Enable) );
    VMW_AO22 U86 ( .A(ScanOut[6]), .B(n363), .C(\count260[6] ), .D(n364), .Z(
        n405) );
    VMW_AO22 U103 ( .A(\count[5] ), .B(n366), .C(\ScanReg[5] ), .D(n365), .Z(
        n397) );
    VMW_BUFIZ U118 ( .A(n376), .E(n377), .Z(\arr[9] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nOut0_1[1] , \nOut0_2[2] , \nScanOut4[1] , \nScanOut7[2] , 
        \nScanOut11[1] , \nScanOut12[2] , \nOut2_0[2] , \nScanOut9[4] , 
        \nOut2_3[1] , \nOut1_1[7] , \nOut1_2[4] , \nScanOut14[5] , 
        \nScanOut1[5] , \nScanOut2[6] , \nOut2_0[6] , \nOut2_3[5] , 
        \nOut0_1[5] , \nScanOut9[0] , \nOut0_2[6] , \nScanOut4[5] , 
        \nScanOut7[6] , \nScanOut11[5] , \nScanOut12[6] , \nScanOut1[1] , 
        \nScanOut2[2] , \nOut1_1[3] , \nScanOut14[1] , \nOut1_2[0] , 
        \nScanOut1[3] , \nOut1_1[1] , \nOut1_2[2] , \nScanOut2[0] , 
        \nScanEnable[0] , \nScanOut14[3] , \nOut0_1[7] , \nOut0_2[4] , 
        \nScanOut4[7] , \nScanOut7[4] , \nScanOut11[7] , \nScanOut12[4] , 
        \nOut2_0[4] , \nOut2_3[7] , \nScanOut1[7] , \nScanOut2[4] , 
        \nScanOut9[2] , \nScanOut14[7] , \nOut1_1[5] , \nOut1_2[6] , 
        \nOut2_0[0] , \nScanOut9[6] , \nOut2_3[3] , \nScanOut0[3] , 
        \nOut0_1[3] , \nScanOut4[3] , \nScanOut11[3] , \nScanOut12[0] , 
        \nScanOut7[0] , \nOut0_2[0] , \nScanOut3[0] , \nOut3_1[2] , 
        \nOut3_2[1] , \nScanOut15[3] , \nScanOut16[0] , \nOut1_0[1] , 
        \nOut1_3[2] , \nOut2_1[4] , \nOut2_2[7] , \nScanOut8[2] , 
        \nScanOut5[7] , \nScanOut6[4] , \nScanOut10[7] , \nScanOut13[4] , 
        \nOut1_0[5] , \nOut1_3[6] , \nScanOut0[7] , \nScanOut15[7] , 
        \nScanOut16[4] , \nScanOut3[4] , \nScanOut5[3] , \nScanOut6[0] , 
        \nOut3_1[6] , \nScanOut10[3] , \nOut3_2[5] , \nScanOut13[0] , 
        \nScanOut8[6] , \nOut2_1[0] , \nOut2_2[3] , \nScanOut8[4] , 
        \nOut2_1[2] , \nOut2_2[1] , \nScanOut5[1] , \nScanOut10[1] , 
        \nScanOut13[2] , \nScanOut6[2] , \nScanOut15[5] , \nScanOut16[6] , 
        \nScanOut0[5] , \nScanOut3[6] , \nOut3_1[4] , \nOut3_2[7] , 
        \nOut1_0[7] , \nOut1_3[4] , \nScanOut5[5] , \nScanOut6[6] , 
        \nOut2_1[6] , \nScanOut10[5] , \nScanOut13[6] , \nOut2_2[5] , 
        \nScanOut8[0] , \nOut1_0[3] , \nOut1_3[0] , \nScanOut0[1] , 
        \nOut3_1[0] , \nOut3_2[3] , \nScanOut3[2] , \nScanOut15[1] , 
        \nScanOut16[2] , \nScanOut5[4] , \nScanOut6[7] , \nOut2_1[7] , 
        \nOut2_2[4] , \nScanOut10[4] , \nScanOut13[7] , \nScanOut8[1] , 
        \nOut1_0[2] , \nOut1_3[1] , \nScanOut0[0] , \nScanOut3[3] , 
        \nOut3_1[1] , \nOut3_2[2] , \nScanOut8[5] , \nScanOut15[0] , 
        \nScanOut16[3] , \nOut2_1[3] , \nOut2_2[0] , \nScanOut10[0] , 
        \nScanOut13[3] , \nScanOut5[0] , \nScanOut6[3] , \nScanOut15[4] , 
        \nScanOut16[7] , \nScanOut0[4] , \nOut3_1[5] , \nOut3_2[6] , 
        \nScanOut3[7] , \nOut1_0[6] , \nOut1_3[5] , \nOut1_0[4] , \nOut1_3[7] , 
        \nScanOut15[6] , \nScanOut16[5] , \nScanOut0[6] , \nScanOut3[5] , 
        \nOut3_1[7] , \nOut3_2[4] , \nScanOut10[2] , \nScanOut13[1] , 
        \nScanOut5[2] , \nScanOut6[1] , \nScanOut8[7] , \nScanOut0[2] , 
        \nOut2_1[1] , \nOut2_2[2] , \nScanOut3[1] , \nOut3_1[3] , \nOut3_2[0] , 
        \nOut1_0[0] , \nOut1_3[3] , \nScanOut15[2] , \nScanOut16[1] , 
        \nOut2_1[5] , \nOut2_2[6] , \nScanOut8[3] , \nScanOut5[6] , 
        \nScanOut6[5] , \nScanOut10[6] , \nScanOut13[5] , \nScanOut14[6] , 
        \nScanOut1[6] , \nScanOut2[5] , \nOut1_1[4] , \nOut1_2[7] , 
        \nOut2_0[1] , \nScanOut9[7] , \nOut2_3[2] , \nScanOut11[2] , 
        \nScanOut12[1] , \nScanOut1[2] , \nOut0_1[2] , \nOut0_2[1] , 
        \nScanOut2[1] , \nScanOut4[2] , \nScanOut7[1] , \nOut1_1[0] , 
        \nOut1_2[3] , \nScanOut14[2] , \nOut0_1[6] , \nScanOut4[6] , 
        \nScanOut7[5] , \nOut0_2[5] , \nOut2_0[5] , \nOut2_3[6] , 
        \nScanOut11[6] , \nScanOut12[5] , \nOut2_0[7] , \nScanOut9[3] , 
        \nOut2_3[4] , \nOut0_1[4] , \nOut0_2[7] , \nScanOut4[4] , 
        \nScanOut7[7] , \nScanOut9[1] , \nScanOut1[0] , \nScanOut11[4] , 
        \nScanOut12[7] , \nScanOut2[3] , \nScanOut14[0] , \nEnable[0] , 
        \nOut1_1[2] , \nOut1_2[1] , \nScanOut11[0] , \nScanOut12[3] , 
        \nOut0_1[0] , \nOut0_2[3] , \nScanOut4[0] , \nScanOut7[3] , 
        \nOut2_0[3] , \nScanOut9[5] , \nOut2_3[0] , \nScanOut1[4] , 
        \nScanOut2[7] , \nOut1_1[6] , \nOut1_2[5] , \nScanOut14[4] ;
    Jacobi_Control_WIDTH8_CWIDTH7_IDWIDTH1_SCAN1 U_Jacobi_Control ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanOut({\nScanOut16[7] , 
        \nScanOut16[6] , \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , 
        \nScanOut16[2] , \nScanOut16[1] , \nScanOut16[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b1), .ScanId(1'b0), .Enable(\nEnable[0] ) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut1[7] , \nScanOut1[6] , 
        \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , 
        \nScanOut1[1] , \nScanOut1[0] }), .ScanOut({\nScanOut0[7] , 
        \nScanOut0[6] , \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , 
        \nScanOut0[2] , \nScanOut0[1] , \nScanOut0[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut3[7] , \nScanOut3[6] , 
        \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , 
        \nScanOut3[1] , \nScanOut3[0] }), .ScanOut({\nScanOut2[7] , 
        \nScanOut2[6] , \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , 
        \nScanOut2[2] , \nScanOut2[1] , \nScanOut2[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_2[7] , \nOut0_2[6] , 
        \nOut0_2[5] , \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , 
        \nOut0_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut4[7] , \nScanOut4[6] , 
        \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , 
        \nScanOut4[1] , \nScanOut4[0] }), .ScanOut({\nScanOut3[7] , 
        \nScanOut3[6] , \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , 
        \nScanOut3[2] , \nScanOut3[1] , \nScanOut3[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut5[7] , \nScanOut5[6] , 
        \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , 
        \nScanOut5[1] , \nScanOut5[0] }), .ScanOut({\nScanOut4[7] , 
        \nScanOut4[6] , \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , 
        \nScanOut4[2] , \nScanOut4[1] , \nScanOut4[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_0[7] , \nOut1_0[6] , 
        \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , 
        \nOut1_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut11[7] , \nScanOut11[6] , 
        \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , 
        \nScanOut11[1] , \nScanOut11[0] }), .ScanOut({\nScanOut10[7] , 
        \nScanOut10[6] , \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , 
        \nScanOut10[2] , \nScanOut10[1] , \nScanOut10[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , 
        \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), .SouthIn({\nOut2_3[7] , 
        \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , 
        \nOut2_3[1] , \nOut2_3[0] }), .EastIn({\nOut3_2[7] , \nOut3_2[6] , 
        \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , 
        \nOut3_2[0] }), .WestIn({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , 
        \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), 
        .Out({\nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , 
        \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut6[7] , \nScanOut6[6] , 
        \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , 
        \nScanOut6[1] , \nScanOut6[0] }), .ScanOut({\nScanOut5[7] , 
        \nScanOut5[6] , \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , 
        \nScanOut5[2] , \nScanOut5[1] , \nScanOut5[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_0[7] , \nOut1_0[6] , \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , 
        \nOut1_0[2] , \nOut1_0[1] , \nOut1_0[0] }), .SouthIn({\nOut1_2[7] , 
        \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , 
        \nOut1_2[1] , \nOut1_2[0] }), .EastIn({\nOut2_1[7] , \nOut2_1[6] , 
        \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , 
        \nOut2_1[0] }), .WestIn({\nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , 
        \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), 
        .Out({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , 
        \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut12[7] , \nScanOut12[6] , 
        \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , 
        \nScanOut12[1] , \nScanOut12[0] }), .ScanOut({\nScanOut11[7] , 
        \nScanOut11[6] , \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , 
        \nScanOut11[2] , \nScanOut11[1] , \nScanOut11[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_3[7] , \nOut2_3[6] , 
        \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , 
        \nOut2_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut8[7] , \nScanOut8[6] , 
        \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , 
        \nScanOut8[1] , \nScanOut8[0] }), .ScanOut({\nScanOut7[7] , 
        \nScanOut7[6] , \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , 
        \nScanOut7[2] , \nScanOut7[1] , \nScanOut7[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut1_3[7] , \nOut1_3[6] , 
        \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , 
        \nOut1_3[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut14[7] , \nScanOut14[6] , 
        \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , 
        \nScanOut14[1] , \nScanOut14[0] }), .ScanOut({\nScanOut13[7] , 
        \nScanOut13[6] , \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , 
        \nScanOut13[2] , \nScanOut13[1] , \nScanOut13[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_1[7] , \nOut3_1[6] , 
        \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , 
        \nOut3_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut15[7] , \nScanOut15[6] , 
        \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , 
        \nScanOut15[1] , \nScanOut15[0] }), .ScanOut({\nScanOut14[7] , 
        \nScanOut14[6] , \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , 
        \nScanOut14[2] , \nScanOut14[1] , \nScanOut14[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut3_2[7] , \nOut3_2[6] , 
        \nOut3_2[5] , \nOut3_2[4] , \nOut3_2[3] , \nOut3_2[2] , \nOut3_2[1] , 
        \nOut3_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut2[7] , \nScanOut2[6] , 
        \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , 
        \nScanOut2[1] , \nScanOut2[0] }), .ScanOut({\nScanOut1[7] , 
        \nScanOut1[6] , \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , 
        \nScanOut1[2] , \nScanOut1[1] , \nScanOut1[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut0_1[7] , \nOut0_1[6] , 
        \nOut0_1[5] , \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , 
        \nOut0_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut10[7] , \nScanOut10[6] , 
        \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , 
        \nScanOut10[1] , \nScanOut10[0] }), .ScanOut({\nScanOut9[7] , 
        \nScanOut9[6] , \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , 
        \nScanOut9[2] , \nScanOut9[1] , \nScanOut9[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut2_0[7] , \nOut2_0[6] , \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , 
        \nOut2_0[2] , \nOut2_0[1] , \nOut2_0[0] }), .SouthIn({\nOut2_2[7] , 
        \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , 
        \nOut2_2[1] , \nOut2_2[0] }), .EastIn({\nOut3_1[7] , \nOut3_1[6] , 
        \nOut3_1[5] , \nOut3_1[4] , \nOut3_1[3] , \nOut3_1[2] , \nOut3_1[1] , 
        \nOut3_1[0] }), .WestIn({\nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , 
        \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), 
        .Out({\nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , 
        \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY0_SCAN1 U_Jacobi_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut7[7] , \nScanOut7[6] , 
        \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , 
        \nScanOut7[1] , \nScanOut7[0] }), .ScanOut({\nScanOut6[7] , 
        \nScanOut6[6] , \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , 
        \nScanOut6[2] , \nScanOut6[1] , \nScanOut6[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Enable(\nEnable[0] ), .NorthIn({
        \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , \nOut1_1[3] , 
        \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), .SouthIn({\nOut1_3[7] , 
        \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , 
        \nOut1_3[1] , \nOut1_3[0] }), .EastIn({\nOut2_2[7] , \nOut2_2[6] , 
        \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , 
        \nOut2_2[0] }), .WestIn({\nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , 
        \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), 
        .Out({\nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , 
        \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut9[7] , \nScanOut9[6] , 
        \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , 
        \nScanOut9[1] , \nScanOut9[0] }), .ScanOut({\nScanOut8[7] , 
        \nScanOut8[6] , \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , 
        \nScanOut8[2] , \nScanOut8[1] , \nScanOut8[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0), .Out({\nOut2_0[7] , \nOut2_0[6] , 
        \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , \nOut2_0[2] , \nOut2_0[1] , 
        \nOut2_0[0] }) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut16[7] , \nScanOut16[6] , 
        \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , 
        \nScanOut16[1] , \nScanOut16[0] }), .ScanOut({\nScanOut15[7] , 
        \nScanOut15[6] , \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , 
        \nScanOut15[2] , \nScanOut15[1] , \nScanOut15[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
    Jacobi_Node_WIDTH8_IDWIDTH1_BOUNDARY1_SCAN1 U_Jacobi_Node_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut13[7] , \nScanOut13[6] , 
        \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , 
        \nScanOut13[1] , \nScanOut13[0] }), .ScanOut({\nScanOut12[7] , 
        \nScanOut12[6] , \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , 
        \nScanOut12[2] , \nScanOut12[1] , \nScanOut12[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b0) );
endmodule

