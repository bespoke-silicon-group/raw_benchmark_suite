
module Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, Load, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  Clk, Reset, RD, WR, ScanEnable, Load;
    wire \Out[31] , \Out[5] , n175, n190, n217, n182, n222, n167, n205, n199, 
        n185, n160, n219, n169, n210, n202, n224, n172, n203, n197, \Out[24] , 
        \Out[17] , n161, n184, \Out[30] , n196, n218, \Out[29] , \Out[22] , 
        \Out[20] , \Out[13] , \Out[8] , \Out[1] , n173, n168, n211, \Out[11] , 
        n216, \Out[2] , n183, \Out[18] , \Out[3] , n174, n191, \Out[26] , 
        \Out[15] , n166, n223, \Out[7] , n204, n198, n193, \Out[27] , 
        \Out[14] , n214, n176, \Out[23] , \Out[10] , \Out[6] , n188, n206, 
        n221, \Out[28] , \Out[19] , n164, n181, \Out[0] , n186, \Out[21] , 
        \Out[12] , \Out[9] , n163, n178, n213, n201, \Out[25] , \Out[16] , 
        \Out[4] , n171, n208, n194, n179, n200, n162, n187, n209, n195, n170, 
        n212, n215, n192, n189, n177, n180, n165, n220, n207;
    assign ScanOut[31] = \Out[31] ;
    assign ScanOut[30] = \Out[30] ;
    assign ScanOut[29] = \Out[29] ;
    assign ScanOut[28] = \Out[28] ;
    assign ScanOut[27] = \Out[27] ;
    assign ScanOut[26] = \Out[26] ;
    assign ScanOut[25] = \Out[25] ;
    assign ScanOut[24] = \Out[24] ;
    assign ScanOut[23] = \Out[23] ;
    assign ScanOut[22] = \Out[22] ;
    assign ScanOut[21] = \Out[21] ;
    assign ScanOut[20] = \Out[20] ;
    assign ScanOut[19] = \Out[19] ;
    assign ScanOut[18] = \Out[18] ;
    assign ScanOut[17] = \Out[17] ;
    assign ScanOut[16] = \Out[16] ;
    assign ScanOut[15] = \Out[15] ;
    assign ScanOut[14] = \Out[14] ;
    assign ScanOut[13] = \Out[13] ;
    assign ScanOut[12] = \Out[12] ;
    assign ScanOut[11] = \Out[11] ;
    assign ScanOut[10] = \Out[10] ;
    assign ScanOut[9] = \Out[9] ;
    assign ScanOut[8] = \Out[8] ;
    assign ScanOut[7] = \Out[7] ;
    assign ScanOut[6] = \Out[6] ;
    assign ScanOut[5] = \Out[5] ;
    assign ScanOut[4] = \Out[4] ;
    assign ScanOut[3] = \Out[3] ;
    assign ScanOut[2] = \Out[2] ;
    assign ScanOut[1] = \Out[1] ;
    assign ScanOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AO21 U54 ( .A(\Out[27] ), .B(n160), .C(n188), .Z(n197) );
    VMW_AO21 U73 ( .A(ScanIn[26]), .B(ScanEnable), .C(Reset), .Z(n187) );
    VMW_AO21 U68 ( .A(ScanIn[30]), .B(ScanEnable), .C(Reset), .Z(n191) );
    VMW_AO21 U28 ( .A(\Out[1] ), .B(n160), .C(n162), .Z(n223) );
    VMW_AO21 U33 ( .A(\Out[6] ), .B(n160), .C(n167), .Z(n218) );
    VMW_AO21 U34 ( .A(\Out[7] ), .B(n160), .C(n168), .Z(n217) );
    VMW_AO21 U41 ( .A(\Out[14] ), .B(n160), .C(n175), .Z(n210) );
    VMW_AO21 U46 ( .A(\Out[19] ), .B(n160), .C(n180), .Z(n205) );
    VMW_AO21 U61 ( .A(ScanIn[8]), .B(ScanEnable), .C(Reset), .Z(n169) );
    VMW_AO21 U84 ( .A(ScanIn[16]), .B(ScanEnable), .C(Reset), .Z(n177) );
    VMW_AO21 U66 ( .A(ScanIn[3]), .B(ScanEnable), .C(Reset), .Z(n164) );
    VMW_AO21 U83 ( .A(ScanIn[17]), .B(ScanEnable), .C(Reset), .Z(n178) );
    VMW_AO21 U35 ( .A(\Out[8] ), .B(n160), .C(n169), .Z(n216) );
    VMW_AO21 U48 ( .A(\Out[21] ), .B(n160), .C(n182), .Z(n203) );
    VMW_AO21 U53 ( .A(\Out[26] ), .B(n160), .C(n187), .Z(n198) );
    VMW_AO21 U91 ( .A(ScanIn[0]), .B(ScanEnable), .C(Reset), .Z(n161) );
    VMW_AO21 U74 ( .A(ScanIn[25]), .B(ScanEnable), .C(Reset), .Z(n186) );
    VMW_FD \Out_reg[25]  ( .D(n199), .CP(Clk), .Q(\Out[25] ) );
    VMW_FD \Out_reg[16]  ( .D(n208), .CP(Clk), .Q(\Out[16] ) );
    VMW_AO21 U27 ( .A(\Out[0] ), .B(n160), .C(n161), .Z(n224) );
    VMW_AO21 U40 ( .A(\Out[13] ), .B(n160), .C(n174), .Z(n211) );
    VMW_AO21 U82 ( .A(ScanIn[18]), .B(ScanEnable), .C(Reset), .Z(n179) );
    VMW_FD \Out_reg[5]  ( .D(n219), .CP(Clk), .Q(\Out[5] ) );
    VMW_AO21 U52 ( .A(\Out[25] ), .B(n160), .C(n186), .Z(n199) );
    VMW_AO21 U67 ( .A(ScanIn[31]), .B(ScanEnable), .C(Reset), .Z(n192) );
    VMW_AO21 U75 ( .A(ScanIn[24]), .B(ScanEnable), .C(Reset), .Z(n185) );
    VMW_FD \Out_reg[12]  ( .D(n212), .CP(Clk), .Q(\Out[12] ) );
    VMW_AO21 U90 ( .A(ScanIn[10]), .B(ScanEnable), .C(Reset), .Z(n171) );
    VMW_FD \Out_reg[21]  ( .D(n203), .CP(Clk), .Q(\Out[21] ) );
    VMW_FD \Out_reg[8]  ( .D(n216), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO21 U29 ( .A(\Out[2] ), .B(n160), .C(n163), .Z(n222) );
    VMW_AO21 U47 ( .A(\Out[20] ), .B(n160), .C(n181), .Z(n204) );
    VMW_AO21 U49 ( .A(\Out[22] ), .B(n160), .C(n183), .Z(n202) );
    VMW_FD \Out_reg[31]  ( .D(n193), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n196), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n223), .CP(Clk), .Q(\Out[1] ) );
    VMW_AO21 U55 ( .A(\Out[28] ), .B(n160), .C(n189), .Z(n196) );
    VMW_AO21 U69 ( .A(ScanIn[2]), .B(ScanEnable), .C(Reset), .Z(n163) );
    VMW_FD \Out_reg[19]  ( .D(n205), .CP(Clk), .Q(\Out[19] ) );
    VMW_AO21 U72 ( .A(ScanIn[27]), .B(ScanEnable), .C(Reset), .Z(n188) );
    VMW_FD \Out_reg[3]  ( .D(n221), .CP(Clk), .Q(\Out[3] ) );
    VMW_FD \Out_reg[23]  ( .D(n201), .CP(Clk), .Q(\Out[23] ) );
    VMW_FD \Out_reg[10]  ( .D(n214), .CP(Clk), .Q(\Out[10] ) );
    VMW_AO21 U60 ( .A(ScanIn[9]), .B(ScanEnable), .C(Reset), .Z(n170) );
    VMW_FD \Out_reg[7]  ( .D(n217), .CP(Clk), .Q(\Out[7] ) );
    VMW_AO21 U32 ( .A(\Out[5] ), .B(n160), .C(n166), .Z(n219) );
    VMW_AO21 U85 ( .A(ScanIn[15]), .B(ScanEnable), .C(Reset), .Z(n176) );
    VMW_FD \Out_reg[27]  ( .D(n197), .CP(Clk), .Q(\Out[27] ) );
    VMW_FD \Out_reg[14]  ( .D(n210), .CP(Clk), .Q(\Out[14] ) );
    VMW_AO21 U30 ( .A(\Out[3] ), .B(n160), .C(n164), .Z(n221) );
    VMW_AO21 U39 ( .A(\Out[12] ), .B(n160), .C(n173), .Z(n212) );
    VMW_AO21 U57 ( .A(\Out[30] ), .B(n160), .C(n191), .Z(n194) );
    VMW_FD \Out_reg[6]  ( .D(n218), .CP(Clk), .Q(\Out[6] ) );
    VMW_AO21 U70 ( .A(ScanIn[29]), .B(ScanEnable), .C(Reset), .Z(n190) );
    VMW_AO21 U79 ( .A(ScanIn[20]), .B(ScanEnable), .C(Reset), .Z(n181) );
    VMW_FD \Out_reg[26]  ( .D(n198), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n209), .CP(Clk), .Q(\Out[15] ) );
    VMW_FD \Out_reg[18]  ( .D(n206), .CP(Clk), .Q(\Out[18] ) );
    VMW_AO21 U31 ( .A(\Out[4] ), .B(n160), .C(n165), .Z(n220) );
    VMW_AO21 U36 ( .A(\Out[9] ), .B(n160), .C(n170), .Z(n215) );
    VMW_AO21 U37 ( .A(\Out[10] ), .B(n160), .C(n171), .Z(n214) );
    VMW_AO21 U42 ( .A(\Out[15] ), .B(n160), .C(n176), .Z(n209) );
    VMW_AO21 U45 ( .A(\Out[18] ), .B(n160), .C(n179), .Z(n206) );
    VMW_AO21 U87 ( .A(ScanIn[13]), .B(ScanEnable), .C(Reset), .Z(n174) );
    VMW_FD \Out_reg[2]  ( .D(n222), .CP(Clk), .Q(\Out[2] ) );
    VMW_FD \Out_reg[11]  ( .D(n213), .CP(Clk), .Q(\Out[11] ) );
    VMW_AO21 U62 ( .A(ScanIn[7]), .B(ScanEnable), .C(Reset), .Z(n168) );
    VMW_FD \Out_reg[22]  ( .D(n202), .CP(Clk), .Q(\Out[22] ) );
    VMW_AO21 U65 ( .A(ScanIn[4]), .B(ScanEnable), .C(Reset), .Z(n165) );
    VMW_FD \Out_reg[20]  ( .D(n204), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n211), .CP(Clk), .Q(\Out[13] ) );
    VMW_AO21 U80 ( .A(ScanIn[1]), .B(ScanEnable), .C(Reset), .Z(n162) );
    VMW_FD \Out_reg[9]  ( .D(n215), .CP(Clk), .Q(\Out[9] ) );
    VMW_AO21 U50 ( .A(\Out[23] ), .B(n160), .C(n184), .Z(n201) );
    VMW_NOR2 U59 ( .A(ScanEnable), .B(Load), .Z(n160) );
    VMW_FD \Out_reg[30]  ( .D(n194), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n224), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n195), .CP(Clk), .Q(\Out[29] ) );
    VMW_AO21 U77 ( .A(ScanIn[22]), .B(ScanEnable), .C(Reset), .Z(n183) );
    VMW_AO21 U89 ( .A(ScanIn[11]), .B(ScanEnable), .C(Reset), .Z(n172) );
    VMW_FD \Out_reg[24]  ( .D(n200), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n207), .CP(Clk), .Q(\Out[17] ) );
    VMW_FD \Out_reg[4]  ( .D(n220), .CP(Clk), .Q(\Out[4] ) );
    VMW_AO21 U58 ( .A(\Out[31] ), .B(n160), .C(n192), .Z(n193) );
    VMW_AO21 U38 ( .A(\Out[11] ), .B(n160), .C(n172), .Z(n213) );
    VMW_AO21 U43 ( .A(\Out[16] ), .B(n160), .C(n177), .Z(n208) );
    VMW_AO21 U64 ( .A(ScanIn[5]), .B(ScanEnable), .C(Reset), .Z(n166) );
    VMW_AO21 U81 ( .A(ScanIn[19]), .B(ScanEnable), .C(Reset), .Z(n180) );
    VMW_AO21 U51 ( .A(\Out[24] ), .B(n160), .C(n185), .Z(n200) );
    VMW_AO21 U76 ( .A(ScanIn[23]), .B(ScanEnable), .C(Reset), .Z(n184) );
    VMW_AO21 U88 ( .A(ScanIn[12]), .B(ScanEnable), .C(Reset), .Z(n173) );
    VMW_AO21 U44 ( .A(\Out[17] ), .B(n160), .C(n178), .Z(n207) );
    VMW_AO21 U56 ( .A(\Out[29] ), .B(n160), .C(n190), .Z(n195) );
    VMW_AO21 U71 ( .A(ScanIn[28]), .B(ScanEnable), .C(Reset), .Z(n189) );
    VMW_AO21 U63 ( .A(ScanIn[6]), .B(ScanEnable), .C(Reset), .Z(n167) );
    VMW_AO21 U86 ( .A(ScanIn[14]), .B(ScanEnable), .C(Reset), .Z(n175) );
    VMW_AO21 U78 ( .A(ScanIn[21]), .B(ScanEnable), .C(Reset), .Z(n182) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n15, n55, n72, n97, n20, n69, n100, n112, n32, n29, n85, n47, n60, 
        n109, n40, n67, n82, n99, n27, n35, n49, n115, n107, n90, n52, n75, 
        n98, n114, n34, n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, 
        n101, n21, n46, n54, n96, n73, n61, n108, n28, n84, n33, n38, n56, n71, 
        n113, n94, n23, n103, n16, n111, n31, n36, n44, n63, n86, n43, n64, 
        n81, n58, n104, n18, n24, n88, n37, n51, n93, n59, n76, n80, n42, n65, 
        n19, n50, n77, n89, n92, n25, n102, n105, n22, n39, n95, n45, n57, n62, 
        n87, n17, n30, n79, n110;
    VMW_AO21 U3 ( .A(n15), .B(A[31]), .C(n16), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n96), .Z(n99) );
    VMW_INV U73 ( .A(B[27]), .Z(n105) );
    VMW_INV U96 ( .A(n115), .Z(n16) );
    VMW_INV U68 ( .A(A[30]), .Z(n110) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n80), .C(n74), .D(n68), .Z(n79) );
    VMW_NAND2 U46 ( .A(n86), .B(A[21]), .Z(n87) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n112), .C(n107), .D(n102), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(A[6]), .Z(n30) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(B[13]), .Z(n58) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n90), .B(B[24]), .Z(n89) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n98), .C(n94), .D(n89), .Z(n97) );
    VMW_INV U91 ( .A(A[28]), .Z(n103) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(A[26]), .Z(n96) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n77), .B(B[20]), .Z(n76) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n96), .B(B[26]), .Z(n95) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n98) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n92), .C(n88), .D(n83), .Z(n91) );
    VMW_INV U69 ( .A(B[17]), .Z(n72) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n84), .C(n87), .D(n85), .Z(n88) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n101), .C(n99), .D(n97), .Z(n100) );
    VMW_INV U72 ( .A(A[27]), .Z(n108) );
    VMW_INV U97 ( .A(A[16]), .Z(n62) );
    VMW_NAND2 U60 ( .A(n110), .B(B[30]), .Z(n109) );
    VMW_INV U100 ( .A(B[23]), .Z(n92) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n90) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n75), .C(n73), .D(n71), .Z(n74) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n105), .C(n100), .D(n95), .Z(n104) );
    VMW_INV U70 ( .A(A[17]), .Z(n75) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n86) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n80), .B(A[19]), .Z(n81) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n86), .C(n82), .D(n76), .Z(n85) );
    VMW_NAND2 U62 ( .A(n112), .B(A[29]), .Z(n113) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U102 ( .A(B[2]), .Z(n21) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n72), .C(n66), .D(n61), .Z(n71) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n108), .C(n106), .D(n104), .Z(n107) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n92), .B(A[23]), .Z(n93) );
    VMW_INV U77 ( .A(A[20]), .Z(n77) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n103), .Z(n106) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n112) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n77), .C(n81), .D(n79), .Z(n82) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n15), .C(n114), .D(n109), .Z(n115) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n90), .C(n93), .D(n91), .Z(n94) );
    VMW_INV U76 ( .A(A[25]), .Z(n101) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n73) );
    VMW_NAND2 U44 ( .A(n84), .B(B[22]), .Z(n83) );
    VMW_NAND2 U56 ( .A(n103), .B(B[28]), .Z(n102) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n84) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n110), .C(n113), .D(n111), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n80) );
endmodule


module Merge_Node_DWIDTH32_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, n182, 
        n129, n185, n147, n160, n120, n132, n202, n169, n210, n155, n172, n197, 
        n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, n211, 
        n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, n193, 
        n198, n151, n176, n124, n188, n206, n136, n143, n158, n144, n163, n164, 
        n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, n138, 
        n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, n170, 
        n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, n165, 
        n159, n137, n207;
    VMW_OAI21 U3 ( .A(A[31]), .B(n116), .C(n117), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n119), .C(B[0]), .Z(n120) );
    VMW_AO22 U6 ( .A(A[2]), .B(n122), .C(n120), .D(A[0]), .Z(n121) );
    VMW_OR2 U14 ( .A(B[6]), .B(n131), .Z(n134) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n147), .C(n142), .D(n137), .Z(n146) );
    VMW_OR2 U54 ( .A(B[26]), .B(n195), .Z(n198) );
    VMW_INV U73 ( .A(B[27]), .Z(n204) );
    VMW_INV U96 ( .A(A[16]), .Z(n163) );
    VMW_INV U68 ( .A(A[30]), .Z(n212) );
    VMW_NAND2 U28 ( .A(n157), .B(B[14]), .Z(n156) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n165), .C(n161), .D(n156), .Z(n164) );
    VMW_OAI22 U7 ( .A(n118), .B(n121), .C(A[2]), .D(n122), .Z(n123) );
    VMW_NAND2 U8 ( .A(n125), .B(B[4]), .Z(n124) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n133), .C(n129), .D(n124), .Z(n132) );
    VMW_OR2 U34 ( .A(B[16]), .B(n163), .Z(n166) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n179), .C(n174), .D(n169), .Z(n178) );
    VMW_NAND2 U46 ( .A(n185), .B(A[21]), .Z(n186) );
    VMW_NAND2 U61 ( .A(n209), .B(A[29]), .Z(n210) );
    VMW_INV U84 ( .A(A[4]), .Z(n125) );
    VMW_INV U101 ( .A(B[2]), .Z(n122) );
    VMW_INV U66 ( .A(B[7]), .Z(n140) );
    VMW_INV U83 ( .A(B[15]), .Z(n165) );
    VMW_INV U98 ( .A(A[26]), .Z(n195) );
    VMW_NAND2 U26 ( .A(n153), .B(A[11]), .Z(n154) );
    VMW_NAND2 U48 ( .A(n189), .B(B[24]), .Z(n188) );
    VMW_AO21 U9 ( .A(B[3]), .B(n127), .C(n123), .Z(n126) );
    VMW_NAND2 U12 ( .A(n131), .B(B[6]), .Z(n130) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n168), .C(n166), .D(n164), .Z(n167) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n197), .C(n193), .D(n188), .Z(n196) );
    VMW_INV U91 ( .A(A[28]), .Z(n202) );
    VMW_INV U74 ( .A(A[3]), .Z(n127) );
    VMW_INV U99 ( .A(B[23]), .Z(n191) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n151), .C(n154), .D(n152), .Z(n155) );
    VMW_NAND2 U40 ( .A(n177), .B(B[20]), .Z(n176) );
    VMW_INV U82 ( .A(A[15]), .Z(n168) );
    VMW_NAND2 U52 ( .A(n195), .B(B[26]), .Z(n194) );
    VMW_INV U67 ( .A(A[7]), .Z(n143) );
    VMW_INV U75 ( .A(B[25]), .Z(n197) );
    VMW_INV U90 ( .A(B[11]), .Z(n153) );
    VMW_NAND2 U20 ( .A(n145), .B(B[10]), .Z(n144) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n191), .C(n187), .D(n182), .Z(n190) );
    VMW_INV U69 ( .A(B[17]), .Z(n172) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n159), .C(n155), .D(n150), .Z(n158) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n183), .C(n186), .D(n184), .Z(n187) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n200), .C(n198), .D(n196), .Z(n199) );
    VMW_INV U72 ( .A(A[27]), .Z(n207) );
    VMW_INV U97 ( .A(B[13]), .Z(n159) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n209), .C(n206), .D(n201), .Z(n208) );
    VMW_INV U100 ( .A(A[6]), .Z(n131) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n136), .C(n134), .D(n132), .Z(n135) );
    VMW_INV U85 ( .A(A[24]), .Z(n189) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n140), .C(n135), .D(n130), .Z(n139) );
    VMW_NAND2 U22 ( .A(n147), .B(A[9]), .Z(n148) );
    VMW_NAND2 U32 ( .A(n163), .B(B[16]), .Z(n162) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n175), .C(n173), .D(n171), .Z(n174) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n204), .C(n199), .D(n194), .Z(n203) );
    VMW_INV U70 ( .A(A[17]), .Z(n175) );
    VMW_INV U95 ( .A(B[31]), .Z(n116) );
    VMW_NAND2 U30 ( .A(n159), .B(A[13]), .Z(n160) );
    VMW_INV U79 ( .A(A[10]), .Z(n145) );
    VMW_INV U87 ( .A(B[21]), .Z(n185) );
    VMW_OR2 U10 ( .A(B[4]), .B(n125), .Z(n128) );
    VMW_NAND2 U42 ( .A(n179), .B(A[19]), .Z(n180) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n185), .C(n181), .D(n176), .Z(n184) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n212), .C(n210), .D(n208), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n151) );
    VMW_INV U80 ( .A(B[9]), .Z(n147) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n127), .C(n128), .D(n126), .Z(n129) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n143), .C(n141), .D(n139), .Z(n142) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n153), .C(n149), .D(n144), .Z(n152) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n172), .C(n167), .D(n162), .Z(n171) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n207), .C(n205), .D(n203), .Z(n206) );
    VMW_INV U89 ( .A(A[14]), .Z(n157) );
    VMW_NAND2 U50 ( .A(n191), .B(A[23]), .Z(n192) );
    VMW_INV U77 ( .A(A[20]), .Z(n177) );
    VMW_INV U92 ( .A(A[5]), .Z(n136) );
    VMW_OR2 U58 ( .A(B[28]), .B(n202), .Z(n205) );
    VMW_NAND2 U36 ( .A(n170), .B(B[18]), .Z(n169) );
    VMW_INV U81 ( .A(B[29]), .Z(n209) );
    VMW_NOR2 U4 ( .A(n119), .B(B[1]), .Z(n118) );
    VMW_OR2 U18 ( .A(B[8]), .B(n138), .Z(n141) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n177), .C(n180), .D(n178), .Z(n181) );
    VMW_AO22 U64 ( .A(n211), .B(n213), .C(A[31]), .D(n116), .Z(n117) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n189), .C(n192), .D(n190), .Z(n193) );
    VMW_INV U76 ( .A(A[25]), .Z(n200) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n145), .C(n148), .D(n146), .Z(n149) );
    VMW_NAND2 U24 ( .A(n151), .B(B[12]), .Z(n150) );
    VMW_INV U88 ( .A(A[18]), .Z(n170) );
    VMW_INV U93 ( .A(B[5]), .Z(n133) );
    VMW_OR2 U38 ( .A(B[18]), .B(n170), .Z(n173) );
    VMW_NAND2 U44 ( .A(n183), .B(B[22]), .Z(n182) );
    VMW_NAND2 U56 ( .A(n202), .B(B[28]), .Z(n201) );
    VMW_INV U94 ( .A(A[1]), .Z(n119) );
    VMW_INV U71 ( .A(A[22]), .Z(n183) );
    VMW_NAND2 U63 ( .A(n212), .B(B[30]), .Z(n213) );
    VMW_INV U86 ( .A(A[8]), .Z(n138) );
    VMW_NAND2 U16 ( .A(n138), .B(B[8]), .Z(n137) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n157), .C(n160), .D(n158), .Z(n161) );
    VMW_INV U78 ( .A(B[19]), .Z(n179) );
endmodule


module Merge_Node_DWIDTH32 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, Load, 
    Out, In1, In2, Read1, Read2 );
input  [14:0] Addr;
input  [31:0] DataIn;
input  [31:0] DataOut;
input  [31:0] In1;
output [31:0] Out;
input  [31:0] In2;
input  Clk, Reset, RD, WR, Load;
output Read1, Read2;
    wire n337, n339, n217, n287, n330, n317, n245, n262, n279, n230, n222, 
        n219, n257, n270, n239, n295, n305, n322, n292, n325, n302, n250, n277, 
        n225, n289, n319, n237, n259, n265, n242, n336, n218, n224, n280, n310, 
        n251, n276, n288, n318, n293, n303, n324, n338, n216, n231, n236, n243, 
        n264, n281, n311, n258, n278, n223, n238, n244, n263, n286, n316, n294, 
        n331, n304, n323, n256, n271, n70, n215, n214, n228, n284, n333, n314, 
        n246, n261, n221, n233, n328, n226, n248, n254, n268, n78, n273, n253, 
        n291, n296, n321, n301, n306, n326, n274, n227, n234, n241, n298, n308, 
        n266, n283, n313, n334, n249, n252, n275, n282, n290, n300, n327, n312, 
        n335, n235, n240, n267, n299, n309, n232, n329, n247, n260, n332, n229, 
        n285, n315, n297, n307, n320, n255, n272, n220, n269;
    VMW_PULLDOWN U36 ( .Z(n337) );
    VMW_PULLUP U37 ( .Z(n336) );
    VMW_PULLUP U39 ( .Z(n338) );
    VMW_OAI21 U40 ( .A(n70), .B(n215), .C(Load), .Z(n214) );
    VMW_AO21 U41 ( .A(n215), .B(n217), .C(Reset), .Z(n216) );
    VMW_AOI211 U46 ( .A(n219), .B(In2[5]), .C(n228), .D(n216), .Z(n227) );
    VMW_AOI211 U54 ( .A(n219), .B(In2[27]), .C(n244), .D(n216), .Z(n243) );
    VMW_AOI211 U73 ( .A(n219), .B(In2[0]), .C(n282), .D(n216), .Z(n281) );
    VMW_AO22 U113 ( .A(Out[22]), .B(n293), .C(n294), .D(In1[22]), .Z(n254) );
    VMW_INV U134 ( .A(n225), .Z(n329) );
    VMW_AOI211 U61 ( .A(n219), .B(In2[20]), .C(n258), .D(n216), .Z(n257) );
    VMW_AOI211 U68 ( .A(n219), .B(In2[14]), .C(n272), .D(n216), .Z(n271) );
    VMW_AO22 U96 ( .A(Out[9]), .B(n293), .C(n294), .D(In1[9]), .Z(n220) );
    VMW_AO22 U108 ( .A(Out[27]), .B(n293), .C(n294), .D(In1[27]), .Z(n244) );
    VMW_INV U141 ( .A(n239), .Z(n306) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_1 r140 ( .A(In1), .B(In2), .LEQ(n338), 
        .TC(n339), .GE_GT(n70) );
    VMW_AND4 U84 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(n285
        ) );
    VMW_INV U148 ( .A(n253), .Z(n313) );
    VMW_INV U153 ( .A(n263), .Z(n317) );
    VMW_AO22 U101 ( .A(Out[4]), .B(n293), .C(n294), .D(In1[4]), .Z(n230) );
    VMW_AO22 U126 ( .A(Out[10]), .B(n293), .C(n294), .D(In1[10]), .Z(n280) );
    VMW_AOI211 U48 ( .A(n219), .B(In2[3]), .C(n232), .D(n216), .Z(n231) );
    VMW_AOI211 U66 ( .A(n219), .B(In2[16]), .C(n268), .D(n216), .Z(n267) );
    VMW_AO22 U106 ( .A(Out[29]), .B(n293), .C(n294), .D(In1[29]), .Z(n240) );
    VMW_AO22 U121 ( .A(Out[15]), .B(n293), .C(n294), .D(In1[15]), .Z(n270) );
    VMW_AND4 U83 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(n286
        ) );
    VMW_AO22 U98 ( .A(Out[7]), .B(n293), .C(n294), .D(In1[7]), .Z(n224) );
    VMW_OAI21 U128 ( .A(n78), .B(n217), .C(Load), .Z(n303) );
    VMW_INV U154 ( .A(n265), .Z(n318) );
    VMW_AOI211 U53 ( .A(n219), .B(In2[28]), .C(n242), .D(n216), .Z(n241) );
    VMW_AND4 U91 ( .A(n302), .B(n301), .C(n300), .D(n299), .Z(n292) );
    VMW_INV U146 ( .A(n249), .Z(n311) );
    VMW_INV U161 ( .A(n279), .Z(n325) );
    VMW_AND5 U74 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(n287), .Z(n217)
         );
    VMW_AO22 U114 ( .A(Out[21]), .B(n293), .C(n294), .D(In1[21]), .Z(n256) );
    VMW_INV U133 ( .A(n223), .Z(n328) );
    VMW_AND4 U82 ( .A(n298), .B(n297), .C(n296), .D(n295), .Z(n287) );
    VMW_AO22 U99 ( .A(Out[6]), .B(n293), .C(n294), .D(In1[6]), .Z(n226) );
    VMW_INV U155 ( .A(n267), .Z(n319) );
    VMW_FD \Out_reg[16]  ( .D(n319), .CP(Clk), .Q(Out[16]) );
    VMW_FD \Out_reg[25]  ( .D(n310), .CP(Clk), .Q(Out[25]) );
    VMW_FD \Out_reg[5]  ( .D(n330), .CP(Clk), .Q(Out[5]) );
    VMW_AOI211 U47 ( .A(n219), .B(In2[4]), .C(n230), .D(n216), .Z(n229) );
    VMW_AOI211 U49 ( .A(n219), .B(In2[31]), .C(n234), .D(n216), .Z(n233) );
    VMW_AOI211 U52 ( .A(n219), .B(In2[29]), .C(n240), .D(n216), .Z(n239) );
    VMW_AOI211 U67 ( .A(n219), .B(In2[15]), .C(n270), .D(n216), .Z(n269) );
    VMW_AO22 U107 ( .A(Out[28]), .B(n293), .C(n294), .D(In1[28]), .Z(n242) );
    VMW_AO22 U120 ( .A(Out[16]), .B(n293), .C(n294), .D(In1[16]), .Z(n268) );
    VMW_AND5 U75 ( .A(n288), .B(n289), .C(n290), .D(n291), .E(n292), .Z(n215)
         );
    VMW_AO22 U115 ( .A(Out[20]), .B(n293), .C(n294), .D(In1[20]), .Z(n258) );
    VMW_INV U132 ( .A(n221), .Z(n327) );
    VMW_FD \Out_reg[12]  ( .D(n323), .CP(Clk), .Q(Out[12]) );
    VMW_AND4 U90 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(n302
        ) );
    VMW_FD \Out_reg[21]  ( .D(n314), .CP(Clk), .Q(Out[21]) );
    VMW_INV U129 ( .A(n214), .Z(Read1) );
    VMW_INV U147 ( .A(n251), .Z(n312) );
    VMW_FD \Out_reg[8]  ( .D(n327), .CP(Clk), .Q(Out[8]) );
    VMW_INV U160 ( .A(n277), .Z(n324) );
    VMW_FD \Out_reg[31]  ( .D(n304), .CP(Clk), .Q(Out[31]) );
    VMW_FD \Out_reg[28]  ( .D(n307), .CP(Clk), .Q(Out[28]) );
    VMW_FD \Out_reg[1]  ( .D(n334), .CP(Clk), .Q(Out[1]) );
    VMW_AOI211 U55 ( .A(n219), .B(In2[26]), .C(n246), .D(n216), .Z(n245) );
    VMW_AOI211 U69 ( .A(n219), .B(In2[13]), .C(n274), .D(n216), .Z(n273) );
    VMW_AO22 U109 ( .A(Out[26]), .B(n293), .C(n294), .D(In1[26]), .Z(n246) );
    VMW_FD \Out_reg[19]  ( .D(n316), .CP(Clk), .Q(Out[19]) );
    VMW_AOI211 U72 ( .A(n219), .B(In2[10]), .C(n280), .D(n216), .Z(n279) );
    VMW_AO22 U97 ( .A(Out[8]), .B(n293), .C(n294), .D(In1[8]), .Z(n222) );
    VMW_INV U140 ( .A(n237), .Z(n333) );
    VMW_FD \Out_reg[3]  ( .D(n332), .CP(Clk), .Q(Out[3]) );
    VMW_AO22 U112 ( .A(Out[23]), .B(n293), .C(n294), .D(In1[23]), .Z(n252) );
    VMW_INV U135 ( .A(n227), .Z(n330) );
    VMW_FD \Out_reg[10]  ( .D(n325), .CP(Clk), .Q(Out[10]) );
    VMW_FD \Out_reg[23]  ( .D(n312), .CP(Clk), .Q(Out[23]) );
    VMW_AOI211 U60 ( .A(n219), .B(In2[21]), .C(n256), .D(n216), .Z(n255) );
    VMW_FD \Out_reg[7]  ( .D(n328), .CP(Clk), .Q(Out[7]) );
    VMW_AO22 U100 ( .A(Out[5]), .B(n293), .C(n294), .D(In1[5]), .Z(n228) );
    VMW_AO22 U127 ( .A(Out[0]), .B(n293), .C(n294), .D(In1[0]), .Z(n282) );
    VMW_AOI211 U57 ( .A(n219), .B(In2[24]), .C(n250), .D(n216), .Z(n249) );
    VMW_AND4 U85 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(n284
        ) );
    VMW_INV U149 ( .A(n255), .Z(n314) );
    VMW_INV U137 ( .A(n231), .Z(n332) );
    VMW_INV U152 ( .A(n261), .Z(n316) );
    VMW_FD \Out_reg[27]  ( .D(n308), .CP(Clk), .Q(Out[27]) );
    VMW_FD \Out_reg[14]  ( .D(n321), .CP(Clk), .Q(Out[14]) );
    VMW_FD \Out_reg[6]  ( .D(n329), .CP(Clk), .Q(Out[6]) );
    VMW_AOI211 U70 ( .A(n219), .B(In2[12]), .C(n276), .D(n216), .Z(n275) );
    VMW_AO22 U110 ( .A(Out[25]), .B(n293), .C(n294), .D(In1[25]), .Z(n248) );
    VMW_INV U159 ( .A(n275), .Z(n323) );
    VMW_AOI211 U42 ( .A(n219), .B(In2[9]), .C(n220), .D(n216), .Z(n218) );
    VMW_AOI211 U45 ( .A(n219), .B(In2[6]), .C(n226), .D(n216), .Z(n225) );
    VMW_AND4 U79 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n296) );
    VMW_AND4 U95 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(n288
        ) );
    VMW_AO22 U119 ( .A(Out[17]), .B(n293), .C(n294), .D(In1[17]), .Z(n266) );
    VMW_INV U142 ( .A(n241), .Z(n307) );
    VMW_FD \Out_reg[26]  ( .D(n309), .CP(Clk), .Q(Out[26]) );
    VMW_FD \Out_reg[15]  ( .D(n320), .CP(Clk), .Q(Out[15]) );
    VMW_FD \Out_reg[18]  ( .D(n317), .CP(Clk), .Q(Out[18]) );
    VMW_AND4 U87 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n299) );
    VMW_INV U150 ( .A(n257), .Z(n315) );
    VMW_FD \Out_reg[2]  ( .D(n333), .CP(Clk), .Q(Out[2]) );
    VMW_AO22 U125 ( .A(Out[11]), .B(n293), .C(n294), .D(In1[11]), .Z(n278) );
    VMW_FD \Out_reg[11]  ( .D(n324), .CP(Clk), .Q(Out[11]) );
    VMW_AOI211 U62 ( .A(n219), .B(In2[1]), .C(n260), .D(n216), .Z(n259) );
    VMW_FD \Out_reg[22]  ( .D(n313), .CP(Clk), .Q(Out[22]) );
    VMW_AOI211 U65 ( .A(n219), .B(In2[17]), .C(n266), .D(n216), .Z(n265) );
    VMW_AO22 U102 ( .A(Out[3]), .B(n293), .C(n294), .D(In1[3]), .Z(n232) );
    VMW_AO22 U105 ( .A(Out[2]), .B(n293), .C(n294), .D(In1[2]), .Z(n238) );
    VMW_FD \Out_reg[20]  ( .D(n315), .CP(Clk), .Q(Out[20]) );
    VMW_FD \Out_reg[13]  ( .D(n322), .CP(Clk), .Q(Out[13]) );
    VMW_AND4 U80 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n297)
         );
    VMW_AO22 U122 ( .A(Out[14]), .B(n293), .C(n294), .D(In1[14]), .Z(n272) );
    VMW_INV U157 ( .A(n271), .Z(n321) );
    VMW_FD \Out_reg[9]  ( .D(n326), .CP(Clk), .Q(Out[9]) );
    VMW_AOI211 U50 ( .A(n219), .B(In2[30]), .C(n236), .D(n216), .Z(n235) );
    VMW_AOI211 U59 ( .A(n219), .B(In2[22]), .C(n254), .D(n216), .Z(n253) );
    VMW_INV U139 ( .A(n235), .Z(n305) );
    VMW_FD \Out_reg[30]  ( .D(n305), .CP(Clk), .Q(Out[30]) );
    VMW_FD \Out_reg[0]  ( .D(n335), .CP(Clk), .Q(Out[0]) );
    VMW_FD \Out_reg[29]  ( .D(n306), .CP(Clk), .Q(Out[29]) );
    VMW_AND2 U77 ( .A(n70), .B(Load), .Z(n294) );
    VMW_AND4 U89 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n301)
         );
    VMW_AND4 U92 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(n291
        ) );
    VMW_INV U145 ( .A(n247), .Z(n310) );
    VMW_INV U162 ( .A(n281), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n311), .CP(Clk), .Q(Out[24]) );
    VMW_FD \Out_reg[17]  ( .D(n318), .CP(Clk), .Q(Out[17]) );
    VMW_AO22 U117 ( .A(Out[19]), .B(n293), .C(n294), .D(In1[19]), .Z(n262) );
    VMW_FD \Out_reg[4]  ( .D(n331), .CP(Clk), .Q(Out[4]) );
    VMW_AOI211 U58 ( .A(n219), .B(In2[23]), .C(n252), .D(n216), .Z(n251) );
    VMW_INV U130 ( .A(Load), .Z(n293) );
    VMW_INV U138 ( .A(n233), .Z(n304) );
    VMW_INV U156 ( .A(n269), .Z(n320) );
    VMW_PULLDOWN U38 ( .Z(n339) );
    VMW_AOI211 U43 ( .A(n219), .B(In2[8]), .C(n222), .D(n216), .Z(n221) );
    VMW_AOI211 U64 ( .A(n219), .B(In2[18]), .C(n264), .D(n216), .Z(n263) );
    VMW_AND4 U81 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(n298
        ) );
    VMW_AO22 U104 ( .A(Out[30]), .B(n293), .C(n294), .D(In1[30]), .Z(n236) );
    VMW_AOI211 U51 ( .A(n219), .B(In2[2]), .C(n238), .D(n216), .Z(n237) );
    VMW_NOR2 U76 ( .A(n293), .B(n70), .Z(n219) );
    VMW_AO22 U116 ( .A(Out[1]), .B(n293), .C(n294), .D(In1[1]), .Z(n260) );
    VMW_AO22 U123 ( .A(Out[13]), .B(n293), .C(n294), .D(In1[13]), .Z(n274) );
    VMW_AND4 U88 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n300) );
    VMW_AND4 U93 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(n290
        ) );
    VMW_INV U131 ( .A(n218), .Z(n326) );
    VMW_INV U143 ( .A(n243), .Z(n308) );
    VMW_INV U144 ( .A(n245), .Z(n309) );
    VMW_INV U163 ( .A(n303), .Z(Read2) );
    VMW_INV U158 ( .A(n273), .Z(n322) );
    VMW_AOI211 U44 ( .A(n219), .B(In2[7]), .C(n224), .D(n216), .Z(n223) );
    VMW_AOI211 U56 ( .A(n219), .B(In2[25]), .C(n248), .D(n216), .Z(n247) );
    VMW_AND4 U94 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(n289
        ) );
    VMW_INV U136 ( .A(n229), .Z(n331) );
    VMW_AOI211 U71 ( .A(n219), .B(In2[11]), .C(n278), .D(n216), .Z(n277) );
    VMW_AO22 U111 ( .A(Out[24]), .B(n293), .C(n294), .D(In1[24]), .Z(n250) );
    VMW_AO22 U124 ( .A(Out[12]), .B(n293), .C(n294), .D(In1[12]), .Z(n276) );
    Merge_Node_DWIDTH32_DW01_cmp2_32_0 lte_86 ( .A(In1), .B(In2), .LEQ(n336), 
        .TC(n337), .LT_LE(n78) );
    VMW_AOI211 U63 ( .A(n219), .B(In2[19]), .C(n262), .D(n216), .Z(n261) );
    VMW_AND4 U78 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n295) );
    VMW_AND4 U86 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(n283
        ) );
    VMW_AO22 U103 ( .A(Out[31]), .B(n293), .C(n294), .D(In1[31]), .Z(n234) );
    VMW_AO22 U118 ( .A(Out[18]), .B(n293), .C(n294), .D(In1[18]), .Z(n264) );
    VMW_INV U151 ( .A(n259), .Z(n334) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n55, n72, n97, n20, n15, n69, n112, n32, n29, n85, n47, n60, n109, 
        n40, n67, n82, n99, n27, n35, n49, n107, n90, n52, n75, n98, n114, n34, 
        n26, n41, n66, n83, n53, n74, n91, n48, n106, n68, n101, n21, n46, n54, 
        n96, n73, n61, n28, n84, n33, n38, n56, n71, n113, n94, n23, n103, n16, 
        n78, n111, n31, n36, n44, n63, n86, n43, n64, n81, n58, n104, n18, n24, 
        n88, n37, n51, n93, n59, n76, n80, n42, n65, n19, n50, n77, n89, n92, 
        n25, n102, n105, n22, n39, n95, n45, n57, n70, n62, n87, n17, n30, n79, 
        n110;
    VMW_OAI21 U3 ( .A(A[31]), .B(n15), .C(n16), .Z(LT_LE) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n18), .C(B[0]), .Z(n19) );
    VMW_AO22 U6 ( .A(A[2]), .B(n21), .C(n19), .D(A[0]), .Z(n20) );
    VMW_OR2 U14 ( .A(B[6]), .B(n30), .Z(n33) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n46), .C(n41), .D(n36), .Z(n45) );
    VMW_OR2 U54 ( .A(B[26]), .B(n94), .Z(n97) );
    VMW_INV U73 ( .A(B[27]), .Z(n104) );
    VMW_INV U96 ( .A(A[16]), .Z(n62) );
    VMW_INV U68 ( .A(A[30]), .Z(n113) );
    VMW_NAND2 U28 ( .A(n56), .B(B[14]), .Z(n55) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n64), .C(n60), .D(n55), .Z(n63) );
    VMW_OAI22 U7 ( .A(n17), .B(n20), .C(A[2]), .D(n21), .Z(n22) );
    VMW_NAND2 U8 ( .A(n24), .B(B[4]), .Z(n23) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n32), .C(n28), .D(n23), .Z(n31) );
    VMW_OR2 U34 ( .A(B[16]), .B(n62), .Z(n65) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n78), .C(n73), .D(n68), .Z(n77) );
    VMW_NAND2 U46 ( .A(n84), .B(A[21]), .Z(n85) );
    VMW_NAND2 U61 ( .A(n110), .B(A[29]), .Z(n111) );
    VMW_INV U84 ( .A(A[4]), .Z(n24) );
    VMW_INV U101 ( .A(B[2]), .Z(n21) );
    VMW_INV U66 ( .A(B[7]), .Z(n39) );
    VMW_INV U83 ( .A(B[15]), .Z(n64) );
    VMW_INV U98 ( .A(A[26]), .Z(n94) );
    VMW_NAND2 U26 ( .A(n52), .B(A[11]), .Z(n53) );
    VMW_NAND2 U48 ( .A(n88), .B(B[24]), .Z(n87) );
    VMW_AO21 U9 ( .A(B[3]), .B(n26), .C(n22), .Z(n25) );
    VMW_NAND2 U12 ( .A(n30), .B(B[6]), .Z(n29) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n67), .C(n65), .D(n63), .Z(n66) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n96), .C(n92), .D(n87), .Z(n95) );
    VMW_INV U91 ( .A(A[28]), .Z(n102) );
    VMW_INV U74 ( .A(A[3]), .Z(n26) );
    VMW_INV U99 ( .A(B[23]), .Z(n90) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n50), .C(n53), .D(n51), .Z(n54) );
    VMW_NAND2 U40 ( .A(n76), .B(B[20]), .Z(n75) );
    VMW_INV U82 ( .A(A[15]), .Z(n67) );
    VMW_NAND2 U52 ( .A(n94), .B(B[26]), .Z(n93) );
    VMW_INV U67 ( .A(A[7]), .Z(n42) );
    VMW_INV U75 ( .A(B[25]), .Z(n96) );
    VMW_INV U90 ( .A(B[11]), .Z(n52) );
    VMW_NAND2 U20 ( .A(n44), .B(B[10]), .Z(n43) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n90), .C(n86), .D(n81), .Z(n89) );
    VMW_INV U69 ( .A(B[17]), .Z(n71) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n58), .C(n54), .D(n49), .Z(n57) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n82), .C(n85), .D(n83), .Z(n86) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n99), .C(n97), .D(n95), .Z(n98) );
    VMW_INV U72 ( .A(A[27]), .Z(n107) );
    VMW_INV U97 ( .A(B[13]), .Z(n58) );
    VMW_OAI211 U60 ( .A(A[29]), .B(n110), .C(n106), .D(n101), .Z(n109) );
    VMW_INV U100 ( .A(A[6]), .Z(n30) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n35), .C(n33), .D(n31), .Z(n34) );
    VMW_INV U85 ( .A(A[24]), .Z(n88) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n39), .C(n34), .D(n29), .Z(n38) );
    VMW_NAND2 U22 ( .A(n46), .B(A[9]), .Z(n47) );
    VMW_NAND2 U32 ( .A(n62), .B(B[16]), .Z(n61) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n74), .C(n72), .D(n70), .Z(n73) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n104), .C(n98), .D(n93), .Z(n103) );
    VMW_INV U70 ( .A(A[17]), .Z(n74) );
    VMW_INV U95 ( .A(B[31]), .Z(n15) );
    VMW_NAND2 U30 ( .A(n58), .B(A[13]), .Z(n59) );
    VMW_INV U79 ( .A(A[10]), .Z(n44) );
    VMW_INV U87 ( .A(B[21]), .Z(n84) );
    VMW_OR2 U10 ( .A(B[4]), .B(n24), .Z(n27) );
    VMW_NAND2 U42 ( .A(n78), .B(A[19]), .Z(n79) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n84), .C(n80), .D(n75), .Z(n83) );
    VMW_OAI211 U62 ( .A(B[30]), .B(n113), .C(n111), .D(n109), .Z(n112) );
    VMW_INV U65 ( .A(A[12]), .Z(n50) );
    VMW_INV U80 ( .A(B[9]), .Z(n46) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n26), .C(n27), .D(n25), .Z(n28) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n42), .C(n40), .D(n38), .Z(n41) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n52), .C(n48), .D(n43), .Z(n51) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n71), .C(n66), .D(n61), .Z(n70) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n107), .C(n105), .D(n103), .Z(n106) );
    VMW_INV U89 ( .A(A[14]), .Z(n56) );
    VMW_NAND2 U50 ( .A(n90), .B(A[23]), .Z(n91) );
    VMW_INV U77 ( .A(A[20]), .Z(n76) );
    VMW_INV U92 ( .A(A[5]), .Z(n35) );
    VMW_OR2 U58 ( .A(B[28]), .B(n102), .Z(n105) );
    VMW_NAND2 U36 ( .A(n69), .B(B[18]), .Z(n68) );
    VMW_INV U81 ( .A(B[29]), .Z(n110) );
    VMW_NOR2 U4 ( .A(n18), .B(B[1]), .Z(n17) );
    VMW_OR2 U18 ( .A(B[8]), .B(n37), .Z(n40) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n76), .C(n79), .D(n77), .Z(n80) );
    VMW_AO22 U64 ( .A(n112), .B(n114), .C(A[31]), .D(n15), .Z(n16) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n88), .C(n91), .D(n89), .Z(n92) );
    VMW_INV U76 ( .A(A[25]), .Z(n99) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n44), .C(n47), .D(n45), .Z(n48) );
    VMW_NAND2 U24 ( .A(n50), .B(B[12]), .Z(n49) );
    VMW_INV U88 ( .A(A[18]), .Z(n69) );
    VMW_INV U93 ( .A(B[5]), .Z(n32) );
    VMW_OR2 U38 ( .A(B[18]), .B(n69), .Z(n72) );
    VMW_NAND2 U44 ( .A(n82), .B(B[22]), .Z(n81) );
    VMW_NAND2 U56 ( .A(n102), .B(B[28]), .Z(n101) );
    VMW_INV U94 ( .A(A[1]), .Z(n18) );
    VMW_INV U71 ( .A(A[22]), .Z(n82) );
    VMW_NAND2 U63 ( .A(n113), .B(B[30]), .Z(n114) );
    VMW_INV U86 ( .A(A[8]), .Z(n37) );
    VMW_NAND2 U16 ( .A(n37), .B(B[8]), .Z(n36) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n56), .C(n59), .D(n57), .Z(n60) );
    VMW_INV U78 ( .A(B[19]), .Z(n78) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 ( A, B, LEQ, TC, 
    LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n115, n190, n149, n152, n175, n127, n135, n205, n199, n140, n167, 
        n182, n129, n185, n147, n160, n132, n202, n120, n169, n210, n155, n172, 
        n197, n133, n203, n146, n161, n121, n128, n184, n154, n196, n168, n173, 
        n211, n126, n148, n153, n174, n183, n191, n166, n141, n118, n134, n204, 
        n193, n198, n151, n176, n124, n188, n206, n136, n144, n143, n158, n164, 
        n163, n181, n186, n178, n116, n123, n131, n201, n213, n171, n156, n117, 
        n138, n194, n208, n130, n179, n200, n145, n162, n187, n195, n139, n209, 
        n170, n157, n122, n125, n212, n189, n150, n177, n192, n119, n142, n180, 
        n165, n159, n137, n207;
    VMW_AO21 U3 ( .A(n115), .B(A[31]), .C(n116), .Z(GE_GT) );
    VMW_AOI21 U5 ( .A(B[1]), .B(n118), .C(B[0]), .Z(n119) );
    VMW_AO22 U6 ( .A(A[2]), .B(n121), .C(n119), .D(A[0]), .Z(n120) );
    VMW_OR2 U14 ( .A(B[6]), .B(n130), .Z(n133) );
    VMW_OAI211 U21 ( .A(A[9]), .B(n146), .C(n141), .D(n136), .Z(n145) );
    VMW_OR2 U54 ( .A(B[26]), .B(n194), .Z(n197) );
    VMW_INV U73 ( .A(B[27]), .Z(n203) );
    VMW_INV U96 ( .A(n213), .Z(n116) );
    VMW_INV U68 ( .A(A[30]), .Z(n208) );
    VMW_NAND2 U28 ( .A(n156), .B(B[14]), .Z(n155) );
    VMW_OAI211 U33 ( .A(A[15]), .B(n164), .C(n160), .D(n155), .Z(n163) );
    VMW_OAI22 U7 ( .A(n117), .B(n120), .C(A[2]), .D(n121), .Z(n122) );
    VMW_NAND2 U8 ( .A(n124), .B(B[4]), .Z(n123) );
    VMW_OAI211 U13 ( .A(A[5]), .B(n132), .C(n128), .D(n123), .Z(n131) );
    VMW_OR2 U34 ( .A(B[16]), .B(n162), .Z(n165) );
    VMW_OAI211 U41 ( .A(A[19]), .B(n178), .C(n173), .D(n168), .Z(n177) );
    VMW_NAND2 U46 ( .A(n184), .B(A[21]), .Z(n185) );
    VMW_OAI211 U61 ( .A(A[29]), .B(n210), .C(n205), .D(n200), .Z(n209) );
    VMW_INV U84 ( .A(A[4]), .Z(n124) );
    VMW_INV U101 ( .A(A[6]), .Z(n130) );
    VMW_INV U66 ( .A(B[7]), .Z(n139) );
    VMW_INV U83 ( .A(B[15]), .Z(n164) );
    VMW_INV U98 ( .A(B[13]), .Z(n158) );
    VMW_NAND2 U26 ( .A(n152), .B(A[11]), .Z(n153) );
    VMW_NAND2 U48 ( .A(n188), .B(B[24]), .Z(n187) );
    VMW_AO21 U9 ( .A(B[3]), .B(n126), .C(n122), .Z(n125) );
    VMW_NAND2 U12 ( .A(n130), .B(B[6]), .Z(n129) );
    VMW_OAI211 U35 ( .A(B[15]), .B(n167), .C(n165), .D(n163), .Z(n166) );
    VMW_OAI211 U53 ( .A(A[25]), .B(n196), .C(n192), .D(n187), .Z(n195) );
    VMW_INV U91 ( .A(A[28]), .Z(n201) );
    VMW_INV U74 ( .A(A[3]), .Z(n126) );
    VMW_INV U99 ( .A(A[26]), .Z(n194) );
    VMW_OAI211 U27 ( .A(B[12]), .B(n150), .C(n153), .D(n151), .Z(n154) );
    VMW_NAND2 U40 ( .A(n176), .B(B[20]), .Z(n175) );
    VMW_INV U82 ( .A(A[15]), .Z(n167) );
    VMW_NAND2 U52 ( .A(n194), .B(B[26]), .Z(n193) );
    VMW_INV U67 ( .A(A[7]), .Z(n142) );
    VMW_INV U75 ( .A(B[25]), .Z(n196) );
    VMW_INV U90 ( .A(B[11]), .Z(n152) );
    VMW_NAND2 U20 ( .A(n144), .B(B[10]), .Z(n143) );
    VMW_OAI211 U49 ( .A(A[23]), .B(n190), .C(n186), .D(n181), .Z(n189) );
    VMW_INV U69 ( .A(B[17]), .Z(n171) );
    VMW_OAI211 U29 ( .A(A[13]), .B(n158), .C(n154), .D(n149), .Z(n157) );
    VMW_OAI211 U47 ( .A(B[22]), .B(n182), .C(n185), .D(n183), .Z(n186) );
    VMW_OAI211 U55 ( .A(B[25]), .B(n199), .C(n197), .D(n195), .Z(n198) );
    VMW_INV U72 ( .A(A[27]), .Z(n206) );
    VMW_INV U97 ( .A(A[16]), .Z(n162) );
    VMW_NAND2 U60 ( .A(n208), .B(B[30]), .Z(n207) );
    VMW_INV U100 ( .A(B[23]), .Z(n190) );
    VMW_OAI211 U15 ( .A(B[5]), .B(n135), .C(n133), .D(n131), .Z(n134) );
    VMW_INV U85 ( .A(A[24]), .Z(n188) );
    VMW_OAI211 U17 ( .A(A[7]), .B(n139), .C(n134), .D(n129), .Z(n138) );
    VMW_NAND2 U22 ( .A(n146), .B(A[9]), .Z(n147) );
    VMW_NAND2 U32 ( .A(n162), .B(B[16]), .Z(n161) );
    VMW_OAI211 U39 ( .A(B[17]), .B(n174), .C(n172), .D(n170), .Z(n173) );
    VMW_OAI211 U57 ( .A(A[27]), .B(n203), .C(n198), .D(n193), .Z(n202) );
    VMW_INV U70 ( .A(A[17]), .Z(n174) );
    VMW_INV U95 ( .A(B[31]), .Z(n115) );
    VMW_NAND2 U30 ( .A(n158), .B(A[13]), .Z(n159) );
    VMW_INV U79 ( .A(A[10]), .Z(n144) );
    VMW_INV U87 ( .A(B[21]), .Z(n184) );
    VMW_OR2 U10 ( .A(B[4]), .B(n124), .Z(n127) );
    VMW_NAND2 U42 ( .A(n178), .B(A[19]), .Z(n179) );
    VMW_OAI211 U45 ( .A(A[21]), .B(n184), .C(n180), .D(n175), .Z(n183) );
    VMW_NAND2 U62 ( .A(n210), .B(A[29]), .Z(n211) );
    VMW_INV U65 ( .A(A[12]), .Z(n150) );
    VMW_INV U102 ( .A(B[2]), .Z(n121) );
    VMW_INV U80 ( .A(B[9]), .Z(n146) );
    VMW_OAI211 U11 ( .A(B[3]), .B(n126), .C(n127), .D(n125), .Z(n128) );
    VMW_OAI211 U19 ( .A(B[7]), .B(n142), .C(n140), .D(n138), .Z(n141) );
    VMW_OAI211 U25 ( .A(A[11]), .B(n152), .C(n148), .D(n143), .Z(n151) );
    VMW_OAI211 U37 ( .A(A[17]), .B(n171), .C(n166), .D(n161), .Z(n170) );
    VMW_OAI211 U59 ( .A(B[27]), .B(n206), .C(n204), .D(n202), .Z(n205) );
    VMW_INV U89 ( .A(A[14]), .Z(n156) );
    VMW_NAND2 U50 ( .A(n190), .B(A[23]), .Z(n191) );
    VMW_INV U77 ( .A(A[20]), .Z(n176) );
    VMW_INV U92 ( .A(A[5]), .Z(n135) );
    VMW_OR2 U58 ( .A(B[28]), .B(n201), .Z(n204) );
    VMW_NAND2 U36 ( .A(n169), .B(B[18]), .Z(n168) );
    VMW_INV U81 ( .A(B[29]), .Z(n210) );
    VMW_NOR2 U4 ( .A(n118), .B(B[1]), .Z(n117) );
    VMW_OR2 U18 ( .A(B[8]), .B(n137), .Z(n140) );
    VMW_OAI211 U43 ( .A(B[20]), .B(n176), .C(n179), .D(n177), .Z(n180) );
    VMW_OAI211 U64 ( .A(A[31]), .B(n115), .C(n212), .D(n207), .Z(n213) );
    VMW_OAI211 U51 ( .A(B[24]), .B(n188), .C(n191), .D(n189), .Z(n192) );
    VMW_INV U76 ( .A(A[25]), .Z(n199) );
    VMW_OAI211 U23 ( .A(B[10]), .B(n144), .C(n147), .D(n145), .Z(n148) );
    VMW_NAND2 U24 ( .A(n150), .B(B[12]), .Z(n149) );
    VMW_INV U88 ( .A(A[18]), .Z(n169) );
    VMW_INV U93 ( .A(B[5]), .Z(n132) );
    VMW_OR2 U38 ( .A(B[18]), .B(n169), .Z(n172) );
    VMW_NAND2 U44 ( .A(n182), .B(B[22]), .Z(n181) );
    VMW_NAND2 U56 ( .A(n201), .B(B[28]), .Z(n200) );
    VMW_INV U94 ( .A(A[1]), .Z(n118) );
    VMW_INV U71 ( .A(A[22]), .Z(n182) );
    VMW_OAI211 U63 ( .A(B[30]), .B(n208), .C(n211), .D(n209), .Z(n212) );
    VMW_INV U86 ( .A(A[8]), .Z(n137) );
    VMW_NAND2 U16 ( .A(n137), .B(B[8]), .Z(n136) );
    VMW_OAI211 U31 ( .A(B[14]), .B(n156), .C(n159), .D(n157), .Z(n160) );
    VMW_INV U78 ( .A(B[19]), .Z(n178) );
endmodule


module Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, ScanId, Id, In1, In2, Read1, 
    Read2, Out );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] In1;
input  [31:0] ScanIn;
output [31:0] Out;
output [31:0] ScanOut;
input  [31:0] In2;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Read1, Read2;
    wire \Out[31] , n100, n245, n287, n317, n330, n262, n279, n362, n345, n357, 
        n339, n270, n257, n295, n305, n322, n292, n325, n302, n250, n277, n350, 
        n289, n319, n259, n342, n365, n265, n359, n356, \Out[5] , n280, n310, 
        n337, n288, n318, n351, \Out[24] , \Out[17] , n276, n251, \Out[30] , 
        n293, n303, n324, n281, n336, n311, \Out[29] , \Out[8] , \Out[1] , 
        n358, n243, n264, n258, n343, n364, \Out[20] , \Out[13] , \Out[26] , 
        \Out[22] , \Out[11] , \Out[18] , \Out[3] , n344, n278, n363, n244, 
        n263, n286, n316, n331, \Out[15] , n294, n304, n323, n256, n108, n271, 
        \Out[27] , \Out[14] , \Out[7] , n338, n284, n314, n333, n246, n261, 
        n361, n346, \Out[6] , n328, \Out[28] , \Out[23] , \Out[10] , \Out[19] , 
        \Out[2] , n268, n354, n368, n254, n273, n321, n306, n296, \Out[9] , 
        \Out[0] , n291, n301, n326, n348, n274, n253, n248, n353, \Out[25] , 
        \Out[21] , \Out[12] , \Out[16] , \Out[4] , n366, n298, n308, n341, 
        n266, n283, n313, n334, n249, n352, n349, n252, n275, n282, n290, n300, 
        n312, n327, n335, n267, n315, n367, n340, n299, n309, n329, n360, n347, 
        n247, n260, n332, n285, n269, n255, n297, n307, n320, n272, n355;
    assign ScanEnable = WR;
    assign DataOut[31] = \Out[31] ;
    assign DataOut[30] = \Out[30] ;
    assign DataOut[29] = \Out[29] ;
    assign DataOut[28] = \Out[28] ;
    assign DataOut[27] = \Out[27] ;
    assign DataOut[26] = \Out[26] ;
    assign DataOut[25] = \Out[25] ;
    assign DataOut[24] = \Out[24] ;
    assign DataOut[23] = \Out[23] ;
    assign DataOut[22] = \Out[22] ;
    assign DataOut[21] = \Out[21] ;
    assign DataOut[20] = \Out[20] ;
    assign DataOut[19] = \Out[19] ;
    assign DataOut[18] = \Out[18] ;
    assign DataOut[17] = \Out[17] ;
    assign DataOut[16] = \Out[16] ;
    assign DataOut[15] = \Out[15] ;
    assign DataOut[14] = \Out[14] ;
    assign DataOut[13] = \Out[13] ;
    assign DataOut[12] = \Out[12] ;
    assign DataOut[11] = \Out[11] ;
    assign DataOut[10] = \Out[10] ;
    assign DataOut[9] = \Out[9] ;
    assign DataOut[8] = \Out[8] ;
    assign DataOut[7] = \Out[7] ;
    assign DataOut[6] = \Out[6] ;
    assign DataOut[5] = \Out[5] ;
    assign DataOut[4] = \Out[4] ;
    assign DataOut[3] = \Out[3] ;
    assign DataOut[2] = \Out[2] ;
    assign DataOut[1] = \Out[1] ;
    assign DataOut[0] = \Out[0] ;
    assign Out[31] = \Out[31] ;
    assign Out[30] = \Out[30] ;
    assign Out[29] = \Out[29] ;
    assign Out[28] = \Out[28] ;
    assign Out[27] = \Out[27] ;
    assign Out[26] = \Out[26] ;
    assign Out[25] = \Out[25] ;
    assign Out[24] = \Out[24] ;
    assign Out[23] = \Out[23] ;
    assign Out[22] = \Out[22] ;
    assign Out[21] = \Out[21] ;
    assign Out[20] = \Out[20] ;
    assign Out[19] = \Out[19] ;
    assign Out[18] = \Out[18] ;
    assign Out[17] = \Out[17] ;
    assign Out[16] = \Out[16] ;
    assign Out[15] = \Out[15] ;
    assign Out[14] = \Out[14] ;
    assign Out[13] = \Out[13] ;
    assign Out[12] = \Out[12] ;
    assign Out[11] = \Out[11] ;
    assign Out[10] = \Out[10] ;
    assign Out[9] = \Out[9] ;
    assign Out[8] = \Out[8] ;
    assign Out[7] = \Out[7] ;
    assign Out[6] = \Out[6] ;
    assign Out[5] = \Out[5] ;
    assign Out[4] = \Out[4] ;
    assign Out[3] = \Out[3] ;
    assign Out[2] = \Out[2] ;
    assign Out[1] = \Out[1] ;
    assign Out[0] = \Out[0] ;
    VMW_AND2 U54 ( .A(DataIn[24]), .B(ScanEnable), .Z(ScanOut[24]) );
    VMW_AND2 U73 ( .A(DataIn[5]), .B(ScanEnable), .Z(ScanOut[5]) );
    VMW_AND5 U113 ( .A(n317), .B(n318), .C(n319), .D(n320), .E(n321), .Z(n246)
         );
    VMW_AO22 U134 ( .A(\Out[9] ), .B(n322), .C(n323), .D(In1[9]), .Z(n249) );
    VMW_AND2 U68 ( .A(DataIn[10]), .B(ScanEnable), .Z(ScanOut[10]) );
    VMW_AOI211 U96 ( .A(n248), .B(In2[23]), .C(n281), .D(n245), .Z(n280) );
    VMW_INV U198 ( .A(n306), .Z(n353) );
    VMW_AOI211 U108 ( .A(n248), .B(In2[12]), .C(n305), .D(n245), .Z(n304) );
    VMW_AO22 U141 ( .A(\Out[31] ), .B(n322), .C(n323), .D(In1[31]), .Z(n263)
         );
    VMW_OAI21 U166 ( .A(n108), .B(n246), .C(RD), .Z(n332) );
    VMW_INV U183 ( .A(n276), .Z(n339) );
    VMW_OAI21 U46 ( .A(n100), .B(n244), .C(RD), .Z(n243) );
    VMW_AND2 U61 ( .A(DataIn[17]), .B(ScanEnable), .Z(ScanOut[17]) );
    VMW_AOI211 U84 ( .A(n248), .B(In2[5]), .C(n257), .D(n245), .Z(n256) );
    VMW_AO22 U148 ( .A(\Out[25] ), .B(n322), .C(n323), .D(In1[25]), .Z(n277)
         );
    VMW_AO22 U153 ( .A(\Out[20] ), .B(n322), .C(n323), .D(In1[20]), .Z(n287)
         );
    VMW_INV U174 ( .A(n258), .Z(n360) );
    VMW_INV U191 ( .A(n292), .Z(n346) );
    VMW_AOI211 U101 ( .A(n248), .B(In2[19]), .C(n291), .D(n245), .Z(n290) );
    VMW_AND4 U126 ( .A(In1[7]), .B(In1[6]), .C(In1[5]), .D(In1[4]), .Z(n329)
         );
    VMW_AND2 U48 ( .A(DataIn[30]), .B(ScanEnable), .Z(ScanOut[30]) );
    VMW_AND2 U66 ( .A(DataIn[12]), .B(ScanEnable), .Z(ScanOut[12]) );
    VMW_AOI211 U106 ( .A(n248), .B(In2[14]), .C(n301), .D(n245), .Z(n300) );
    VMW_AND4 U121 ( .A(In2[19]), .B(In2[18]), .C(In2[17]), .D(In2[16]), .Z(
        n320) );
    VMW_AOI211 U83 ( .A(n248), .B(In2[6]), .C(n255), .D(n245), .Z(n254) );
    VMW_INV U168 ( .A(RD), .Z(n322) );
    VMW_AOI211 U98 ( .A(n248), .B(In2[21]), .C(n285), .D(n245), .Z(n284) );
    VMW_AND4 U128 ( .A(In1[15]), .B(In1[14]), .C(In1[13]), .D(In1[12]), .Z(
        n331) );
    VMW_AO22 U154 ( .A(\Out[1] ), .B(n322), .C(n323), .D(In1[1]), .Z(n289) );
    VMW_INV U173 ( .A(n256), .Z(n359) );
    VMW_INV U184 ( .A(n278), .Z(n340) );
    VMW_INV U196 ( .A(n302), .Z(n351) );
    VMW_AND2 U53 ( .A(DataIn[25]), .B(ScanEnable), .Z(ScanOut[25]) );
    VMW_AOI211 U91 ( .A(n248), .B(In2[28]), .C(n271), .D(n245), .Z(n270) );
    VMW_AO22 U146 ( .A(\Out[27] ), .B(n322), .C(n323), .D(In1[27]), .Z(n273)
         );
    VMW_AO22 U161 ( .A(\Out[13] ), .B(n322), .C(n323), .D(In1[13]), .Z(n303)
         );
    VMW_AND2 U74 ( .A(DataIn[4]), .B(ScanEnable), .Z(ScanOut[4]) );
    VMW_NOR2 U114 ( .A(n322), .B(n100), .Z(n248) );
    VMW_AND4 U133 ( .A(In1[31]), .B(In1[30]), .C(In1[29]), .D(In1[28]), .Z(
        n312) );
    VMW_AOI211 U99 ( .A(n248), .B(In2[20]), .C(n287), .D(n245), .Z(n286) );
    VMW_INV U197 ( .A(n304), .Z(n352) );
    VMW_AO22 U155 ( .A(\Out[19] ), .B(n322), .C(n323), .D(In1[19]), .Z(n291)
         );
    VMW_FD \Out_reg[16]  ( .D(n348), .CP(Clk), .Q(\Out[16] ) );
    VMW_INV U172 ( .A(n254), .Z(n358) );
    VMW_FD \Out_reg[25]  ( .D(n339), .CP(Clk), .Q(\Out[25] ) );
    VMW_AND2 U47 ( .A(DataIn[31]), .B(ScanEnable), .Z(ScanOut[31]) );
    VMW_AND2 U49 ( .A(DataIn[29]), .B(ScanEnable), .Z(ScanOut[29]) );
    VMW_AND2 U52 ( .A(DataIn[26]), .B(ScanEnable), .Z(ScanOut[26]) );
    VMW_AND2 U67 ( .A(DataIn[11]), .B(ScanEnable), .Z(ScanOut[11]) );
    VMW_AOI211 U82 ( .A(n248), .B(In2[7]), .C(n253), .D(n245), .Z(n252) );
    VMW_INV U169 ( .A(n247), .Z(n355) );
    VMW_AOI211 U107 ( .A(n248), .B(In2[13]), .C(n303), .D(n245), .Z(n302) );
    VMW_AND4 U120 ( .A(n327), .B(n326), .C(n325), .D(n324), .Z(n321) );
    VMW_FD \Out_reg[5]  ( .D(n359), .CP(Clk), .Q(\Out[5] ) );
    VMW_AND2 U75 ( .A(DataIn[3]), .B(ScanEnable), .Z(ScanOut[3]) );
    VMW_AND2 U115 ( .A(n100), .B(RD), .Z(n323) );
    VMW_AND4 U132 ( .A(In1[27]), .B(In1[26]), .C(In1[25]), .D(In1[24]), .Z(
        n313) );
    VMW_FD \Out_reg[12]  ( .D(n352), .CP(Clk), .Q(\Out[12] ) );
    VMW_AOI211 U90 ( .A(n248), .B(In2[29]), .C(n269), .D(n245), .Z(n268) );
    VMW_FD \Out_reg[21]  ( .D(n343), .CP(Clk), .Q(\Out[21] ) );
    VMW_AND4 U129 ( .A(n331), .B(n330), .C(n329), .D(n328), .Z(n316) );
    VMW_AO22 U147 ( .A(\Out[26] ), .B(n322), .C(n323), .D(In1[26]), .Z(n275)
         );
    VMW_FD \Out_reg[8]  ( .D(n356), .CP(Clk), .Q(\Out[8] ) );
    VMW_AO22 U160 ( .A(\Out[14] ), .B(n322), .C(n323), .D(In1[14]), .Z(n301)
         );
    VMW_INV U185 ( .A(n280), .Z(n341) );
    VMW_FD \Out_reg[31]  ( .D(n333), .CP(Clk), .Q(\Out[31] ) );
    VMW_FD \Out_reg[28]  ( .D(n336), .CP(Clk), .Q(\Out[28] ) );
    VMW_FD \Out_reg[1]  ( .D(n363), .CP(Clk), .Q(\Out[1] ) );
    VMW_AND2 U55 ( .A(DataIn[23]), .B(ScanEnable), .Z(ScanOut[23]) );
    VMW_AND2 U69 ( .A(ScanEnable), .B(DataIn[9]), .Z(ScanOut[9]) );
    VMW_AOI211 U109 ( .A(n248), .B(In2[11]), .C(n307), .D(n245), .Z(n306) );
    VMW_INV U182 ( .A(n274), .Z(n338) );
    VMW_FD \Out_reg[19]  ( .D(n345), .CP(Clk), .Q(\Out[19] ) );
    VMW_AND2 U72 ( .A(DataIn[6]), .B(ScanEnable), .Z(ScanOut[6]) );
    VMW_AOI211 U97 ( .A(n248), .B(In2[22]), .C(n283), .D(n245), .Z(n282) );
    VMW_AO22 U140 ( .A(\Out[3] ), .B(n322), .C(n323), .D(In1[3]), .Z(n261) );
    VMW_INV U167 ( .A(n243), .Z(Read1) );
    VMW_FD \Out_reg[3]  ( .D(n361), .CP(Clk), .Q(\Out[3] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_0 r141 ( .A(In1), .B(
        In2), .LEQ(n365), .TC(n366), .GE_GT(n100) );
    VMW_AND5 U112 ( .A(n312), .B(n313), .C(n314), .D(n315), .E(n316), .Z(n244)
         );
    VMW_AO22 U135 ( .A(\Out[8] ), .B(n322), .C(n323), .D(In1[8]), .Z(n251) );
    VMW_FD \Out_reg[10]  ( .D(n354), .CP(Clk), .Q(\Out[10] ) );
    VMW_FD \Out_reg[23]  ( .D(n341), .CP(Clk), .Q(\Out[23] ) );
    VMW_AND2 U60 ( .A(DataIn[18]), .B(ScanEnable), .Z(ScanOut[18]) );
    VMW_INV U199 ( .A(n308), .Z(n354) );
    VMW_FD \Out_reg[7]  ( .D(n357), .CP(Clk), .Q(\Out[7] ) );
    VMW_AOI211 U100 ( .A(n248), .B(In2[1]), .C(n289), .D(n245), .Z(n288) );
    VMW_AND4 U127 ( .A(In1[11]), .B(In1[10]), .C(In1[9]), .D(In1[8]), .Z(n330)
         );
    VMW_AOI211 U85 ( .A(n248), .B(In2[4]), .C(n259), .D(n245), .Z(n258) );
    VMW_AO22 U149 ( .A(\Out[24] ), .B(n322), .C(n323), .D(In1[24]), .Z(n279)
         );
    VMW_AO22 U152 ( .A(\Out[21] ), .B(n322), .C(n323), .D(In1[21]), .Z(n285)
         );
    VMW_INV U175 ( .A(n260), .Z(n361) );
    VMW_FD \Out_reg[14]  ( .D(n350), .CP(Clk), .Q(\Out[14] ) );
    VMW_FD \Out_reg[27]  ( .D(n337), .CP(Clk), .Q(\Out[27] ) );
    VMW_PULLDOWN U42 ( .Z(n366) );
    VMW_PULLUP U45 ( .Z(n367) );
    VMW_AND2 U57 ( .A(DataIn[21]), .B(ScanEnable), .Z(ScanOut[21]) );
    VMW_AO22 U137 ( .A(\Out[6] ), .B(n322), .C(n323), .D(In1[6]), .Z(n255) );
    VMW_INV U190 ( .A(n290), .Z(n345) );
    VMW_FD \Out_reg[6]  ( .D(n358), .CP(Clk), .Q(\Out[6] ) );
    VMW_AND2 U70 ( .A(DataIn[8]), .B(ScanEnable), .Z(ScanOut[8]) );
    VMW_AO21 U79 ( .A(n246), .B(n244), .C(Reset), .Z(n245) );
    VMW_AOI211 U95 ( .A(n248), .B(In2[24]), .C(n279), .D(n245), .Z(n278) );
    VMW_AOI211 U110 ( .A(n248), .B(In2[10]), .C(n309), .D(n245), .Z(n308) );
    VMW_AO22 U159 ( .A(\Out[15] ), .B(n322), .C(n323), .D(In1[15]), .Z(n299)
         );
    VMW_AND4 U119 ( .A(In2[15]), .B(In2[14]), .C(In2[13]), .D(In2[12]), .Z(
        n327) );
    VMW_AO22 U142 ( .A(\Out[30] ), .B(n322), .C(n323), .D(In1[30]), .Z(n265)
         );
    VMW_AO22 U165 ( .A(\Out[0] ), .B(n322), .C(n323), .D(In1[0]), .Z(n311) );
    VMW_INV U180 ( .A(n270), .Z(n336) );
    VMW_FD \Out_reg[26]  ( .D(n338), .CP(Clk), .Q(\Out[26] ) );
    VMW_FD \Out_reg[15]  ( .D(n349), .CP(Clk), .Q(\Out[15] ) );
    VMW_INV U192 ( .A(n294), .Z(n347) );
    VMW_FD \Out_reg[18]  ( .D(n346), .CP(Clk), .Q(\Out[18] ) );
    VMW_AOI211 U87 ( .A(n248), .B(In2[31]), .C(n263), .D(n245), .Z(n262) );
    VMW_AO22 U150 ( .A(\Out[23] ), .B(n322), .C(n323), .D(In1[23]), .Z(n281)
         );
    VMW_INV U177 ( .A(n264), .Z(n334) );
    VMW_FD \Out_reg[2]  ( .D(n362), .CP(Clk), .Q(\Out[2] ) );
    VMW_AND4 U125 ( .A(In1[3]), .B(In1[2]), .C(In1[1]), .D(In1[0]), .Z(n328)
         );
    VMW_FD \Out_reg[11]  ( .D(n353), .CP(Clk), .Q(\Out[11] ) );
    VMW_AND2 U62 ( .A(DataIn[16]), .B(ScanEnable), .Z(ScanOut[16]) );
    VMW_FD \Out_reg[22]  ( .D(n342), .CP(Clk), .Q(\Out[22] ) );
    VMW_AND2 U65 ( .A(DataIn[13]), .B(ScanEnable), .Z(ScanOut[13]) );
    VMW_AOI211 U102 ( .A(n248), .B(In2[18]), .C(n293), .D(n245), .Z(n292) );
    VMW_AOI211 U105 ( .A(n248), .B(In2[15]), .C(n299), .D(n245), .Z(n298) );
    VMW_INV U189 ( .A(n288), .Z(n363) );
    VMW_FD \Out_reg[20]  ( .D(n344), .CP(Clk), .Q(\Out[20] ) );
    VMW_FD \Out_reg[13]  ( .D(n351), .CP(Clk), .Q(\Out[13] ) );
    VMW_PULLUP U43 ( .Z(n365) );
    VMW_AND2 U50 ( .A(DataIn[28]), .B(ScanEnable), .Z(ScanOut[28]) );
    VMW_AND2 U59 ( .A(DataIn[19]), .B(ScanEnable), .Z(ScanOut[19]) );
    VMW_AOI211 U80 ( .A(n248), .B(In2[9]), .C(n249), .D(n245), .Z(n247) );
    VMW_AND4 U122 ( .A(In2[23]), .B(In2[22]), .C(In2[21]), .D(In2[20]), .Z(
        n319) );
    VMW_AO22 U139 ( .A(\Out[4] ), .B(n322), .C(n323), .D(In1[4]), .Z(n259) );
    VMW_AO22 U157 ( .A(\Out[17] ), .B(n322), .C(n323), .D(In1[17]), .Z(n295)
         );
    VMW_INV U170 ( .A(n250), .Z(n356) );
    VMW_FD \Out_reg[9]  ( .D(n355), .CP(Clk), .Q(\Out[9] ) );
    VMW_INV U195 ( .A(n300), .Z(n350) );
    VMW_FD \Out_reg[30]  ( .D(n334), .CP(Clk), .Q(\Out[30] ) );
    VMW_FD \Out_reg[0]  ( .D(n364), .CP(Clk), .Q(\Out[0] ) );
    VMW_FD \Out_reg[29]  ( .D(n335), .CP(Clk), .Q(\Out[29] ) );
    VMW_AND2 U77 ( .A(DataIn[1]), .B(ScanEnable), .Z(ScanOut[1]) );
    VMW_AOI211 U89 ( .A(n248), .B(In2[2]), .C(n267), .D(n245), .Z(n266) );
    VMW_INV U187 ( .A(n284), .Z(n343) );
    VMW_AOI211 U92 ( .A(n248), .B(In2[27]), .C(n273), .D(n245), .Z(n272) );
    VMW_AO22 U145 ( .A(\Out[28] ), .B(n322), .C(n323), .D(In1[28]), .Z(n271)
         );
    VMW_AO22 U162 ( .A(\Out[12] ), .B(n322), .C(n323), .D(In1[12]), .Z(n305)
         );
    VMW_INV U179 ( .A(n268), .Z(n335) );
    VMW_FD \Out_reg[24]  ( .D(n340), .CP(Clk), .Q(\Out[24] ) );
    VMW_FD \Out_reg[17]  ( .D(n347), .CP(Clk), .Q(\Out[17] ) );
    VMW_AND4 U117 ( .A(In2[7]), .B(In2[6]), .C(In2[5]), .D(In2[4]), .Z(n325)
         );
    VMW_FD \Out_reg[4]  ( .D(n360), .CP(Clk), .Q(\Out[4] ) );
    VMW_INV U200 ( .A(n310), .Z(n364) );
    VMW_AND2 U58 ( .A(DataIn[20]), .B(ScanEnable), .Z(ScanOut[20]) );
    VMW_AND4 U130 ( .A(In1[19]), .B(In1[18]), .C(In1[17]), .D(In1[16]), .Z(
        n315) );
    VMW_AO22 U138 ( .A(\Out[5] ), .B(n322), .C(n323), .D(In1[5]), .Z(n257) );
    VMW_INV U194 ( .A(n298), .Z(n349) );
    VMW_AND2 U64 ( .A(DataIn[14]), .B(ScanEnable), .Z(ScanOut[14]) );
    VMW_AOI211 U81 ( .A(n248), .B(In2[8]), .C(n251), .D(n245), .Z(n250) );
    VMW_AO22 U156 ( .A(\Out[18] ), .B(n322), .C(n323), .D(In1[18]), .Z(n293)
         );
    VMW_INV U171 ( .A(n252), .Z(n357) );
    VMW_AOI211 U104 ( .A(n248), .B(In2[16]), .C(n297), .D(n245), .Z(n296) );
    VMW_PULLDOWN U44 ( .Z(n368) );
    VMW_AND2 U51 ( .A(DataIn[27]), .B(ScanEnable), .Z(ScanOut[27]) );
    VMW_AND2 U76 ( .A(DataIn[2]), .B(ScanEnable), .Z(ScanOut[2]) );
    VMW_AND4 U116 ( .A(In2[3]), .B(In2[2]), .C(In2[1]), .D(In2[0]), .Z(n324)
         );
    VMW_AND4 U123 ( .A(In2[27]), .B(In2[26]), .C(In2[25]), .D(In2[24]), .Z(
        n318) );
    VMW_AND2 U56 ( .A(DataIn[22]), .B(ScanEnable), .Z(ScanOut[22]) );
    VMW_AOI211 U88 ( .A(n248), .B(In2[30]), .C(n265), .D(n245), .Z(n264) );
    VMW_AOI211 U93 ( .A(n248), .B(In2[26]), .C(n275), .D(n245), .Z(n274) );
    VMW_AND4 U131 ( .A(In1[23]), .B(In1[22]), .C(In1[21]), .D(In1[20]), .Z(
        n314) );
    VMW_INV U201 ( .A(n332), .Z(Read2) );
    VMW_INV U178 ( .A(n266), .Z(n362) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1_DW01_cmp2_32_1 lte_43 ( .A(In1), 
        .B(In2), .LEQ(n367), .TC(n368), .LT_LE(n108) );
    VMW_AOI211 U94 ( .A(n248), .B(In2[25]), .C(n277), .D(n245), .Z(n276) );
    VMW_AO22 U143 ( .A(\Out[2] ), .B(n322), .C(n323), .D(In1[2]), .Z(n267) );
    VMW_AO22 U144 ( .A(\Out[29] ), .B(n322), .C(n323), .D(In1[29]), .Z(n269)
         );
    VMW_AO22 U163 ( .A(\Out[11] ), .B(n322), .C(n323), .D(In1[11]), .Z(n307)
         );
    VMW_INV U181 ( .A(n272), .Z(n337) );
    VMW_INV U186 ( .A(n282), .Z(n342) );
    VMW_AO22 U158 ( .A(\Out[16] ), .B(n322), .C(n323), .D(In1[16]), .Z(n297)
         );
    VMW_AO22 U164 ( .A(\Out[10] ), .B(n322), .C(n323), .D(In1[10]), .Z(n309)
         );
    VMW_AO22 U136 ( .A(\Out[7] ), .B(n322), .C(n323), .D(In1[7]), .Z(n253) );
    VMW_AND2 U71 ( .A(DataIn[7]), .B(ScanEnable), .Z(ScanOut[7]) );
    VMW_AOI211 U111 ( .A(n248), .B(In2[0]), .C(n311), .D(n245), .Z(n310) );
    VMW_AND4 U124 ( .A(In2[31]), .B(In2[30]), .C(In2[29]), .D(In2[28]), .Z(
        n317) );
    VMW_AND2 U63 ( .A(DataIn[15]), .B(ScanEnable), .Z(ScanOut[15]) );
    VMW_AND2 U78 ( .A(DataIn[0]), .B(ScanEnable), .Z(ScanOut[0]) );
    VMW_AOI211 U86 ( .A(n248), .B(In2[3]), .C(n261), .D(n245), .Z(n260) );
    VMW_AOI211 U103 ( .A(n248), .B(In2[17]), .C(n295), .D(n245), .Z(n294) );
    VMW_INV U188 ( .A(n286), .Z(n344) );
    VMW_AND4 U118 ( .A(In2[11]), .B(In2[10]), .C(In2[9]), .D(In2[8]), .Z(n326)
         );
    VMW_AO22 U151 ( .A(\Out[22] ), .B(n322), .C(n323), .D(In1[22]), .Z(n283)
         );
    VMW_INV U176 ( .A(n262), .Z(n333) );
    VMW_INV U193 ( .A(n296), .Z(n348) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \Level1Out10[15] , \Level1Out33[24] , \Level1Out46[14] , 
        \Level2Out8[24] , \Level1Out53[20] , \ScanLink0[13] , \Level1Out11[2] , 
        \ScanLink24[18] , \Level1Out26[10] , \ScanLink50[8] , \ScanLink51[31] , 
        \ScanLink51[28] , \Level4Out0[18] , \Level1Out12[1] , 
        \Level1Out26[23] , \ScanLink29[3] , \ScanLink0[20] , \Level1Out10[26] , 
        \Level1Out33[17] , \Level1Out53[13] , \Level1Out46[27] , 
        \Level2Out8[17] , \ScanLink1[19] , \Level1Out1[7] , \Level1Out2[23] , 
        \ScanLink19[22] , \Level1Load28[0] , \Level8Out8[6] , 
        \Level2Out52[15] , \Level2Out32[11] , \Level1Out2[10] , \ScanLink9[6] , 
        \ScanLink55[5] , \ScanLink56[6] , \Level2Load44[0] , \Level4Out48[1] , 
        \Level32Out32[30] , \Level32Out32[29] , \ScanLink32[2] , 
        \Level1Out38[31] , \Level1Out38[28] , \Level2Out60[0] , 
        \Level1Out6[21] , \ScanLink15[7] , \ScanLink19[11] , \Level2Out32[22] , 
        \Level4Out32[9] , \Level2Out52[26] , \ScanLink31[1] , 
        \Level8Out16[31] , \Level8Out16[28] , \Level8Out40[29] , 
        \Level8Out40[30] , \Level1Out49[2] , \Level2Out0[0] , \Level2Out20[2] , 
        \Level16Out48[19] , \Level1Out49[30] , \Level1Out49[29] , 
        \ScanLink16[4] , \Level1Out30[9] , \Level2Out36[13] , 
        \Level2Out60[12] , \Level2Out44[6] , \Level2Out56[17] , 
        \Level1Out2[4] , \ScanLink4[22] , \ScanLink4[11] , \Level1Out6[12] , 
        \Level2Out36[20] , \Level2Out56[24] , \Level2Out60[21] , 
        \Level1Load7[0] , \Level1Out52[3] , \Level16Out32[27] , 
        \Level1Out7[9] , \ScanLink13[9] , \Level1Out14[17] , \Level1Out22[12] , 
        \Level1Out51[0] , \Level1Out57[22] , \Level2Out28[18] , 
        \Level2Out38[0] , \Level8Load16[0] , \Level4Out4[6] , 
        \Level1Out37[26] , \Level1Out42[16] , \Level1Out61[27] , 
        \Level4Out4[30] , \Level4Out4[29] , \Level2Out42[8] , \ScanLink5[31] , 
        \ScanLink5[28] , \Level1Out7[18] , \Level1Out14[24] , \Level1Out35[4] , 
        \Level1Out36[7] , \Level1Out37[15] , \Level16Out32[14] , 
        \Level1Out42[25] , \ScanLink20[30] , \Level1Out22[21] , 
        \Level1Out61[14] , \Level1Out57[11] , \ScanLink20[29] , 
        \Level1Out28[14] , \ScanLink55[19] , \ScanLink17[26] , \ScanLink18[2] , 
        \Level1Out20[3] , \Level1Out23[0] , \Level1Out48[10] , 
        \Level2Out6[20] , \Level1Out28[27] , \Level1Out47[4] , \ScanLink61[9] , 
        \Level2Out14[31] , \Level2Out42[29] , \Level2Out42[30] , 
        \Level1Out48[23] , \Level2Out6[13] , \Level2Out14[28] , 
        \Level1Out44[7] , \Level1Out59[8] , \Level4Out52[29] , 
        \Level2Out30[8] , \Level4Out52[30] , \ScanLink21[23] , 
        \Level1Out38[1] , \ScanLink54[13] , \ScanLink34[17] , \ScanLink62[16] , 
        \ScanLink41[27] , \ScanLink64[4] , \Level2Out52[2] , \Level1Out8[25] , 
        \ScanLink17[15] , \Level1Out23[18] , \Level1Out56[28] , 
        \Level1Out56[31] , \ScanLink62[25] , \Level2Out8[8] , \ScanLink21[10] , 
        \ScanLink34[24] , \ScanLink41[14] , \ScanLink54[20] , \ScanLink27[5] , 
        \Level1Out42[9] , \Level2Out36[6] , \Level1Out27[29] , 
        \Level2Out12[0] , \Level2Load36[0] , \Level4Out48[13] , 
        \Level4Out28[17] , \Level1Out52[19] , \ScanLink13[24] , 
        \Level1Out27[30] , \ScanLink39[9] , \ScanLink24[6] , \ScanLink30[15] , 
        \ScanLink45[25] , \Level2Out58[13] , \ScanLink25[21] , 
        \ScanLink50[11] , \Level2Out38[17] , \Level4Out28[24] , 
        \Level8Out8[10] , \Level1Out8[16] , \ScanLink13[17] , \ScanLink25[12] , 
        \ScanLink40[2] , \ScanLink43[1] , \Level4Out48[20] , \ScanLink50[22] , 
        \Level2Out38[24] , \Level8Out8[23] , \ScanLink30[26] , 
        \ScanLink45[16] , \Level16Out0[6] , \Level2Out58[20] , 
        \Level4Out40[9] , \ScanLink22[8] , \Level1Out60[1] , \Level4Out56[18] , 
        \Level1Out63[2] , \Level2Out10[19] , \Level2Out46[18] , 
        \Level2Out2[22] , \Level1Out39[22] , \ScanLink58[0] , 
        \Level1Out59[26] , \ScanLink0[30] , \ScanLink1[23] , \ScanLink1[10] , 
        \Level1Out3[30] , \ScanLink4[3] , \ScanLink7[0] , \Level32Out0[31] , 
        \Level32Out0[28] , \Level1Out3[29] , \Level1Out59[15] , 
        \Level1Out3[20] , \ScanLink5[21] , \ScanLink5[12] , \Level1Out15[14] , 
        \ScanLink18[31] , \ScanLink18[28] , \Level1Out39[11] , 
        \Level2Out2[11] , \Level1Out60[24] , \ScanLink21[19] , 
        \Level1Out23[11] , \Level1Out36[25] , \Level1Out43[15] , 
        \Level1Out41[3] , \Level1Out56[21] , \ScanLink54[29] , 
        \Level1Load63[0] , \Level2Out8[1] , \ScanLink54[30] , \Level2Out28[3] , 
        \Level1Out9[6] , \Level1Out42[0] , \Level1Out15[27] , 
        \Level1Out23[22] , \Level1Out38[8] , \Level1Out56[12] , 
        \Level1Out25[7] , \Level1Out36[16] , \Level1Out60[17] , 
        \Level1Out43[26] , \ScanLink7[9] , \Level1Out7[22] , \Level1Out26[4] , 
        \Level2Out14[21] , \Level2Out22[24] , \Level2Out42[20] , 
        \Level1Out7[11] , \Level1Out48[19] , \Level1Out59[1] , 
        \Level4Out32[24] , \Level4Out52[20] , \ScanLink62[3] , 
        \Level2Out6[29] , \Level2Out30[1] , \Level2Out6[30] , \Level1Out19[3] , 
        \Level1Out23[9] , \Level2Out14[12] , \Level2Out42[13] , 
        \ScanLink58[9] , \ScanLink61[0] , \Level2Out22[17] , \Level2Out54[5] , 
        \Level4Out52[13] , \Level4Out32[17] , \Level4Out56[22] , 
        \Level1Out39[18] , \ScanLink45[6] , \Level4Out60[27] , 
        \Level32Out0[21] , \Level2Out2[18] , \Level4Out36[26] , 
        \Level1Out3[13] , \ScanLink18[21] , \ScanLink46[5] , \Level2Out10[23] , 
        \Level2Out46[22] , \ScanLink18[12] , \ScanLink21[2] , 
        \Level2Out26[26] , \Level4Out36[15] , \Level4Load60[0] , 
        \Level4Out60[14] , \Level4Out56[11] , \Level1Out60[8] , 
        \Level2Out14[7] , \Level32Out0[12] , \Level2Out10[10] , 
        \Level2Out26[15] , \Level2Out46[11] , \Level8Out0[7] , \ScanLink22[1] , 
        \Level4Out48[30] , \Level4Out48[29] , \ScanLink1[7] , \ScanLink2[4] , 
        \ScanLink43[8] , \Level2Out58[30] , \Level2Out58[29] , 
        \Level1Out11[16] , \Level1Out27[13] , \Level1Out52[23] , 
        \Level1Out32[27] , \Level1Out47[17] , \Level4Out40[0] , 
        \Level2Out12[9] , \Level32Out32[3] , \Level1Out2[19] , 
        \Level1Out11[25] , \ScanLink25[31] , \ScanLink25[28] , 
        \Level1Out27[20] , \Level1Out32[14] , \Level1Out47[24] , 
        \ScanLink39[0] , \Level1Out52[10] , \Level4Out24[4] , \ScanLink50[18] , 
        \Level8Out8[19] , \Level1Out9[26] , \ScanLink12[27] , \Level1Out14[6] , 
        \Level1Out17[5] , \ScanLink19[18] , \Level1Out38[21] , 
        \Level1Out58[25] , \ScanLink31[8] , \Level4Out32[0] , 
        \Level8Out16[21] , \Level8Out40[20] , \Level32Out32[13] , 
        \Level16Out48[10] , \Level1Out38[12] , \Level2Out32[18] , 
        \Level4Out56[4] , \Level1Out58[16] , \Level2Out60[9] , 
        \Level4Out48[8] , \Level16Out48[23] , \Level8Out40[13] , 
        \Level32Out32[20] , \ScanLink24[22] , \ScanLink48[3] , 
        \Level8Out16[12] , \ScanLink31[16] , \ScanLink51[12] , \ScanLink34[5] , 
        \ScanLink44[26] , \Level4Load12[0] , \ScanLink0[29] , \ScanLink4[18] , 
        \Level1Out4[3] , \Level1Out7[0] , \Level1Out9[15] , \ScanLink37[6] , 
        \Level1Load49[0] , \Level4Out0[22] , \Level1Out53[30] , 
        \ScanLink12[14] , \Level1Out26[19] , \Level1Out53[29] , 
        \ScanLink31[25] , \ScanLink44[15] , \Level1Out12[8] , \ScanLink24[11] , 
        \ScanLink50[1] , \ScanLink51[21] , \ScanLink53[2] , \Level4Out0[11] , 
        \Level4Out4[20] , \Level1Out22[31] , \Level2Out42[1] , 
        \Level1Out22[28] , \Level1Out57[18] , \ScanLink16[25] , 
        \ScanLink35[14] , \ScanLink40[24] , \Level2Out28[22] , 
        \ScanLink20[20] , \Level1Out28[2] , \ScanLink63[15] , 
        \Level2Out48[26] , \ScanLink55[10] , \Level2Out26[5] , 
        \Level4Out4[13] , \Level1Out6[31] , \Level1Out6[28] , \ScanLink10[3] , 
        \ScanLink13[0] , \ScanLink55[23] , \Level2Out6[7] , \Level2Out48[15] , 
        \Level1Load11[0] , \ScanLink16[16] , \ScanLink20[13] , 
        \ScanLink35[27] , \ScanLink40[17] , \Level2Out28[11] , 
        \ScanLink63[26] , \Level2Out38[9] , \Level1Out30[0] , \Level1Out51[9] , 
        \Level1Out33[3] , \Level2Out36[30] , \Level8Out24[26] , 
        \Level2Out36[29] , \Level2Out60[28] , \Level2Out60[31] , 
        \Level1Out49[13] , \Level1Out29[17] , \Level1Out54[4] , 
        \Level8Out24[15] , \Level2Out0[9] , \ScanLink7[4] , \Level1Out29[24] , 
        \Level1Out39[26] , \Level1Out49[20] , \Level1Out57[7] , 
        \Level4Out16[6] , \Level1Out59[22] , \Level1Out39[15] , 
        \Level1Out60[5] , \Level1Out63[6] , \Level2Out2[26] , 
        \Level2Out26[18] , \Level4Out36[18] , \Level4Out60[19] , 
        \ScanLink46[8] , \Level2Out2[15] , \Level1Out59[11] , \ScanLink4[7] , 
        \ScanLink58[4] , \ScanLink0[17] , \ScanEnable[0] , \ScanLink2[9] , 
        \Level1Out8[21] , \Level1Out11[31] , \ScanLink13[20] , \ScanLink24[2] , 
        \ScanLink25[25] , \Level8Out8[14] , \ScanLink30[11] , \ScanLink50[15] , 
        \Level2Out38[13] , \ScanLink45[21] , \Level2Out58[17] , 
        \Level1Out32[19] , \Level1Out11[28] , \Level1Out47[29] , 
        \Level1Out47[30] , \Level1Out8[12] , \ScanLink27[1] , \Level2Out12[4] , 
        \Level4Out24[9] , \Level4Out28[13] , \Level4Out48[17] , 
        \ScanLink13[13] , \ScanLink30[22] , \ScanLink45[12] , 
        \Level2Out58[24] , \Level16Out0[2] , \ScanLink25[16] , \ScanLink40[6] , 
        \ScanLink50[26] , \Level2Out38[20] , \Level8Out8[27] , \ScanLink43[5] , 
        \ScanLink4[26] , \ScanLink4[15] , \Level1Out14[13] , \Level1Out15[19] , 
        \ScanLink17[22] , \Level1Out26[9] , \Level2Load52[0] , 
        \Level2Out52[6] , \Level4Out28[20] , \Level4Out48[24] , 
        \ScanLink34[13] , \ScanLink41[23] , \ScanLink64[0] , \ScanLink17[11] , 
        \ScanLink21[27] , \Level1Out38[5] , \ScanLink62[12] , \ScanLink21[14] , 
        \ScanLink54[24] , \ScanLink54[17] , \Level2Out36[2] , \ScanLink34[20] , 
        \ScanLink41[10] , \ScanLink62[21] , \Level1Out36[28] , 
        \Level1Out43[18] , \Level1Out60[30] , \Level1Out60[29] , 
        \ScanLink18[6] , \Level1Out20[7] , \Level1Out36[31] , \Level2Out54[8] , 
        \Level1Out23[4] , \Level1Out28[10] , \Level1Out48[14] , 
        \Level2Out6[24] , \Level1Out28[23] , \Level1Out44[3] , 
        \Level4Out32[30] , \Level4Out32[29] , \Level1Out47[0] , 
        \Level1Out48[27] , \Level2Out6[17] , \Level2Out22[30] , 
        \Level2Out22[29] , \Level1Out61[23] , \Level1Out22[16] , 
        \Level1Out37[22] , \Level1Out42[12] , \Level1Out51[4] , 
        \Level1Out57[26] , \Level4Out4[2] , \Level2Out38[4] , 
        \Level2Out48[18] , \Level16Out32[23] , \Level1Out14[20] , 
        \ScanLink16[31] , \ScanLink16[28] , \Level1Out52[7] , \Level2Out26[8] , 
        \ScanLink35[19] , \ScanLink40[30] , \ScanLink63[18] , 
        \Level1Out22[25] , \ScanLink40[29] , \Level1Out57[15] , 
        \Level1Out35[0] , \Level1Out37[11] , \Level1Out61[10] , 
        \Level1Out42[21] , \Level1Out6[25] , \Level1Load14[0] , 
        \Level1Out36[3] , \Level16Out32[10] , \Level1Out29[30] , 
        \Level1Out29[29] , \Level2Out36[17] , \Level2Out56[13] , 
        \Level2Out60[16] , \ScanLink15[3] , \ScanLink16[0] , \Level1Out49[6] , 
        \Level1Out1[3] , \Level1Out2[0] , \Level1Out6[16] , \Level1Out54[9] , 
        \Level2Out0[4] , \Level2Out20[6] , \Level8Out24[18] , 
        \Level2Out36[24] , \Level2Out60[25] , \Level2Out56[20] , 
        \Level1Out2[27] , \ScanLink9[2] , \Level2Out44[2] , \Level2Out60[4] , 
        \ScanLink55[1] , \Level4Out48[5] , \Level1Out2[14] , \Level1Out17[8] , 
        \ScanLink56[2] , \Level2Out32[15] , \ScanLink19[26] , \Level4Out56[9] , 
        \ScanLink19[15] , \ScanLink31[5] , \Level2Load20[0] , 
        \Level2Out52[11] , \Level1Out58[31] , \Level1Out58[28] , 
        \Level2Out32[26] , \Level2Out52[22] , \Level1Out12[5] , 
        \ScanLink32[6] , \ScanLink12[19] , \ScanLink31[31] , \ScanLink31[28] , 
        \ScanLink44[18] , \Level1Out53[24] , \ScanLink0[24] , \Level1Out9[18] , 
        \Level1Out11[6] , \Level1Out26[14] , \Level1Out10[11] , 
        \Level2Out8[20] , \Level1Out33[20] , \Level1Out46[10] , 
        \Level1Out10[22] , \Level8Out8[2] , \Level1Out26[27] , 
        \Level1Out33[13] , \Level2Out8[13] , \Level1Out46[23] , 
        \Level1Load2[0] , \Level1Out2[9] , \ScanLink29[7] , \Level1Out53[17] , 
        \Level1Out29[13] , \ScanLink34[8] , \Level1Out33[7] , 
        \Level1Out49[17] , \Level2Out56[30] , \Level1Out30[4] , 
        \Level2Out56[29] , \Level8Out24[22] , \Level1Out4[7] , 
        \Level1Out14[29] , \ScanLink16[21] , \ScanLink16[9] , 
        \Level1Out29[20] , \Level1Out49[24] , \Level1Out57[3] , 
        \Level4Out16[2] , \ScanLink20[24] , \Level1Out54[0] , 
        \Level2Out48[22] , \Level8Out24[11] , \Level1Out28[6] , 
        \ScanLink55[14] , \ScanLink35[10] , \ScanLink63[11] , \ScanLink40[20] , 
        \Level2Out28[26] , \Level1Out7[4] , \Level1Out14[30] , 
        \Level1Out37[18] , \Level1Out42[31] , \Level1Out61[19] , 
        \Level1Out35[9] , \Level1Out42[28] , \Level2Out42[5] , 
        \Level16Out32[19] , \ScanLink10[7] , \ScanLink16[12] , 
        \ScanLink63[22] , \Level4Out4[24] , \ScanLink35[23] , \ScanLink40[13] , 
        \Level2Out28[15] , \ScanLink55[27] , \Level2Out48[11] , 
        \ScanLink13[4] , \ScanLink20[17] , \Level2Out6[3] , \Level4Out4[17] , 
        \ScanLink37[2] , \Level2Out26[1] , \Level4Out0[26] , \ScanLink1[27] , 
        \ScanLink1[14] , \ScanLink1[3] , \Level1Out9[22] , \Level1Out9[11] , 
        \Level1Out10[18] , \ScanLink12[23] , \ScanLink12[10] , 
        \ScanLink24[26] , \ScanLink31[12] , \ScanLink34[1] , \ScanLink44[22] , 
        \ScanLink24[15] , \ScanLink50[5] , \ScanLink51[25] , \ScanLink51[16] , 
        \ScanLink53[6] , \Level4Out0[15] , \ScanLink31[21] , \ScanLink44[11] , 
        \Level1Out33[30] , \Level1Out33[29] , \Level1Out46[19] , 
        \Level2Out8[29] , \Level2Out8[30] , \Level1Out11[12] , 
        \Level1Out14[2] , \Level1Out38[25] , \Level4Out32[4] , 
        \Level8Out16[25] , \Level16Out48[14] , \Level32Out32[17] , 
        \Level8Out40[24] , \ScanLink48[7] , \Level1Out58[21] , 
        \Level4Load0[0] , \Level8Out16[16] , \Level1Out17[1] , 
        \Level1Out38[16] , \ScanLink55[8] , \Level8Out40[17] , 
        \Level1Out58[12] , \Level16Out48[27] , \Level32Out32[24] , 
        \Level2Out52[18] , \Level4Out56[0] , \Level1Out32[23] , 
        \Level1Out47[13] , \Level4Out40[4] , \Level32Out32[7] , 
        \Level1Out27[17] , \Level1Out52[27] , \Level2Out38[30] , 
        \ScanLink2[0] , \Level2Out38[29] , \Level4Out28[30] , 
        \Level4Out28[29] , \Level1Out8[31] , \Level1Out8[28] , 
        \ScanLink13[30] , \ScanLink30[18] , \ScanLink13[29] , \ScanLink45[28] , 
        \ScanLink45[31] , \Level1Out27[24] , \ScanLink39[4] , 
        \Level1Out11[21] , \Level1Out32[10] , \Level1Out52[14] , 
        \Level4Out24[0] , \Level1Out47[20] , \Level1Out3[24] , 
        \ScanLink18[25] , \ScanLink27[8] , \Level2Out26[22] , 
        \Level2Out10[27] , \Level2Out46[26] , \ScanLink46[1] , 
        \Level1Out59[18] , \ScanLink1[25] , \ScanLink1[16] , \Level1Out3[17] , 
        \Level1Out19[7] , \ScanLink45[2] , \Level4Out36[22] , 
        \Level4Out60[23] , \Level4Out56[26] , \Level32Out0[25] , 
        \ScanLink22[5] , \ScanLink5[25] , \ScanLink5[16] , \Level1Out7[26] , 
        \ScanLink18[16] , \Level2Out10[14] , \Level8Out0[3] , 
        \Level2Out26[11] , \Level2Out46[15] , \ScanLink21[6] , 
        \Level2Out14[3] , \Level1Out59[5] , \Level2Out30[5] , 
        \Level4Out36[11] , \Level4Out56[15] , \Level32Out0[16] , 
        \Level4Out60[10] , \Level4Out52[24] , \Level4Out32[20] , 
        \Level1Out7[15] , \Level1Out47[9] , \Level2Out14[25] , \ScanLink61[4] , 
        \Level2Out22[20] , \Level2Out42[24] , \Level4Out32[13] , 
        \Level2Out14[16] , \Level2Out22[13] , \Level2Out54[1] , 
        \Level4Out52[17] , \Level2Out42[17] , \Level1Out28[19] , 
        \Level1Out42[4] , \ScanLink62[7] , \Level1Out15[10] , \ScanLink17[18] , 
        \ScanLink34[29] , \ScanLink41[19] , \ScanLink62[31] , \ScanLink62[28] , 
        \Level2Out28[7] , \Level1Out23[15] , \ScanLink34[30] , 
        \Level1Out41[7] , \Level1Out56[25] , \Level2Out8[5] , 
        \Level1Out36[21] , \Level1Out43[11] , \Level1Out60[20] , 
        \Level1Out9[2] , \Level1Out15[23] , \Level1Out25[3] , \Level1Out26[0] , 
        \Level1Out36[12] , \Level1Out43[22] , \Level1Out23[26] , 
        \Level1Out60[13] , \Level1Out56[16] , \ScanLink64[9] , \ScanLink1[1] , 
        \ScanLink2[2] , \ScanLink13[18] , \ScanLink30[30] , \ScanLink30[29] , 
        \ScanLink45[19] , \Level16Out0[9] , \Level1Out8[19] , 
        \Level1Out11[10] , \Level1Out27[15] , \Level1Out32[21] , 
        \Level1Out52[25] , \Level1Out47[11] , \Level32Out32[5] , 
        \Level4Out40[6] , \Level4Out28[18] , \Level1Out1[8] , \Level1Out3[26] , 
        \Level1Out11[23] , \Level1Out32[12] , \Level1Out47[22] , 
        \Level1Out19[5] , \ScanLink24[9] , \Level1Out27[26] , \ScanLink39[6] , 
        \Level1Out52[16] , \Level4Out24[2] , \Level2Out38[18] , 
        \Level1Load47[0] , \Level4Out56[24] , \Level32Out0[27] , 
        \ScanLink45[0] , \Level4Out36[20] , \ScanLink46[3] , \Level4Out60[21] , 
        \Level1Out3[15] , \ScanLink18[27] , \Level2Out10[25] , 
        \Level2Out26[20] , \Level2Out46[24] , \ScanLink18[14] , 
        \ScanLink21[4] , \Level4Out36[13] , \Level4Out60[12] , 
        \Level2Out14[1] , \Level4Out56[17] , \Level32Out0[14] , 
        \Level2Out26[13] , \Level2Out10[16] , \Level2Out46[17] , 
        \ScanLink5[27] , \ScanLink5[14] , \Level1Out7[24] , \ScanLink22[7] , 
        \Level1Out59[30] , \Level1Out59[29] , \Level8Out0[1] , 
        \Level2Out14[27] , \Level2Out22[22] , \Level2Out42[26] , 
        \Level1Out7[17] , \Level1Out28[31] , \Level1Out28[28] , 
        \Level1Out44[8] , \Level1Out59[7] , \Level4Out32[22] , 
        \Level4Out52[26] , \ScanLink62[5] , \Level2Out30[7] , 
        \Level1Out15[12] , \Level1Out36[23] , \ScanLink61[6] , 
        \Level2Out14[14] , \Level2Out22[11] , \Level2Out42[15] , 
        \Level4Load44[0] , \Level2Out54[3] , \Level4Out32[11] , 
        \Level4Out52[15] , \Level1Out43[13] , \Level1Out23[17] , 
        \Level1Out41[5] , \Level1Out60[22] , \Level2Out8[7] , 
        \Level1Out56[27] , \Level2Out28[5] , \Level1Out9[0] , \ScanLink17[30] , 
        \ScanLink41[28] , \Level1Out42[6] , \Level2Out36[9] , \ScanLink17[29] , 
        \ScanLink34[18] , \ScanLink41[31] , \ScanLink62[19] , 
        \Level1Out15[21] , \Level1Out23[24] , \Level1Out56[14] , 
        \Level1Out25[1] , \Level1Out43[20] , \Level1Out36[10] , 
        \Level1Out60[11] , \Level1Out26[2] , \Level8Out24[20] , 
        \Level1Out4[5] , \Level1Out7[6] , \ScanLink15[8] , \Level1Out29[11] , 
        \Level1Out30[6] , \Level1Out33[5] , \Level2Out44[9] , 
        \Level1Out49[15] , \Level1Out54[2] , \Level8Out24[13] , 
        \Level1Out29[22] , \Level1Out36[8] , \Level1Out49[26] , 
        \Level1Out57[1] , \Level2Out56[18] , \Level4Out16[0] , 
        \Level4Out4[26] , \Level2Out42[7] , \Level1Out9[20] , \ScanLink10[5] , 
        \ScanLink13[6] , \ScanLink16[23] , \ScanLink63[13] , \ScanLink20[26] , 
        \ScanLink35[12] , \ScanLink40[22] , \Level2Out28[24] , 
        \ScanLink55[16] , \Level2Out48[20] , \Level1Out28[4] , 
        \Level2Out26[3] , \Level16Out32[31] , \Level16Out32[28] , 
        \Level2Out6[1] , \Level4Out4[15] , \Level1Out10[30] , 
        \Level1Out10[29] , \ScanLink12[21] , \Level1Out14[18] , 
        \ScanLink16[10] , \ScanLink20[15] , \Level2Out48[13] , 
        \ScanLink55[25] , \ScanLink35[21] , \ScanLink63[20] , 
        \Level1Out37[30] , \ScanLink40[11] , \Level2Out28[17] , 
        \ScanLink24[24] , \Level1Out37[29] , \Level1Out61[28] , 
        \Level4Load36[0] , \Level1Out42[19] , \Level1Out61[31] , 
        \ScanLink51[14] , \Level4Out4[9] , \ScanLink31[10] , \ScanLink34[3] , 
        \ScanLink44[20] , \Level1Out46[31] , \Level1Out46[28] , 
        \Level2Out8[18] , \Level1Out33[18] , \ScanLink37[0] , \Level4Out0[24] , 
        \Level8Out8[9] , \Level1Out9[13] , \Level1Out1[1] , \ScanLink4[24] , 
        \ScanLink4[17] , \ScanLink9[9] , \ScanLink12[12] , \Level1Out14[0] , 
        \Level1Out17[3] , \ScanLink24[17] , \ScanLink31[23] , \ScanLink44[13] , 
        \ScanLink50[7] , \Level1Out38[27] , \ScanLink51[27] , \ScanLink53[4] , 
        \Level1Out58[23] , \Level4Out0[17] , \Level2Out52[30] , 
        \Level2Out52[29] , \Level4Out32[6] , \Level8Out16[27] , 
        \Level8Out40[26] , \Level16Out48[16] , \Level32Out32[15] , 
        \Level1Load35[0] , \Level1Out38[14] , \Level4Out56[2] , 
        \ScanLink56[9] , \Level1Out58[10] , \Level16Out48[25] , 
        \Level32Out32[26] , \ScanLink48[5] , \Level8Out16[14] , 
        \Level8Out40[15] , \Level1Out52[5] , \Level1Out14[11] , 
        \ScanLink16[19] , \ScanLink35[31] , \Level2Out6[8] , 
        \Level16Out32[21] , \Level1Out22[14] , \ScanLink35[28] , 
        \ScanLink63[29] , \Level2Out38[6] , \ScanLink40[18] , \ScanLink63[30] , 
        \Level1Out51[6] , \Level1Out57[24] , \Level4Out4[0] , \Level1Out36[1] , 
        \Level1Out37[20] , \Level1Out61[21] , \Level1Out42[10] , 
        \Level16Out32[12] , \Level1Out6[27] , \Level1Out14[22] , 
        \Level1Out61[12] , \ScanLink15[1] , \Level1Out22[27] , 
        \Level1Out35[2] , \Level1Out42[23] , \Level1Out37[13] , 
        \Level1Out57[17] , \Level1Out49[4] , \Level2Out20[4] , 
        \Level2Out48[30] , \Level2Out48[29] , \Level2Out0[6] , \ScanLink16[2] , 
        \Level1Out57[8] , \Level2Out36[15] , \Level2Out56[11] , 
        \Level2Out60[14] , \Level4Out16[9] , \Level2Load60[0] , 
        \Level8Out24[29] , \Level1Out2[25] , \Level1Out2[2] , \Level2Out44[0] , 
        \Level8Out24[30] , \Level2Out56[22] , \Level1Out6[14] , 
        \Level1Out29[18] , \Level2Out36[26] , \Level2Out60[27] , 
        \ScanLink19[24] , \ScanLink56[0] , \Level1Out58[19] , 
        \Level2Out32[17] , \Level2Out52[13] , \Level1Out2[16] , \ScanLink9[0] , 
        \ScanLink55[3] , \Level4Out48[7] , \Level1Out14[9] , \ScanLink32[4] , 
        \Level2Out60[6] , \Level1Out10[13] , \ScanLink19[17] , 
        \Level2Out32[24] , \ScanLink31[7] , \Level2Out52[20] , 
        \Level1Out11[4] , \Level1Out33[22] , \Level2Out8[22] , 
        \Level1Out46[12] , \Level1Out26[16] , \ScanLink0[15] , 
        \Level1Out53[26] , \ScanLink12[31] , \ScanLink12[28] , 
        \Level1Out12[7] , \ScanLink44[30] , \ScanLink44[29] , \ScanLink31[19] , 
        \Level1Out53[15] , \Level8Load32[0] , \ScanLink0[26] , 
        \Level1Out9[30] , \Level2Load38[0] , \Level1Out9[29] , 
        \Level1Out26[25] , \ScanLink29[5] , \Level1Out10[20] , 
        \Level2Out8[11] , \Level1Out33[11] , \Level1Out46[21] , 
        \Level8Out8[0] , \ScanLink37[9] , \Level1Out39[24] , \Level1Load54[0] , 
        \Level1Out60[7] , \Level1Out63[4] , \Level2Out14[8] , \ScanLink58[6] , 
        \Level1Out59[20] , \Level2Out2[24] , \Level8Out0[8] , 
        \Level4Out60[31] , \ScanLink0[18] , \ScanLink1[8] , \ScanLink4[5] , 
        \ScanLink7[6] , \Level1Load26[0] , \ScanLink45[9] , \Level4Out36[29] , 
        \Level4Out60[28] , \Level1Out59[13] , \Level4Out36[30] , 
        \Level1Out8[23] , \ScanLink27[3] , \Level1Out39[17] , \Level2Out2[17] , 
        \Level8Load40[0] , \Level2Out26[30] , \Level2Out26[29] , 
        \Level2Out12[6] , \Level4Out28[11] , \Level4Out48[15] , 
        \ScanLink13[22] , \ScanLink24[0] , \ScanLink45[23] , \ScanLink30[13] , 
        \Level2Out58[15] , \ScanLink25[27] , \ScanLink50[17] , 
        \Level2Out38[11] , \Level8Out8[16] , \ScanLink43[7] , 
        \Level4Out28[22] , \Level4Out48[26] , \Level1Out2[31] , 
        \Level1Out2[28] , \Level1Out8[10] , \Level1Out11[19] , 
        \ScanLink13[11] , \ScanLink25[14] , \ScanLink40[4] , \Level8Out8[25] , 
        \ScanLink30[20] , \ScanLink50[24] , \Level2Out38[22] , 
        \Level16Out0[0] , \ScanLink45[10] , \Level2Out58[26] , 
        \Level1Out32[31] , \Level1Out32[28] , \Level1Out47[18] , 
        \Level1Load9[0] , \Level1Out9[9] , \Level1Out38[7] , \ScanLink54[15] , 
        \Level1Out15[31] , \ScanLink17[20] , \ScanLink21[25] , 
        \ScanLink34[11] , \ScanLink41[21] , \ScanLink64[2] , \ScanLink62[10] , 
        \Level1Out25[8] , \Level1Out43[29] , \Level1Out15[28] , 
        \Level1Out36[19] , \Level1Out43[30] , \Level1Out60[18] , 
        \ScanLink17[13] , \ScanLink34[22] , \Level2Out52[4] , \ScanLink41[12] , 
        \ScanLink62[23] , \Level1Out14[4] , \ScanLink18[4] , \Level1Out20[5] , 
        \ScanLink21[16] , \Level1Out23[6] , \Level1Out28[12] , 
        \ScanLink54[26] , \Level2Load12[0] , \Level2Out36[0] , 
        \Level1Out48[16] , \Level2Out6[26] , \Level2Out22[18] , 
        \Level1Out28[21] , \Level1Out47[2] , \Level4Out32[18] , 
        \Level1Out48[25] , \Level2Out6[15] , \Level1Out44[1] , \ScanLink32[9] , 
        \Level1Out38[23] , \Level2Out32[30] , \Level8Out16[23] , 
        \Level8Out40[22] , \Level16Out48[12] , \Level32Out32[11] , 
        \Level2Out32[29] , \Level4Out32[2] , \ScanLink48[1] , 
        \Level1Load51[0] , \Level1Out58[27] , \Level8Out16[10] , 
        \Level8Out40[11] , \Level16Out48[21] , \Level32Out32[22] , 
        \Level1Out58[14] , \Level1Out9[24] , \Level1Out17[7] , 
        \ScanLink19[30] , \Level1Out38[10] , \ScanLink19[29] , 
        \Level4Out56[6] , \Level1Out26[31] , \ScanLink29[8] , \ScanLink37[4] , 
        \Level4Out0[20] , \ScanLink12[25] , \Level1Out26[28] , 
        \Level1Out53[18] , \ScanLink31[14] , \ScanLink34[7] , \ScanLink44[24] , 
        \ScanLink24[20] , \ScanLink51[10] , \ScanLink4[30] , \Level1Out4[1] , 
        \Level1Out9[17] , \ScanLink12[16] , \ScanLink24[13] , \ScanLink50[3] , 
        \ScanLink53[0] , \Level4Out0[13] , \ScanLink31[27] , \ScanLink51[23] , 
        \ScanLink44[17] , \Level1Out11[9] , \ScanLink16[27] , \ScanLink20[22] , 
        \Level1Out28[0] , \ScanLink55[12] , \Level2Out48[24] , 
        \ScanLink35[16] , \ScanLink40[26] , \Level2Out28[20] , 
        \ScanLink63[17] , \Level1Out7[2] , \Level4Load52[0] , \ScanLink4[29] , 
        \Level2Out42[3] , \ScanLink10[1] , \ScanLink16[14] , \Level1Out22[19] , 
        \Level1Out57[30] , \Level4Out4[22] , \ScanLink35[25] , 
        \Level1Out57[29] , \ScanLink40[15] , \Level2Out28[13] , 
        \ScanLink63[24] , \ScanLink13[2] , \ScanLink20[11] , \Level2Out48[17] , 
        \ScanLink55[21] , \Level2Out6[5] , \ScanLink1[31] , \ScanLink1[28] , 
        \ScanLink1[21] , \ScanLink1[12] , \ScanLink1[5] , \Level1Out3[22] , 
        \ScanLink5[23] , \ScanLink5[10] , \Level1Out6[19] , \Level1Out52[8] , 
        \Level4Out4[11] , \Level2Out26[7] , \Level1Out29[26] , 
        \Level1Out29[15] , \Level1Out30[2] , \Level1Out33[1] , 
        \Level1Out49[11] , \Level1Out49[22] , \Level1Out57[5] , 
        \Level8Out24[24] , \Level2Out36[18] , \Level2Out60[19] , 
        \Level4Out16[4] , \Level1Out42[2] , \Level1Out49[9] , \Level1Out54[6] , 
        \Level2Out20[9] , \Level8Out24[17] , \Level1Out15[16] , 
        \Level1Out23[13] , \Level1Out41[1] , \Level2Out28[1] , 
        \Level1Out56[23] , \Level2Out8[3] , \Level1Out26[6] , 
        \Level1Out36[27] , \Level1Out60[26] , \Level1Out43[17] , 
        \Level2Out52[9] , \Level1Out7[20] , \Level1Out9[4] , \Level1Out15[25] , 
        \Level1Out60[15] , \Level1Out23[20] , \Level1Out25[5] , 
        \Level1Out43[24] , \Level1Out36[14] , \Level1Out56[10] , 
        \ScanLink54[18] , \ScanLink18[9] , \ScanLink21[31] , \ScanLink21[28] , 
        \Level2Out30[3] , \Level1Out48[31] , \Level1Out59[3] , 
        \Level4Out52[22] , \Level4Out32[26] , \Level1Out48[28] , 
        \Level2Out6[18] , \Level1Out7[13] , \Level1Out20[8] , \ScanLink61[2] , 
        \Level2Out14[23] , \Level2Out42[22] , \Level2Out22[26] , 
        \Level4Load20[0] , \Level4Out32[15] , \Level4Out52[11] , 
        \Level2Out14[10] , \Level2Out22[15] , \Level2Out54[7] , 
        \Level2Out42[11] , \ScanLink18[23] , \ScanLink62[1] , \ScanLink46[7] , 
        \Level2Out10[21] , \Level2Out26[24] , \Level2Out46[20] , 
        \Level1Out3[11] , \ScanLink4[8] , \ScanLink45[4] , \Level4Out36[24] , 
        \Level4Out60[25] , \Level1Out19[1] , \Level4Out56[20] , 
        \ScanLink22[3] , \Level1Out39[30] , \Level32Out0[23] , 
        \Level2Out2[29] , \Level1Out39[29] , \Level2Out2[30] , \Level8Out0[5] , 
        \Level1Out11[14] , \ScanLink18[10] , \Level2Out10[12] , 
        \Level2Out46[13] , \ScanLink21[0] , \Level1Out63[9] , \Level2Out14[5] , 
        \Level2Out26[17] , \Level4Out56[13] , \Level4Out36[17] , 
        \Level4Out60[16] , \Level32Out0[10] , \Level1Load23[0] , 
        \ScanLink25[19] , \Level1Out27[11] , \Level1Out32[25] , 
        \Level1Out47[15] , \Level32Out32[1] , \Level4Out40[2] , 
        \ScanLink40[9] , \Level1Out52[21] , \ScanLink50[29] , \Level8Out8[31] , 
        \ScanLink2[6] , \ScanLink50[30] , \Level8Out8[28] , \Level1Out11[27] , 
        \Level1Out27[22] , \Level1Out52[12] , \Level2Out58[18] , 
        \Level4Out24[6] , \ScanLink39[2] , \Level1Out32[16] , 
        \Level1Out47[26] , \Level4Out48[18] , \ScanLink5[19] , 
        \Level1Out7[30] , \ScanLink18[0] , \Level1Out20[1] , \Level4Out52[18] , 
        \Level1Out23[2] , \Level2Out14[19] , \Level2Out42[18] , 
        \Level1Out28[16] , \Level1Out48[12] , \ScanLink62[8] , 
        \Level2Out6[22] , \Level1Out28[25] , \Level1Out44[5] , 
        \Level1Out7[29] , \ScanLink17[24] , \Level1Out23[30] , 
        \Level1Out23[29] , \Level1Out47[6] , \Level1Out48[21] , 
        \Level2Out6[11] , \Level1Out56[19] , \Level2Out52[0] , 
        \ScanLink62[14] , \Level2Load4[0] , \ScanLink21[21] , \ScanLink34[15] , 
        \ScanLink41[25] , \ScanLink64[6] , \ScanLink54[11] , \Level1Out38[3] , 
        \Level1Out8[27] , \ScanLink13[26] , \ScanLink17[17] , \ScanLink21[12] , 
        \Level2Out36[4] , \ScanLink54[22] , \ScanLink25[23] , \ScanLink34[26] , 
        \ScanLink62[27] , \Level2Out28[8] , \ScanLink41[16] , \Level1Out41[8] , 
        \ScanLink50[13] , \Level2Out38[15] , \Level8Out8[12] , \ScanLink24[4] , 
        \ScanLink45[27] , \ScanLink30[17] , \Level2Out58[11] , 
        \Level2Out12[2] , \Level4Out28[15] , \Level1Out3[18] , 
        \Level1Out8[14] , \ScanLink27[7] , \Level4Out48[11] , 
        \Level1Out27[18] , \Level1Out52[28] , \ScanLink13[15] , 
        \Level1Out52[31] , \Level32Out32[8] , \ScanLink25[10] , 
        \ScanLink30[24] , \ScanLink40[0] , \ScanLink45[14] , \Level2Out58[22] , 
        \Level16Out0[4] , \ScanLink43[3] , \ScanLink50[20] , \Level2Out38[26] , 
        \Level8Out8[21] , \Level1Out59[24] , \Level4Out28[26] , 
        \Level4Out48[22] , \Level8Load24[0] , \ScanLink7[2] , \ScanLink18[19] , 
        \Level1Out39[20] , \Level2Out2[20] , \ScanLink21[9] , \Level1Out60[3] , 
        \Level1Out63[0] , \Level1Out39[13] , \Level1Load42[0] , 
        \Level32Out0[19] , \Level2Out2[13] , \Level2Out10[31] , 
        \Level2Out10[28] , \Level2Out46[29] , \Level2Out46[30] , 
        \Level1Out59[17] , \Level1Out19[8] , \Level4Out56[29] , 
        \Level4Out56[30] , \ScanLink0[11] , \ScanLink4[1] , \Level1Out12[3] , 
        \ScanLink58[2] , \Level1Out11[0] , \Level1Load30[0] , \ScanLink53[9] , 
        \Level8Load56[0] , \Level1Out26[12] , \ScanLink0[22] , 
        \Level1Out10[17] , \Level1Out33[26] , \Level1Out53[22] , 
        \Level1Out46[16] , \Level2Out8[26] , \Level4Out0[30] , 
        \Level4Out0[29] , \Level8Out8[4] , \Level1Out10[24] , 
        \Level1Out33[15] , \Level1Out46[25] , \Level2Out8[15] , 
        \ScanLink29[1] , \Level1Out53[11] , \Level1Out0[27] , \Level1Out0[14] , 
        \Level1Out0[8] , \Level1Out1[5] , \Level1Out2[21] , \ScanLink9[4] , 
        \ScanLink24[30] , \Level1Out26[21] , \ScanLink24[29] , 
        \ScanLink51[19] , \Level2Out60[2] , \Level8Out16[19] , 
        \Level8Out40[18] , \Level1Out38[19] , \ScanLink48[8] , \ScanLink55[7] , 
        \Level4Out48[3] , \Level16Out48[31] , \Level16Out48[28] , 
        \ScanLink56[4] , \Level1Out2[12] , \ScanLink19[20] , \Level2Out32[13] , 
        \Level2Out52[17] , \ScanLink19[13] , \ScanLink31[3] , 
        \Level32Out32[18] , \Level2Out52[24] , \Level2Out32[20] , 
        \Level1Out2[6] , \Level1Out6[23] , \ScanLink16[6] , \ScanLink32[0] , 
        \Level2Out36[11] , \Level2Out56[15] , \Level2Out60[10] , 
        \Level1Out6[10] , \ScanLink15[5] , \Level1Out49[18] , \Level1Out49[0] , 
        \Level2Out0[2] , \Level2Out20[0] , \Level2Out36[22] , 
        \Level2Out60[23] , \Level2Out56[26] , \Level1Out33[8] , 
        \Level2Out44[4] , \ScanLink2[24] , \ScanLink4[20] , \ScanLink4[13] , 
        \ScanLink10[8] , \Level1Out14[15] , \Level1Out37[24] , 
        \Level1Out42[14] , \Level1Out22[10] , \Level1Out51[2] , 
        \Level1Out61[25] , \ScanLink55[31] , \Level1Out57[20] , 
        \Level4Out4[4] , \ScanLink20[18] , \ScanLink55[28] , \Level2Out38[2] , 
        \Level4Out4[18] , \Level1Out4[8] , \Level1Out14[26] , 
        \Level1Out22[23] , \Level1Out28[9] , \Level1Out52[1] , 
        \Level16Out32[25] , \Level2Out28[30] , \Level2Out28[29] , 
        \Level1Out57[13] , \Level1Out35[6] , \Level1Out42[27] , 
        \Level1Out37[17] , \Level1Out61[16] , \Level1Out36[5] , 
        \Level16Out32[16] , \Level1Out56[1] , \Level8Out32[3] , 
        \ScanLink2[17] , \Level1Out12[22] , \Level1Out24[27] , 
        \Level1Out51[17] , \Level1Out31[13] , \Level1Out44[23] , 
        \Level1Out55[2] , \Level4Out0[4] , \ScanLink14[8] , \Level2Out18[31] , 
        \Level2Out18[28] , \ScanLink10[19] , \Level1Out32[5] , 
        \ScanLink33[28] , \Level8Out56[7] , \ScanLink46[18] , 
        \Level1Out12[11] , \Level1Out31[20] , \ScanLink33[31] , 
        \Level2Out58[6] , \Level1Out44[10] , \ScanLink11[5] , 
        \Level1Out24[14] , \Level1Out31[6] , \Level1Out51[24] , 
        \ScanLink12[6] , \ScanLink38[24] , \ScanLink58[20] , \Level2Out4[2] , 
        \Level4Out16[23] , \Level4Out20[26] , \Level4Out40[22] , 
        \Level2Out24[0] , \Level8Out0[21] , \Level2Out30[26] , 
        \Level2Out50[22] , \Level1Out5[5] , \ScanLink9[31] , \Level2Out40[4] , 
        \Level4Out16[10] , \Level4Out40[11] , \ScanLink9[28] , 
        \Level1Out29[4] , \Level4Out20[15] , \Level1Out4[25] , 
        \Level1Out4[16] , \Level1Out6[6] , \Level1Out37[8] , \ScanLink38[17] , 
        \Level2Out50[11] , \Level8Out0[12] , \ScanLink58[13] , 
        \Level2Out30[15] , \ScanLink29[21] , \ScanLink29[12] , 
        \ScanLink49[16] , \ScanLink52[4] , \Level2Out54[20] , 
        \Level2Out62[25] , \ScanLink51[7] , \Level2Out34[24] , 
        \Level4Out12[21] , \Level4Out44[20] , \Level2Out34[17] , 
        \Level2Out62[16] , \Level4Out24[24] , \ScanLink36[0] , 
        \ScanLink49[25] , \Level2Out54[13] , \ScanLink6[26] , \ScanLink8[9] , 
        \ScanLink14[31] , \ScanLink35[3] , \Level4Out24[17] , \Level4Out28[7] , 
        \Level4Out44[13] , \ScanLink37[19] , \ScanLink42[29] , 
        \Level4Out12[12] , \ScanLink14[28] , \ScanLink42[30] , 
        \ScanLink61[18] , \Level1Out15[0] , \Level1Out16[20] , 
        \Level1Out35[11] , \Level1Out40[21] , \Level1Out63[10] , 
        \Level1Out20[25] , \ScanLink49[5] , \Level1Out55[15] , 
        \Level2Load58[0] , \Level1Out16[3] , \Level1Out16[13] , 
        \Level1Out20[16] , \Level1Load34[0] , \ScanLink57[9] , 
        \Level1Out35[22] , \Level1Out55[26] , \Level1Out40[12] , 
        \Level1Out63[23] , \Level2Out18[4] , \ScanLink0[1] , \ScanLink6[15] , 
        \Level8Out16[5] , \ScanLink25[9] , \ScanLink38[6] , \Level8Out32[26] , 
        \Level1Load46[0] , \Level2Out4[17] , \Level2Out20[30] , 
        \Level16Out16[8] , \Level2Out20[29] , \ScanLink3[2] , \ScanLink28[18] , 
        \Level8Out32[15] , \Level2Out4[24] , \ScanLink15[11] , \ScanLink23[7] , 
        \Level2Out16[2] , \Level1Out17[19] , \ScanLink20[4] , \ScanLink23[14] , 
        \ScanLink36[20] , \ScanLink60[21] , \ScanLink43[10] , \ScanLink56[24] , 
        \Level1Out34[31] , \Level1Out34[28] , \Level1Out62[29] , 
        \Level1Out41[18] , \ScanLink47[3] , \Level1Out62[30] , 
        \ScanLink15[22] , \Level1Out18[5] , \ScanLink23[27] , \ScanLink56[17] , 
        \ScanLink60[12] , \ScanLink36[13] , \ScanLink43[23] , \ScanLink44[0] , 
        \Level2Load0[0] , \ScanLink11[20] , \ScanLink11[13] , \ScanLink27[16] , 
        \ScanLink52[26] , \ScanLink60[6] , \ScanLink32[22] , \ScanLink64[23] , 
        \ScanLink47[12] , \ScanLink63[5] , \ScanLink64[10] , \Level2Out56[0] , 
        \ScanLink27[25] , \ScanLink32[11] , \ScanLink47[21] , \ScanLink52[15] , 
        \Level1Out58[7] , \ScanLink0[8] , \ScanLink5[5] , \ScanLink6[6] , 
        \ScanLink8[22] , \Level1Out13[31] , \Level1Out13[28] , 
        \Level1Out45[30] , \Level1Out30[19] , \Level1Out45[29] , 
        \Level1Out45[8] , \Level1Out18[24] , \Level1Out27[2] , 
        \ScanLink59[19] , \Level2Out32[4] , \Level16Out16[30] , 
        \Level8Out48[18] , \Level16Out16[29] , \Level2Out0[15] , 
        \ScanLink8[11] , \Level1Out8[0] , \Level8Out40[3] , \Level16Out48[6] , 
        \Level1Out18[17] , \Level1Out24[1] , \Level4Out8[30] , 
        \Level8Out56[20] , \Level4Out8[29] , \Level1Out40[5] , 
        \Level1Out43[6] , \Level2Out0[26] , \Level2Out24[18] , 
        \Level8Out56[13] , \Level8Out24[7] , \ScanLink7[25] , 
        \Level1Out17[23] , \Level1Out21[26] , \Level1Out54[16] , 
        \ScanLink59[6] , \Level4Out44[2] , \Level32Load32[0] , 
        \Level1Out62[13] , \Level1Out34[12] , \Level1Out41[22] , 
        \ScanLink7[16] , \Level1Load27[0] , \ScanLink44[9] , \ScanLink15[18] , 
        \Level1Out62[4] , \Level1Out17[10] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink60[28] , \ScanLink43[19] , \ScanLink60[31] , 
        \Level1Out21[15] , \Level1Out34[21] , \Level1Out62[20] , 
        \Level1Out41[11] , \Level4Out20[6] , \Level1Out54[25] , 
        \Level1Out61[7] , \Level1Out1[24] , \Level1Out1[17] , \Level1Out5[26] , 
        \Level1Out5[15] , \ScanLink28[11] , \ScanLink41[4] , \ScanLink42[7] , 
        \ScanLink48[15] , \Level2Out16[16] , \Level2Out40[17] , 
        \Level2Out20[13] , \ScanLink25[0] , \Level2Out10[5] , \ScanLink26[3] , 
        \ScanLink28[22] , \ScanLink48[26] , \Level2Out20[20] , 
        \Level16Out16[1] , \Level2Out16[25] , \Level2Out40[24] , 
        \ScanLink8[18] , \Level1Load8[0] , \ScanLink39[27] , \ScanLink59[23] , 
        \Level2Out24[11] , \Level2Out44[15] , \Level4Load24[0] , 
        \Level16Out32[7] , \Level2Out12[14] , \Level2Out34[3] , 
        \Level4Out8[13] , \Level4Out8[5] , \ScanLink39[14] , \ScanLink59[10] , 
        \Level2Out12[27] , \Level2Out44[26] , \Level2Out24[22] , 
        \Level1Out8[9] , \Level1Out39[7] , \ScanLink11[30] , \ScanLink11[29] , 
        \Level1Out24[8] , \ScanLink47[31] , \ScanLink64[19] , \Level2Out50[7] , 
        \Level4Out8[20] , \Level8Out56[30] , \Level8Out56[29] , 
        \ScanLink32[18] , \ScanLink47[28] , \Level1Out13[21] , \ScanLink19[4] , 
        \Level1Out25[24] , \Level1Out30[10] , \Level1Out45[20] , 
        \Level1Out45[1] , \Level1Out50[14] , \ScanLink3[27] , \Level1Out46[2] , 
        \Level1Out13[12] , \Level1Out21[5] , \Level1Out25[17] , 
        \Level8Out48[11] , \Level16Out16[20] , \Level16Out0[25] , 
        \Level1Out50[27] , \Level32Out0[4] , \Level1Out30[23] , 
        \Level1Out45[13] , \Level4Out60[4] , \Level2Out48[5] , \Level1Out0[1] , 
        \ScanLink3[14] , \Level1Out22[6] , \Level8Out48[22] , 
        \Level16Out0[16] , \Level2Out56[9] , \Level1Out3[2] , \ScanLink9[21] , 
        \Level1Out34[2] , \Level16Out16[13] , \ScanLink9[12] , 
        \Level1Out19[27] , \Level4Out16[19] , \Level4Out40[18] , 
        \Level1Out37[1] , \Level2Out50[18] , \Level1Out19[14] , 
        \Level1Out50[6] , \Level1Out53[5] , \Level2Out24[9] , \ScanLink58[30] , 
        \ScanLink58[29] , \Level4Out12[4] , \Level8Out0[28] , \Level8Out0[31] , 
        \Level2Out46[3] , \ScanLink10[10] , \ScanLink33[21] , \ScanLink46[11] , 
        \ScanLink26[15] , \Level2Out18[12] , \ScanLink53[25] , 
        \Level8Out48[2] , \Level1Out1[30] , \Level1Out1[29] , \ScanLink8[26] , 
        \ScanLink8[0] , \ScanLink10[23] , \Level1Out12[18] , \Level1Out31[29] , 
        \Level1Out44[19] , \Level4Load56[0] , \ScanLink14[1] , \ScanLink17[2] , 
        \Level1Out31[30] , \Level2Out2[5] , \ScanLink26[26] , \Level1Out48[4] , 
        \Level1Out56[8] , \Level2Out22[7] , \ScanLink53[16] , 
        \Level2Out18[21] , \ScanLink33[12] , \ScanLink46[22] , 
        \ScanLink14[21] , \ScanLink14[12] , \ScanLink22[17] , \ScanLink30[7] , 
        \ScanLink37[23] , \ScanLink57[27] , \ScanLink42[13] , \ScanLink33[4] , 
        \ScanLink61[22] , \ScanLink37[10] , \ScanLink42[20] , \ScanLink54[3] , 
        \ScanLink61[11] , \ScanLink22[24] , \ScanLink57[14] , \Level1Out8[4] , 
        \Level1Out10[4] , \Level1Out13[7] , \Level1Out15[9] , 
        \Level1Out16[30] , \Level1Out35[18] , \Level1Out40[28] , 
        \Level1Out16[29] , \Level1Out40[31] , \Level1Out63[19] , 
        \ScanLink28[5] , \ScanLink29[31] , \ScanLink57[0] , \Level2Out62[5] , 
        \Level4Out36[2] , \ScanLink29[28] , \ScanLink36[9] , \Level1Load55[0] , 
        \Level2Out54[29] , \Level4Out52[6] , \Level2Out54[30] , 
        \Level1Out24[5] , \Level4Out12[31] , \Level4Out12[28] , 
        \Level4Out44[29] , \Level4Out44[30] , \Level8Out40[7] , 
        \Level8Out56[24] , \Level16Out48[2] , \Level1Out18[20] , 
        \Level2Out0[11] , \ScanLink3[19] , \ScanLink8[15] , \Level1Out27[6] , 
        \ScanLink39[19] , \Level4Out8[8] , \Level8Out24[3] , \Level1Out18[13] , 
        \Level1Out40[1] , \Level1Out43[2] , \Level8Out56[17] , 
        \Level2Out12[19] , \Level2Out44[18] , \Level2Out0[22] , 
        \Level2Out56[4] , \ScanLink11[17] , \ScanLink32[26] , \ScanLink63[1] , 
        \ScanLink47[16] , \ScanLink27[12] , \ScanLink64[27] , \Level2Out48[8] , 
        \ScanLink52[22] , \ScanLink60[2] , \Level32Out0[9] , \ScanLink19[9] , 
        \Level1Out21[8] , \Level2Load16[0] , \Level4Out60[9] , 
        \Level2Out32[0] , \Level16Out0[31] , \Level16Out0[28] , \ScanLink0[5] , 
        \ScanLink3[6] , \ScanLink5[8] , \ScanLink11[24] , \Level1Out25[30] , 
        \Level1Out25[29] , \Level1Out50[19] , \ScanLink27[21] , 
        \ScanLink52[11] , \Level1Out58[3] , \ScanLink32[15] , \ScanLink47[25] , 
        \ScanLink64[14] , \ScanLink15[15] , \ScanLink20[0] , \Level1Out21[18] , 
        \Level1Out54[31] , \ScanLink23[10] , \Level1Out54[28] , 
        \ScanLink36[24] , \ScanLink56[20] , \ScanLink43[14] , \ScanLink23[3] , 
        \ScanLink60[25] , \ScanLink36[17] , \ScanLink43[27] , \ScanLink44[4] , 
        \Level1Out62[9] , \Level2Out16[6] , \ScanLink60[16] , \ScanLink7[31] , 
        \ScanLink15[26] , \Level1Out18[1] , \ScanLink23[23] , \ScanLink56[13] , 
        \ScanLink7[28] , \ScanLink38[2] , \ScanLink47[7] , \Level2Out4[13] , 
        \Level2Out16[31] , \Level2Out16[28] , \Level2Out40[30] , 
        \Level2Out40[29] , \Level2Out10[8] , \Level8Out32[22] , 
        \Level1Out5[18] , \Level2Out4[20] , \Level1Load22[0] , \ScanLink41[9] , 
        \ScanLink48[18] , \Level8Out32[11] , \ScanLink6[22] , \Level1Out16[7] , 
        \ScanLink6[11] , \Level1Out15[4] , \Level1Out16[24] , 
        \Level1Out20[21] , \Level1Out55[11] , \Level2Out62[8] , 
        \ScanLink49[1] , \Level1Out63[14] , \ScanLink22[30] , \ScanLink22[29] , 
        \Level1Out35[15] , \Level1Out40[25] , \ScanLink57[19] , 
        \ScanLink33[9] , \Level1Load50[0] , \Level8Out16[1] , \Level1Out0[23] , 
        \Level1Out0[10] , \Level1Out4[21] , \Level1Out4[12] , \Level1Out10[9] , 
        \Level1Out16[17] , \Level2Out18[0] , \Level1Out20[12] , 
        \Level1Out35[26] , \Level1Out63[27] , \Level1Out40[16] , 
        \ScanLink51[3] , \Level1Out55[22] , \Level4Out24[20] , 
        \Level4Out12[25] , \Level4Out44[24] , \ScanLink29[16] , 
        \ScanLink49[12] , \Level2Out34[20] , \Level2Out54[24] , 
        \Level2Out62[21] , \ScanLink52[0] , \ScanLink28[8] , \ScanLink35[7] , 
        \ScanLink36[4] , \Level4Out12[16] , \Level4Out24[13] , 
        \Level4Out28[3] , \Level4Out44[17] , \ScanLink29[25] , 
        \ScanLink49[21] , \Level2Out34[13] , \Level2Out54[17] , 
        \Level2Out62[12] , \Level1Out6[2] , \ScanLink11[1] , \ScanLink12[2] , 
        \Level1Out19[19] , \ScanLink38[20] , \Level1Out53[8] , 
        \Level2Out50[26] , \ScanLink58[24] , \Level2Out4[6] , \Level2Out24[4] , 
        \Level2Out30[22] , \Level4Out12[9] , \Level8Out0[25] , 
        \Level4Out16[27] , \Level4Out20[22] , \Level4Out40[26] , 
        \ScanLink58[17] , \Level2Out30[11] , \ScanLink38[13] , 
        \Level2Out50[15] , \Level8Out0[16] , \Level1Out0[19] , \Level1Out0[5] , 
        \ScanLink2[20] , \Level1Out5[1] , \Level1Out29[0] , \Level2Out40[0] , 
        \Level4Out16[14] , \Level4Out20[11] , \Level4Out40[15] , 
        \Level1Out12[26] , \Level1Out48[9] , \Level1Out24[23] , 
        \Level1Out31[17] , \Level1Out44[27] , \Level1Out55[6] , 
        \Level1Out51[13] , \Level4Out0[0] , \Level1Out56[5] , \ScanLink2[13] , 
        \Level1Out12[15] , \Level1Out24[10] , \Level2Out2[8] , 
        \Level8Out32[7] , \Level1Out31[2] , \Level1Out51[20] , 
        \ScanLink26[18] , \Level1Out31[24] , \Level1Out44[14] , 
        \Level2Out58[2] , \Level1Out32[1] , \ScanLink53[31] , \ScanLink53[28] , 
        \Level8Out56[3] , \Level1Out4[31] , \ScanLink28[1] , \Level1Out4[28] , 
        \ScanLink6[18] , \Level1Out10[0] , \ScanLink49[31] , \ScanLink49[28] , 
        \Level4Out36[6] , \Level4Out24[30] , \Level4Out24[29] , 
        \Level1Out13[3] , \Level1Load31[0] , \ScanLink52[9] , 
        \Level2Out34[30] , \Level2Out34[29] , \Level2Out62[31] , 
        \Level2Out62[28] , \Level4Out52[2] , \ScanLink8[4] , \ScanLink14[16] , 
        \ScanLink33[0] , \Level8Out16[8] , \ScanLink22[13] , \ScanLink37[27] , 
        \ScanLink61[26] , \Level2Out18[9] , \ScanLink42[17] , \ScanLink30[3] , 
        \Level1Out55[18] , \ScanLink57[23] , \ScanLink57[4] , \Level2Out62[1] , 
        \ScanLink14[25] , \Level1Out20[31] , \Level1Out20[28] , 
        \ScanLink49[8] , \ScanLink22[20] , \ScanLink57[10] , \ScanLink61[15] , 
        \Level1Out24[19] , \ScanLink37[14] , \ScanLink42[24] , \ScanLink54[7] , 
        \Level1Out51[29] , \Level8Out48[6] , \ScanLink2[30] , \ScanLink2[29] , 
        \Level1Out3[6] , \ScanLink10[14] , \ScanLink26[11] , \Level1Out51[30] , 
        \ScanLink53[21] , \Level2Out18[16] , \ScanLink33[25] , 
        \ScanLink46[15] , \ScanLink10[27] , \Level1Out32[8] , \Level2Out46[7] , 
        \ScanLink14[5] , \ScanLink26[22] , \ScanLink33[16] , \ScanLink46[26] , 
        \ScanLink53[12] , \Level1Out48[0] , \Level2Out18[25] , \Level4Out0[9] , 
        \Level4Load32[0] , \Level2Out22[3] , \Level1Out5[8] , \ScanLink9[25] , 
        \ScanLink17[6] , \Level1Out19[23] , \Level1Out37[5] , \Level2Out2[1] , 
        \Level2Out30[18] , \Level1Out29[9] , \Level1Out34[6] , 
        \Level4Out20[18] , \Level2Out40[9] , \Level1Out19[10] , 
        \ScanLink3[23] , \ScanLink9[16] , \ScanLink38[30] , \Level1Out53[1] , 
        \Level4Out12[0] , \ScanLink38[29] , \Level1Out50[2] , \ScanLink11[8] , 
        \Level1Out46[6] , \Level8Out48[15] , \Level16Out0[21] , 
        \Level16Out16[24] , \ScanLink3[10] , \Level1Out13[25] , 
        \ScanLink19[0] , \Level2Out32[9] , \Level1Out25[20] , 
        \Level1Out50[10] , \Level1Out30[14] , \Level1Out45[24] , 
        \Level1Out45[5] , \ScanLink27[31] , \ScanLink27[28] , \ScanLink52[18] , 
        \Level16Out16[17] , \Level1Out22[2] , \ScanLink63[8] , 
        \Level8Out48[26] , \Level1Out1[20] , \Level1Out1[13] , 
        \Level1Out13[16] , \Level1Out30[27] , \Level2Out48[1] , 
        \Level16Out0[12] , \Level1Out45[17] , \Level4Out60[0] , 
        \Level1Out21[1] , \Level1Out25[13] , \Level32Out0[0] , 
        \ScanLink39[23] , \Level1Out40[8] , \Level1Out50[23] , 
        \Level4Out8[17] , \Level4Out8[1] , \ScanLink59[27] , \Level2Out12[10] , 
        \Level2Out34[7] , \Level2Out44[11] , \Level2Out24[15] , 
        \Level16Out32[3] , \Level1Out39[3] , \Level2Out50[3] , 
        \Level4Out8[24] , \Level1Out5[11] , \Level1Out18[30] , 
        \Level1Out18[29] , \ScanLink39[10] , \Level2Out0[18] , 
        \Level2Out24[26] , \Level4Load40[0] , \ScanLink59[14] , 
        \Level2Out12[23] , \Level2Out44[22] , \ScanLink42[3] , 
        \Level2Out4[30] , \ScanLink48[11] , \Level2Out4[29] , 
        \Level2Out20[17] , \ScanLink3[21] , \ScanLink5[1] , \Level1Out5[22] , 
        \ScanLink26[7] , \ScanLink28[26] , \ScanLink28[15] , \Level2Out16[12] , 
        \ScanLink41[0] , \Level2Out40[13] , \Level8Out32[18] , 
        \Level2Out16[21] , \Level16Out16[5] , \ScanLink48[22] , 
        \Level2Out20[24] , \Level2Out40[20] , \Level1Out18[8] , 
        \ScanLink25[4] , \Level2Out10[1] , \ScanLink6[2] , \ScanLink7[21] , 
        \Level1Out17[27] , \Level1Out34[16] , \Level1Out41[26] , 
        \Level1Out62[17] , \Level1Out21[22] , \Level1Out54[12] , 
        \ScanLink59[2] , \Level4Out44[6] , \ScanLink7[12] , \Level1Out17[14] , 
        \Level1Out21[11] , \Level1Out34[25] , \Level1Out54[21] , 
        \Level1Out61[3] , \Level1Out41[15] , \Level4Out20[2] , \ScanLink20[9] , 
        \ScanLink23[19] , \ScanLink56[30] , \Level1Out62[24] , 
        \Level1Load43[0] , \ScanLink56[29] , \Level1Out62[0] , 
        \Level1Out13[27] , \Level1Out30[16] , \Level1Out58[8] , 
        \Level1Out45[26] , \Level1Out45[7] , \ScanLink19[2] , 
        \Level1Out25[22] , \Level1Out50[12] , \Level16Out16[26] , 
        \Level1Out13[14] , \Level1Out21[3] , \Level1Out25[11] , 
        \Level1Out46[4] , \Level1Out50[21] , \Level8Out48[17] , 
        \Level16Out0[23] , \Level32Out0[2] , \Level1Out30[25] , 
        \Level1Out45[15] , \Level4Out60[2] , \ScanLink27[19] , 
        \ScanLink52[30] , \Level2Out48[3] , \ScanLink52[29] , \ScanLink60[9] , 
        \Level16Out0[10] , \Level1Out1[22] , \Level1Out1[11] , \ScanLink3[12] , 
        \Level1Out22[0] , \Level8Out48[24] , \Level16Out16[15] , 
        \Level1Out18[18] , \Level2Out0[30] , \ScanLink39[21] , 
        \Level2Out0[29] , \Level2Out24[17] , \Level16Out32[1] , 
        \ScanLink39[12] , \Level1Out43[9] , \ScanLink59[25] , 
        \Level2Out12[12] , \ScanLink59[16] , \Level2Out12[21] , 
        \Level2Out34[5] , \Level2Out44[13] , \Level4Out8[15] , \Level4Out8[3] , 
        \Level8Out24[8] , \Level2Out44[20] , \Level2Out24[24] , 
        \Level1Out4[19] , \ScanLink5[3] , \Level1Out5[20] , \Level1Out5[13] , 
        \ScanLink28[17] , \Level1Out39[1] , \Level16Out48[9] , \ScanLink41[2] , 
        \Level2Out50[1] , \Level4Out8[26] , \Level8Load8[0] , 
        \Level16Load48[0] , \Level2Out16[10] , \ScanLink42[1] , 
        \ScanLink48[13] , \Level2Out20[15] , \Level2Out40[11] , 
        \ScanLink25[6] , \ScanLink38[9] , \Level2Out10[3] , \Level8Out32[29] , 
        \Level8Out32[30] , \ScanLink6[0] , \ScanLink26[5] , \ScanLink28[24] , 
        \ScanLink48[20] , \Level2Out4[18] , \Level2Out20[26] , 
        \Level2Out16[23] , \Level2Out40[22] , \Level16Out16[7] , 
        \ScanLink7[23] , \Level1Out17[25] , \Level1Out21[20] , \ScanLink59[0] , 
        \Level4Out44[4] , \Level1Out34[14] , \Level1Out54[10] , 
        \Level1Out41[24] , \Level1Out62[15] , \ScanLink7[10] , 
        \ScanLink23[31] , \ScanLink23[28] , \ScanLink56[18] , 
        \Level1Out17[16] , \ScanLink23[8] , \Level1Out62[2] , 
        \Level1Out34[27] , \Level1Out41[17] , \Level4Out20[0] , 
        \Level1Out62[26] , \Level1Out21[13] , \Level1Out54[23] , 
        \ScanLink28[3] , \Level1Out61[1] , \Level2Out34[18] , \Level4Out36[4] , 
        \Level2Out62[19] , \Level4Out24[18] , \Level4Out28[8] , 
        \Level1Out10[2] , \Level1Out13[1] , \Level4Out52[0] , \ScanLink49[19] , 
        \Level4Load4[0] , \Level1Out20[19] , \ScanLink51[8] , 
        \Level1Out55[29] , \Level1Out55[30] , \Level1Out0[31] , 
        \Level1Out0[7] , \ScanLink2[18] , \Level1Out3[4] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink8[6] , \ScanLink14[27] , \ScanLink14[14] , 
        \ScanLink22[11] , \ScanLink57[21] , \ScanLink30[1] , \ScanLink61[24] , 
        \ScanLink33[2] , \ScanLink37[25] , \ScanLink42[15] , \ScanLink22[22] , 
        \ScanLink37[16] , \ScanLink61[17] , \ScanLink42[26] , \ScanLink54[5] , 
        \ScanLink57[12] , \Level1Load29[0] , \Level2Out62[3] , \ScanLink57[6] , 
        \Level2Out46[5] , \ScanLink10[16] , \Level2Out58[9] , \Level8Out56[8] , 
        \ScanLink26[13] , \ScanLink33[27] , \ScanLink46[17] , \ScanLink53[23] , 
        \Level1Out31[9] , \Level2Out18[14] , \ScanLink9[27] , \ScanLink10[25] , 
        \ScanLink17[4] , \Level2Out2[3] , \Level8Out48[4] , \Level1Out24[31] , 
        \Level1Out24[28] , \Level2Out22[1] , \Level1Out51[18] , 
        \ScanLink26[20] , \Level1Out48[2] , \ScanLink53[10] , 
        \Level2Out18[27] , \ScanLink14[7] , \ScanLink33[14] , \Level1Out34[4] , 
        \ScanLink46[24] , \Level1Out19[21] , \Level1Out0[28] , \ScanLink6[20] , 
        \Level1Load6[0] , \Level1Out6[9] , \ScanLink9[14] , \Level1Out37[7] , 
        \ScanLink38[18] , \Level1Out50[0] , \Level4Out20[30] , 
        \Level4Out20[29] , \ScanLink12[9] , \Level1Out53[3] , 
        \Level2Out30[30] , \Level2Out30[29] , \Level4Out12[2] , 
        \Level1Out15[6] , \Level1Out16[26] , \Level1Out19[12] , 
        \Level1Out35[17] , \Level1Out63[16] , \Level1Out20[23] , 
        \Level1Out40[27] , \ScanLink49[3] , \Level1Out55[13] , 
        \Level1Out16[15] , \Level1Out16[5] , \Level1Out20[10] , 
        \Level1Out55[20] , \Level1Out63[25] , \Level1Out35[24] , 
        \Level1Out40[14] , \ScanLink57[28] , \Level2Out18[2] , 
        \Level1Out4[10] , \ScanLink6[13] , \ScanLink22[18] , \ScanLink30[8] , 
        \ScanLink57[31] , \Level8Out16[3] , \Level1Out13[8] , \ScanLink52[2] , 
        \ScanLink29[27] , \ScanLink29[14] , \ScanLink49[10] , 
        \Level2Out34[22] , \Level2Out54[26] , \ScanLink51[1] , 
        \Level2Out62[23] , \Level4Out52[9] , \Level4Out12[27] , 
        \Level4Out24[22] , \Level4Out44[26] , \Level2Out34[11] , 
        \Level2Out62[10] , \Level1Out0[21] , \Level1Out0[12] , 
        \Level1Out4[23] , \Level1Load48[0] , \Level2Out54[15] , 
        \ScanLink49[23] , \ScanLink11[3] , \ScanLink35[5] , \ScanLink36[6] , 
        \Level4Out12[14] , \Level4Out24[11] , \Level2Load24[0] , 
        \Level4Out28[1] , \Level4Out20[20] , \Level4Out44[15] , 
        \ScanLink12[0] , \ScanLink38[22] , \Level1Out50[9] , \Level2Out4[4] , 
        \Level4Out16[25] , \Level2Out24[6] , \Level4Out40[24] , 
        \ScanLink58[26] , \Level2Out30[20] , \Level2Out50[24] , 
        \Level8Out0[27] , \Level1Out5[3] , \Level2Out40[2] , \Level1Out29[2] , 
        \Level4Out16[16] , \Level4Out20[13] , \Level4Out40[17] , 
        \Level1Out1[18] , \ScanLink2[22] , \Level1Out6[0] , \Level1Out19[31] , 
        \Level1Out19[28] , \ScanLink38[11] , \Level2Out50[17] , 
        \ScanLink58[15] , \Level2Out30[13] , \Level8Out0[14] , 
        \Level8Out32[5] , \ScanLink2[11] , \Level1Out12[24] , 
        \Level1Out24[21] , \Level1Out56[7] , \Level2Out22[8] , 
        \Level1Out51[11] , \ScanLink26[30] , \ScanLink26[29] , 
        \Level1Out31[15] , \Level4Out0[2] , \Level1Out44[25] , 
        \Level1Out55[4] , \ScanLink53[19] , \ScanLink8[24] , \Level1Out8[6] , 
        \Level1Load10[0] , \Level1Out32[3] , \Level1Out12[17] , 
        \Level2Out58[0] , \Level8Out56[1] , \Level1Out18[22] , 
        \Level1Out24[12] , \Level1Out31[26] , \Level1Out44[16] , 
        \Level1Out51[22] , \Level1Out27[4] , \Level1Out31[0] , 
        \Level2Out12[28] , \Level2Out44[30] , \Level2Out12[31] , 
        \Level2Out44[29] , \Level2Out0[13] , \Level8Out40[5] , 
        \Level16Out48[0] , \Level1Out18[11] , \Level1Out24[7] , 
        \Level1Out39[8] , \Level2Out50[8] , \Level8Out56[26] , 
        \Level2Out0[20] , \ScanLink8[17] , \ScanLink39[31] , \ScanLink39[28] , 
        \Level16Out32[8] , \Level1Out43[0] , \Level1Out40[3] , 
        \Level1Load62[0] , \Level8Out56[15] , \Level1Out50[31] , 
        \Level8Out24[1] , \ScanLink11[26] , \ScanLink11[15] , 
        \Level1Out25[18] , \Level1Out50[28] , \ScanLink27[10] , 
        \ScanLink52[20] , \ScanLink32[24] , \ScanLink47[14] , \ScanLink60[0] , 
        \ScanLink64[25] , \Level1Out22[9] , \ScanLink63[3] , \Level2Out56[6] , 
        \Level16Out0[19] , \ScanLink32[17] , \ScanLink47[27] , 
        \ScanLink27[23] , \Level1Out58[1] , \ScanLink64[16] , \ScanLink52[13] , 
        \Level1Out0[3] , \ScanLink0[7] , \ScanLink3[31] , \ScanLink3[28] , 
        \Level1Out5[30] , \Level1Out5[29] , \ScanLink6[9] , \ScanLink7[19] , 
        \Level2Out16[4] , \Level2Out32[2] , \ScanLink15[17] , \ScanLink23[1] , 
        \ScanLink36[26] , \ScanLink43[16] , \ScanLink60[27] , \ScanLink20[2] , 
        \ScanLink23[12] , \ScanLink56[22] , \Level1Out61[8] , \Level4Out20[9] , 
        \ScanLink15[24] , \Level1Out18[3] , \Level1Out21[30] , \ScanLink47[5] , 
        \Level2Load56[0] , \Level1Out21[29] , \ScanLink59[9] , 
        \Level1Out54[19] , \ScanLink23[21] , \ScanLink36[15] , 
        \ScanLink56[11] , \ScanLink43[25] , \ScanLink44[6] , \ScanLink38[0] , 
        \ScanLink60[14] , \Level8Out32[20] , \Level2Out4[11] , 
        \ScanLink48[30] , \ScanLink48[29] , \ScanLink3[4] , \Level2Out16[19] , 
        \Level8Out32[13] , \Level2Out40[18] , \ScanLink9[23] , 
        \Level1Load15[0] , \Level1Out37[3] , \ScanLink42[8] , \Level2Out4[22] , 
        \Level8Out0[19] , \ScanLink58[18] , \Level1Out19[25] , \ScanLink9[10] , 
        \Level1Out19[16] , \Level1Out34[0] , \Level1Out50[4] , 
        \Level1Out53[7] , \Level2Out50[29] , \Level4Out12[6] , 
        \Level2Out50[30] , \Level2Out4[9] , \Level4Out16[31] , 
        \Level4Out40[29] , \Level4Out16[28] , \Level4Out40[30] , 
        \Level1Out1[26] , \Level1Out1[15] , \ScanLink3[9] , \Level1Out3[0] , 
        \ScanLink10[12] , \ScanLink26[17] , \ScanLink53[27] , 
        \Level2Out18[10] , \Level8Out48[0] , \ScanLink33[23] , 
        \ScanLink46[13] , \Level2Out46[1] , \ScanLink5[7] , \ScanLink8[2] , 
        \ScanLink10[21] , \ScanLink14[3] , \ScanLink33[10] , \ScanLink46[20] , 
        \Level1Out12[30] , \ScanLink26[24] , \Level1Out48[6] , 
        \Level2Out18[23] , \ScanLink53[14] , \Level1Out12[29] , 
        \Level1Out31[18] , \Level1Out44[28] , \Level1Out55[9] , 
        \ScanLink14[10] , \ScanLink17[0] , \Level1Out44[31] , \Level2Out22[5] , 
        \ScanLink33[6] , \Level2Out2[7] , \Level8Out32[8] , \ScanLink37[21] , 
        \ScanLink42[11] , \ScanLink61[20] , \Level1Out16[18] , 
        \ScanLink22[15] , \ScanLink57[25] , \ScanLink30[5] , \Level1Out35[30] , 
        \Level1Out35[29] , \Level1Out40[19] , \Level1Out63[31] , 
        \Level1Out63[28] , \Level4Load16[0] , \Level1Out16[8] , 
        \ScanLink57[2] , \Level2Out62[7] , \Level1Out10[6] , \ScanLink14[23] , 
        \ScanLink22[26] , \ScanLink37[12] , \ScanLink57[16] , \ScanLink42[22] , 
        \ScanLink54[1] , \ScanLink28[7] , \ScanLink61[13] , \ScanLink35[8] , 
        \Level4Out12[19] , \Level4Out44[18] , \Level2Out54[18] , 
        \Level4Out36[0] , \Level1Out13[5] , \ScanLink29[19] , \Level4Out52[4] , 
        \Level1Out5[17] , \ScanLink6[4] , \ScanLink7[27] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink43[31] , \ScanLink60[19] , 
        \Level1Out17[21] , \ScanLink36[18] , \ScanLink43[28] , 
        \Level1Out21[24] , \Level1Out34[10] , \Level1Out62[11] , 
        \Level1Out41[20] , \Level4Out44[0] , \Level1Out54[14] , 
        \ScanLink59[4] , \ScanLink47[8] , \ScanLink7[14] , \Level1Out17[12] , 
        \Level1Out21[17] , \Level1Out54[27] , \Level1Out61[5] , 
        \Level1Out62[22] , \Level1Out34[23] , \Level1Out41[13] , 
        \Level4Out20[4] , \Level1Out62[6] , \Level2Out16[9] , \ScanLink42[5] , 
        \Level1Out5[24] , \ScanLink28[20] , \ScanLink28[13] , \ScanLink48[17] , 
        \Level2Out20[11] , \ScanLink41[6] , \Level2Out16[14] , 
        \Level2Out40[15] , \ScanLink48[24] , \Level2Out16[27] , 
        \Level2Out40[26] , \Level16Out16[3] , \Level2Out20[22] , 
        \ScanLink25[2] , \ScanLink26[1] , \ScanLink39[25] , \ScanLink59[21] , 
        \Level2Out10[7] , \Level2Out34[1] , \Level4Out8[11] , \Level4Out8[7] , 
        \Level8Out56[18] , \Level2Out12[16] , \Level2Out44[17] , 
        \Level2Out24[13] , \Level16Out32[5] , \ScanLink8[30] , \ScanLink8[29] , 
        \Level2Out50[5] , \Level4Out8[22] , \Level1Out39[5] , \Level8Out40[8] , 
        \ScanLink3[25] , \Level1Out27[9] , \ScanLink39[16] , \ScanLink59[12] , 
        \Level2Out24[20] , \Level2Out44[24] , \Level2Out12[25] , 
        \Level8Out48[13] , \Level16Out0[27] , \ScanLink3[16] , 
        \Level1Out13[23] , \ScanLink19[6] , \Level1Out25[26] , 
        \Level1Out46[0] , \Level16Out16[22] , \Level1Out50[16] , 
        \Level1Out30[12] , \Level1Out45[22] , \Level1Out45[3] , 
        \Level1Out22[4] , \Level16Out16[11] , \Level8Out48[20] , 
        \Level16Out0[14] , \ScanLink11[18] , \ScanLink32[30] , 
        \ScanLink64[28] , \Level2Out48[7] , \Level1Out13[10] , 
        \ScanLink32[29] , \ScanLink47[19] , \ScanLink64[31] , 
        \Level1Out30[21] , \Level1Out45[11] , \Level4Out60[6] , 
        \Level1Out50[25] , \Level1Out21[7] , \Level1Out25[15] , 
        \Level32Out0[6] , \ScanLink0[3] , \ScanLink3[0] , \ScanLink26[8] , 
        \ScanLink28[30] , \ScanLink28[29] , \ScanLink38[4] , \Level2Out4[15] , 
        \Level2Out4[26] , \Level8Out32[24] , \Level2Out20[18] , 
        \Level8Out32[17] , \ScanLink15[20] , \ScanLink15[13] , \ScanLink20[6] , 
        \ScanLink23[16] , \ScanLink56[26] , \ScanLink60[23] , \ScanLink23[5] , 
        \ScanLink36[22] , \ScanLink43[12] , \Level2Load32[0] , 
        \Level2Out16[0] , \Level1Out17[31] , \Level1Out17[28] , 
        \Level1Out18[7] , \ScanLink23[25] , \ScanLink36[11] , \ScanLink60[10] , 
        \ScanLink43[21] , \ScanLink44[2] , \ScanLink56[15] , \Level4Out44[9] , 
        \Level1Out41[30] , \Level1Out62[18] , \Level1Out34[19] , 
        \Level1Out41[29] , \ScanLink47[1] , \Level2Out56[2] , 
        \Level16Out16[18] , \ScanLink11[11] , \ScanLink63[7] , 
        \Level8Out48[30] , \ScanLink64[21] , \Level8Out48[29] , 
        \ScanLink27[14] , \ScanLink32[20] , \ScanLink47[10] , \ScanLink52[24] , 
        \ScanLink60[4] , \Level1Out13[19] , \Level1Out30[31] , 
        \Level1Out30[28] , \Level1Out45[18] , \Level1Out46[9] , 
        \Level2Out32[6] , \Level1Out0[25] , \Level1Out0[16] , \ScanLink2[26] , 
        \ScanLink8[20] , \ScanLink11[22] , \ScanLink27[27] , \ScanLink52[17] , 
        \Level1Out58[5] , \Level1Out24[3] , \ScanLink32[13] , \ScanLink64[12] , 
        \ScanLink47[23] , \Level8Out56[22] , \ScanLink8[13] , \Level1Out8[2] , 
        \Level1Out18[26] , \Level8Out40[1] , \Level16Out48[4] , 
        \Level1Out27[0] , \Level2Out0[17] , \Level2Out24[30] , 
        \Level2Out24[29] , \Level8Out24[5] , \ScanLink10[31] , 
        \Level1Out18[15] , \Level1Out40[7] , \Level2Out34[8] , 
        \Level8Out56[11] , \Level1Out43[4] , \Level4Out8[18] , 
        \ScanLink59[31] , \ScanLink59[28] , \Level2Out0[24] , \ScanLink10[28] , 
        \ScanLink33[19] , \ScanLink46[29] , \Level1Out12[20] , 
        \Level1Out31[11] , \ScanLink46[30] , \Level1Out44[21] , 
        \Level1Out55[0] , \Level4Out0[6] , \Level1Out24[25] , 
        \Level1Out51[15] , \Level2Load18[0] , \ScanLink2[15] , 
        \Level1Load3[0] , \Level1Out3[9] , \Level1Out12[13] , \ScanLink17[9] , 
        \Level1Out56[3] , \Level8Out32[1] , \Level1Out24[16] , 
        \Level1Out51[26] , \Level8Out48[9] , \Level1Out31[22] , 
        \Level1Out31[4] , \Level1Out44[12] , \Level1Out32[7] , 
        \Level2Out18[19] , \Level2Out58[4] , \Level2Out46[8] , 
        \Level8Out56[5] , \ScanLink12[4] , \ScanLink38[26] , \Level2Out50[20] , 
        \ScanLink58[22] , \Level8Out0[23] , \Level2Out24[2] , 
        \Level2Out30[24] , \Level1Out6[4] , \ScanLink9[19] , \ScanLink11[7] , 
        \Level2Out4[0] , \Level4Out16[21] , \Level4Out40[20] , 
        \Level4Out20[24] , \Level8Out0[10] , \ScanLink38[15] , 
        \ScanLink58[11] , \Level2Out30[17] , \Level2Out50[13] , 
        \Level1Out4[27] , \Level1Out4[14] , \Level1Out5[7] , \Level1Out29[6] , 
        \Level4Out20[17] , \Level4Out16[12] , \Level4Out40[13] , 
        \ScanLink29[10] , \Level1Out34[9] , \Level2Out40[6] , \ScanLink51[5] , 
        \Level2Out34[26] , \Level2Load40[0] , \Level4Out24[26] , 
        \Level2Out62[27] , \Level4Out12[23] , \Level4Out44[22] , 
        \ScanLink49[14] , \ScanLink52[6] , \Level2Out54[22] , \ScanLink35[1] , 
        \Level4Out12[10] , \Level4Out28[5] , \Level4Out44[11] , 
        \Level4Out24[15] , \ScanLink6[24] , \ScanLink29[23] , \ScanLink36[2] , 
        \ScanLink49[27] , \Level2Out54[11] , \Level2Out62[14] , 
        \Level4Out36[9] , \Level2Out34[15] , \ScanLink6[17] , \Level1Out15[2] , 
        \Level1Out16[1] , \Level1Out20[27] , \ScanLink49[7] , 
        \Level1Out35[13] , \Level1Out55[17] , \Level1Out16[22] , 
        \Level1Out40[23] , \ScanLink54[8] , \Level1Out63[12] , 
        \Level8Out16[7] , \Level1Out0[2] , \Level1Out3[1] , \ScanLink14[19] , 
        \ScanLink37[31] , \ScanLink37[28] , \ScanLink42[18] , \ScanLink61[30] , 
        \ScanLink61[29] , \Level2Out18[6] , \Level1Out16[11] , 
        \Level1Out35[20] , \Level1Out40[10] , \Level1Out63[21] , 
        \Level1Out20[14] , \Level1Out55[24] , \Level2Load62[0] , 
        \Level2Out46[0] , \ScanLink3[24] , \ScanLink3[8] , \ScanLink8[3] , 
        \ScanLink9[22] , \ScanLink10[20] , \ScanLink10[13] , \Level8Out48[1] , 
        \ScanLink17[1] , \ScanLink26[16] , \ScanLink33[22] , \ScanLink46[12] , 
        \ScanLink53[26] , \Level2Out2[6] , \Level2Out18[11] , \Level2Out22[4] , 
        \Level8Out32[9] , \ScanLink26[25] , \Level1Out48[7] , \ScanLink53[15] , 
        \Level2Out18[22] , \Level1Out12[31] , \Level1Out12[28] , 
        \ScanLink14[2] , \ScanLink33[11] , \ScanLink46[21] , \Level1Out44[30] , 
        \Level1Out31[19] , \Level1Out44[29] , \Level1Out55[8] , 
        \ScanLink9[11] , \Level1Out19[24] , \Level1Out34[1] , \Level1Out37[2] , 
        \ScanLink58[19] , \Level8Out0[18] , \Level1Out50[5] , \Level2Out4[8] , 
        \Level4Out40[31] , \Level4Out16[30] , \Level4Out16[29] , 
        \Level4Out40[28] , \Level1Out10[7] , \Level1Out13[4] , 
        \Level1Out19[17] , \ScanLink28[6] , \Level1Out53[6] , 
        \Level2Out50[31] , \Level2Out50[28] , \Level2Out54[19] , 
        \Level4Out12[7] , \Level4Out36[1] , \ScanLink29[18] , \ScanLink35[9] , 
        \Level1Load56[0] , \Level4Out12[18] , \Level4Out44[19] , 
        \Level4Out52[5] , \ScanLink14[11] , \ScanLink22[14] , \ScanLink30[4] , 
        \ScanLink57[24] , \ScanLink61[21] , \Level1Out16[19] , 
        \Level1Out35[31] , \ScanLink37[20] , \ScanLink42[10] , 
        \Level1Out63[29] , \ScanLink33[7] , \Level1Out35[28] , 
        \Level1Out40[18] , \Level1Out63[30] , \ScanLink14[22] , 
        \Level1Out16[9] , \ScanLink22[27] , \ScanLink37[13] , \ScanLink61[12] , 
        \ScanLink42[23] , \ScanLink54[0] , \ScanLink57[17] , \ScanLink57[3] , 
        \Level2Out62[6] , \ScanLink41[7] , \ScanLink5[6] , \Level1Out5[25] , 
        \Level1Out5[16] , \ScanLink42[4] , \ScanLink25[3] , \ScanLink28[12] , 
        \Level2Out16[15] , \Level2Out40[14] , \ScanLink48[16] , 
        \Level2Out20[10] , \ScanLink28[21] , \ScanLink48[25] , 
        \Level2Out10[6] , \Level2Out16[26] , \Level2Out20[23] , 
        \Level2Out40[27] , \Level16Out16[2] , \ScanLink6[5] , \ScanLink7[26] , 
        \ScanLink26[0] , \ScanLink15[31] , \Level1Load24[0] , \ScanLink47[9] , 
        \ScanLink15[28] , \ScanLink36[19] , \ScanLink43[29] , \ScanLink7[15] , 
        \Level1Out17[20] , \Level1Out21[25] , \ScanLink43[30] , 
        \ScanLink59[5] , \ScanLink60[18] , \Level4Out44[1] , \Level1Out34[11] , 
        \Level1Out54[15] , \Level2Load48[0] , \Level1Out41[21] , 
        \Level1Out62[10] , \Level1Out13[22] , \Level1Out17[13] , 
        \Level1Out34[22] , \Level1Out41[12] , \Level1Out62[7] , 
        \Level2Out16[8] , \Level4Out20[5] , \Level1Out62[23] , 
        \Level1Out21[16] , \Level1Out54[26] , \Level1Out61[4] , 
        \Level1Out30[13] , \Level1Out45[23] , \Level1Out45[2] , 
        \ScanLink19[7] , \Level1Out25[27] , \Level1Out50[17] , 
        \Level8Out48[12] , \Level16Out0[26] , \Level16Out16[23] , 
        \ScanLink11[19] , \ScanLink32[31] , \ScanLink32[28] , \Level1Out46[1] , 
        \ScanLink47[18] , \ScanLink64[30] , \ScanLink64[29] , \Level2Out48[6] , 
        \Level32Out0[7] , \ScanLink3[17] , \Level1Out13[11] , \Level1Out21[6] , 
        \Level1Out50[24] , \Level1Out25[14] , \Level1Out30[20] , 
        \Level1Out45[10] , \Level4Out60[7] , \Level1Out22[5] , 
        \Level16Out16[10] , \Level16Out0[15] , \ScanLink0[2] , 
        \Level1Out1[27] , \Level1Out1[14] , \ScanLink39[24] , 
        \Level2Out24[12] , \Level8Out48[21] , \Level16Out32[4] , 
        \ScanLink59[20] , \Level2Out12[17] , \Level2Out44[16] , 
        \Level2Load10[0] , \Level4Out8[6] , \Level2Out34[0] , \Level4Out8[10] , 
        \Level8Out56[19] , \ScanLink8[31] , \Level1Out27[8] , \ScanLink39[17] , 
        \ScanLink59[13] , \Level2Out12[24] , \Level2Out44[25] , 
        \Level2Out24[21] , \Level2Out50[4] , \Level4Out8[23] , 
        \Level16Load0[0] , \ScanLink8[28] , \Level8Out40[9] , \ScanLink15[21] , 
        \ScanLink15[12] , \ScanLink23[4] , \Level1Out39[4] , \ScanLink36[23] , 
        \ScanLink43[13] , \Level2Out16[1] , \ScanLink60[22] , \Level1Out18[6] , 
        \ScanLink20[7] , \ScanLink56[27] , \ScanLink23[17] , \ScanLink47[0] , 
        \ScanLink23[24] , \ScanLink36[10] , \ScanLink56[14] , \ScanLink43[20] , 
        \ScanLink44[3] , \Level1Out17[30] , \ScanLink60[11] , 
        \Level1Out17[29] , \Level1Out34[18] , \Level1Out41[28] , 
        \ScanLink26[9] , \ScanLink28[31] , \ScanLink38[5] , \Level1Out41[31] , 
        \Level1Out62[19] , \Level4Out44[8] , \Level8Out32[25] , 
        \ScanLink28[28] , \Level1Load45[0] , \Level2Out4[14] , 
        \Level8Out32[16] , \ScanLink3[1] , \ScanLink8[21] , \Level1Out8[3] , 
        \Level1Out18[27] , \Level2Out4[27] , \Level2Out20[19] , 
        \Level1Out24[2] , \Level1Out27[1] , \Level2Out0[16] , 
        \Level2Out24[31] , \Level2Out24[28] , \Level8Out56[23] , 
        \Level16Out48[5] , \Level8Out40[0] , \ScanLink8[12] , 
        \Level1Out18[14] , \Level1Out43[5] , \ScanLink59[30] , 
        \ScanLink59[29] , \Level2Out0[25] , \ScanLink11[10] , \ScanLink27[15] , 
        \Level1Out40[6] , \Level2Out34[9] , \Level4Out8[19] , \Level8Out24[4] , 
        \ScanLink52[25] , \Level8Out56[10] , \ScanLink60[5] , \ScanLink32[21] , 
        \ScanLink47[11] , \ScanLink64[20] , \Level1Out13[18] , 
        \Level1Out30[30] , \Level1Out30[29] , \Level1Out45[19] , 
        \ScanLink63[6] , \Level2Out56[3] , \Level16Out16[19] , 
        \Level8Out48[28] , \Level8Out48[31] , \Level1Out0[24] , 
        \Level1Out0[17] , \ScanLink9[18] , \ScanLink11[23] , \ScanLink32[12] , 
        \ScanLink47[22] , \ScanLink27[26] , \Level1Out58[4] , \ScanLink64[13] , 
        \Level1Out46[8] , \ScanLink52[16] , \Level2Out32[7] , \Level2Out24[3] , 
        \Level4Out20[25] , \ScanLink11[6] , \ScanLink12[5] , \Level2Out4[1] , 
        \Level4Out16[20] , \Level4Out40[21] , \Level1Out5[6] , 
        \Level1Out29[7] , \ScanLink38[27] , \ScanLink58[23] , 
        \Level2Out30[25] , \Level8Out0[22] , \Level2Out50[21] , 
        \Level4Out16[13] , \Level4Out20[16] , \Level4Out40[12] , 
        \Level1Out34[8] , \Level2Out40[7] , \Level1Out6[5] , \ScanLink38[14] , 
        \Level2Out50[12] , \ScanLink58[10] , \Level2Out30[16] , 
        \Level8Out0[11] , \ScanLink2[27] , \ScanLink2[14] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink17[8] , \Level1Out56[2] , \Level8Out32[0] , 
        \ScanLink46[31] , \Level1Out12[21] , \Level1Out24[24] , 
        \ScanLink33[18] , \ScanLink46[28] , \Level1Out51[14] , 
        \Level1Out31[10] , \Level4Out0[7] , \Level1Out44[20] , 
        \Level1Out55[1] , \Level8Out56[4] , \Level1Out3[8] , \ScanLink6[25] , 
        \Level1Out12[12] , \Level1Out32[6] , \Level2Out46[9] , 
        \Level1Out15[3] , \Level1Out16[23] , \Level1Out24[17] , 
        \Level1Out31[23] , \Level1Out44[13] , \Level1Out31[5] , 
        \Level1Out51[27] , \Level2Out18[18] , \Level8Out48[8] , 
        \Level2Out58[5] , \Level1Out35[12] , \Level1Out63[13] , 
        \Level1Out40[22] , \Level1Out20[26] , \Level1Load37[0] , 
        \ScanLink49[6] , \Level1Out55[16] , \ScanLink54[9] , \ScanLink14[18] , 
        \Level1Out16[0] , \ScanLink37[30] , \ScanLink61[28] , \Level2Out18[7] , 
        \ScanLink37[29] , \ScanLink42[19] , \ScanLink61[31] , \Level1Out1[23] , 
        \Level1Out1[10] , \Level1Out4[26] , \Level1Out4[15] , \ScanLink6[16] , 
        \Level1Out16[10] , \Level1Out20[15] , \Level1Out55[25] , 
        \Level1Out63[20] , \Level1Out35[21] , \Level1Out40[11] , 
        \ScanLink29[11] , \ScanLink49[15] , \Level8Out16[6] , 
        \Level2Out34[27] , \Level2Out54[23] , \Level2Out62[26] , 
        \ScanLink51[4] , \ScanLink52[7] , \Level4Out12[22] , \Level4Out24[27] , 
        \Level4Out44[23] , \Level1Out18[19] , \ScanLink29[22] , 
        \ScanLink36[3] , \ScanLink35[0] , \ScanLink49[26] , \Level2Out34[14] , 
        \Level2Out54[10] , \Level2Out62[15] , \Level4Out36[8] , 
        \Level4Out12[11] , \Level4Out24[14] , \Level2Out34[4] , 
        \Level4Out8[14] , \Level4Out28[4] , \Level4Out44[10] , \Level4Out8[2] , 
        \Level8Out24[9] , \Level2Out0[31] , \Level2Out0[28] , 
        \Level1Load18[0] , \ScanLink39[20] , \Level1Out43[8] , 
        \ScanLink59[24] , \Level2Out12[13] , \Level2Out44[12] , 
        \Level2Out24[16] , \Level16Out32[0] , \ScanLink39[13] , 
        \Level1Out39[0] , \Level2Out50[0] , \Level16Out48[8] , 
        \Level4Out8[27] , \ScanLink59[17] , \Level2Out24[25] , 
        \Level2Out44[21] , \Level2Load6[0] , \Level2Out12[20] , 
        \ScanLink3[20] , \Level1Out13[26] , \ScanLink19[3] , \Level1Out25[23] , 
        \Level1Out46[5] , \Level1Out58[9] , \Level8Out48[16] , 
        \Level16Out0[22] , \Level16Out16[27] , \Level1Out50[13] , 
        \Level1Out30[17] , \Level1Out45[27] , \Level1Out45[6] , 
        \Level8Out48[25] , \Level16Out0[11] , \ScanLink3[13] , \ScanLink5[2] , 
        \Level1Out13[15] , \Level1Out22[1] , \Level16Out16[14] , 
        \Level1Out17[24] , \Level1Out21[2] , \Level1Out30[24] , 
        \Level1Out45[14] , \Level4Out60[3] , \Level1Out50[20] , 
        \Level1Out25[10] , \ScanLink27[18] , \ScanLink52[28] , 
        \Level32Out0[3] , \ScanLink60[8] , \ScanLink52[31] , \Level2Out48[2] , 
        \Level1Out21[21] , \Level1Out34[15] , \Level1Out62[14] , 
        \Level1Out41[25] , \Level4Out44[5] , \ScanLink23[30] , 
        \ScanLink23[29] , \Level1Out54[11] , \ScanLink59[1] , \ScanLink56[19] , 
        \Level1Out5[21] , \Level1Out5[12] , \ScanLink6[1] , \ScanLink7[22] , 
        \ScanLink7[11] , \Level1Out17[17] , \Level1Out21[12] , 
        \Level1Out54[22] , \Level1Out61[0] , \Level1Out62[27] , 
        \Level1Out34[26] , \Level1Out41[16] , \Level4Out20[1] , 
        \Level1Out62[3] , \ScanLink23[9] , \Level1Load40[0] , \ScanLink28[16] , 
        \ScanLink48[12] , \Level2Out20[14] , \Level2Out40[10] , 
        \Level2Out16[11] , \ScanLink41[3] , \ScanLink42[0] , \Level2Out4[19] , 
        \ScanLink14[15] , \Level1Out20[18] , \ScanLink25[7] , \ScanLink26[4] , 
        \ScanLink28[25] , \Level2Out40[23] , \ScanLink38[8] , \ScanLink48[21] , 
        \Level2Out16[22] , \Level16Out16[6] , \Level2Out10[2] , 
        \Level2Out20[27] , \Level8Out32[31] , \Level8Out32[28] , 
        \ScanLink33[3] , \Level1Out55[31] , \Level1Out55[28] , 
        \ScanLink37[24] , \ScanLink42[14] , \ScanLink61[25] , \Level1Out0[30] , 
        \Level1Out0[29] , \Level1Out4[18] , \ScanLink6[31] , \ScanLink22[10] , 
        \ScanLink30[0] , \ScanLink57[20] , \ScanLink6[28] , \Level2Out62[2] , 
        \ScanLink8[7] , \ScanLink14[26] , \ScanLink22[23] , \ScanLink57[7] , 
        \ScanLink37[17] , \ScanLink57[13] , \ScanLink42[27] , \ScanLink54[4] , 
        \ScanLink61[16] , \Level1Out10[3] , \ScanLink28[2] , \Level4Out24[19] , 
        \Level4Out28[9] , \Level2Out34[19] , \Level2Out62[18] , 
        \Level4Out36[5] , \Level1Load32[0] , \ScanLink51[9] , \Level1Out13[0] , 
        \ScanLink49[18] , \Level4Out52[1] , \Level1Out0[6] , \Level1Out6[8] , 
        \Level1Out19[20] , \Level1Out37[6] , \ScanLink38[19] , \ScanLink9[26] , 
        \Level1Out34[5] , \ScanLink9[15] , \ScanLink12[8] , \Level1Out19[13] , 
        \Level1Out53[2] , \Level2Out30[31] , \Level2Out30[28] , 
        \Level4Out12[3] , \Level4Out20[31] , \Level4Out20[28] , 
        \ScanLink10[17] , \ScanLink26[12] , \Level1Out50[1] , \ScanLink53[22] , 
        \Level2Out18[15] , \ScanLink33[26] , \ScanLink46[16] , 
        \Level2Out58[8] , \ScanLink2[19] , \Level1Out31[8] , \Level8Out48[5] , 
        \Level1Out3[5] , \Level2Out46[4] , \Level1Out4[22] , \Level1Out4[11] , 
        \ScanLink10[24] , \ScanLink14[6] , \Level1Out24[30] , \Level8Out56[9] , 
        \Level1Out24[29] , \ScanLink33[15] , \Level1Out51[19] , 
        \ScanLink46[25] , \ScanLink17[5] , \ScanLink26[21] , \Level1Out48[3] , 
        \Level2Out18[26] , \ScanLink53[11] , \ScanLink51[0] , \Level2Out2[2] , 
        \Level2Out22[0] , \ScanLink52[3] , \Level4Out12[26] , 
        \Level4Out24[23] , \Level4Out44[27] , \Level1Out13[9] , 
        \ScanLink29[15] , \Level2Out34[23] , \Level2Out62[22] , 
        \Level4Out52[8] , \ScanLink49[11] , \Level2Out54[27] , 
        \ScanLink29[26] , \ScanLink35[4] , \Level4Out12[15] , \Level4Out28[0] , 
        \Level4Out44[14] , \ScanLink49[22] , \Level2Out54[14] , 
        \Level4Out24[10] , \Level2Out62[11] , \Level2Out34[10] , 
        \ScanLink6[21] , \ScanLink36[7] , \ScanLink6[12] , \Level1Out15[7] , 
        \Level1Out16[4] , \Level1Out20[22] , \ScanLink49[2] , 
        \Level1Out35[16] , \Level1Out55[12] , \Level1Out40[26] , 
        \Level1Out16[27] , \Level1Out63[17] , \Level8Out16[2] , 
        \Level1Out16[14] , \Level1Out35[25] , \Level1Out40[15] , 
        \Level1Out63[24] , \Level1Out20[11] , \Level1Out55[21] , 
        \ScanLink57[30] , \ScanLink57[29] , \Level1Out0[20] , \Level1Out0[13] , 
        \ScanLink2[23] , \Level1Out12[25] , \ScanLink22[19] , \ScanLink30[9] , 
        \Level1Load53[0] , \Level1Out31[14] , \Level2Out18[3] , 
        \Level1Out44[24] , \Level4Out0[3] , \Level1Out55[5] , 
        \Level1Out24[20] , \ScanLink26[31] , \Level1Out51[10] , 
        \ScanLink26[28] , \ScanLink53[18] , \Level2Out22[9] , \Level8Out32[4] , 
        \ScanLink2[10] , \Level1Out12[16] , \Level1Out24[13] , 
        \Level1Out31[1] , \Level1Out51[23] , \Level1Out56[6] , 
        \Level2Out58[1] , \Level8Load0[0] , \Level1Out31[27] , 
        \Level1Out44[17] , \Level1Out32[2] , \ScanLink38[23] , 
        \Level8Out56[0] , \ScanLink58[27] , \Level2Out30[21] , 
        \Level2Out50[25] , \Level8Out0[26] , \ScanLink11[2] , \ScanLink12[1] , 
        \Level2Out4[5] , \Level4Out40[25] , \Level4Out16[24] , 
        \Level1Out19[30] , \Level1Out50[8] , \Level2Out24[7] , 
        \Level4Out20[21] , \Level1Out19[29] , \Level1Out5[2] , \Level1Out6[1] , 
        \Level8Out0[15] , \ScanLink38[10] , \ScanLink58[14] , 
        \Level2Out30[12] , \Level2Out50[16] , \Level1Out22[8] , 
        \Level1Out29[3] , \Level2Out40[3] , \Level4Out20[12] , \ScanLink63[2] , 
        \Level4Out16[17] , \Level4Out40[16] , \Level16Out0[18] , 
        \Level2Out56[7] , \Level1Out25[19] , \Level1Out50[29] , 
        \ScanLink3[30] , \ScanLink3[29] , \ScanLink11[14] , \Level1Out50[30] , 
        \ScanLink64[24] , \ScanLink27[11] , \ScanLink32[25] , \ScanLink47[15] , 
        \ScanLink52[21] , \ScanLink60[1] , \Level2Out32[3] , \ScanLink11[27] , 
        \ScanLink27[22] , \ScanLink52[12] , \Level1Out58[0] , \ScanLink32[16] , 
        \ScanLink64[17] , \ScanLink47[26] , \ScanLink0[6] , \Level1Out1[19] , 
        \ScanLink8[25] , \ScanLink8[16] , \Level1Out8[7] , \Level1Out39[9] , 
        \Level16Out48[1] , \Level1Out18[23] , \Level1Out24[6] , 
        \Level2Out50[9] , \Level8Out40[4] , \Level1Out27[5] , 
        \Level2Out12[30] , \Level2Out44[28] , \Level8Out56[27] , 
        \Level2Out12[29] , \Level2Out44[31] , \Level1Out40[2] , 
        \Level2Out0[12] , \Level8Out56[14] , \Level8Out24[0] , \ScanLink3[5] , 
        \Level1Out5[31] , \Level1Out18[10] , \Level2Out0[21] , 
        \Level16Load32[0] , \ScanLink39[30] , \ScanLink39[29] , 
        \Level1Out43[1] , \Level16Out32[9] , \Level1Out5[28] , 
        \Level1Load21[0] , \ScanLink38[1] , \ScanLink48[31] , \Level2Out4[10] , 
        \ScanLink48[28] , \Level2Out16[18] , \Level2Out40[19] , 
        \Level8Out32[21] , \ScanLink42[9] , \Level2Out4[23] , \ScanLink6[8] , 
        \ScanLink7[18] , \ScanLink15[16] , \ScanLink20[3] , \ScanLink56[23] , 
        \Level8Out32[12] , \ScanLink23[13] , \ScanLink60[26] , 
        \ScanLink36[27] , \ScanLink43[17] , \Level1Out61[9] , \Level4Out20[8] , 
        \ScanLink15[25] , \Level1Out21[31] , \Level1Out21[28] , 
        \ScanLink23[0] , \Level2Out16[5] , \Level1Out54[18] , \ScanLink59[8] , 
        \Level1Out18[2] , \ScanLink23[20] , \ScanLink36[14] , \ScanLink60[15] , 
        \ScanLink43[24] , \ScanLink44[7] , \ScanLink56[10] , \ScanLink47[4] , 
        \ScanLink11[16] , \ScanLink27[13] , \ScanLink60[3] , \ScanLink52[23] , 
        \Level1Out21[9] , \ScanLink32[27] , \ScanLink64[26] , \Level2Out48[9] , 
        \ScanLink47[17] , \Level4Out60[8] , \ScanLink3[18] , \Level32Out0[8] , 
        \Level1Out25[28] , \Level1Out50[18] , \ScanLink63[0] , 
        \Level2Out56[5] , \ScanLink0[4] , \Level1Out1[31] , \ScanLink11[25] , 
        \ScanLink19[8] , \Level1Out25[31] , \ScanLink64[15] , \ScanLink27[20] , 
        \ScanLink32[14] , \ScanLink47[24] , \ScanLink52[10] , \Level1Out58[2] , 
        \Level2Out32[1] , \Level16Out0[30] , \Level16Out0[29] , 
        \Level1Out1[28] , \ScanLink8[27] , \Level1Out18[21] , \Level2Out0[10] , 
        \Level1Out24[4] , \Level1Out27[7] , \ScanLink39[18] , 
        \Level8Out56[25] , \ScanLink8[14] , \Level1Out8[5] , \Level8Out40[6] , 
        \Level1Out18[12] , \Level1Out43[3] , \Level2Out12[18] , 
        \Level2Out44[19] , \Level16Out48[3] , \Level1Load61[0] , 
        \Level2Out0[23] , \ScanLink38[3] , \Level1Out40[0] , \Level4Out8[9] , 
        \Level8Out24[2] , \Level8Out56[16] , \Level2Out10[9] , 
        \Level8Out32[23] , \Level2Out4[12] , \Level2Out16[30] , 
        \Level2Out16[29] , \Level2Out40[28] , \Level2Out40[31] , 
        \Level8Out32[10] , \ScanLink3[7] , \Level1Out5[19] , \ScanLink41[8] , 
        \Level2Out4[21] , \Level1Out4[20] , \Level1Out4[13] , \ScanLink5[9] , 
        \ScanLink7[30] , \ScanLink7[29] , \ScanLink15[14] , \Level1Out21[19] , 
        \ScanLink23[2] , \ScanLink48[19] , \Level1Out62[8] , \Level2Out16[7] , 
        \Level1Out54[30] , \Level1Out54[29] , \ScanLink20[1] , 
        \ScanLink36[25] , \ScanLink60[24] , \ScanLink43[15] , \ScanLink23[11] , 
        \ScanLink56[21] , \ScanLink15[27] , \Level1Out18[0] , \ScanLink23[22] , 
        \Level1Load39[0] , \ScanLink47[6] , \ScanLink56[12] , \ScanLink60[17] , 
        \ScanLink29[17] , \ScanLink36[16] , \ScanLink43[26] , \ScanLink44[5] , 
        \ScanLink49[13] , \Level2Out54[25] , \Level2Out62[20] , 
        \Level2Out34[21] , \Level1Out10[8] , \ScanLink51[2] , \ScanLink52[1] , 
        \Level4Out12[24] , \Level4Out44[25] , \Level4Out24[21] , 
        \ScanLink36[5] , \ScanLink6[23] , \Level1Out15[5] , \ScanLink28[9] , 
        \ScanLink29[24] , \Level2Out34[12] , \Level2Out62[13] , 
        \ScanLink49[20] , \Level2Out54[16] , \ScanLink35[6] , 
        \Level4Out24[12] , \Level4Out28[2] , \Level4Out44[16] , 
        \Level1Out40[24] , \Level4Out12[17] , \Level1Out16[25] , 
        \Level1Out35[14] , \Level1Out63[15] , \Level1Out16[6] , 
        \Level1Out20[20] , \ScanLink49[0] , \Level1Out55[10] , 
        \ScanLink22[31] , \ScanLink22[28] , \ScanLink57[18] , \Level2Out62[9] , 
        \Level2Out18[1] , \Level1Out0[22] , \Level1Out0[11] , \ScanLink2[21] , 
        \ScanLink6[10] , \Level1Out16[16] , \Level1Out20[13] , 
        \Level1Out35[27] , \Level1Out55[23] , \Level1Out40[17] , 
        \Level1Out63[26] , \ScanLink33[8] , \Level8Out16[0] , \Level1Out56[4] , 
        \ScanLink2[12] , \Level1Out12[27] , \Level1Out24[22] , 
        \Level1Out48[8] , \Level2Out2[9] , \Level8Out32[6] , \Level1Out51[12] , 
        \Level1Out31[16] , \Level1Out44[26] , \Level1Out55[7] , 
        \Level4Out0[1] , \Level4Load48[0] , \Level8Out56[2] , \ScanLink11[0] , 
        \Level1Out12[14] , \Level1Out31[25] , \Level1Out32[0] , 
        \Level1Out44[15] , \Level1Load13[0] , \Level1Out24[11] , 
        \Level1Out31[3] , \ScanLink26[19] , \Level1Out51[21] , 
        \ScanLink53[30] , \ScanLink53[29] , \Level2Out24[5] , \Level2Out58[3] , 
        \ScanLink12[3] , \Level1Out19[18] , \Level2Out4[7] , \Level4Out20[23] , 
        \Level4Out40[27] , \Level4Out16[26] , \Level1Out5[0] , 
        \Level1Out29[1] , \ScanLink38[21] , \ScanLink58[25] , 
        \Level2Out30[23] , \Level4Out12[8] , \Level8Out0[24] , 
        \Level1Out53[9] , \Level2Out50[27] , \Level4Out16[15] , 
        \Level4Out40[14] , \Level4Out20[10] , \Level1Out6[3] , 
        \ScanLink38[12] , \Level2Out40[1] , \ScanLink58[16] , 
        \Level2Out30[10] , \Level2Out50[14] , \Level8Out0[17] , 
        \Level1Out0[18] , \Level1Out4[30] , \Level1Out4[29] , \ScanLink6[19] , 
        \ScanLink14[17] , \ScanLink22[12] , \ScanLink30[2] , \ScanLink37[26] , 
        \ScanLink57[22] , \ScanLink42[16] , \ScanLink61[27] , \Level2Out18[8] , 
        \ScanLink8[5] , \Level1Out20[30] , \ScanLink33[1] , \ScanLink49[9] , 
        \Level8Out16[9] , \Level1Out55[19] , \ScanLink14[24] , 
        \Level1Out20[29] , \ScanLink37[15] , \ScanLink42[25] , \ScanLink54[6] , 
        \ScanLink61[14] , \ScanLink22[21] , \ScanLink57[11] , \ScanLink57[5] , 
        \Level2Load46[0] , \Level2Out62[0] , \Level1Load5[0] , \Level1Out5[9] , 
        \ScanLink9[24] , \Level1Out10[1] , \Level1Out13[2] , \ScanLink28[0] , 
        \ScanLink49[30] , \ScanLink49[29] , \Level4Out36[7] , 
        \Level2Out34[31] , \Level2Out62[29] , \Level2Out34[28] , 
        \Level2Out62[30] , \Level4Out52[3] , \ScanLink52[8] , 
        \Level4Out24[31] , \Level4Out24[28] , \Level1Out29[8] , 
        \Level4Out20[19] , \Level1Out19[22] , \Level1Out34[7] , 
        \Level1Out37[4] , \Level2Out40[8] , \Level2Out30[19] , 
        \Level1Out50[3] , \ScanLink9[17] , \ScanLink11[9] , \Level1Out0[4] , 
        \Level1Out3[7] , \Level1Out19[11] , \Level1Out32[9] , \ScanLink38[31] , 
        \ScanLink38[28] , \Level1Out53[0] , \Level4Out12[1] , \Level2Out46[6] , 
        \Level8Out48[7] , \Level1Out1[12] , \ScanLink2[31] , \ScanLink10[15] , 
        \Level1Out24[18] , \Level1Out51[31] , \ScanLink33[24] , 
        \Level1Out51[28] , \ScanLink46[14] , \ScanLink26[10] , 
        \Level2Out18[17] , \ScanLink53[20] , \ScanLink2[28] , \Level2Out22[2] , 
        \ScanLink10[26] , \ScanLink14[4] , \ScanLink17[7] , \Level2Out2[0] , 
        \ScanLink26[23] , \Level1Out48[1] , \Level2Out18[24] , 
        \ScanLink53[13] , \ScanLink46[27] , \ScanLink33[17] , \ScanLink39[22] , 
        \Level4Out0[8] , \ScanLink59[26] , \Level2Out24[14] , 
        \Level16Out32[2] , \Level2Out44[10] , \Level2Out12[11] , 
        \Level4Out8[0] , \Level1Out1[21] , \Level1Out18[31] , 
        \Level1Out18[28] , \Level1Out40[9] , \Level2Out34[6] , 
        \Level4Out8[16] , \Level2Out0[19] , \ScanLink3[22] , \Level1Out13[24] , 
        \ScanLink39[11] , \ScanLink59[15] , \Level2Out12[22] , 
        \Level2Out44[23] , \Level2Out24[27] , \Level1Out39[2] , 
        \Level2Out50[2] , \Level4Out8[25] , \ScanLink19[1] , \Level1Out25[21] , 
        \Level1Out30[15] , \Level1Out45[25] , \Level1Out45[4] , 
        \Level1Out50[11] , \ScanLink27[30] , \ScanLink27[29] , 
        \ScanLink52[19] , \Level1Out46[7] , \Level8Out48[14] , 
        \Level16Out0[20] , \Level2Out32[8] , \ScanLink3[11] , 
        \Level1Out13[17] , \Level1Out21[0] , \Level2Out48[0] , 
        \Level16Out16[25] , \Level1Out25[12] , \Level1Out50[22] , 
        \Level32Out0[1] , \Level1Out22[3] , \Level1Out30[26] , 
        \Level1Out45[16] , \Level4Out60[1] , \Level16Out16[16] , 
        \Level1Load0[0] , \Level1Out0[26] , \Level1Out0[15] , \ScanLink5[0] , 
        \ScanLink6[3] , \ScanLink7[20] , \ScanLink63[9] , \Level8Out48[27] , 
        \Level16Out0[13] , \Level1Out5[23] , \Level1Out5[10] , \ScanLink7[13] , 
        \Level1Out17[26] , \Level1Out18[9] , \Level1Out21[23] , 
        \Level1Out54[13] , \ScanLink59[3] , \Level4Out44[7] , 
        \Level1Out62[16] , \Level1Out34[17] , \Level1Out41[27] , 
        \Level1Out17[15] , \Level1Out62[1] , \ScanLink20[8] , 
        \Level1Out21[10] , \Level1Out34[24] , \Level1Out62[25] , 
        \Level1Out41[14] , \Level4Out20[3] , \Level1Out61[2] , 
        \Level1Out54[20] , \ScanLink23[18] , \ScanLink41[1] , \ScanLink56[31] , 
        \ScanLink56[28] , \Level8Out32[19] , \ScanLink42[2] , \Level2Out4[28] , 
        \Level2Out4[31] , \ScanLink25[5] , \ScanLink28[14] , \Level2Out40[12] , 
        \ScanLink48[10] , \Level2Out16[13] , \Level2Out20[16] , 
        \ScanLink26[6] , \ScanLink28[27] , \ScanLink48[23] , \Level2Out10[0] , 
        \Level2Load34[0] , \Level1Load58[0] , \Level2Out20[25] , 
        \Level2Out40[21] , \Level16Out16[4] , \Level2Out16[20] , 
        \ScanLink38[25] , \ScanLink58[21] , \Level2Out30[27] , 
        \Level2Out50[23] , \Level8Out0[20] , \ScanLink11[4] , \ScanLink12[7] , 
        \Level2Out4[3] , \Level4Out16[22] , \Level4Out20[27] , 
        \Level4Out40[23] , \Level2Out24[1] , \Level1Out5[4] , \Level1Out6[7] , 
        \ScanLink58[12] , \Level2Out30[14] , \Level1Out37[9] , 
        \ScanLink38[16] , \Level8Out0[13] , \Level2Out40[5] , 
        \Level2Out50[10] , \ScanLink9[30] , \ScanLink9[29] , \Level1Out29[5] , 
        \Level4Out20[14] , \Level1Out12[23] , \Level4Out16[11] , 
        \Level4Out40[10] , \Level1Out31[12] , \Level1Out44[22] , 
        \Level1Out55[3] , \Level4Out0[5] , \Level1Out0[9] , \ScanLink2[25] , 
        \ScanLink14[9] , \Level1Out24[26] , \Level1Out51[16] , 
        \Level2Out18[30] , \Level2Out18[29] , \Level1Out56[0] , 
        \Level8Out32[2] , \ScanLink10[18] , \Level1Out24[15] , 
        \Level1Out31[7] , \ScanLink33[30] , \ScanLink33[29] , \Level2Out58[7] , 
        \ScanLink46[19] , \Level1Out51[25] , \ScanLink2[16] , 
        \Level1Out12[10] , \Level1Out31[21] , \Level1Out32[4] , 
        \Level1Out44[11] , \ScanLink6[27] , \Level1Out16[2] , \Level8Out56[6] , 
        \ScanLink6[14] , \ScanLink8[8] , \ScanLink14[30] , \ScanLink14[29] , 
        \ScanLink42[31] , \ScanLink57[8] , \ScanLink61[19] , \ScanLink37[18] , 
        \ScanLink42[28] , \Level1Out20[24] , \Level1Out55[14] , 
        \Level1Out15[1] , \Level1Out16[21] , \ScanLink49[4] , 
        \Level1Out63[11] , \Level1Out40[20] , \Level1Out35[10] , 
        \Level8Out16[4] , \Level1Out16[12] , \Level1Out20[17] , 
        \Level1Out35[23] , \Level1Out63[22] , \Level1Out40[13] , 
        \Level1Out55[27] , \ScanLink0[0] , \ScanLink3[3] , \Level1Out4[24] , 
        \Level1Out4[17] , \ScanLink51[6] , \Level2Out18[5] , \Level4Out24[25] , 
        \ScanLink52[5] , \Level4Out12[20] , \Level4Out44[21] , 
        \ScanLink29[20] , \ScanLink29[13] , \ScanLink35[2] , \ScanLink49[17] , 
        \Level2Out34[25] , \Level2Out54[21] , \Level2Out62[24] , 
        \ScanLink49[24] , \Level4Out12[13] , \Level4Out24[16] , 
        \Level4Out28[6] , \Level4Out44[12] , \Level2Out34[16] , 
        \Level2Out54[12] , \ScanLink36[1] , \Level2Out62[17] , 
        \ScanLink15[23] , \ScanLink15[10] , \ScanLink20[5] , \ScanLink23[15] , 
        \ScanLink36[21] , \ScanLink56[25] , \ScanLink43[11] , 
        \Level1Out17[18] , \Level1Out34[29] , \ScanLink60[20] , 
        \Level1Out41[19] , \Level1Out62[31] , \ScanLink23[6] , 
        \Level1Out34[30] , \Level1Out62[28] , \Level2Out16[3] , 
        \ScanLink36[12] , \ScanLink43[22] , \ScanLink44[1] , \ScanLink60[13] , 
        \Level1Out18[4] , \ScanLink23[26] , \ScanLink56[16] , \ScanLink25[8] , 
        \ScanLink38[7] , \ScanLink47[2] , \Level2Out4[16] , \Level16Load16[0] , 
        \Level2Out20[31] , \Level2Out20[28] , \Level16Out16[9] , 
        \Level8Out32[27] , \ScanLink28[19] , \Level2Out4[25] , \ScanLink8[23] , 
        \Level1Out8[1] , \Level8Out32[14] , \Level8Out40[2] , 
        \Level16Out48[7] , \ScanLink8[10] , \Level1Out18[25] , 
        \Level1Out24[0] , \Level4Out8[28] , \Level1Out27[3] , \Level4Out8[31] , 
        \Level8Out56[21] , \ScanLink59[18] , \Level2Out0[14] , 
        \Level1Out40[4] , \Level8Out24[6] , \Level8Out56[12] , 
        \Level1Out18[16] , \Level1Out43[7] , \Level2Out0[27] , 
        \Level2Out24[19] , \ScanLink63[4] , \Level2Out56[1] , \ScanLink11[21] , 
        \ScanLink11[12] , \ScanLink32[23] , \ScanLink47[13] , \ScanLink27[24] , 
        \ScanLink27[17] , \ScanLink60[7] , \ScanLink64[22] , \ScanLink52[27] , 
        \ScanLink52[14] , \Level1Out58[6] , \Level2Out32[5] , 
        \Level16Out16[31] , \Level16Out16[28] , \Level8Out48[19] , 
        \ScanLink32[10] , \ScanLink47[20] , \ScanLink64[11] , 
        \Level1Out13[30] , \Level1Out30[18] , \Level1Out45[28] , 
        \Level1Out45[9] , \Level1Out13[29] , \Level1Out45[31] , \ScanLink0[9] , 
        \Level1Out5[14] , \ScanLink28[10] , \ScanLink48[14] , 
        \Level2Out16[17] , \Level2Out20[12] , \Level2Out40[16] , 
        \ScanLink41[5] , \ScanLink42[6] , \Level2Load50[0] , \ScanLink3[26] , 
        \ScanLink5[4] , \Level1Out5[27] , \ScanLink26[2] , \Level1Out17[22] , 
        \ScanLink25[1] , \ScanLink28[23] , \Level2Out16[24] , 
        \Level2Out40[25] , \Level16Out16[0] , \ScanLink48[27] , 
        \Level2Out10[4] , \Level2Out20[21] , \Level1Out34[13] , 
        \Level1Out41[23] , \Level1Out62[12] , \Level1Out21[27] , 
        \Level1Out54[17] , \ScanLink59[7] , \ScanLink44[8] , \Level4Out44[3] , 
        \ScanLink6[7] , \ScanLink7[24] , \ScanLink7[17] , \ScanLink15[19] , 
        \ScanLink36[28] , \ScanLink43[18] , \ScanLink60[30] , 
        \Level1Out17[11] , \Level1Out21[14] , \ScanLink36[31] , 
        \ScanLink60[29] , \Level1Out61[6] , \Level1Out34[20] , 
        \Level1Out54[24] , \Level1Out41[10] , \Level4Out20[7] , 
        \Level1Out62[21] , \Level1Out62[5] , \Level1Out46[3] , 
        \Level16Out16[21] , \ScanLink11[31] , \ScanLink32[19] , 
        \ScanLink47[29] , \Level8Out48[10] , \Level16Out0[24] , 
        \ScanLink11[28] , \ScanLink47[30] , \ScanLink64[18] , 
        \Level1Out13[20] , \ScanLink19[5] , \Level1Out25[25] , 
        \Level1Out50[15] , \Level1Out30[11] , \Level1Out45[21] , 
        \Level1Out45[0] , \Level8Out48[23] , \Level1Out0[0] , \Level1Out1[25] , 
        \Level1Out1[16] , \ScanLink3[15] , \Level16Out0[17] , 
        \Level16Out16[12] , \ScanLink8[19] , \Level1Out13[13] , 
        \Level1Out22[7] , \Level1Out30[22] , \Level2Out56[8] , 
        \Level1Out45[12] , \Level4Out60[5] , \Level1Out21[4] , 
        \Level32Out0[5] , \Level1Out25[16] , \Level1Out50[26] , 
        \Level2Out34[2] , \Level2Out48[4] , \Level4Out8[12] , \Level4Out8[4] , 
        \Level1Out8[8] , \ScanLink39[26] , \ScanLink59[22] , \Level2Out12[15] , 
        \Level2Out44[14] , \Level2Out24[10] , \Level16Out32[6] , 
        \Level1Out24[9] , \Level1Out39[6] , \Level4Out8[21] , 
        \Level8Out56[31] , \Level8Out56[28] , \ScanLink39[15] , 
        \Level2Out24[23] , \Level2Out50[6] , \ScanLink59[11] , 
        \Level2Out12[26] , \Level2Out44[27] , \ScanLink10[11] , 
        \ScanLink26[14] , \ScanLink53[24] , \Level2Out18[13] , 
        \Level1Out12[19] , \ScanLink33[20] , \ScanLink46[10] , 
        \Level1Out31[31] , \Level1Out31[28] , \Level1Out44[18] , 
        \Level8Out48[3] , \ScanLink0[19] , \Level1Out3[3] , \ScanLink8[1] , 
        \ScanLink9[20] , \ScanLink10[22] , \Level2Out46[2] , \ScanLink14[0] , 
        \ScanLink46[23] , \Level1Load16[0] , \ScanLink17[3] , \ScanLink26[27] , 
        \ScanLink33[13] , \ScanLink53[17] , \Level1Out48[5] , 
        \Level2Out18[20] , \Level1Out19[26] , \Level1Out56[9] , 
        \Level2Out2[4] , \Level2Out22[6] , \Level1Out34[3] , \Level1Out37[0] , 
        \Level2Out50[19] , \Level2Load8[0] , \Level4Out16[18] , 
        \Level4Out40[19] , \ScanLink9[13] , \Level1Out19[15] , 
        \Level1Out53[4] , \ScanLink58[31] , \ScanLink58[28] , \Level8Out0[30] , 
        \Level4Out12[5] , \Level8Out0[29] , \Level1Out10[5] , \ScanLink28[4] , 
        \Level1Out50[7] , \Level2Out24[8] , \ScanLink29[30] , \ScanLink29[29] , 
        \ScanLink36[8] , \Level4Out36[3] , \Level1Out13[6] , \Level2Out54[31] , 
        \Level4Out12[30] , \Level4Out12[29] , \Level4Out44[31] , 
        \Level4Out44[28] , \ScanLink14[20] , \ScanLink14[13] , \ScanLink33[5] , 
        \Level2Load22[0] , \Level2Out54[28] , \Level4Out52[7] , 
        \ScanLink22[25] , \ScanLink22[16] , \ScanLink30[6] , \ScanLink37[22] , 
        \ScanLink61[23] , \ScanLink42[12] , \ScanLink57[26] , \ScanLink57[15] , 
        \ScanLink57[1] , \Level2Out62[4] , \ScanLink61[10] , \Level1Out15[8] , 
        \Level1Out16[28] , \ScanLink37[11] , \ScanLink42[21] , \ScanLink54[2] , 
        \Level1Out40[30] , \Level1Out63[18] , \Level1Out40[29] , 
        \Level1Out16[31] , \Level1Out35[19] , \Level1Out9[25] , 
        \Level1Out26[30] , \Level1Out26[29] , \Level1Out53[19] , 
        \ScanLink29[9] , \Level1Out9[16] , \Level1Out11[8] , \ScanLink12[24] , 
        \ScanLink24[21] , \ScanLink51[11] , \ScanLink12[17] , \ScanLink31[15] , 
        \ScanLink34[6] , \ScanLink44[25] , \ScanLink37[5] , \Level4Out0[21] , 
        \Level2Load26[0] , \ScanLink24[12] , \ScanLink31[26] , 
        \ScanLink44[16] , \ScanLink50[2] , \ScanLink51[22] , \Level1Out2[30] , 
        \ScanLink32[8] , \ScanLink53[1] , \Level1Out58[26] , \Level2Out32[31] , 
        \Level2Out32[28] , \Level4Out0[12] , \Level4Out32[3] , 
        \Level1Out38[22] , \Level1Out38[11] , \Level8Out16[22] , 
        \Level16Out48[13] , \Level32Out32[10] , \Level8Out40[23] , 
        \Level1Out58[15] , \Level1Out2[29] , \ScanLink4[31] , \ScanLink4[28] , 
        \Level1Out6[18] , \Level1Load12[0] , \Level1Out14[5] , 
        \Level1Out17[6] , \ScanLink19[31] , \ScanLink19[28] , \Level4Out56[7] , 
        \Level1Out30[3] , \ScanLink48[0] , \Level8Out16[11] , 
        \Level8Out40[10] , \Level8Out24[25] , \Level16Out48[20] , 
        \Level32Out32[23] , \Level1Out29[14] , \Level1Out49[10] , 
        \Level1Out29[27] , \Level1Out33[0] , \Level1Out49[8] , 
        \Level1Out54[7] , \Level8Out24[16] , \Level1Out57[4] , 
        \Level2Out20[8] , \Level2Out36[19] , \Level4Out16[5] , 
        \Level2Out60[18] , \Level1Out49[23] , \Level1Out7[3] , 
        \Level2Out42[2] , \Level1Out4[0] , \ScanLink16[26] , \ScanLink63[16] , 
        \Level4Out4[23] , \ScanLink20[23] , \ScanLink35[17] , \ScanLink40[27] , 
        \Level2Out28[21] , \ScanLink55[13] , \Level1Out28[1] , 
        \Level2Out48[25] , \ScanLink13[3] , \ScanLink1[20] , \ScanLink1[13] , 
        \ScanLink2[7] , \ScanLink5[22] , \ScanLink5[11] , \Level1Out7[21] , 
        \ScanLink10[0] , \ScanLink20[10] , \Level1Out22[18] , \Level1Out52[9] , 
        \Level2Out6[4] , \Level4Out4[10] , \Level2Out26[6] , \Level1Out57[31] , 
        \Level1Out57[28] , \ScanLink16[15] , \ScanLink55[20] , 
        \Level2Out48[16] , \ScanLink35[24] , \ScanLink63[25] , 
        \ScanLink40[14] , \Level2Out28[12] , \Level1Out7[12] , \ScanLink18[8] , 
        \Level1Out48[30] , \Level1Out48[29] , \Level2Out6[19] , 
        \Level2Out14[22] , \Level2Out22[27] , \Level2Out42[23] , 
        \Level1Out59[2] , \Level2Out30[2] , \Level4Out32[27] , \ScanLink62[0] , 
        \Level2Out14[11] , \Level4Out52[23] , \Level2Out22[14] , 
        \Level2Out42[10] , \Level1Out15[17] , \Level1Out20[9] , 
        \ScanLink61[3] , \Level4Out32[14] , \Level4Out52[10] , 
        \Level1Out36[26] , \Level2Out28[0] , \Level2Out54[6] , 
        \Level1Out43[16] , \Level1Out23[12] , \Level1Out60[27] , 
        \Level2Out8[2] , \Level1Out41[0] , \Level1Out56[22] , \Level1Out9[5] , 
        \Level1Out15[24] , \Level1Out23[21] , \Level1Out42[3] , 
        \Level1Out56[11] , \Level1Load60[0] , \Level1Out25[4] , 
        \Level1Out36[15] , \Level1Out43[25] , \Level1Out60[14] , 
        \ScanLink21[30] , \ScanLink21[29] , \ScanLink54[19] , \Level1Out26[7] , 
        \Level2Out52[8] , \ScanLink1[4] , \Level1Out11[15] , \Level1Out27[10] , 
        \Level1Out32[24] , \Level1Out52[20] , \Level32Out32[0] , 
        \Level1Out47[14] , \Level4Out40[3] , \ScanLink50[31] , 
        \Level8Out8[29] , \ScanLink25[18] , \ScanLink40[8] , \ScanLink50[28] , 
        \Level8Out8[30] , \Level1Out3[23] , \ScanLink4[9] , \Level1Out11[26] , 
        \Level1Out32[17] , \Level1Out47[27] , \Level2Out58[19] , 
        \Level4Out48[19] , \Level1Out19[0] , \Level1Out27[23] , 
        \ScanLink39[3] , \Level1Out52[13] , \Level4Out24[7] , 
        \Level32Out0[22] , \Level2Load54[0] , \Level4Out56[21] , 
        \Level4Out36[25] , \ScanLink18[22] , \Level1Load38[0] , 
        \ScanLink45[5] , \Level4Out60[24] , \Level2Out10[20] , 
        \Level2Out26[25] , \Level2Out46[21] , \ScanLink46[6] , 
        \Level1Out3[19] , \Level1Out3[10] , \ScanLink21[1] , \Level2Out14[4] , 
        \Level4Out36[16] , \Level4Out60[17] , \Level32Out0[11] , 
        \Level4Out56[12] , \ScanLink5[18] , \ScanLink17[25] , \ScanLink18[11] , 
        \ScanLink22[2] , \Level1Out39[28] , \Level2Out2[31] , \Level8Out0[4] , 
        \Level1Out39[31] , \Level2Out2[28] , \Level1Out63[8] , 
        \Level2Out26[16] , \ScanLink21[20] , \Level1Out23[31] , 
        \Level2Out10[13] , \Level2Out46[12] , \Level1Out23[28] , 
        \Level1Out56[18] , \Level1Out38[2] , \ScanLink54[10] , 
        \ScanLink34[14] , \ScanLink41[24] , \ScanLink64[7] , \ScanLink62[15] , 
        \ScanLink17[16] , \ScanLink34[27] , \Level2Out52[1] , \ScanLink41[17] , 
        \ScanLink21[13] , \ScanLink62[26] , \Level2Out28[9] , \Level1Out41[9] , 
        \ScanLink54[23] , \Level2Out36[5] , \Level1Out7[31] , \Level1Out7[28] , 
        \Level1Out20[0] , \Level1Out23[3] , \Level1Out28[17] , 
        \Level2Out14[18] , \Level2Out42[19] , \Level1Out48[13] , 
        \ScanLink62[9] , \Level2Out6[23] , \Level4Out52[19] , 
        \Level1Out48[20] , \Level2Out6[10] , \Level1Out28[24] , 
        \ScanLink18[1] , \Level1Out44[4] , \Level1Out47[7] , \ScanLink21[8] , 
        \Level1Out60[2] , \Level32Out0[18] , \Level1Out39[21] , 
        \Level2Out2[21] , \ScanLink4[0] , \ScanLink18[18] , \Level1Out59[25] , 
        \Level1Out63[1] , \ScanLink1[30] , \ScanLink7[3] , \Level1Out19[9] , 
        \Level4Out56[31] , \ScanLink58[3] , \Level4Out56[28] , 
        \Level1Out59[16] , \Level2Out10[30] , \Level2Out10[29] , 
        \Level2Out46[31] , \Level2Out46[28] , \Level1Out39[12] , 
        \Level1Load59[0] , \Level2Out2[12] , \Level4Out48[10] , 
        \ScanLink1[29] , \Level1Out2[20] , \Level1Out8[26] , \ScanLink13[27] , 
        \ScanLink24[5] , \ScanLink27[6] , \Level2Out12[3] , \Level4Out28[14] , 
        \ScanLink30[16] , \ScanLink45[26] , \Level2Out58[10] , 
        \ScanLink25[22] , \ScanLink50[12] , \Level8Out8[13] , 
        \Level2Out38[14] , \Level1Out8[15] , \ScanLink43[2] , 
        \Level4Out28[27] , \Level4Out48[23] , \Level32Out32[9] , 
        \ScanLink13[14] , \ScanLink25[11] , \Level1Out27[19] , 
        \Level1Out52[30] , \Level1Out52[29] , \Level8Out8[20] , 
        \ScanLink30[25] , \ScanLink40[1] , \ScanLink50[21] , \Level2Out38[27] , 
        \Level2Out58[23] , \Level16Out0[5] , \ScanLink45[15] , \ScanLink56[5] , 
        \Level1Out2[13] , \ScanLink9[5] , \ScanLink19[21] , \Level1Out38[18] , 
        \ScanLink48[9] , \Level2Out32[12] , \Level2Out52[16] , 
        \ScanLink19[12] , \ScanLink55[6] , \Level2Out60[3] , \Level8Out16[18] , 
        \Level8Out40[19] , \Level2Out32[21] , \Level4Out48[2] , 
        \Level16Out48[30] , \Level16Out48[29] , \ScanLink32[1] , 
        \Level2Out52[25] , \Level1Out10[16] , \ScanLink31[2] , 
        \Level32Out32[19] , \Level1Out11[1] , \Level1Out26[13] , 
        \Level1Out33[27] , \Level2Out8[27] , \Level1Out46[17] , 
        \ScanLink0[10] , \Level1Out53[23] , \Level1Out12[2] , \ScanLink53[8] , 
        \Level1Out53[10] , \ScanLink0[23] , \Level1Out10[25] , 
        \Level1Out26[20] , \ScanLink29[0] , \Level2Out8[14] , \ScanLink24[31] , 
        \ScanLink24[28] , \Level1Out33[14] , \Level1Out46[24] , 
        \ScanLink51[18] , \Level4Out0[31] , \Level4Out0[28] , \Level8Out8[5] , 
        \ScanLink1[24] , \ScanLink1[17] , \ScanLink1[0] , \Level1Out1[4] , 
        \ScanLink4[21] , \ScanLink4[12] , \Level1Out52[0] , \Level4Out4[19] , 
        \Level4Load28[0] , \Level1Load4[0] , \Level1Out22[11] , 
        \Level16Out32[24] , \Level1Out51[3] , \Level1Out57[21] , 
        \ScanLink10[9] , \Level1Out14[14] , \Level4Out4[5] , \ScanLink20[19] , 
        \Level1Out37[25] , \Level1Out61[24] , \Level1Out42[15] , 
        \Level2Out38[3] , \Level1Out36[4] , \ScanLink55[30] , \ScanLink55[29] , 
        \Level16Out32[17] , \Level1Out4[9] , \Level1Out28[8] , 
        \Level1Out61[17] , \Level2Out28[31] , \Level2Out28[28] , 
        \Level1Out6[22] , \Level1Out14[27] , \ScanLink15[4] , 
        \Level1Out22[22] , \Level1Out35[7] , \Level1Out37[16] , 
        \Level1Out42[26] , \Level1Out57[12] , \Level1Out49[1] , 
        \Level2Out0[3] , \ScanLink16[7] , \Level2Out20[1] , \Level2Out36[10] , 
        \Level2Out56[14] , \Level2Out60[11] , \Level1Out2[7] , 
        \Level1Out6[11] , \Level2Out44[5] , \Level1Out33[9] , 
        \Level1Out49[19] , \Level2Out56[27] , \Level1Out3[27] , 
        \ScanLink46[2] , \Level2Out36[23] , \Level2Out60[22] , 
        \Level1Out3[14] , \ScanLink18[26] , \ScanLink18[15] , \Level1Out19[4] , 
        \ScanLink45[1] , \Level2Out10[24] , \Level2Out26[21] , 
        \Level2Out46[25] , \Level4Out60[20] , \Level4Out36[21] , 
        \Level2Out10[17] , \Level2Out46[16] , \Level4Out56[25] , 
        \Level32Out0[26] , \ScanLink22[6] , \Level2Out26[12] , 
        \Level1Out59[28] , \Level8Out0[0] , \ScanLink21[5] , \Level1Out59[31] , 
        \Level2Load30[0] , \Level4Out56[16] , \Level32Out0[15] , 
        \Level2Out14[0] , \Level4Out36[12] , \Level4Out60[13] , 
        \Level1Out8[18] , \Level1Out11[11] , \ScanLink13[19] , 
        \ScanLink30[31] , \ScanLink30[28] , \Level16Out0[8] , \ScanLink45[18] , 
        \Level1Out27[14] , \Level1Out32[20] , \Level32Out32[4] , 
        \Level1Out47[10] , \Level4Out40[7] , \Level1Out52[24] , \ScanLink2[3] , 
        \Level1Out11[22] , \Level1Out27[27] , \Level1Out52[17] , 
        \Level4Out24[3] , \ScanLink39[7] , \ScanLink24[8] , \Level1Out32[13] , 
        \Level1Out47[23] , \Level2Out38[19] , \Level32Load0[0] , 
        \Level1Out4[4] , \ScanLink5[26] , \ScanLink5[15] , \Level1Out42[7] , 
        \Level4Out28[19] , \Level2Out36[8] , \Level1Out15[13] , 
        \Level1Out23[16] , \Level1Out41[4] , \Level1Out56[26] , 
        \Level2Out8[6] , \Level1Out26[3] , \Level1Out36[22] , 
        \Level1Out60[23] , \Level1Out43[12] , \Level2Out28[4] , 
        \Level1Out7[25] , \Level1Out9[1] , \Level1Out15[20] , \ScanLink17[31] , 
        \ScanLink17[28] , \ScanLink41[30] , \ScanLink62[18] , \ScanLink41[29] , 
        \ScanLink34[19] , \Level1Out60[10] , \Level1Out23[25] , 
        \Level1Out25[0] , \Level1Out36[11] , \Level1Out43[21] , 
        \Level1Out56[15] , \Level1Out28[29] , \Level1Out44[9] , 
        \Level1Out59[6] , \Level4Out32[23] , \Level4Out52[27] , 
        \Level2Out14[26] , \Level2Out30[6] , \Level2Out42[27] , 
        \Level2Out22[23] , \Level1Out7[16] , \Level1Out28[30] , 
        \ScanLink61[7] , \Level2Out54[2] , \Level4Out32[10] , 
        \Level4Out52[14] , \ScanLink62[4] , \Level2Out14[15] , 
        \Level2Out22[10] , \Level2Out42[14] , \Level1Out7[7] , 
        \ScanLink16[22] , \ScanLink20[27] , \Level1Out28[5] , \ScanLink55[17] , 
        \ScanLink35[13] , \ScanLink40[23] , \Level2Out28[25] , 
        \Level2Out48[21] , \ScanLink63[12] , \Level4Out4[27] , \ScanLink10[4] , 
        \ScanLink16[11] , \ScanLink35[20] , \Level1Out36[9] , \Level2Out42[6] , 
        \ScanLink40[10] , \Level2Out28[16] , \ScanLink20[14] , 
        \ScanLink63[21] , \ScanLink13[7] , \Level1Out14[19] , 
        \Level1Out37[31] , \Level1Out37[28] , \ScanLink55[24] , 
        \Level2Out48[12] , \Level4Out4[8] , \Level1Out42[18] , 
        \Level1Out61[30] , \Level1Out61[29] , \Level2Out6[0] , 
        \Level2Out26[2] , \Level16Out32[30] , \Level16Out32[29] , 
        \Level1Load1[0] , \Level1Out1[9] , \Level1Out29[10] , \Level1Out33[4] , 
        \Level4Out4[14] , \Level1Out30[7] , \Level1Out49[14] , 
        \Level2Out44[8] , \Level1Out29[23] , \Level1Out49[27] , 
        \Level8Out24[21] , \Level1Out54[3] , \Level1Out57[0] , 
        \Level2Out56[19] , \Level4Out16[1] , \ScanLink9[8] , \ScanLink15[9] , 
        \Level8Out24[12] , \Level1Out38[26] , \Level8Out16[26] , 
        \Level8Out40[27] , \Level16Out48[17] , \Level32Out32[14] , 
        \Level1Out58[22] , \Level2Out52[31] , \Level2Out52[28] , 
        \Level4Out32[7] , \Level16Out48[24] , \Level32Out32[27] , 
        \Level1Out9[21] , \ScanLink12[20] , \Level1Out14[1] , \ScanLink48[4] , 
        \Level8Out16[15] , \Level8Out40[14] , \Level1Out17[2] , 
        \Level4Out56[3] , \ScanLink31[11] , \ScanLink34[2] , \ScanLink37[1] , 
        \Level1Out38[15] , \ScanLink56[8] , \Level1Out58[11] , \Level8Out8[8] , 
        \Level4Out0[25] , \ScanLink44[21] , \ScanLink24[25] , \ScanLink51[15] , 
        \Level1Out9[12] , \Level1Out10[31] , \Level1Out46[29] , 
        \Level1Out10[28] , \Level1Out33[19] , \Level1Out46[30] , 
        \ScanLink53[5] , \Level2Out8[19] , \Level2Load42[0] , \Level4Out0[16] , 
        \Level8Load48[0] , \ScanLink0[14] , \Level1Out1[0] , \Level1Out2[3] , 
        \Level1Out6[26] , \ScanLink12[13] , \ScanLink24[16] , \ScanLink31[22] , 
        \ScanLink50[6] , \ScanLink51[26] , \ScanLink44[12] , \ScanLink16[3] , 
        \ScanLink15[0] , \Level1Out57[9] , \Level2Out56[10] , \Level4Out16[8] , 
        \Level2Out20[5] , \Level2Out36[14] , \Level2Out60[15] , 
        \Level1Out49[5] , \Level2Out0[7] , \Level2Out36[27] , 
        \Level2Out60[26] , \Level2Out56[23] , \Level1Out6[15] , 
        \Level1Out29[19] , \Level2Out44[1] , \Level8Out24[31] , 
        \ScanLink4[25] , \ScanLink4[16] , \Level1Out14[10] , \ScanLink16[18] , 
        \ScanLink35[30] , \ScanLink35[29] , \Level8Out24[28] , 
        \ScanLink40[19] , \ScanLink63[31] , \Level1Out37[21] , 
        \ScanLink63[28] , \Level2Out38[7] , \Level1Out42[11] , 
        \Level1Out22[15] , \Level1Out61[20] , \Level1Out51[7] , 
        \Level1Out57[25] , \Level4Out4[1] , \Level1Out14[23] , 
        \Level1Out22[26] , \Level1Out52[4] , \Level16Out32[20] , 
        \Level1Out57[16] , \Level2Out6[9] , \Level1Out35[3] , 
        \Level1Out37[12] , \Level1Out42[22] , \Level1Out61[13] , 
        \Level1Load17[0] , \Level1Out36[0] , \Level2Out48[31] , 
        \Level2Out48[28] , \Level16Out32[13] , \Level1Out12[6] , 
        \Level1Out11[5] , \Level1Out26[17] , \ScanLink0[27] , 
        \Level1Out10[12] , \Level1Out33[23] , \Level1Out53[27] , 
        \Level1Out46[13] , \Level2Out8[23] , \Level8Out8[1] , \Level1Out9[28] , 
        \Level1Out10[21] , \ScanLink12[30] , \ScanLink37[8] , \ScanLink44[28] , 
        \ScanLink12[29] , \ScanLink31[18] , \ScanLink44[31] , 
        \Level1Out33[10] , \Level1Out46[20] , \Level2Out8[10] , 
        \ScanLink29[4] , \Level1Out53[14] , \ScanLink1[9] , \Level1Out2[24] , 
        \ScanLink9[1] , \Level1Out9[31] , \Level1Out14[8] , \Level1Out26[24] , 
        \ScanLink55[2] , \Level4Out48[6] , \Level2Out60[7] , \ScanLink19[25] , 
        \Level2Out32[16] , \Level2Out52[12] , \ScanLink56[1] , 
        \Level1Out2[17] , \ScanLink31[6] , \Level1Out58[18] , \Level1Out8[22] , 
        \ScanLink19[16] , \ScanLink32[5] , \Level2Out52[21] , 
        \Level2Out32[25] , \ScanLink13[23] , \ScanLink25[26] , 
        \ScanLink50[16] , \Level2Out38[10] , \Level8Out8[17] , 
        \ScanLink13[10] , \ScanLink24[1] , \ScanLink27[2] , \ScanLink30[12] , 
        \ScanLink45[22] , \Level2Out58[14] , \Level2Out12[7] , 
        \Level4Out28[10] , \Level4Out48[14] , \ScanLink25[15] , 
        \ScanLink30[21] , \Level2Out58[27] , \ScanLink45[11] , 
        \Level16Out0[1] , \ScanLink40[5] , \ScanLink50[25] , \Level2Out38[23] , 
        \Level8Out8[24] , \ScanLink4[4] , \ScanLink7[7] , \Level1Out8[11] , 
        \Level1Out11[18] , \Level1Out32[30] , \Level1Out32[29] , 
        \Level1Out39[25] , \ScanLink43[6] , \Level1Out47[19] , 
        \Level4Out28[23] , \Level4Out48[27] , \Level1Out59[21] , 
        \Level1Out63[5] , \Level8Out0[9] , \Level2Out2[25] , \Level1Out39[16] , 
        \Level1Out60[6] , \Level2Out2[16] , \Level2Out14[9] , 
        \Level1Out59[12] , \ScanLink45[8] , \ScanLink58[7] , \Level2Out26[31] , 
        \Level2Out26[28] , \Level4Out36[31] , \Level4Out60[29] , 
        \Level4Out60[30] , \Level4Out36[28] , \ScanLink2[8] , \Level1Out8[20] , 
        \Level1Out9[8] , \ScanLink17[21] , \ScanLink18[5] , \Level1Out20[4] , 
        \Level1Out23[7] , \Level1Out28[13] , \Level1Out48[17] , 
        \Level2Out6[27] , \Level4Out32[19] , \Level2Out22[19] , 
        \Level1Out28[20] , \Level1Out44[0] , \Level1Out47[3] , 
        \Level1Out48[24] , \Level2Out6[14] , \ScanLink62[11] , 
        \Level2Out52[5] , \ScanLink21[24] , \ScanLink34[10] , \ScanLink41[20] , 
        \ScanLink64[3] , \ScanLink54[14] , \ScanLink13[21] , \Level1Out15[30] , 
        \Level1Out15[29] , \Level1Out38[6] , \Level1Out43[31] , 
        \Level1Out60[19] , \Level1Out25[9] , \Level1Out43[28] , 
        \ScanLink17[12] , \ScanLink21[17] , \Level1Out36[18] , 
        \Level2Out36[1] , \ScanLink54[27] , \ScanLink27[0] , \ScanLink34[23] , 
        \ScanLink62[22] , \ScanLink41[13] , \Level2Out12[5] , 
        \Level4Out48[16] , \Level4Out28[12] , \ScanLink24[3] , 
        \ScanLink30[10] , \Level2Out58[16] , \ScanLink25[24] , 
        \ScanLink45[20] , \ScanLink50[14] , \Level2Out38[12] , 
        \Level4Out24[8] , \Level8Out8[15] , \Level1Out11[30] , 
        \Level1Out11[29] , \Level1Out32[18] , \Level1Out47[31] , 
        \Level1Out47[28] , \ScanLink4[6] , \Level1Out8[13] , \ScanLink43[4] , 
        \Level4Out28[21] , \Level4Out48[25] , \ScanLink13[12] , 
        \ScanLink25[17] , \ScanLink50[27] , \Level2Out38[21] , \ScanLink40[7] , 
        \Level4Load8[0] , \Level8Out8[26] , \ScanLink30[23] , \ScanLink45[13] , 
        \Level2Out58[25] , \Level16Out0[3] , \Level1Out39[27] , 
        \Level1Out60[4] , \Level2Out2[27] , \Level4Out36[19] , 
        \Level4Out60[18] , \Level1Out59[23] , \Level1Out63[7] , 
        \Level2Out26[19] , \Level1Out1[2] , \Level1Out6[24] , \ScanLink7[5] , 
        \ScanLink58[5] , \ScanLink15[2] , \Level1Out15[18] , \ScanLink17[23] , 
        \ScanLink18[7] , \Level1Out20[6] , \Level1Out23[5] , \Level1Load25[0] , 
        \Level1Out59[10] , \Level1Out39[14] , \ScanLink46[9] , 
        \Level2Out2[14] , \Level1Out28[11] , \Level1Out48[15] , 
        \Level2Out6[25] , \Level2Out54[9] , \Level1Out28[22] , 
        \Level1Out48[26] , \Level2Out6[16] , \Level1Out44[2] , 
        \Level1Out47[1] , \Level2Out22[31] , \Level2Out22[28] , 
        \ScanLink21[26] , \Level4Out32[31] , \Level4Out32[28] , 
        \Level1Out38[4] , \ScanLink54[16] , \ScanLink17[10] , \Level1Out26[8] , 
        \ScanLink34[12] , \ScanLink62[13] , \ScanLink41[22] , \ScanLink64[1] , 
        \Level2Out52[7] , \ScanLink62[20] , \ScanLink21[15] , \ScanLink34[21] , 
        \ScanLink41[11] , \ScanLink54[25] , \Level1Out60[28] , 
        \Level1Out36[30] , \Level1Out36[29] , \Level1Out43[19] , 
        \Level1Out60[31] , \Level1Out49[7] , \Level2Out0[5] , \Level2Out36[3] , 
        \Level1Out29[31] , \Level1Out54[8] , \Level2Out20[7] , 
        \Level2Out36[16] , \Level2Out60[17] , \Level8Out24[19] , 
        \Level2Out56[12] , \ScanLink16[1] , \Level1Out29[28] , 
        \Level2Out44[3] , \Level1Out2[1] , \Level1Out6[17] , \ScanLink4[27] , 
        \ScanLink4[14] , \Level1Out52[6] , \Level2Out26[9] , \Level2Out36[25] , 
        \Level2Out56[21] , \Level2Out60[24] , \Level16Out32[22] , 
        \Level1Out14[12] , \Level1Out22[17] , \Level1Out57[27] , 
        \Level4Out4[3] , \Level1Out37[23] , \Level1Out42[13] , 
        \Level1Out51[5] , \Level1Out61[22] , \Level2Out38[5] , 
        \Level2Out48[19] , \Level1Out9[19] , \Level1Out10[10] , 
        \ScanLink12[18] , \Level1Out14[21] , \ScanLink16[30] , 
        \ScanLink35[18] , \Level1Out36[2] , \Level16Out32[11] , 
        \ScanLink16[29] , \ScanLink40[28] , \Level1Out35[1] , 
        \Level1Out37[10] , \ScanLink40[31] , \ScanLink63[19] , 
        \Level1Out42[20] , \Level1Out22[24] , \Level1Out61[11] , 
        \ScanLink31[29] , \ScanLink44[19] , \Level1Out57[14] , 
        \ScanLink31[30] , \Level1Out33[21] , \Level1Out46[11] , 
        \Level2Out8[21] , \Level1Out53[25] , \ScanLink0[16] , \Level1Out11[7] , 
        \Level1Out26[15] , \Level1Out12[4] , \Level1Out26[26] , 
        \ScanLink29[6] , \ScanLink0[25] , \Level1Out10[23] , \Level1Out33[12] , 
        \Level1Out53[16] , \Level1Out46[22] , \ScanLink34[9] , 
        \Level1Load57[0] , \Level2Out8[12] , \Level1Out2[26] , \Level8Out8[3] , 
        \Level1Out2[15] , \ScanLink9[3] , \Level1Out17[9] , \ScanLink19[27] , 
        \ScanLink56[3] , \Level2Out52[10] , \Level4Out56[8] , 
        \Level2Out32[14] , \ScanLink19[14] , \ScanLink55[0] , \Level2Out60[5] , 
        \Level4Out48[4] , \Level2Out32[27] , \Level2Out52[23] , 
        \ScanLink32[7] , \Level1Out58[30] , \Level1Out2[8] , \Level1Out4[6] , 
        \Level1Out7[5] , \ScanLink31[4] , \Level1Out58[29] , \Level1Out14[31] , 
        \ScanLink16[20] , \ScanLink35[11] , \Level2Out42[4] , \Level4Out4[25] , 
        \Level16Out32[18] , \ScanLink40[21] , \Level2Out28[27] , 
        \ScanLink20[25] , \Level1Out28[7] , \ScanLink63[10] , 
        \Level1Out37[19] , \ScanLink55[15] , \Level2Out48[23] , 
        \Level1Out35[8] , \Level1Out42[29] , \ScanLink10[6] , \ScanLink13[5] , 
        \Level1Out14[28] , \Level1Out42[30] , \Level1Out61[18] , 
        \Level4Out4[16] , \ScanLink20[16] , \ScanLink55[26] , \Level2Out6[2] , 
        \Level2Out26[0] , \Level2Out48[10] , \ScanLink16[13] , 
        \ScanLink35[22] , \ScanLink40[12] , \Level2Out28[14] , 
        \ScanLink63[23] , \Level1Out29[12] , \Level1Out30[5] , 
        \Level1Out49[16] , \Level8Out24[23] , \Level1Out9[23] , 
        \Level1Out14[3] , \ScanLink16[8] , \Level1Out33[6] , \Level2Out56[31] , 
        \Level2Out56[28] , \Level1Out54[1] , \Level8Out24[10] , 
        \Level1Out57[2] , \Level4Out16[3] , \Level1Out17[0] , 
        \Level1Out29[21] , \Level1Out38[24] , \Level1Out49[25] , 
        \Level1Out58[20] , \Level4Out32[5] , \Level1Out38[17] , 
        \Level8Out16[24] , \Level8Out40[25] , \Level16Out48[15] , 
        \Level32Out32[16] , \Level1Out58[13] , \Level2Out52[19] , 
        \Level4Out56[1] , \Level8Out40[16] , \Level1Load36[0] , 
        \ScanLink48[6] , \Level8Out16[17] , \Level16Out48[26] , 
        \ScanLink55[9] , \Level32Out32[25] , \Level1Out9[10] , 
        \ScanLink12[22] , \ScanLink24[27] , \ScanLink31[13] , \ScanLink51[17] , 
        \ScanLink34[0] , \ScanLink44[23] , \ScanLink12[11] , \ScanLink31[20] , 
        \ScanLink37[3] , \Level4Out0[27] , \ScanLink44[10] , \ScanLink24[14] , 
        \ScanLink51[24] , \ScanLink50[4] , \Level1Out10[19] , 
        \Level1Out33[28] , \Level1Out46[18] , \Level2Out8[31] , 
        \Level1Out19[6] , \Level1Out33[31] , \Level2Out8[28] , \ScanLink53[7] , 
        \Level4Out0[14] , \ScanLink45[3] , \Level4Out56[27] , 
        \Level32Out0[24] , \Level4Out36[23] , \Level4Out60[22] , 
        \ScanLink0[12] , \ScanLink1[26] , \ScanLink1[15] , \ScanLink2[1] , 
        \Level1Out3[25] , \ScanLink18[24] , \Level2Out10[26] , 
        \Level2Out46[27] , \Level1Out59[19] , \Level2Out26[23] , 
        \Level1Out3[16] , \ScanLink21[7] , \ScanLink46[0] , \Level2Out14[2] , 
        \Level4Out36[10] , \Level4Out60[11] , \Level4Out56[14] , 
        \Level32Out0[17] , \Level8Out0[2] , \ScanLink18[17] , \ScanLink22[4] , 
        \Level2Out10[15] , \Level2Out26[10] , \Level2Out46[14] , 
        \ScanLink1[2] , \Level1Out11[13] , \Level1Out27[16] , 
        \Level1Out52[26] , \Level4Out28[31] , \Level4Out28[28] , 
        \Level1Out32[22] , \Level1Out47[12] , \Level4Out40[5] , 
        \Level32Out32[6] , \Level2Out38[31] , \Level2Out38[28] , 
        \Level1Out2[22] , \ScanLink5[24] , \ScanLink5[17] , \Level1Out8[30] , 
        \Level1Out11[20] , \ScanLink13[31] , \ScanLink13[28] , \ScanLink27[9] , 
        \Level1Load44[0] , \ScanLink30[19] , \ScanLink45[30] , 
        \ScanLink45[29] , \Level1Out27[25] , \Level1Out32[11] , 
        \Level1Out47[21] , \Level4Out24[1] , \Level1Out8[29] , 
        \Level1Out52[15] , \Level2Load28[0] , \Level1Out15[11] , 
        \ScanLink17[19] , \ScanLink39[5] , \ScanLink62[29] , \Level2Out28[6] , 
        \ScanLink34[31] , \ScanLink34[28] , \ScanLink41[18] , \ScanLink62[30] , 
        \Level1Out60[21] , \Level1Out23[14] , \Level1Out36[20] , 
        \Level1Out43[10] , \Level1Out56[24] , \Level1Out41[6] , 
        \Level2Out8[4] , \Level1Out9[3] , \Level1Out15[22] , \Level1Out23[27] , 
        \Level1Out42[5] , \Level1Out56[17] , \Level1Out25[2] , 
        \Level1Out36[13] , \Level1Out60[12] , \Level1Out43[23] , 
        \ScanLink64[8] , \Level1Out7[27] , \Level1Out26[1] , \Level1Out7[14] , 
        \Level1Out28[18] , \Level1Out47[8] , \Level2Out14[24] , 
        \Level2Out22[21] , \Level2Out42[25] , \Level1Out59[4] , 
        \Level2Out30[4] , \Level4Out32[21] , \ScanLink62[6] , \Level2Load2[0] , 
        \Level2Out14[17] , \Level2Out42[16] , \Level4Out52[25] , 
        \Level2Out22[12] , \ScanLink9[7] , \ScanLink55[4] , \ScanLink61[5] , 
        \Level4Out52[16] , \Level2Out54[0] , \Level4Out32[12] , 
        \Level2Out60[1] , \Level4Out48[0] , \Level32Out32[28] , 
        \Level32Out32[31] , \ScanLink19[23] , \Level2Out32[10] , 
        \Level2Out52[14] , \Level1Out2[11] , \ScanLink31[0] , \ScanLink56[7] , 
        \Level8Out16[30] , \Level8Out16[29] , \Level8Out40[31] , 
        \Level8Out40[28] , \Level16Out48[18] , \Level1Out12[0] , 
        \ScanLink19[10] , \ScanLink32[3] , \Level1Out38[30] , 
        \Level1Out38[29] , \Level2Out32[23] , \Level2Out52[27] , 
        \Level4Out0[19] , \Level4Out32[8] , \Level1Out53[21] , \ScanLink0[21] , 
        \Level1Out10[14] , \Level1Out11[3] , \Level1Out26[11] , 
        \Level2Out8[25] , \ScanLink24[19] , \Level1Load33[0] , 
        \Level1Out33[25] , \Level1Out46[15] , \ScanLink51[29] , 
        \ScanLink50[9] , \ScanLink51[30] , \Level1Out10[27] , \Level8Out8[7] , 
        \Level1Out26[22] , \Level1Out33[16] , \Level2Out8[16] , 
        \Level1Out46[26] , \Level1Out1[6] , \Level1Out2[5] , \ScanLink4[23] , 
        \ScanLink4[10] , \Level1Out14[16] , \ScanLink29[2] , \Level1Out53[12] , 
        \Level1Out61[26] , \Level2Out28[19] , \Level2Out38[1] , 
        \Level1Out22[13] , \Level1Out37[27] , \Level1Out42[17] , 
        \Level1Out57[23] , \Level4Out4[7] , \Level1Out51[1] , 
        \Level16Out32[26] , \ScanLink13[8] , \Level1Out52[2] , 
        \Level1Out14[25] , \Level1Out22[20] , \Level1Out57[10] , 
        \ScanLink20[31] , \ScanLink20[28] , \Level1Out35[5] , 
        \Level1Out37[14] , \Level1Out61[15] , \Level1Out42[24] , 
        \ScanLink55[18] , \Level4Out4[31] , \Level4Out4[28] , \Level1Out6[20] , 
        \Level1Out7[8] , \Level1Out36[6] , \Level2Out42[9] , 
        \Level16Out32[15] , \ScanLink15[6] , \ScanLink16[5] , 
        \Level1Out49[31] , \Level1Out49[28] , \Level2Out20[3] , 
        \Level2Out36[12] , \Level2Out56[16] , \Level2Out60[13] , 
        \Level1Out49[3] , \Level2Out0[1] , \Level2Out36[21] , 
        \Level2Out60[20] , \Level1Out6[13] , \Level2Out56[25] , 
        \Level1Out3[31] , \Level1Out3[28] , \ScanLink5[30] , \Level1Load19[0] , 
        \Level1Out30[8] , \Level2Out44[7] , \ScanLink5[29] , \Level1Out7[19] , 
        \ScanLink17[27] , \ScanLink34[16] , \Level2Out52[3] , \ScanLink41[26] , 
        \ScanLink64[5] , \ScanLink17[14] , \ScanLink21[22] , \Level1Out38[0] , 
        \ScanLink62[17] , \ScanLink21[11] , \Level1Out23[19] , 
        \Level1Out42[8] , \ScanLink54[12] , \Level2Out36[7] , 
        \Level1Out56[30] , \Level1Out56[29] , \Level2Out8[9] , 
        \ScanLink54[21] , \ScanLink34[25] , \ScanLink41[15] , \ScanLink62[24] , 
        \Level1Out20[2] , \Level1Out48[11] , \ScanLink61[8] , \Level2Out6[21] , 
        \ScanLink18[3] , \Level1Out23[1] , \Level1Out28[15] , \Level1Out59[9] , 
        \Level4Out52[31] , \Level4Out52[28] , \ScanLink22[9] , 
        \Level1Out28[26] , \Level1Out44[6] , \Level2Out30[9] , 
        \Level1Out47[5] , \Level2Out42[31] , \Level2Out14[30] , 
        \Level2Out14[29] , \Level2Out42[28] , \Level1Out39[23] , 
        \Level1Out48[22] , \Level1Out59[27] , \Level1Out63[3] , 
        \Level2Out6[12] , \Level2Out10[18] , \Level2Out46[19] , 
        \Level1Load41[0] , \Level1Out39[10] , \Level1Out60[0] , 
        \Level2Out2[23] , \Level4Out56[19] , \Level2Out2[10] , \ScanLink4[2] , 
        \ScanLink7[1] , \ScanLink18[30] , \Level1Out59[14] , \ScanLink18[29] , 
        \ScanLink58[1] , \Level32Out0[30] , \Level32Out0[29] , \ScanLink0[31] , 
        \ScanLink0[28] , \ScanLink1[22] , \ScanLink1[18] , \Level1Out8[24] , 
        \Level1Out8[17] , \ScanLink13[25] , \ScanLink24[7] , \ScanLink25[20] , 
        \Level1Out27[31] , \Level1Out27[28] , \ScanLink39[8] , 
        \Level1Out52[18] , \Level8Out8[11] , \ScanLink30[14] , 
        \ScanLink50[10] , \Level2Out38[16] , \Level2Out58[12] , 
        \ScanLink45[24] , \ScanLink13[16] , \ScanLink27[4] , \ScanLink30[27] , 
        \ScanLink45[17] , \Level2Out12[1] , \Level4Out28[16] , 
        \Level4Out48[12] , \Level2Out58[21] , \Level16Out0[7] , 
        \ScanLink25[13] , \ScanLink50[23] , \Level8Out8[22] , 
        \Level2Out38[25] , \ScanLink40[3] , \Level4Out40[8] , 
        \Level4Out48[21] , \ScanLink1[11] , \ScanLink1[6] , \ScanLink5[20] , 
        \ScanLink5[13] , \Level1Out7[23] , \ScanLink43[0] , \Level4Out28[25] , 
        \Level1Out59[0] , \Level2Load14[0] , \Level4Out32[25] , 
        \Level4Out52[21] , \Level2Out14[20] , \Level2Out30[0] , 
        \Level2Out22[25] , \Level2Out42[21] , \Level1Out7[10] , 
        \ScanLink61[1] , \Level2Out54[4] , \Level4Out32[16] , 
        \Level4Out52[12] , \Level1Out23[8] , \Level1Out48[18] , 
        \ScanLink62[2] , \Level2Out6[31] , \Level2Out6[28] , \Level2Out22[16] , 
        \Level1Out42[1] , \Level2Out14[13] , \Level2Out42[12] , 
        \Level1Out15[15] , \Level1Out23[10] , \Level1Out56[20] , 
        \Level2Out8[0] , \Level1Out36[24] , \Level1Out41[2] , 
        \Level1Out43[14] , \Level1Out60[25] , \ScanLink21[18] , 
        \ScanLink54[31] , \Level2Out28[2] , \ScanLink54[28] , \Level1Out9[7] , 
        \Level1Out26[5] , \Level1Out38[9] , \Level1Out15[26] , 
        \Level1Out25[6] , \Level1Out36[17] , \Level1Out43[27] , 
        \Level1Out23[23] , \Level1Out60[16] , \Level1Out56[13] , 
        \Level1Out11[17] , \Level1Out32[26] , \Level1Out47[16] , 
        \Level2Out58[31] , \Level2Out58[28] , \Level4Out40[1] , 
        \Level32Out32[2] , \Level1Out27[12] , \Level1Out52[22] , 
        \ScanLink2[5] , \Level1Load20[0] , \Level4Out48[31] , 
        \Level4Out48[28] , \ScanLink43[9] , \Level1Out11[24] , 
        \Level1Out27[21] , \ScanLink39[1] , \Level1Out32[15] , 
        \Level1Out52[11] , \Level4Out24[5] , \Level1Out47[25] , 
        \ScanLink25[30] , \ScanLink25[29] , \Level8Out8[18] , \ScanLink50[19] , 
        \Level1Out3[21] , \Level2Out12[8] , \Level1Out3[12] , \ScanLink7[8] , 
        \ScanLink46[4] , \ScanLink18[20] , \Level1Out39[19] , \Level2Out2[19] , 
        \Level2Out26[27] , \ScanLink18[13] , \Level1Out19[2] , \ScanLink45[7] , 
        \ScanLink58[8] , \Level2Out10[22] , \Level2Out46[23] , 
        \Level4Out36[27] , \Level4Out60[26] , \Level32Out0[20] , 
        \Level2Out10[11] , \Level4Out56[23] , \Level2Out26[14] , 
        \Level2Out46[10] , \ScanLink22[0] , \ScanLink21[3] , \Level8Out0[6] , 
        \Level32Out0[13] , \Level1Out60[9] , \Level2Out14[6] , 
        \Level4Out36[14] , \Level4Out56[10] , \Level4Out60[15] , 
        \Level1Out2[18] , \Level1Out9[27] , \ScanLink12[26] , \ScanLink37[7] , 
        \Level4Out0[23] , \ScanLink24[23] , \ScanLink31[17] , \ScanLink34[4] , 
        \ScanLink44[27] , \ScanLink51[13] , \Level1Out9[14] , \Level1Out12[9] , 
        \ScanLink53[3] , \Level4Out0[10] , \Level1Out26[18] , 
        \Level1Out53[28] , \Level1Out53[31] , \ScanLink12[15] , 
        \ScanLink24[10] , \ScanLink51[20] , \ScanLink50[0] , \ScanLink31[24] , 
        \ScanLink44[14] , \ScanLink31[9] , \Level1Load52[0] , 
        \Level8Out16[20] , \Level8Out40[21] , \Level16Out48[11] , 
        \Level1Out38[20] , \Level32Out32[12] , \Level1Out58[24] , 
        \ScanLink4[19] , \Level1Out4[2] , \Level1Out6[30] , \Level1Out14[7] , 
        \ScanLink19[19] , \Level4Out32[1] , \ScanLink48[2] , \Level4Out48[9] , 
        \Level32Out32[21] , \Level16Out48[22] , \Level2Out60[8] , 
        \Level8Out16[13] , \Level1Out17[4] , \Level2Out32[19] , 
        \Level4Out56[5] , \Level8Out40[12] , \Level1Out29[16] , 
        \Level1Out33[2] , \Level1Out38[13] , \Level1Out58[17] , 
        \Level2Out36[31] , \Level2Out36[28] , \Level2Out60[30] , 
        \Level2Out60[29] , \Level1Out30[1] , \Level1Out49[12] , 
        \Level8Out24[27] , \Level1Out49[21] , \Level1Out6[29] , 
        \Level1Out29[25] , \Level1Out54[5] , \Level1Out57[6] , 
        \Level4Out16[7] , \Level2Out0[8] , \Level8Out24[14] , \Level1Out7[1] , 
        \ScanLink16[24] , \ScanLink20[21] , \Level1Out22[30] , 
        \Level1Out22[29] , \Level1Out57[19] , \Level1Out28[3] , 
        \ScanLink55[11] , \Level2Out48[27] , \ScanLink35[15] , 
        \ScanLink63[14] , \ScanLink40[25] , \Level2Out28[23] , 
        \Level2Out42[0] , \Level4Out4[21] , \ScanLink10[2] , \ScanLink16[17] , 
        \ScanLink63[27] , \Level2Out38[8] , \ScanLink20[12] , \ScanLink35[26] , 
        \ScanLink40[16] , \Level2Out28[10] , \ScanLink55[22] , 
        \Level2Out48[14] , \Level1Out51[8] , \Level2Out26[4] , \Level2Out6[6] , 
        \Level4Out4[12] , \ScanLink13[1] ;
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_1 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink1[31] , \ScanLink1[30] , 
        \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , \ScanLink1[26] , 
        \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , \ScanLink1[22] , 
        \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , \ScanLink1[18] , 
        \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , \ScanLink1[14] , 
        \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , \ScanLink1[10] , 
        \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , \ScanLink1[6] , 
        \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , \ScanLink1[2] , 
        \ScanLink1[1] , \ScanLink1[0] }), .ScanOut({\ScanLink2[31] , 
        \ScanLink2[30] , \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , 
        \ScanLink2[26] , \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , 
        \ScanLink2[22] , \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , 
        \ScanLink2[18] , \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , 
        \ScanLink2[14] , \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , 
        \ScanLink2[10] , \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , 
        \ScanLink2[6] , \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , 
        \ScanLink2[2] , \ScanLink2[1] , \ScanLink2[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load1[0] ), .Out({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_21 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink21[31] , \ScanLink21[30] , 
        \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , \ScanLink21[26] , 
        \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , \ScanLink21[22] , 
        \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , \ScanLink21[18] , 
        \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , \ScanLink21[14] , 
        \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , \ScanLink21[10] , 
        \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , \ScanLink21[6] , 
        \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , \ScanLink21[2] , 
        \ScanLink21[1] , \ScanLink21[0] }), .ScanOut({\ScanLink22[31] , 
        \ScanLink22[30] , \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , 
        \ScanLink22[26] , \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , 
        \ScanLink22[22] , \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , 
        \ScanLink22[18] , \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , 
        \ScanLink22[14] , \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , 
        \ScanLink22[10] , \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , 
        \ScanLink22[6] , \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , 
        \ScanLink22[2] , \ScanLink22[1] , \ScanLink22[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load21[0] ), .Out({
        \Level1Out21[31] , \Level1Out21[30] , \Level1Out21[29] , 
        \Level1Out21[28] , \Level1Out21[27] , \Level1Out21[26] , 
        \Level1Out21[25] , \Level1Out21[24] , \Level1Out21[23] , 
        \Level1Out21[22] , \Level1Out21[21] , \Level1Out21[20] , 
        \Level1Out21[19] , \Level1Out21[18] , \Level1Out21[17] , 
        \Level1Out21[16] , \Level1Out21[15] , \Level1Out21[14] , 
        \Level1Out21[13] , \Level1Out21[12] , \Level1Out21[11] , 
        \Level1Out21[10] , \Level1Out21[9] , \Level1Out21[8] , 
        \Level1Out21[7] , \Level1Out21[6] , \Level1Out21[5] , \Level1Out21[4] , 
        \Level1Out21[3] , \Level1Out21[2] , \Level1Out21[1] , \Level1Out21[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_36_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load36[0] ), .Out({\Level2Out36[31] , \Level2Out36[30] , 
        \Level2Out36[29] , \Level2Out36[28] , \Level2Out36[27] , 
        \Level2Out36[26] , \Level2Out36[25] , \Level2Out36[24] , 
        \Level2Out36[23] , \Level2Out36[22] , \Level2Out36[21] , 
        \Level2Out36[20] , \Level2Out36[19] , \Level2Out36[18] , 
        \Level2Out36[17] , \Level2Out36[16] , \Level2Out36[15] , 
        \Level2Out36[14] , \Level2Out36[13] , \Level2Out36[12] , 
        \Level2Out36[11] , \Level2Out36[10] , \Level2Out36[9] , 
        \Level2Out36[8] , \Level2Out36[7] , \Level2Out36[6] , \Level2Out36[5] , 
        \Level2Out36[4] , \Level2Out36[3] , \Level2Out36[2] , \Level2Out36[1] , 
        \Level2Out36[0] }), .In1({\Level1Out36[31] , \Level1Out36[30] , 
        \Level1Out36[29] , \Level1Out36[28] , \Level1Out36[27] , 
        \Level1Out36[26] , \Level1Out36[25] , \Level1Out36[24] , 
        \Level1Out36[23] , \Level1Out36[22] , \Level1Out36[21] , 
        \Level1Out36[20] , \Level1Out36[19] , \Level1Out36[18] , 
        \Level1Out36[17] , \Level1Out36[16] , \Level1Out36[15] , 
        \Level1Out36[14] , \Level1Out36[13] , \Level1Out36[12] , 
        \Level1Out36[11] , \Level1Out36[10] , \Level1Out36[9] , 
        \Level1Out36[8] , \Level1Out36[7] , \Level1Out36[6] , \Level1Out36[5] , 
        \Level1Out36[4] , \Level1Out36[3] , \Level1Out36[2] , \Level1Out36[1] , 
        \Level1Out36[0] }), .In2({\Level1Out37[31] , \Level1Out37[30] , 
        \Level1Out37[29] , \Level1Out37[28] , \Level1Out37[27] , 
        \Level1Out37[26] , \Level1Out37[25] , \Level1Out37[24] , 
        \Level1Out37[23] , \Level1Out37[22] , \Level1Out37[21] , 
        \Level1Out37[20] , \Level1Out37[19] , \Level1Out37[18] , 
        \Level1Out37[17] , \Level1Out37[16] , \Level1Out37[15] , 
        \Level1Out37[14] , \Level1Out37[13] , \Level1Out37[12] , 
        \Level1Out37[11] , \Level1Out37[10] , \Level1Out37[9] , 
        \Level1Out37[8] , \Level1Out37[7] , \Level1Out37[6] , \Level1Out37[5] , 
        \Level1Out37[4] , \Level1Out37[3] , \Level1Out37[2] , \Level1Out37[1] , 
        \Level1Out37[0] }), .Read1(\Level1Load36[0] ), .Read2(
        \Level1Load37[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_54 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink54[31] , \ScanLink54[30] , 
        \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , \ScanLink54[26] , 
        \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , \ScanLink54[22] , 
        \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , \ScanLink54[18] , 
        \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , \ScanLink54[14] , 
        \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , \ScanLink54[10] , 
        \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , \ScanLink54[6] , 
        \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , \ScanLink54[2] , 
        \ScanLink54[1] , \ScanLink54[0] }), .ScanOut({\ScanLink55[31] , 
        \ScanLink55[30] , \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , 
        \ScanLink55[26] , \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , 
        \ScanLink55[22] , \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , 
        \ScanLink55[18] , \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , 
        \ScanLink55[14] , \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , 
        \ScanLink55[10] , \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , 
        \ScanLink55[6] , \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , 
        \ScanLink55[2] , \ScanLink55[1] , \ScanLink55[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load54[0] ), .Out({
        \Level1Out54[31] , \Level1Out54[30] , \Level1Out54[29] , 
        \Level1Out54[28] , \Level1Out54[27] , \Level1Out54[26] , 
        \Level1Out54[25] , \Level1Out54[24] , \Level1Out54[23] , 
        \Level1Out54[22] , \Level1Out54[21] , \Level1Out54[20] , 
        \Level1Out54[19] , \Level1Out54[18] , \Level1Out54[17] , 
        \Level1Out54[16] , \Level1Out54[15] , \Level1Out54[14] , 
        \Level1Out54[13] , \Level1Out54[12] , \Level1Out54[11] , 
        \Level1Out54[10] , \Level1Out54[9] , \Level1Out54[8] , 
        \Level1Out54[7] , \Level1Out54[6] , \Level1Out54[5] , \Level1Out54[4] , 
        \Level1Out54[3] , \Level1Out54[2] , \Level1Out54[1] , \Level1Out54[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load32[0] ), .Out({\Level4Out32[31] , \Level4Out32[30] , 
        \Level4Out32[29] , \Level4Out32[28] , \Level4Out32[27] , 
        \Level4Out32[26] , \Level4Out32[25] , \Level4Out32[24] , 
        \Level4Out32[23] , \Level4Out32[22] , \Level4Out32[21] , 
        \Level4Out32[20] , \Level4Out32[19] , \Level4Out32[18] , 
        \Level4Out32[17] , \Level4Out32[16] , \Level4Out32[15] , 
        \Level4Out32[14] , \Level4Out32[13] , \Level4Out32[12] , 
        \Level4Out32[11] , \Level4Out32[10] , \Level4Out32[9] , 
        \Level4Out32[8] , \Level4Out32[7] , \Level4Out32[6] , \Level4Out32[5] , 
        \Level4Out32[4] , \Level4Out32[3] , \Level4Out32[2] , \Level4Out32[1] , 
        \Level4Out32[0] }), .In1({\Level2Out32[31] , \Level2Out32[30] , 
        \Level2Out32[29] , \Level2Out32[28] , \Level2Out32[27] , 
        \Level2Out32[26] , \Level2Out32[25] , \Level2Out32[24] , 
        \Level2Out32[23] , \Level2Out32[22] , \Level2Out32[21] , 
        \Level2Out32[20] , \Level2Out32[19] , \Level2Out32[18] , 
        \Level2Out32[17] , \Level2Out32[16] , \Level2Out32[15] , 
        \Level2Out32[14] , \Level2Out32[13] , \Level2Out32[12] , 
        \Level2Out32[11] , \Level2Out32[10] , \Level2Out32[9] , 
        \Level2Out32[8] , \Level2Out32[7] , \Level2Out32[6] , \Level2Out32[5] , 
        \Level2Out32[4] , \Level2Out32[3] , \Level2Out32[2] , \Level2Out32[1] , 
        \Level2Out32[0] }), .In2({\Level2Out34[31] , \Level2Out34[30] , 
        \Level2Out34[29] , \Level2Out34[28] , \Level2Out34[27] , 
        \Level2Out34[26] , \Level2Out34[25] , \Level2Out34[24] , 
        \Level2Out34[23] , \Level2Out34[22] , \Level2Out34[21] , 
        \Level2Out34[20] , \Level2Out34[19] , \Level2Out34[18] , 
        \Level2Out34[17] , \Level2Out34[16] , \Level2Out34[15] , 
        \Level2Out34[14] , \Level2Out34[13] , \Level2Out34[12] , 
        \Level2Out34[11] , \Level2Out34[10] , \Level2Out34[9] , 
        \Level2Out34[8] , \Level2Out34[7] , \Level2Out34[6] , \Level2Out34[5] , 
        \Level2Out34[4] , \Level2Out34[3] , \Level2Out34[2] , \Level2Out34[1] , 
        \Level2Out34[0] }), .Read1(\Level2Load32[0] ), .Read2(
        \Level2Load34[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_0 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink0[31] , \ScanLink0[30] , 
        \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , \ScanLink0[26] , 
        \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , \ScanLink0[22] , 
        \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , \ScanLink0[18] , 
        \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , \ScanLink0[14] , 
        \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , \ScanLink0[10] , 
        \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , \ScanLink0[6] , 
        \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , \ScanLink0[2] , 
        \ScanLink0[1] , \ScanLink0[0] }), .ScanOut({\ScanLink1[31] , 
        \ScanLink1[30] , \ScanLink1[29] , \ScanLink1[28] , \ScanLink1[27] , 
        \ScanLink1[26] , \ScanLink1[25] , \ScanLink1[24] , \ScanLink1[23] , 
        \ScanLink1[22] , \ScanLink1[21] , \ScanLink1[20] , \ScanLink1[19] , 
        \ScanLink1[18] , \ScanLink1[17] , \ScanLink1[16] , \ScanLink1[15] , 
        \ScanLink1[14] , \ScanLink1[13] , \ScanLink1[12] , \ScanLink1[11] , 
        \ScanLink1[10] , \ScanLink1[9] , \ScanLink1[8] , \ScanLink1[7] , 
        \ScanLink1[6] , \ScanLink1[5] , \ScanLink1[4] , \ScanLink1[3] , 
        \ScanLink1[2] , \ScanLink1[1] , \ScanLink1[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load0[0] ), .Out({
        \Level1Out0[31] , \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , 
        \Level1Out0[27] , \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , 
        \Level1Out0[23] , \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , 
        \Level1Out0[19] , \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , 
        \Level1Out0[15] , \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , 
        \Level1Out0[11] , \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , 
        \Level1Out0[7] , \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , 
        \Level1Out0[3] , \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_6 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink6[31] , \ScanLink6[30] , 
        \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , \ScanLink6[26] , 
        \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , \ScanLink6[22] , 
        \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , \ScanLink6[18] , 
        \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , \ScanLink6[14] , 
        \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , \ScanLink6[10] , 
        \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , \ScanLink6[6] , 
        \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , \ScanLink6[2] , 
        \ScanLink6[1] , \ScanLink6[0] }), .ScanOut({\ScanLink7[31] , 
        \ScanLink7[30] , \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , 
        \ScanLink7[26] , \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , 
        \ScanLink7[22] , \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , 
        \ScanLink7[18] , \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , 
        \ScanLink7[14] , \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , 
        \ScanLink7[10] , \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , 
        \ScanLink7[6] , \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , 
        \ScanLink7[2] , \ScanLink7[1] , \ScanLink7[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load6[0] ), .Out({
        \Level1Out6[31] , \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , 
        \Level1Out6[27] , \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , 
        \Level1Out6[23] , \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , 
        \Level1Out6[19] , \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , 
        \Level1Out6[15] , \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , 
        \Level1Out6[11] , \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , 
        \Level1Out6[7] , \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , 
        \Level1Out6[3] , \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_8 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink8[31] , \ScanLink8[30] , 
        \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , \ScanLink8[26] , 
        \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , \ScanLink8[22] , 
        \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , \ScanLink8[18] , 
        \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , \ScanLink8[14] , 
        \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , \ScanLink8[10] , 
        \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , \ScanLink8[6] , 
        \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , \ScanLink8[2] , 
        \ScanLink8[1] , \ScanLink8[0] }), .ScanOut({\ScanLink9[31] , 
        \ScanLink9[30] , \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , 
        \ScanLink9[26] , \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , 
        \ScanLink9[22] , \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , 
        \ScanLink9[18] , \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , 
        \ScanLink9[14] , \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , 
        \ScanLink9[10] , \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , 
        \ScanLink9[6] , \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , 
        \ScanLink9[2] , \ScanLink9[1] , \ScanLink9[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load8[0] ), .Out({
        \Level1Out8[31] , \Level1Out8[30] , \Level1Out8[29] , \Level1Out8[28] , 
        \Level1Out8[27] , \Level1Out8[26] , \Level1Out8[25] , \Level1Out8[24] , 
        \Level1Out8[23] , \Level1Out8[22] , \Level1Out8[21] , \Level1Out8[20] , 
        \Level1Out8[19] , \Level1Out8[18] , \Level1Out8[17] , \Level1Out8[16] , 
        \Level1Out8[15] , \Level1Out8[14] , \Level1Out8[13] , \Level1Out8[12] , 
        \Level1Out8[11] , \Level1Out8[10] , \Level1Out8[9] , \Level1Out8[8] , 
        \Level1Out8[7] , \Level1Out8[6] , \Level1Out8[5] , \Level1Out8[4] , 
        \Level1Out8[3] , \Level1Out8[2] , \Level1Out8[1] , \Level1Out8[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_28 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink28[31] , \ScanLink28[30] , 
        \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , \ScanLink28[26] , 
        \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , \ScanLink28[22] , 
        \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , \ScanLink28[18] , 
        \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , \ScanLink28[14] , 
        \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , \ScanLink28[10] , 
        \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , \ScanLink28[6] , 
        \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , \ScanLink28[2] , 
        \ScanLink28[1] , \ScanLink28[0] }), .ScanOut({\ScanLink29[31] , 
        \ScanLink29[30] , \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , 
        \ScanLink29[26] , \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , 
        \ScanLink29[22] , \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , 
        \ScanLink29[18] , \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , 
        \ScanLink29[14] , \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , 
        \ScanLink29[10] , \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , 
        \ScanLink29[6] , \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , 
        \ScanLink29[2] , \ScanLink29[1] , \ScanLink29[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load28[0] ), .Out({
        \Level1Out28[31] , \Level1Out28[30] , \Level1Out28[29] , 
        \Level1Out28[28] , \Level1Out28[27] , \Level1Out28[26] , 
        \Level1Out28[25] , \Level1Out28[24] , \Level1Out28[23] , 
        \Level1Out28[22] , \Level1Out28[21] , \Level1Out28[20] , 
        \Level1Out28[19] , \Level1Out28[18] , \Level1Out28[17] , 
        \Level1Out28[16] , \Level1Out28[15] , \Level1Out28[14] , 
        \Level1Out28[13] , \Level1Out28[12] , \Level1Out28[11] , 
        \Level1Out28[10] , \Level1Out28[9] , \Level1Out28[8] , 
        \Level1Out28[7] , \Level1Out28[6] , \Level1Out28[5] , \Level1Out28[4] , 
        \Level1Out28[3] , \Level1Out28[2] , \Level1Out28[1] , \Level1Out28[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load48[0] ), .Out({\Level4Out48[31] , \Level4Out48[30] , 
        \Level4Out48[29] , \Level4Out48[28] , \Level4Out48[27] , 
        \Level4Out48[26] , \Level4Out48[25] , \Level4Out48[24] , 
        \Level4Out48[23] , \Level4Out48[22] , \Level4Out48[21] , 
        \Level4Out48[20] , \Level4Out48[19] , \Level4Out48[18] , 
        \Level4Out48[17] , \Level4Out48[16] , \Level4Out48[15] , 
        \Level4Out48[14] , \Level4Out48[13] , \Level4Out48[12] , 
        \Level4Out48[11] , \Level4Out48[10] , \Level4Out48[9] , 
        \Level4Out48[8] , \Level4Out48[7] , \Level4Out48[6] , \Level4Out48[5] , 
        \Level4Out48[4] , \Level4Out48[3] , \Level4Out48[2] , \Level4Out48[1] , 
        \Level4Out48[0] }), .In1({\Level2Out48[31] , \Level2Out48[30] , 
        \Level2Out48[29] , \Level2Out48[28] , \Level2Out48[27] , 
        \Level2Out48[26] , \Level2Out48[25] , \Level2Out48[24] , 
        \Level2Out48[23] , \Level2Out48[22] , \Level2Out48[21] , 
        \Level2Out48[20] , \Level2Out48[19] , \Level2Out48[18] , 
        \Level2Out48[17] , \Level2Out48[16] , \Level2Out48[15] , 
        \Level2Out48[14] , \Level2Out48[13] , \Level2Out48[12] , 
        \Level2Out48[11] , \Level2Out48[10] , \Level2Out48[9] , 
        \Level2Out48[8] , \Level2Out48[7] , \Level2Out48[6] , \Level2Out48[5] , 
        \Level2Out48[4] , \Level2Out48[3] , \Level2Out48[2] , \Level2Out48[1] , 
        \Level2Out48[0] }), .In2({\Level2Out50[31] , \Level2Out50[30] , 
        \Level2Out50[29] , \Level2Out50[28] , \Level2Out50[27] , 
        \Level2Out50[26] , \Level2Out50[25] , \Level2Out50[24] , 
        \Level2Out50[23] , \Level2Out50[22] , \Level2Out50[21] , 
        \Level2Out50[20] , \Level2Out50[19] , \Level2Out50[18] , 
        \Level2Out50[17] , \Level2Out50[16] , \Level2Out50[15] , 
        \Level2Out50[14] , \Level2Out50[13] , \Level2Out50[12] , 
        \Level2Out50[11] , \Level2Out50[10] , \Level2Out50[9] , 
        \Level2Out50[8] , \Level2Out50[7] , \Level2Out50[6] , \Level2Out50[5] , 
        \Level2Out50[4] , \Level2Out50[3] , \Level2Out50[2] , \Level2Out50[1] , 
        \Level2Out50[0] }), .Read1(\Level2Load48[0] ), .Read2(
        \Level2Load50[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_46 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink46[31] , \ScanLink46[30] , 
        \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , \ScanLink46[26] , 
        \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , \ScanLink46[22] , 
        \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , \ScanLink46[18] , 
        \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , \ScanLink46[14] , 
        \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , \ScanLink46[10] , 
        \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , \ScanLink46[6] , 
        \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , \ScanLink46[2] , 
        \ScanLink46[1] , \ScanLink46[0] }), .ScanOut({\ScanLink47[31] , 
        \ScanLink47[30] , \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , 
        \ScanLink47[26] , \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , 
        \ScanLink47[22] , \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , 
        \ScanLink47[18] , \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , 
        \ScanLink47[14] , \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , 
        \ScanLink47[10] , \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , 
        \ScanLink47[6] , \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , 
        \ScanLink47[2] , \ScanLink47[1] , \ScanLink47[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load46[0] ), .Out({
        \Level1Out46[31] , \Level1Out46[30] , \Level1Out46[29] , 
        \Level1Out46[28] , \Level1Out46[27] , \Level1Out46[26] , 
        \Level1Out46[25] , \Level1Out46[24] , \Level1Out46[23] , 
        \Level1Out46[22] , \Level1Out46[21] , \Level1Out46[20] , 
        \Level1Out46[19] , \Level1Out46[18] , \Level1Out46[17] , 
        \Level1Out46[16] , \Level1Out46[15] , \Level1Out46[14] , 
        \Level1Out46[13] , \Level1Out46[12] , \Level1Out46[11] , 
        \Level1Out46[10] , \Level1Out46[9] , \Level1Out46[8] , 
        \Level1Out46[7] , \Level1Out46[6] , \Level1Out46[5] , \Level1Out46[4] , 
        \Level1Out46[3] , \Level1Out46[2] , \Level1Out46[1] , \Level1Out46[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_61 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink61[31] , \ScanLink61[30] , 
        \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , \ScanLink61[26] , 
        \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , \ScanLink61[22] , 
        \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , \ScanLink61[18] , 
        \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , \ScanLink61[14] , 
        \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , \ScanLink61[10] , 
        \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , \ScanLink61[6] , 
        \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , \ScanLink61[2] , 
        \ScanLink61[1] , \ScanLink61[0] }), .ScanOut({\ScanLink62[31] , 
        \ScanLink62[30] , \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , 
        \ScanLink62[26] , \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , 
        \ScanLink62[22] , \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , 
        \ScanLink62[18] , \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , 
        \ScanLink62[14] , \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , 
        \ScanLink62[10] , \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , 
        \ScanLink62[6] , \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , 
        \ScanLink62[2] , \ScanLink62[1] , \ScanLink62[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load61[0] ), .Out({
        \Level1Out61[31] , \Level1Out61[30] , \Level1Out61[29] , 
        \Level1Out61[28] , \Level1Out61[27] , \Level1Out61[26] , 
        \Level1Out61[25] , \Level1Out61[24] , \Level1Out61[23] , 
        \Level1Out61[22] , \Level1Out61[21] , \Level1Out61[20] , 
        \Level1Out61[19] , \Level1Out61[18] , \Level1Out61[17] , 
        \Level1Out61[16] , \Level1Out61[15] , \Level1Out61[14] , 
        \Level1Out61[13] , \Level1Out61[12] , \Level1Out61[11] , 
        \Level1Out61[10] , \Level1Out61[9] , \Level1Out61[8] , 
        \Level1Out61[7] , \Level1Out61[6] , \Level1Out61[5] , \Level1Out61[4] , 
        \Level1Out61[3] , \Level1Out61[2] , \Level1Out61[1] , \Level1Out61[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_54_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load54[0] ), .Out({\Level2Out54[31] , \Level2Out54[30] , 
        \Level2Out54[29] , \Level2Out54[28] , \Level2Out54[27] , 
        \Level2Out54[26] , \Level2Out54[25] , \Level2Out54[24] , 
        \Level2Out54[23] , \Level2Out54[22] , \Level2Out54[21] , 
        \Level2Out54[20] , \Level2Out54[19] , \Level2Out54[18] , 
        \Level2Out54[17] , \Level2Out54[16] , \Level2Out54[15] , 
        \Level2Out54[14] , \Level2Out54[13] , \Level2Out54[12] , 
        \Level2Out54[11] , \Level2Out54[10] , \Level2Out54[9] , 
        \Level2Out54[8] , \Level2Out54[7] , \Level2Out54[6] , \Level2Out54[5] , 
        \Level2Out54[4] , \Level2Out54[3] , \Level2Out54[2] , \Level2Out54[1] , 
        \Level2Out54[0] }), .In1({\Level1Out54[31] , \Level1Out54[30] , 
        \Level1Out54[29] , \Level1Out54[28] , \Level1Out54[27] , 
        \Level1Out54[26] , \Level1Out54[25] , \Level1Out54[24] , 
        \Level1Out54[23] , \Level1Out54[22] , \Level1Out54[21] , 
        \Level1Out54[20] , \Level1Out54[19] , \Level1Out54[18] , 
        \Level1Out54[17] , \Level1Out54[16] , \Level1Out54[15] , 
        \Level1Out54[14] , \Level1Out54[13] , \Level1Out54[12] , 
        \Level1Out54[11] , \Level1Out54[10] , \Level1Out54[9] , 
        \Level1Out54[8] , \Level1Out54[7] , \Level1Out54[6] , \Level1Out54[5] , 
        \Level1Out54[4] , \Level1Out54[3] , \Level1Out54[2] , \Level1Out54[1] , 
        \Level1Out54[0] }), .In2({\Level1Out55[31] , \Level1Out55[30] , 
        \Level1Out55[29] , \Level1Out55[28] , \Level1Out55[27] , 
        \Level1Out55[26] , \Level1Out55[25] , \Level1Out55[24] , 
        \Level1Out55[23] , \Level1Out55[22] , \Level1Out55[21] , 
        \Level1Out55[20] , \Level1Out55[19] , \Level1Out55[18] , 
        \Level1Out55[17] , \Level1Out55[16] , \Level1Out55[15] , 
        \Level1Out55[14] , \Level1Out55[13] , \Level1Out55[12] , 
        \Level1Out55[11] , \Level1Out55[10] , \Level1Out55[9] , 
        \Level1Out55[8] , \Level1Out55[7] , \Level1Out55[6] , \Level1Out55[5] , 
        \Level1Out55[4] , \Level1Out55[3] , \Level1Out55[2] , \Level1Out55[1] , 
        \Level1Out55[0] }), .Read1(\Level1Load54[0] ), .Read2(
        \Level1Load55[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_13 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink13[31] , \ScanLink13[30] , 
        \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , \ScanLink13[26] , 
        \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , \ScanLink13[22] , 
        \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , \ScanLink13[18] , 
        \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , \ScanLink13[14] , 
        \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , \ScanLink13[10] , 
        \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , \ScanLink13[6] , 
        \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , \ScanLink13[2] , 
        \ScanLink13[1] , \ScanLink13[0] }), .ScanOut({\ScanLink14[31] , 
        \ScanLink14[30] , \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , 
        \ScanLink14[26] , \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , 
        \ScanLink14[22] , \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , 
        \ScanLink14[18] , \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , 
        \ScanLink14[14] , \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , 
        \ScanLink14[10] , \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , 
        \ScanLink14[6] , \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , 
        \ScanLink14[2] , \ScanLink14[1] , \ScanLink14[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load13[0] ), .Out({
        \Level1Out13[31] , \Level1Out13[30] , \Level1Out13[29] , 
        \Level1Out13[28] , \Level1Out13[27] , \Level1Out13[26] , 
        \Level1Out13[25] , \Level1Out13[24] , \Level1Out13[23] , 
        \Level1Out13[22] , \Level1Out13[21] , \Level1Out13[20] , 
        \Level1Out13[19] , \Level1Out13[18] , \Level1Out13[17] , 
        \Level1Out13[16] , \Level1Out13[15] , \Level1Out13[14] , 
        \Level1Out13[13] , \Level1Out13[12] , \Level1Out13[11] , 
        \Level1Out13[10] , \Level1Out13[9] , \Level1Out13[8] , 
        \Level1Out13[7] , \Level1Out13[6] , \Level1Out13[5] , \Level1Out13[4] , 
        \Level1Out13[3] , \Level1Out13[2] , \Level1Out13[1] , \Level1Out13[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_14 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink14[31] , \ScanLink14[30] , 
        \ScanLink14[29] , \ScanLink14[28] , \ScanLink14[27] , \ScanLink14[26] , 
        \ScanLink14[25] , \ScanLink14[24] , \ScanLink14[23] , \ScanLink14[22] , 
        \ScanLink14[21] , \ScanLink14[20] , \ScanLink14[19] , \ScanLink14[18] , 
        \ScanLink14[17] , \ScanLink14[16] , \ScanLink14[15] , \ScanLink14[14] , 
        \ScanLink14[13] , \ScanLink14[12] , \ScanLink14[11] , \ScanLink14[10] , 
        \ScanLink14[9] , \ScanLink14[8] , \ScanLink14[7] , \ScanLink14[6] , 
        \ScanLink14[5] , \ScanLink14[4] , \ScanLink14[3] , \ScanLink14[2] , 
        \ScanLink14[1] , \ScanLink14[0] }), .ScanOut({\ScanLink15[31] , 
        \ScanLink15[30] , \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , 
        \ScanLink15[26] , \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , 
        \ScanLink15[22] , \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , 
        \ScanLink15[18] , \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , 
        \ScanLink15[14] , \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , 
        \ScanLink15[10] , \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , 
        \ScanLink15[6] , \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , 
        \ScanLink15[2] , \ScanLink15[1] , \ScanLink15[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load14[0] ), .Out({
        \Level1Out14[31] , \Level1Out14[30] , \Level1Out14[29] , 
        \Level1Out14[28] , \Level1Out14[27] , \Level1Out14[26] , 
        \Level1Out14[25] , \Level1Out14[24] , \Level1Out14[23] , 
        \Level1Out14[22] , \Level1Out14[21] , \Level1Out14[20] , 
        \Level1Out14[19] , \Level1Out14[18] , \Level1Out14[17] , 
        \Level1Out14[16] , \Level1Out14[15] , \Level1Out14[14] , 
        \Level1Out14[13] , \Level1Out14[12] , \Level1Out14[11] , 
        \Level1Out14[10] , \Level1Out14[9] , \Level1Out14[8] , 
        \Level1Out14[7] , \Level1Out14[6] , \Level1Out14[5] , \Level1Out14[4] , 
        \Level1Out14[3] , \Level1Out14[2] , \Level1Out14[1] , \Level1Out14[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load8[0] ), .Out({\Level4Out8[31] , \Level4Out8[30] , 
        \Level4Out8[29] , \Level4Out8[28] , \Level4Out8[27] , \Level4Out8[26] , 
        \Level4Out8[25] , \Level4Out8[24] , \Level4Out8[23] , \Level4Out8[22] , 
        \Level4Out8[21] , \Level4Out8[20] , \Level4Out8[19] , \Level4Out8[18] , 
        \Level4Out8[17] , \Level4Out8[16] , \Level4Out8[15] , \Level4Out8[14] , 
        \Level4Out8[13] , \Level4Out8[12] , \Level4Out8[11] , \Level4Out8[10] , 
        \Level4Out8[9] , \Level4Out8[8] , \Level4Out8[7] , \Level4Out8[6] , 
        \Level4Out8[5] , \Level4Out8[4] , \Level4Out8[3] , \Level4Out8[2] , 
        \Level4Out8[1] , \Level4Out8[0] }), .In1({\Level2Out8[31] , 
        \Level2Out8[30] , \Level2Out8[29] , \Level2Out8[28] , \Level2Out8[27] , 
        \Level2Out8[26] , \Level2Out8[25] , \Level2Out8[24] , \Level2Out8[23] , 
        \Level2Out8[22] , \Level2Out8[21] , \Level2Out8[20] , \Level2Out8[19] , 
        \Level2Out8[18] , \Level2Out8[17] , \Level2Out8[16] , \Level2Out8[15] , 
        \Level2Out8[14] , \Level2Out8[13] , \Level2Out8[12] , \Level2Out8[11] , 
        \Level2Out8[10] , \Level2Out8[9] , \Level2Out8[8] , \Level2Out8[7] , 
        \Level2Out8[6] , \Level2Out8[5] , \Level2Out8[4] , \Level2Out8[3] , 
        \Level2Out8[2] , \Level2Out8[1] , \Level2Out8[0] }), .In2({
        \Level2Out10[31] , \Level2Out10[30] , \Level2Out10[29] , 
        \Level2Out10[28] , \Level2Out10[27] , \Level2Out10[26] , 
        \Level2Out10[25] , \Level2Out10[24] , \Level2Out10[23] , 
        \Level2Out10[22] , \Level2Out10[21] , \Level2Out10[20] , 
        \Level2Out10[19] , \Level2Out10[18] , \Level2Out10[17] , 
        \Level2Out10[16] , \Level2Out10[15] , \Level2Out10[14] , 
        \Level2Out10[13] , \Level2Out10[12] , \Level2Out10[11] , 
        \Level2Out10[10] , \Level2Out10[9] , \Level2Out10[8] , 
        \Level2Out10[7] , \Level2Out10[6] , \Level2Out10[5] , \Level2Out10[4] , 
        \Level2Out10[3] , \Level2Out10[2] , \Level2Out10[1] , \Level2Out10[0] 
        }), .Read1(\Level2Load8[0] ), .Read2(\Level2Load10[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_33 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink33[31] , \ScanLink33[30] , 
        \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , \ScanLink33[26] , 
        \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , \ScanLink33[22] , 
        \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , \ScanLink33[18] , 
        \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , \ScanLink33[14] , 
        \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , \ScanLink33[10] , 
        \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , \ScanLink33[6] , 
        \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , \ScanLink33[2] , 
        \ScanLink33[1] , \ScanLink33[0] }), .ScanOut({\ScanLink34[31] , 
        \ScanLink34[30] , \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , 
        \ScanLink34[26] , \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , 
        \ScanLink34[22] , \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , 
        \ScanLink34[18] , \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , 
        \ScanLink34[14] , \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , 
        \ScanLink34[10] , \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , 
        \ScanLink34[6] , \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , 
        \ScanLink34[2] , \ScanLink34[1] , \ScanLink34[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load33[0] ), .Out({
        \Level1Out33[31] , \Level1Out33[30] , \Level1Out33[29] , 
        \Level1Out33[28] , \Level1Out33[27] , \Level1Out33[26] , 
        \Level1Out33[25] , \Level1Out33[24] , \Level1Out33[23] , 
        \Level1Out33[22] , \Level1Out33[21] , \Level1Out33[20] , 
        \Level1Out33[19] , \Level1Out33[18] , \Level1Out33[17] , 
        \Level1Out33[16] , \Level1Out33[15] , \Level1Out33[14] , 
        \Level1Out33[13] , \Level1Out33[12] , \Level1Out33[11] , 
        \Level1Out33[10] , \Level1Out33[9] , \Level1Out33[8] , 
        \Level1Out33[7] , \Level1Out33[6] , \Level1Out33[5] , \Level1Out33[4] , 
        \Level1Out33[3] , \Level1Out33[2] , \Level1Out33[1] , \Level1Out33[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_34 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink34[31] , \ScanLink34[30] , 
        \ScanLink34[29] , \ScanLink34[28] , \ScanLink34[27] , \ScanLink34[26] , 
        \ScanLink34[25] , \ScanLink34[24] , \ScanLink34[23] , \ScanLink34[22] , 
        \ScanLink34[21] , \ScanLink34[20] , \ScanLink34[19] , \ScanLink34[18] , 
        \ScanLink34[17] , \ScanLink34[16] , \ScanLink34[15] , \ScanLink34[14] , 
        \ScanLink34[13] , \ScanLink34[12] , \ScanLink34[11] , \ScanLink34[10] , 
        \ScanLink34[9] , \ScanLink34[8] , \ScanLink34[7] , \ScanLink34[6] , 
        \ScanLink34[5] , \ScanLink34[4] , \ScanLink34[3] , \ScanLink34[2] , 
        \ScanLink34[1] , \ScanLink34[0] }), .ScanOut({\ScanLink35[31] , 
        \ScanLink35[30] , \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , 
        \ScanLink35[26] , \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , 
        \ScanLink35[22] , \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , 
        \ScanLink35[18] , \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , 
        \ScanLink35[14] , \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , 
        \ScanLink35[10] , \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , 
        \ScanLink35[6] , \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , 
        \ScanLink35[2] , \ScanLink35[1] , \ScanLink35[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load34[0] ), .Out({
        \Level1Out34[31] , \Level1Out34[30] , \Level1Out34[29] , 
        \Level1Out34[28] , \Level1Out34[27] , \Level1Out34[26] , 
        \Level1Out34[25] , \Level1Out34[24] , \Level1Out34[23] , 
        \Level1Out34[22] , \Level1Out34[21] , \Level1Out34[20] , 
        \Level1Out34[19] , \Level1Out34[18] , \Level1Out34[17] , 
        \Level1Out34[16] , \Level1Out34[15] , \Level1Out34[14] , 
        \Level1Out34[13] , \Level1Out34[12] , \Level1Out34[11] , 
        \Level1Out34[10] , \Level1Out34[9] , \Level1Out34[8] , 
        \Level1Out34[7] , \Level1Out34[6] , \Level1Out34[5] , \Level1Out34[4] , 
        \Level1Out34[3] , \Level1Out34[2] , \Level1Out34[1] , \Level1Out34[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load0[0] ), .Out({\Level32Out0[31] , \Level32Out0[30] , 
        \Level32Out0[29] , \Level32Out0[28] , \Level32Out0[27] , 
        \Level32Out0[26] , \Level32Out0[25] , \Level32Out0[24] , 
        \Level32Out0[23] , \Level32Out0[22] , \Level32Out0[21] , 
        \Level32Out0[20] , \Level32Out0[19] , \Level32Out0[18] , 
        \Level32Out0[17] , \Level32Out0[16] , \Level32Out0[15] , 
        \Level32Out0[14] , \Level32Out0[13] , \Level32Out0[12] , 
        \Level32Out0[11] , \Level32Out0[10] , \Level32Out0[9] , 
        \Level32Out0[8] , \Level32Out0[7] , \Level32Out0[6] , \Level32Out0[5] , 
        \Level32Out0[4] , \Level32Out0[3] , \Level32Out0[2] , \Level32Out0[1] , 
        \Level32Out0[0] }), .In1({\Level16Out0[31] , \Level16Out0[30] , 
        \Level16Out0[29] , \Level16Out0[28] , \Level16Out0[27] , 
        \Level16Out0[26] , \Level16Out0[25] , \Level16Out0[24] , 
        \Level16Out0[23] , \Level16Out0[22] , \Level16Out0[21] , 
        \Level16Out0[20] , \Level16Out0[19] , \Level16Out0[18] , 
        \Level16Out0[17] , \Level16Out0[16] , \Level16Out0[15] , 
        \Level16Out0[14] , \Level16Out0[13] , \Level16Out0[12] , 
        \Level16Out0[11] , \Level16Out0[10] , \Level16Out0[9] , 
        \Level16Out0[8] , \Level16Out0[7] , \Level16Out0[6] , \Level16Out0[5] , 
        \Level16Out0[4] , \Level16Out0[3] , \Level16Out0[2] , \Level16Out0[1] , 
        \Level16Out0[0] }), .In2({\Level16Out16[31] , \Level16Out16[30] , 
        \Level16Out16[29] , \Level16Out16[28] , \Level16Out16[27] , 
        \Level16Out16[26] , \Level16Out16[25] , \Level16Out16[24] , 
        \Level16Out16[23] , \Level16Out16[22] , \Level16Out16[21] , 
        \Level16Out16[20] , \Level16Out16[19] , \Level16Out16[18] , 
        \Level16Out16[17] , \Level16Out16[16] , \Level16Out16[15] , 
        \Level16Out16[14] , \Level16Out16[13] , \Level16Out16[12] , 
        \Level16Out16[11] , \Level16Out16[10] , \Level16Out16[9] , 
        \Level16Out16[8] , \Level16Out16[7] , \Level16Out16[6] , 
        \Level16Out16[5] , \Level16Out16[4] , \Level16Out16[3] , 
        \Level16Out16[2] , \Level16Out16[1] , \Level16Out16[0] }), .Read1(
        \Level16Load0[0] ), .Read2(\Level16Load16[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_41 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink41[31] , \ScanLink41[30] , 
        \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , \ScanLink41[26] , 
        \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , \ScanLink41[22] , 
        \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , \ScanLink41[18] , 
        \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , \ScanLink41[14] , 
        \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , \ScanLink41[10] , 
        \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , \ScanLink41[6] , 
        \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , \ScanLink41[2] , 
        \ScanLink41[1] , \ScanLink41[0] }), .ScanOut({\ScanLink42[31] , 
        \ScanLink42[30] , \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , 
        \ScanLink42[26] , \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , 
        \ScanLink42[22] , \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , 
        \ScanLink42[18] , \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , 
        \ScanLink42[14] , \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , 
        \ScanLink42[10] , \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , 
        \ScanLink42[6] , \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , 
        \ScanLink42[2] , \ScanLink42[1] , \ScanLink42[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load41[0] ), .Out({
        \Level1Out41[31] , \Level1Out41[30] , \Level1Out41[29] , 
        \Level1Out41[28] , \Level1Out41[27] , \Level1Out41[26] , 
        \Level1Out41[25] , \Level1Out41[24] , \Level1Out41[23] , 
        \Level1Out41[22] , \Level1Out41[21] , \Level1Out41[20] , 
        \Level1Out41[19] , \Level1Out41[18] , \Level1Out41[17] , 
        \Level1Out41[16] , \Level1Out41[15] , \Level1Out41[14] , 
        \Level1Out41[13] , \Level1Out41[12] , \Level1Out41[11] , 
        \Level1Out41[10] , \Level1Out41[9] , \Level1Out41[8] , 
        \Level1Out41[7] , \Level1Out41[6] , \Level1Out41[5] , \Level1Out41[4] , 
        \Level1Out41[3] , \Level1Out41[2] , \Level1Out41[1] , \Level1Out41[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load0[0] ), .Out({\Level2Out0[31] , \Level2Out0[30] , 
        \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , \Level2Out0[26] , 
        \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , \Level2Out0[22] , 
        \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , \Level2Out0[18] , 
        \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , \Level2Out0[14] , 
        \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , \Level2Out0[10] , 
        \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , \Level2Out0[6] , 
        \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , \Level2Out0[2] , 
        \Level2Out0[1] , \Level2Out0[0] }), .In1({\Level1Out0[31] , 
        \Level1Out0[30] , \Level1Out0[29] , \Level1Out0[28] , \Level1Out0[27] , 
        \Level1Out0[26] , \Level1Out0[25] , \Level1Out0[24] , \Level1Out0[23] , 
        \Level1Out0[22] , \Level1Out0[21] , \Level1Out0[20] , \Level1Out0[19] , 
        \Level1Out0[18] , \Level1Out0[17] , \Level1Out0[16] , \Level1Out0[15] , 
        \Level1Out0[14] , \Level1Out0[13] , \Level1Out0[12] , \Level1Out0[11] , 
        \Level1Out0[10] , \Level1Out0[9] , \Level1Out0[8] , \Level1Out0[7] , 
        \Level1Out0[6] , \Level1Out0[5] , \Level1Out0[4] , \Level1Out0[3] , 
        \Level1Out0[2] , \Level1Out0[1] , \Level1Out0[0] }), .In2({
        \Level1Out1[31] , \Level1Out1[30] , \Level1Out1[29] , \Level1Out1[28] , 
        \Level1Out1[27] , \Level1Out1[26] , \Level1Out1[25] , \Level1Out1[24] , 
        \Level1Out1[23] , \Level1Out1[22] , \Level1Out1[21] , \Level1Out1[20] , 
        \Level1Out1[19] , \Level1Out1[18] , \Level1Out1[17] , \Level1Out1[16] , 
        \Level1Out1[15] , \Level1Out1[14] , \Level1Out1[13] , \Level1Out1[12] , 
        \Level1Out1[11] , \Level1Out1[10] , \Level1Out1[9] , \Level1Out1[8] , 
        \Level1Out1[7] , \Level1Out1[6] , \Level1Out1[5] , \Level1Out1[4] , 
        \Level1Out1[3] , \Level1Out1[2] , \Level1Out1[1] , \Level1Out1[0] }), 
        .Read1(\Level1Load0[0] ), .Read2(\Level1Load1[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_58_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load58[0] ), .Out({\Level2Out58[31] , \Level2Out58[30] , 
        \Level2Out58[29] , \Level2Out58[28] , \Level2Out58[27] , 
        \Level2Out58[26] , \Level2Out58[25] , \Level2Out58[24] , 
        \Level2Out58[23] , \Level2Out58[22] , \Level2Out58[21] , 
        \Level2Out58[20] , \Level2Out58[19] , \Level2Out58[18] , 
        \Level2Out58[17] , \Level2Out58[16] , \Level2Out58[15] , 
        \Level2Out58[14] , \Level2Out58[13] , \Level2Out58[12] , 
        \Level2Out58[11] , \Level2Out58[10] , \Level2Out58[9] , 
        \Level2Out58[8] , \Level2Out58[7] , \Level2Out58[6] , \Level2Out58[5] , 
        \Level2Out58[4] , \Level2Out58[3] , \Level2Out58[2] , \Level2Out58[1] , 
        \Level2Out58[0] }), .In1({\Level1Out58[31] , \Level1Out58[30] , 
        \Level1Out58[29] , \Level1Out58[28] , \Level1Out58[27] , 
        \Level1Out58[26] , \Level1Out58[25] , \Level1Out58[24] , 
        \Level1Out58[23] , \Level1Out58[22] , \Level1Out58[21] , 
        \Level1Out58[20] , \Level1Out58[19] , \Level1Out58[18] , 
        \Level1Out58[17] , \Level1Out58[16] , \Level1Out58[15] , 
        \Level1Out58[14] , \Level1Out58[13] , \Level1Out58[12] , 
        \Level1Out58[11] , \Level1Out58[10] , \Level1Out58[9] , 
        \Level1Out58[8] , \Level1Out58[7] , \Level1Out58[6] , \Level1Out58[5] , 
        \Level1Out58[4] , \Level1Out58[3] , \Level1Out58[2] , \Level1Out58[1] , 
        \Level1Out58[0] }), .In2({\Level1Out59[31] , \Level1Out59[30] , 
        \Level1Out59[29] , \Level1Out59[28] , \Level1Out59[27] , 
        \Level1Out59[26] , \Level1Out59[25] , \Level1Out59[24] , 
        \Level1Out59[23] , \Level1Out59[22] , \Level1Out59[21] , 
        \Level1Out59[20] , \Level1Out59[19] , \Level1Out59[18] , 
        \Level1Out59[17] , \Level1Out59[16] , \Level1Out59[15] , 
        \Level1Out59[14] , \Level1Out59[13] , \Level1Out59[12] , 
        \Level1Out59[11] , \Level1Out59[10] , \Level1Out59[9] , 
        \Level1Out59[8] , \Level1Out59[7] , \Level1Out59[6] , \Level1Out59[5] , 
        \Level1Out59[4] , \Level1Out59[3] , \Level1Out59[2] , \Level1Out59[1] , 
        \Level1Out59[0] }), .Read1(\Level1Load58[0] ), .Read2(
        \Level1Load59[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_44_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load44[0] ), .Out({\Level4Out44[31] , \Level4Out44[30] , 
        \Level4Out44[29] , \Level4Out44[28] , \Level4Out44[27] , 
        \Level4Out44[26] , \Level4Out44[25] , \Level4Out44[24] , 
        \Level4Out44[23] , \Level4Out44[22] , \Level4Out44[21] , 
        \Level4Out44[20] , \Level4Out44[19] , \Level4Out44[18] , 
        \Level4Out44[17] , \Level4Out44[16] , \Level4Out44[15] , 
        \Level4Out44[14] , \Level4Out44[13] , \Level4Out44[12] , 
        \Level4Out44[11] , \Level4Out44[10] , \Level4Out44[9] , 
        \Level4Out44[8] , \Level4Out44[7] , \Level4Out44[6] , \Level4Out44[5] , 
        \Level4Out44[4] , \Level4Out44[3] , \Level4Out44[2] , \Level4Out44[1] , 
        \Level4Out44[0] }), .In1({\Level2Out44[31] , \Level2Out44[30] , 
        \Level2Out44[29] , \Level2Out44[28] , \Level2Out44[27] , 
        \Level2Out44[26] , \Level2Out44[25] , \Level2Out44[24] , 
        \Level2Out44[23] , \Level2Out44[22] , \Level2Out44[21] , 
        \Level2Out44[20] , \Level2Out44[19] , \Level2Out44[18] , 
        \Level2Out44[17] , \Level2Out44[16] , \Level2Out44[15] , 
        \Level2Out44[14] , \Level2Out44[13] , \Level2Out44[12] , 
        \Level2Out44[11] , \Level2Out44[10] , \Level2Out44[9] , 
        \Level2Out44[8] , \Level2Out44[7] , \Level2Out44[6] , \Level2Out44[5] , 
        \Level2Out44[4] , \Level2Out44[3] , \Level2Out44[2] , \Level2Out44[1] , 
        \Level2Out44[0] }), .In2({\Level2Out46[31] , \Level2Out46[30] , 
        \Level2Out46[29] , \Level2Out46[28] , \Level2Out46[27] , 
        \Level2Out46[26] , \Level2Out46[25] , \Level2Out46[24] , 
        \Level2Out46[23] , \Level2Out46[22] , \Level2Out46[21] , 
        \Level2Out46[20] , \Level2Out46[19] , \Level2Out46[18] , 
        \Level2Out46[17] , \Level2Out46[16] , \Level2Out46[15] , 
        \Level2Out46[14] , \Level2Out46[13] , \Level2Out46[12] , 
        \Level2Out46[11] , \Level2Out46[10] , \Level2Out46[9] , 
        \Level2Out46[8] , \Level2Out46[7] , \Level2Out46[6] , \Level2Out46[5] , 
        \Level2Out46[4] , \Level2Out46[3] , \Level2Out46[2] , \Level2Out46[1] , 
        \Level2Out46[0] }), .Read1(\Level2Load44[0] ), .Read2(
        \Level2Load46[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_48 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink48[31] , \ScanLink48[30] , 
        \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , \ScanLink48[26] , 
        \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , \ScanLink48[22] , 
        \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , \ScanLink48[18] , 
        \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , \ScanLink48[14] , 
        \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , \ScanLink48[10] , 
        \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , \ScanLink48[6] , 
        \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , \ScanLink48[2] , 
        \ScanLink48[1] , \ScanLink48[0] }), .ScanOut({\ScanLink49[31] , 
        \ScanLink49[30] , \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , 
        \ScanLink49[26] , \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , 
        \ScanLink49[22] , \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , 
        \ScanLink49[18] , \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , 
        \ScanLink49[14] , \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , 
        \ScanLink49[10] , \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , 
        \ScanLink49[6] , \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , 
        \ScanLink49[2] , \ScanLink49[1] , \ScanLink49[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load48[0] ), .Out({
        \Level1Out48[31] , \Level1Out48[30] , \Level1Out48[29] , 
        \Level1Out48[28] , \Level1Out48[27] , \Level1Out48[26] , 
        \Level1Out48[25] , \Level1Out48[24] , \Level1Out48[23] , 
        \Level1Out48[22] , \Level1Out48[21] , \Level1Out48[20] , 
        \Level1Out48[19] , \Level1Out48[18] , \Level1Out48[17] , 
        \Level1Out48[16] , \Level1Out48[15] , \Level1Out48[14] , 
        \Level1Out48[13] , \Level1Out48[12] , \Level1Out48[11] , 
        \Level1Out48[10] , \Level1Out48[9] , \Level1Out48[8] , 
        \Level1Out48[7] , \Level1Out48[6] , \Level1Out48[5] , \Level1Out48[4] , 
        \Level1Out48[3] , \Level1Out48[2] , \Level1Out48[1] , \Level1Out48[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_53 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink53[31] , \ScanLink53[30] , 
        \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , \ScanLink53[26] , 
        \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , \ScanLink53[22] , 
        \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , \ScanLink53[18] , 
        \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , \ScanLink53[14] , 
        \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , \ScanLink53[10] , 
        \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , \ScanLink53[6] , 
        \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , \ScanLink53[2] , 
        \ScanLink53[1] , \ScanLink53[0] }), .ScanOut({\ScanLink54[31] , 
        \ScanLink54[30] , \ScanLink54[29] , \ScanLink54[28] , \ScanLink54[27] , 
        \ScanLink54[26] , \ScanLink54[25] , \ScanLink54[24] , \ScanLink54[23] , 
        \ScanLink54[22] , \ScanLink54[21] , \ScanLink54[20] , \ScanLink54[19] , 
        \ScanLink54[18] , \ScanLink54[17] , \ScanLink54[16] , \ScanLink54[15] , 
        \ScanLink54[14] , \ScanLink54[13] , \ScanLink54[12] , \ScanLink54[11] , 
        \ScanLink54[10] , \ScanLink54[9] , \ScanLink54[8] , \ScanLink54[7] , 
        \ScanLink54[6] , \ScanLink54[5] , \ScanLink54[4] , \ScanLink54[3] , 
        \ScanLink54[2] , \ScanLink54[1] , \ScanLink54[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load53[0] ), .Out({
        \Level1Out53[31] , \Level1Out53[30] , \Level1Out53[29] , 
        \Level1Out53[28] , \Level1Out53[27] , \Level1Out53[26] , 
        \Level1Out53[25] , \Level1Out53[24] , \Level1Out53[23] , 
        \Level1Out53[22] , \Level1Out53[21] , \Level1Out53[20] , 
        \Level1Out53[19] , \Level1Out53[18] , \Level1Out53[17] , 
        \Level1Out53[16] , \Level1Out53[15] , \Level1Out53[14] , 
        \Level1Out53[13] , \Level1Out53[12] , \Level1Out53[11] , 
        \Level1Out53[10] , \Level1Out53[9] , \Level1Out53[8] , 
        \Level1Out53[7] , \Level1Out53[6] , \Level1Out53[5] , \Level1Out53[4] , 
        \Level1Out53[3] , \Level1Out53[2] , \Level1Out53[1] , \Level1Out53[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_10_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load10[0] ), .Out({\Level2Out10[31] , \Level2Out10[30] , 
        \Level2Out10[29] , \Level2Out10[28] , \Level2Out10[27] , 
        \Level2Out10[26] , \Level2Out10[25] , \Level2Out10[24] , 
        \Level2Out10[23] , \Level2Out10[22] , \Level2Out10[21] , 
        \Level2Out10[20] , \Level2Out10[19] , \Level2Out10[18] , 
        \Level2Out10[17] , \Level2Out10[16] , \Level2Out10[15] , 
        \Level2Out10[14] , \Level2Out10[13] , \Level2Out10[12] , 
        \Level2Out10[11] , \Level2Out10[10] , \Level2Out10[9] , 
        \Level2Out10[8] , \Level2Out10[7] , \Level2Out10[6] , \Level2Out10[5] , 
        \Level2Out10[4] , \Level2Out10[3] , \Level2Out10[2] , \Level2Out10[1] , 
        \Level2Out10[0] }), .In1({\Level1Out10[31] , \Level1Out10[30] , 
        \Level1Out10[29] , \Level1Out10[28] , \Level1Out10[27] , 
        \Level1Out10[26] , \Level1Out10[25] , \Level1Out10[24] , 
        \Level1Out10[23] , \Level1Out10[22] , \Level1Out10[21] , 
        \Level1Out10[20] , \Level1Out10[19] , \Level1Out10[18] , 
        \Level1Out10[17] , \Level1Out10[16] , \Level1Out10[15] , 
        \Level1Out10[14] , \Level1Out10[13] , \Level1Out10[12] , 
        \Level1Out10[11] , \Level1Out10[10] , \Level1Out10[9] , 
        \Level1Out10[8] , \Level1Out10[7] , \Level1Out10[6] , \Level1Out10[5] , 
        \Level1Out10[4] , \Level1Out10[3] , \Level1Out10[2] , \Level1Out10[1] , 
        \Level1Out10[0] }), .In2({\Level1Out11[31] , \Level1Out11[30] , 
        \Level1Out11[29] , \Level1Out11[28] , \Level1Out11[27] , 
        \Level1Out11[26] , \Level1Out11[25] , \Level1Out11[24] , 
        \Level1Out11[23] , \Level1Out11[22] , \Level1Out11[21] , 
        \Level1Out11[20] , \Level1Out11[19] , \Level1Out11[18] , 
        \Level1Out11[17] , \Level1Out11[16] , \Level1Out11[15] , 
        \Level1Out11[14] , \Level1Out11[13] , \Level1Out11[12] , 
        \Level1Out11[11] , \Level1Out11[10] , \Level1Out11[9] , 
        \Level1Out11[8] , \Level1Out11[7] , \Level1Out11[6] , \Level1Out11[5] , 
        \Level1Out11[4] , \Level1Out11[3] , \Level1Out11[2] , \Level1Out11[1] , 
        \Level1Out11[0] }), .Read1(\Level1Load10[0] ), .Read2(
        \Level1Load11[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load40[0] ), .Out({\Level2Out40[31] , \Level2Out40[30] , 
        \Level2Out40[29] , \Level2Out40[28] , \Level2Out40[27] , 
        \Level2Out40[26] , \Level2Out40[25] , \Level2Out40[24] , 
        \Level2Out40[23] , \Level2Out40[22] , \Level2Out40[21] , 
        \Level2Out40[20] , \Level2Out40[19] , \Level2Out40[18] , 
        \Level2Out40[17] , \Level2Out40[16] , \Level2Out40[15] , 
        \Level2Out40[14] , \Level2Out40[13] , \Level2Out40[12] , 
        \Level2Out40[11] , \Level2Out40[10] , \Level2Out40[9] , 
        \Level2Out40[8] , \Level2Out40[7] , \Level2Out40[6] , \Level2Out40[5] , 
        \Level2Out40[4] , \Level2Out40[3] , \Level2Out40[2] , \Level2Out40[1] , 
        \Level2Out40[0] }), .In1({\Level1Out40[31] , \Level1Out40[30] , 
        \Level1Out40[29] , \Level1Out40[28] , \Level1Out40[27] , 
        \Level1Out40[26] , \Level1Out40[25] , \Level1Out40[24] , 
        \Level1Out40[23] , \Level1Out40[22] , \Level1Out40[21] , 
        \Level1Out40[20] , \Level1Out40[19] , \Level1Out40[18] , 
        \Level1Out40[17] , \Level1Out40[16] , \Level1Out40[15] , 
        \Level1Out40[14] , \Level1Out40[13] , \Level1Out40[12] , 
        \Level1Out40[11] , \Level1Out40[10] , \Level1Out40[9] , 
        \Level1Out40[8] , \Level1Out40[7] , \Level1Out40[6] , \Level1Out40[5] , 
        \Level1Out40[4] , \Level1Out40[3] , \Level1Out40[2] , \Level1Out40[1] , 
        \Level1Out40[0] }), .In2({\Level1Out41[31] , \Level1Out41[30] , 
        \Level1Out41[29] , \Level1Out41[28] , \Level1Out41[27] , 
        \Level1Out41[26] , \Level1Out41[25] , \Level1Out41[24] , 
        \Level1Out41[23] , \Level1Out41[22] , \Level1Out41[21] , 
        \Level1Out41[20] , \Level1Out41[19] , \Level1Out41[18] , 
        \Level1Out41[17] , \Level1Out41[16] , \Level1Out41[15] , 
        \Level1Out41[14] , \Level1Out41[13] , \Level1Out41[12] , 
        \Level1Out41[11] , \Level1Out41[10] , \Level1Out41[9] , 
        \Level1Out41[8] , \Level1Out41[7] , \Level1Out41[6] , \Level1Out41[5] , 
        \Level1Out41[4] , \Level1Out41[3] , \Level1Out41[2] , \Level1Out41[1] , 
        \Level1Out41[0] }), .Read1(\Level1Load40[0] ), .Read2(
        \Level1Load41[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load4[0] ), .Out({\Level4Out4[31] , \Level4Out4[30] , 
        \Level4Out4[29] , \Level4Out4[28] , \Level4Out4[27] , \Level4Out4[26] , 
        \Level4Out4[25] , \Level4Out4[24] , \Level4Out4[23] , \Level4Out4[22] , 
        \Level4Out4[21] , \Level4Out4[20] , \Level4Out4[19] , \Level4Out4[18] , 
        \Level4Out4[17] , \Level4Out4[16] , \Level4Out4[15] , \Level4Out4[14] , 
        \Level4Out4[13] , \Level4Out4[12] , \Level4Out4[11] , \Level4Out4[10] , 
        \Level4Out4[9] , \Level4Out4[8] , \Level4Out4[7] , \Level4Out4[6] , 
        \Level4Out4[5] , \Level4Out4[4] , \Level4Out4[3] , \Level4Out4[2] , 
        \Level4Out4[1] , \Level4Out4[0] }), .In1({\Level2Out4[31] , 
        \Level2Out4[30] , \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , 
        \Level2Out4[26] , \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , 
        \Level2Out4[22] , \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , 
        \Level2Out4[18] , \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , 
        \Level2Out4[14] , \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , 
        \Level2Out4[10] , \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , 
        \Level2Out4[6] , \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , 
        \Level2Out4[2] , \Level2Out4[1] , \Level2Out4[0] }), .In2({
        \Level2Out6[31] , \Level2Out6[30] , \Level2Out6[29] , \Level2Out6[28] , 
        \Level2Out6[27] , \Level2Out6[26] , \Level2Out6[25] , \Level2Out6[24] , 
        \Level2Out6[23] , \Level2Out6[22] , \Level2Out6[21] , \Level2Out6[20] , 
        \Level2Out6[19] , \Level2Out6[18] , \Level2Out6[17] , \Level2Out6[16] , 
        \Level2Out6[15] , \Level2Out6[14] , \Level2Out6[13] , \Level2Out6[12] , 
        \Level2Out6[11] , \Level2Out6[10] , \Level2Out6[9] , \Level2Out6[8] , 
        \Level2Out6[7] , \Level2Out6[6] , \Level2Out6[5] , \Level2Out6[4] , 
        \Level2Out6[3] , \Level2Out6[2] , \Level2Out6[1] , \Level2Out6[0] }), 
        .Read1(\Level2Load4[0] ), .Read2(\Level2Load6[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load24[0] ), .Out({\Level8Out24[31] , \Level8Out24[30] , 
        \Level8Out24[29] , \Level8Out24[28] , \Level8Out24[27] , 
        \Level8Out24[26] , \Level8Out24[25] , \Level8Out24[24] , 
        \Level8Out24[23] , \Level8Out24[22] , \Level8Out24[21] , 
        \Level8Out24[20] , \Level8Out24[19] , \Level8Out24[18] , 
        \Level8Out24[17] , \Level8Out24[16] , \Level8Out24[15] , 
        \Level8Out24[14] , \Level8Out24[13] , \Level8Out24[12] , 
        \Level8Out24[11] , \Level8Out24[10] , \Level8Out24[9] , 
        \Level8Out24[8] , \Level8Out24[7] , \Level8Out24[6] , \Level8Out24[5] , 
        \Level8Out24[4] , \Level8Out24[3] , \Level8Out24[2] , \Level8Out24[1] , 
        \Level8Out24[0] }), .In1({\Level4Out24[31] , \Level4Out24[30] , 
        \Level4Out24[29] , \Level4Out24[28] , \Level4Out24[27] , 
        \Level4Out24[26] , \Level4Out24[25] , \Level4Out24[24] , 
        \Level4Out24[23] , \Level4Out24[22] , \Level4Out24[21] , 
        \Level4Out24[20] , \Level4Out24[19] , \Level4Out24[18] , 
        \Level4Out24[17] , \Level4Out24[16] , \Level4Out24[15] , 
        \Level4Out24[14] , \Level4Out24[13] , \Level4Out24[12] , 
        \Level4Out24[11] , \Level4Out24[10] , \Level4Out24[9] , 
        \Level4Out24[8] , \Level4Out24[7] , \Level4Out24[6] , \Level4Out24[5] , 
        \Level4Out24[4] , \Level4Out24[3] , \Level4Out24[2] , \Level4Out24[1] , 
        \Level4Out24[0] }), .In2({\Level4Out28[31] , \Level4Out28[30] , 
        \Level4Out28[29] , \Level4Out28[28] , \Level4Out28[27] , 
        \Level4Out28[26] , \Level4Out28[25] , \Level4Out28[24] , 
        \Level4Out28[23] , \Level4Out28[22] , \Level4Out28[21] , 
        \Level4Out28[20] , \Level4Out28[19] , \Level4Out28[18] , 
        \Level4Out28[17] , \Level4Out28[16] , \Level4Out28[15] , 
        \Level4Out28[14] , \Level4Out28[13] , \Level4Out28[12] , 
        \Level4Out28[11] , \Level4Out28[10] , \Level4Out28[9] , 
        \Level4Out28[8] , \Level4Out28[7] , \Level4Out28[6] , \Level4Out28[5] , 
        \Level4Out28[4] , \Level4Out28[3] , \Level4Out28[2] , \Level4Out28[1] , 
        \Level4Out28[0] }), .Read1(\Level4Load24[0] ), .Read2(
        \Level4Load28[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_7 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink7[31] , \ScanLink7[30] , 
        \ScanLink7[29] , \ScanLink7[28] , \ScanLink7[27] , \ScanLink7[26] , 
        \ScanLink7[25] , \ScanLink7[24] , \ScanLink7[23] , \ScanLink7[22] , 
        \ScanLink7[21] , \ScanLink7[20] , \ScanLink7[19] , \ScanLink7[18] , 
        \ScanLink7[17] , \ScanLink7[16] , \ScanLink7[15] , \ScanLink7[14] , 
        \ScanLink7[13] , \ScanLink7[12] , \ScanLink7[11] , \ScanLink7[10] , 
        \ScanLink7[9] , \ScanLink7[8] , \ScanLink7[7] , \ScanLink7[6] , 
        \ScanLink7[5] , \ScanLink7[4] , \ScanLink7[3] , \ScanLink7[2] , 
        \ScanLink7[1] , \ScanLink7[0] }), .ScanOut({\ScanLink8[31] , 
        \ScanLink8[30] , \ScanLink8[29] , \ScanLink8[28] , \ScanLink8[27] , 
        \ScanLink8[26] , \ScanLink8[25] , \ScanLink8[24] , \ScanLink8[23] , 
        \ScanLink8[22] , \ScanLink8[21] , \ScanLink8[20] , \ScanLink8[19] , 
        \ScanLink8[18] , \ScanLink8[17] , \ScanLink8[16] , \ScanLink8[15] , 
        \ScanLink8[14] , \ScanLink8[13] , \ScanLink8[12] , \ScanLink8[11] , 
        \ScanLink8[10] , \ScanLink8[9] , \ScanLink8[8] , \ScanLink8[7] , 
        \ScanLink8[6] , \ScanLink8[5] , \ScanLink8[4] , \ScanLink8[3] , 
        \ScanLink8[2] , \ScanLink8[1] , \ScanLink8[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load7[0] ), .Out({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_12 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink12[31] , \ScanLink12[30] , 
        \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , \ScanLink12[26] , 
        \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , \ScanLink12[22] , 
        \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , \ScanLink12[18] , 
        \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , \ScanLink12[14] , 
        \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , \ScanLink12[10] , 
        \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , \ScanLink12[6] , 
        \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , \ScanLink12[2] , 
        \ScanLink12[1] , \ScanLink12[0] }), .ScanOut({\ScanLink13[31] , 
        \ScanLink13[30] , \ScanLink13[29] , \ScanLink13[28] , \ScanLink13[27] , 
        \ScanLink13[26] , \ScanLink13[25] , \ScanLink13[24] , \ScanLink13[23] , 
        \ScanLink13[22] , \ScanLink13[21] , \ScanLink13[20] , \ScanLink13[19] , 
        \ScanLink13[18] , \ScanLink13[17] , \ScanLink13[16] , \ScanLink13[15] , 
        \ScanLink13[14] , \ScanLink13[13] , \ScanLink13[12] , \ScanLink13[11] , 
        \ScanLink13[10] , \ScanLink13[9] , \ScanLink13[8] , \ScanLink13[7] , 
        \ScanLink13[6] , \ScanLink13[5] , \ScanLink13[4] , \ScanLink13[3] , 
        \ScanLink13[2] , \ScanLink13[1] , \ScanLink13[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load12[0] ), .Out({
        \Level1Out12[31] , \Level1Out12[30] , \Level1Out12[29] , 
        \Level1Out12[28] , \Level1Out12[27] , \Level1Out12[26] , 
        \Level1Out12[25] , \Level1Out12[24] , \Level1Out12[23] , 
        \Level1Out12[22] , \Level1Out12[21] , \Level1Out12[20] , 
        \Level1Out12[19] , \Level1Out12[18] , \Level1Out12[17] , 
        \Level1Out12[16] , \Level1Out12[15] , \Level1Out12[14] , 
        \Level1Out12[13] , \Level1Out12[12] , \Level1Out12[11] , 
        \Level1Out12[10] , \Level1Out12[9] , \Level1Out12[8] , 
        \Level1Out12[7] , \Level1Out12[6] , \Level1Out12[5] , \Level1Out12[4] , 
        \Level1Out12[3] , \Level1Out12[2] , \Level1Out12[1] , \Level1Out12[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_26 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink26[31] , \ScanLink26[30] , 
        \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , \ScanLink26[26] , 
        \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , \ScanLink26[22] , 
        \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , \ScanLink26[18] , 
        \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , \ScanLink26[14] , 
        \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , \ScanLink26[10] , 
        \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , \ScanLink26[6] , 
        \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , \ScanLink26[2] , 
        \ScanLink26[1] , \ScanLink26[0] }), .ScanOut({\ScanLink27[31] , 
        \ScanLink27[30] , \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , 
        \ScanLink27[26] , \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , 
        \ScanLink27[22] , \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , 
        \ScanLink27[18] , \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , 
        \ScanLink27[14] , \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , 
        \ScanLink27[10] , \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , 
        \ScanLink27[6] , \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , 
        \ScanLink27[2] , \ScanLink27[1] , \ScanLink27[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load26[0] ), .Out({
        \Level1Out26[31] , \Level1Out26[30] , \Level1Out26[29] , 
        \Level1Out26[28] , \Level1Out26[27] , \Level1Out26[26] , 
        \Level1Out26[25] , \Level1Out26[24] , \Level1Out26[23] , 
        \Level1Out26[22] , \Level1Out26[21] , \Level1Out26[20] , 
        \Level1Out26[19] , \Level1Out26[18] , \Level1Out26[17] , 
        \Level1Out26[16] , \Level1Out26[15] , \Level1Out26[14] , 
        \Level1Out26[13] , \Level1Out26[12] , \Level1Out26[11] , 
        \Level1Out26[10] , \Level1Out26[9] , \Level1Out26[8] , 
        \Level1Out26[7] , \Level1Out26[6] , \Level1Out26[5] , \Level1Out26[4] , 
        \Level1Out26[3] , \Level1Out26[2] , \Level1Out26[1] , \Level1Out26[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_22_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load22[0] ), .Out({\Level2Out22[31] , \Level2Out22[30] , 
        \Level2Out22[29] , \Level2Out22[28] , \Level2Out22[27] , 
        \Level2Out22[26] , \Level2Out22[25] , \Level2Out22[24] , 
        \Level2Out22[23] , \Level2Out22[22] , \Level2Out22[21] , 
        \Level2Out22[20] , \Level2Out22[19] , \Level2Out22[18] , 
        \Level2Out22[17] , \Level2Out22[16] , \Level2Out22[15] , 
        \Level2Out22[14] , \Level2Out22[13] , \Level2Out22[12] , 
        \Level2Out22[11] , \Level2Out22[10] , \Level2Out22[9] , 
        \Level2Out22[8] , \Level2Out22[7] , \Level2Out22[6] , \Level2Out22[5] , 
        \Level2Out22[4] , \Level2Out22[3] , \Level2Out22[2] , \Level2Out22[1] , 
        \Level2Out22[0] }), .In1({\Level1Out22[31] , \Level1Out22[30] , 
        \Level1Out22[29] , \Level1Out22[28] , \Level1Out22[27] , 
        \Level1Out22[26] , \Level1Out22[25] , \Level1Out22[24] , 
        \Level1Out22[23] , \Level1Out22[22] , \Level1Out22[21] , 
        \Level1Out22[20] , \Level1Out22[19] , \Level1Out22[18] , 
        \Level1Out22[17] , \Level1Out22[16] , \Level1Out22[15] , 
        \Level1Out22[14] , \Level1Out22[13] , \Level1Out22[12] , 
        \Level1Out22[11] , \Level1Out22[10] , \Level1Out22[9] , 
        \Level1Out22[8] , \Level1Out22[7] , \Level1Out22[6] , \Level1Out22[5] , 
        \Level1Out22[4] , \Level1Out22[3] , \Level1Out22[2] , \Level1Out22[1] , 
        \Level1Out22[0] }), .In2({\Level1Out23[31] , \Level1Out23[30] , 
        \Level1Out23[29] , \Level1Out23[28] , \Level1Out23[27] , 
        \Level1Out23[26] , \Level1Out23[25] , \Level1Out23[24] , 
        \Level1Out23[23] , \Level1Out23[22] , \Level1Out23[21] , 
        \Level1Out23[20] , \Level1Out23[19] , \Level1Out23[18] , 
        \Level1Out23[17] , \Level1Out23[16] , \Level1Out23[15] , 
        \Level1Out23[14] , \Level1Out23[13] , \Level1Out23[12] , 
        \Level1Out23[11] , \Level1Out23[10] , \Level1Out23[9] , 
        \Level1Out23[8] , \Level1Out23[7] , \Level1Out23[6] , \Level1Out23[5] , 
        \Level1Out23[4] , \Level1Out23[3] , \Level1Out23[2] , \Level1Out23[1] , 
        \Level1Out23[0] }), .Read1(\Level1Load22[0] ), .Read2(
        \Level1Load23[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level32Load32[0] ), .Out({\Level32Out32[31] , \Level32Out32[30] , 
        \Level32Out32[29] , \Level32Out32[28] , \Level32Out32[27] , 
        \Level32Out32[26] , \Level32Out32[25] , \Level32Out32[24] , 
        \Level32Out32[23] , \Level32Out32[22] , \Level32Out32[21] , 
        \Level32Out32[20] , \Level32Out32[19] , \Level32Out32[18] , 
        \Level32Out32[17] , \Level32Out32[16] , \Level32Out32[15] , 
        \Level32Out32[14] , \Level32Out32[13] , \Level32Out32[12] , 
        \Level32Out32[11] , \Level32Out32[10] , \Level32Out32[9] , 
        \Level32Out32[8] , \Level32Out32[7] , \Level32Out32[6] , 
        \Level32Out32[5] , \Level32Out32[4] , \Level32Out32[3] , 
        \Level32Out32[2] , \Level32Out32[1] , \Level32Out32[0] }), .In1({
        \Level16Out32[31] , \Level16Out32[30] , \Level16Out32[29] , 
        \Level16Out32[28] , \Level16Out32[27] , \Level16Out32[26] , 
        \Level16Out32[25] , \Level16Out32[24] , \Level16Out32[23] , 
        \Level16Out32[22] , \Level16Out32[21] , \Level16Out32[20] , 
        \Level16Out32[19] , \Level16Out32[18] , \Level16Out32[17] , 
        \Level16Out32[16] , \Level16Out32[15] , \Level16Out32[14] , 
        \Level16Out32[13] , \Level16Out32[12] , \Level16Out32[11] , 
        \Level16Out32[10] , \Level16Out32[9] , \Level16Out32[8] , 
        \Level16Out32[7] , \Level16Out32[6] , \Level16Out32[5] , 
        \Level16Out32[4] , \Level16Out32[3] , \Level16Out32[2] , 
        \Level16Out32[1] , \Level16Out32[0] }), .In2({\Level16Out48[31] , 
        \Level16Out48[30] , \Level16Out48[29] , \Level16Out48[28] , 
        \Level16Out48[27] , \Level16Out48[26] , \Level16Out48[25] , 
        \Level16Out48[24] , \Level16Out48[23] , \Level16Out48[22] , 
        \Level16Out48[21] , \Level16Out48[20] , \Level16Out48[19] , 
        \Level16Out48[18] , \Level16Out48[17] , \Level16Out48[16] , 
        \Level16Out48[15] , \Level16Out48[14] , \Level16Out48[13] , 
        \Level16Out48[12] , \Level16Out48[11] , \Level16Out48[10] , 
        \Level16Out48[9] , \Level16Out48[8] , \Level16Out48[7] , 
        \Level16Out48[6] , \Level16Out48[5] , \Level16Out48[4] , 
        \Level16Out48[3] , \Level16Out48[2] , \Level16Out48[1] , 
        \Level16Out48[0] }), .Read1(\Level16Load32[0] ), .Read2(
        \Level16Load48[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_35 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink35[31] , \ScanLink35[30] , 
        \ScanLink35[29] , \ScanLink35[28] , \ScanLink35[27] , \ScanLink35[26] , 
        \ScanLink35[25] , \ScanLink35[24] , \ScanLink35[23] , \ScanLink35[22] , 
        \ScanLink35[21] , \ScanLink35[20] , \ScanLink35[19] , \ScanLink35[18] , 
        \ScanLink35[17] , \ScanLink35[16] , \ScanLink35[15] , \ScanLink35[14] , 
        \ScanLink35[13] , \ScanLink35[12] , \ScanLink35[11] , \ScanLink35[10] , 
        \ScanLink35[9] , \ScanLink35[8] , \ScanLink35[7] , \ScanLink35[6] , 
        \ScanLink35[5] , \ScanLink35[4] , \ScanLink35[3] , \ScanLink35[2] , 
        \ScanLink35[1] , \ScanLink35[0] }), .ScanOut({\ScanLink36[31] , 
        \ScanLink36[30] , \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , 
        \ScanLink36[26] , \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , 
        \ScanLink36[22] , \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , 
        \ScanLink36[18] , \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , 
        \ScanLink36[14] , \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , 
        \ScanLink36[10] , \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , 
        \ScanLink36[6] , \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , 
        \ScanLink36[2] , \ScanLink36[1] , \ScanLink36[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load35[0] ), .Out({
        \Level1Out35[31] , \Level1Out35[30] , \Level1Out35[29] , 
        \Level1Out35[28] , \Level1Out35[27] , \Level1Out35[26] , 
        \Level1Out35[25] , \Level1Out35[24] , \Level1Out35[23] , 
        \Level1Out35[22] , \Level1Out35[21] , \Level1Out35[20] , 
        \Level1Out35[19] , \Level1Out35[18] , \Level1Out35[17] , 
        \Level1Out35[16] , \Level1Out35[15] , \Level1Out35[14] , 
        \Level1Out35[13] , \Level1Out35[12] , \Level1Out35[11] , 
        \Level1Out35[10] , \Level1Out35[9] , \Level1Out35[8] , 
        \Level1Out35[7] , \Level1Out35[6] , \Level1Out35[5] , \Level1Out35[4] , 
        \Level1Out35[3] , \Level1Out35[2] , \Level1Out35[1] , \Level1Out35[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_40 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink40[31] , \ScanLink40[30] , 
        \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , \ScanLink40[26] , 
        \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , \ScanLink40[22] , 
        \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , \ScanLink40[18] , 
        \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , \ScanLink40[14] , 
        \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , \ScanLink40[10] , 
        \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , \ScanLink40[6] , 
        \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , \ScanLink40[2] , 
        \ScanLink40[1] , \ScanLink40[0] }), .ScanOut({\ScanLink41[31] , 
        \ScanLink41[30] , \ScanLink41[29] , \ScanLink41[28] , \ScanLink41[27] , 
        \ScanLink41[26] , \ScanLink41[25] , \ScanLink41[24] , \ScanLink41[23] , 
        \ScanLink41[22] , \ScanLink41[21] , \ScanLink41[20] , \ScanLink41[19] , 
        \ScanLink41[18] , \ScanLink41[17] , \ScanLink41[16] , \ScanLink41[15] , 
        \ScanLink41[14] , \ScanLink41[13] , \ScanLink41[12] , \ScanLink41[11] , 
        \ScanLink41[10] , \ScanLink41[9] , \ScanLink41[8] , \ScanLink41[7] , 
        \ScanLink41[6] , \ScanLink41[5] , \ScanLink41[4] , \ScanLink41[3] , 
        \ScanLink41[2] , \ScanLink41[1] , \ScanLink41[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load40[0] ), .Out({
        \Level1Out40[31] , \Level1Out40[30] , \Level1Out40[29] , 
        \Level1Out40[28] , \Level1Out40[27] , \Level1Out40[26] , 
        \Level1Out40[25] , \Level1Out40[24] , \Level1Out40[23] , 
        \Level1Out40[22] , \Level1Out40[21] , \Level1Out40[20] , 
        \Level1Out40[19] , \Level1Out40[18] , \Level1Out40[17] , 
        \Level1Out40[16] , \Level1Out40[15] , \Level1Out40[14] , 
        \Level1Out40[13] , \Level1Out40[12] , \Level1Out40[11] , 
        \Level1Out40[10] , \Level1Out40[9] , \Level1Out40[8] , 
        \Level1Out40[7] , \Level1Out40[6] , \Level1Out40[5] , \Level1Out40[4] , 
        \Level1Out40[3] , \Level1Out40[2] , \Level1Out40[1] , \Level1Out40[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load48[0] ), .Out({\Level2Out48[31] , \Level2Out48[30] , 
        \Level2Out48[29] , \Level2Out48[28] , \Level2Out48[27] , 
        \Level2Out48[26] , \Level2Out48[25] , \Level2Out48[24] , 
        \Level2Out48[23] , \Level2Out48[22] , \Level2Out48[21] , 
        \Level2Out48[20] , \Level2Out48[19] , \Level2Out48[18] , 
        \Level2Out48[17] , \Level2Out48[16] , \Level2Out48[15] , 
        \Level2Out48[14] , \Level2Out48[13] , \Level2Out48[12] , 
        \Level2Out48[11] , \Level2Out48[10] , \Level2Out48[9] , 
        \Level2Out48[8] , \Level2Out48[7] , \Level2Out48[6] , \Level2Out48[5] , 
        \Level2Out48[4] , \Level2Out48[3] , \Level2Out48[2] , \Level2Out48[1] , 
        \Level2Out48[0] }), .In1({\Level1Out48[31] , \Level1Out48[30] , 
        \Level1Out48[29] , \Level1Out48[28] , \Level1Out48[27] , 
        \Level1Out48[26] , \Level1Out48[25] , \Level1Out48[24] , 
        \Level1Out48[23] , \Level1Out48[22] , \Level1Out48[21] , 
        \Level1Out48[20] , \Level1Out48[19] , \Level1Out48[18] , 
        \Level1Out48[17] , \Level1Out48[16] , \Level1Out48[15] , 
        \Level1Out48[14] , \Level1Out48[13] , \Level1Out48[12] , 
        \Level1Out48[11] , \Level1Out48[10] , \Level1Out48[9] , 
        \Level1Out48[8] , \Level1Out48[7] , \Level1Out48[6] , \Level1Out48[5] , 
        \Level1Out48[4] , \Level1Out48[3] , \Level1Out48[2] , \Level1Out48[1] , 
        \Level1Out48[0] }), .In2({\Level1Out49[31] , \Level1Out49[30] , 
        \Level1Out49[29] , \Level1Out49[28] , \Level1Out49[27] , 
        \Level1Out49[26] , \Level1Out49[25] , \Level1Out49[24] , 
        \Level1Out49[23] , \Level1Out49[22] , \Level1Out49[21] , 
        \Level1Out49[20] , \Level1Out49[19] , \Level1Out49[18] , 
        \Level1Out49[17] , \Level1Out49[16] , \Level1Out49[15] , 
        \Level1Out49[14] , \Level1Out49[13] , \Level1Out49[12] , 
        \Level1Out49[11] , \Level1Out49[10] , \Level1Out49[9] , 
        \Level1Out49[8] , \Level1Out49[7] , \Level1Out49[6] , \Level1Out49[5] , 
        \Level1Out49[4] , \Level1Out49[3] , \Level1Out49[2] , \Level1Out49[1] , 
        \Level1Out49[0] }), .Read1(\Level1Load48[0] ), .Read2(
        \Level1Load49[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_62_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load62[0] ), .Out({\Level2Out62[31] , \Level2Out62[30] , 
        \Level2Out62[29] , \Level2Out62[28] , \Level2Out62[27] , 
        \Level2Out62[26] , \Level2Out62[25] , \Level2Out62[24] , 
        \Level2Out62[23] , \Level2Out62[22] , \Level2Out62[21] , 
        \Level2Out62[20] , \Level2Out62[19] , \Level2Out62[18] , 
        \Level2Out62[17] , \Level2Out62[16] , \Level2Out62[15] , 
        \Level2Out62[14] , \Level2Out62[13] , \Level2Out62[12] , 
        \Level2Out62[11] , \Level2Out62[10] , \Level2Out62[9] , 
        \Level2Out62[8] , \Level2Out62[7] , \Level2Out62[6] , \Level2Out62[5] , 
        \Level2Out62[4] , \Level2Out62[3] , \Level2Out62[2] , \Level2Out62[1] , 
        \Level2Out62[0] }), .In1({\Level1Out62[31] , \Level1Out62[30] , 
        \Level1Out62[29] , \Level1Out62[28] , \Level1Out62[27] , 
        \Level1Out62[26] , \Level1Out62[25] , \Level1Out62[24] , 
        \Level1Out62[23] , \Level1Out62[22] , \Level1Out62[21] , 
        \Level1Out62[20] , \Level1Out62[19] , \Level1Out62[18] , 
        \Level1Out62[17] , \Level1Out62[16] , \Level1Out62[15] , 
        \Level1Out62[14] , \Level1Out62[13] , \Level1Out62[12] , 
        \Level1Out62[11] , \Level1Out62[10] , \Level1Out62[9] , 
        \Level1Out62[8] , \Level1Out62[7] , \Level1Out62[6] , \Level1Out62[5] , 
        \Level1Out62[4] , \Level1Out62[3] , \Level1Out62[2] , \Level1Out62[1] , 
        \Level1Out62[0] }), .In2({\Level1Out63[31] , \Level1Out63[30] , 
        \Level1Out63[29] , \Level1Out63[28] , \Level1Out63[27] , 
        \Level1Out63[26] , \Level1Out63[25] , \Level1Out63[24] , 
        \Level1Out63[23] , \Level1Out63[22] , \Level1Out63[21] , 
        \Level1Out63[20] , \Level1Out63[19] , \Level1Out63[18] , 
        \Level1Out63[17] , \Level1Out63[16] , \Level1Out63[15] , 
        \Level1Out63[14] , \Level1Out63[13] , \Level1Out63[12] , 
        \Level1Out63[11] , \Level1Out63[10] , \Level1Out63[9] , 
        \Level1Out63[8] , \Level1Out63[7] , \Level1Out63[6] , \Level1Out63[5] , 
        \Level1Out63[4] , \Level1Out63[3] , \Level1Out63[2] , \Level1Out63[1] , 
        \Level1Out63[0] }), .Read1(\Level1Load62[0] ), .Read2(
        \Level1Load63[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load16[0] ), .Out({\Level8Out16[31] , \Level8Out16[30] , 
        \Level8Out16[29] , \Level8Out16[28] , \Level8Out16[27] , 
        \Level8Out16[26] , \Level8Out16[25] , \Level8Out16[24] , 
        \Level8Out16[23] , \Level8Out16[22] , \Level8Out16[21] , 
        \Level8Out16[20] , \Level8Out16[19] , \Level8Out16[18] , 
        \Level8Out16[17] , \Level8Out16[16] , \Level8Out16[15] , 
        \Level8Out16[14] , \Level8Out16[13] , \Level8Out16[12] , 
        \Level8Out16[11] , \Level8Out16[10] , \Level8Out16[9] , 
        \Level8Out16[8] , \Level8Out16[7] , \Level8Out16[6] , \Level8Out16[5] , 
        \Level8Out16[4] , \Level8Out16[3] , \Level8Out16[2] , \Level8Out16[1] , 
        \Level8Out16[0] }), .In1({\Level4Out16[31] , \Level4Out16[30] , 
        \Level4Out16[29] , \Level4Out16[28] , \Level4Out16[27] , 
        \Level4Out16[26] , \Level4Out16[25] , \Level4Out16[24] , 
        \Level4Out16[23] , \Level4Out16[22] , \Level4Out16[21] , 
        \Level4Out16[20] , \Level4Out16[19] , \Level4Out16[18] , 
        \Level4Out16[17] , \Level4Out16[16] , \Level4Out16[15] , 
        \Level4Out16[14] , \Level4Out16[13] , \Level4Out16[12] , 
        \Level4Out16[11] , \Level4Out16[10] , \Level4Out16[9] , 
        \Level4Out16[8] , \Level4Out16[7] , \Level4Out16[6] , \Level4Out16[5] , 
        \Level4Out16[4] , \Level4Out16[3] , \Level4Out16[2] , \Level4Out16[1] , 
        \Level4Out16[0] }), .In2({\Level4Out20[31] , \Level4Out20[30] , 
        \Level4Out20[29] , \Level4Out20[28] , \Level4Out20[27] , 
        \Level4Out20[26] , \Level4Out20[25] , \Level4Out20[24] , 
        \Level4Out20[23] , \Level4Out20[22] , \Level4Out20[21] , 
        \Level4Out20[20] , \Level4Out20[19] , \Level4Out20[18] , 
        \Level4Out20[17] , \Level4Out20[16] , \Level4Out20[15] , 
        \Level4Out20[14] , \Level4Out20[13] , \Level4Out20[12] , 
        \Level4Out20[11] , \Level4Out20[10] , \Level4Out20[9] , 
        \Level4Out20[8] , \Level4Out20[7] , \Level4Out20[6] , \Level4Out20[5] , 
        \Level4Out20[4] , \Level4Out20[3] , \Level4Out20[2] , \Level4Out20[1] , 
        \Level4Out20[0] }), .Read1(\Level4Load16[0] ), .Read2(
        \Level4Load20[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load56[0] ), .Out({\Level8Out56[31] , \Level8Out56[30] , 
        \Level8Out56[29] , \Level8Out56[28] , \Level8Out56[27] , 
        \Level8Out56[26] , \Level8Out56[25] , \Level8Out56[24] , 
        \Level8Out56[23] , \Level8Out56[22] , \Level8Out56[21] , 
        \Level8Out56[20] , \Level8Out56[19] , \Level8Out56[18] , 
        \Level8Out56[17] , \Level8Out56[16] , \Level8Out56[15] , 
        \Level8Out56[14] , \Level8Out56[13] , \Level8Out56[12] , 
        \Level8Out56[11] , \Level8Out56[10] , \Level8Out56[9] , 
        \Level8Out56[8] , \Level8Out56[7] , \Level8Out56[6] , \Level8Out56[5] , 
        \Level8Out56[4] , \Level8Out56[3] , \Level8Out56[2] , \Level8Out56[1] , 
        \Level8Out56[0] }), .In1({\Level4Out56[31] , \Level4Out56[30] , 
        \Level4Out56[29] , \Level4Out56[28] , \Level4Out56[27] , 
        \Level4Out56[26] , \Level4Out56[25] , \Level4Out56[24] , 
        \Level4Out56[23] , \Level4Out56[22] , \Level4Out56[21] , 
        \Level4Out56[20] , \Level4Out56[19] , \Level4Out56[18] , 
        \Level4Out56[17] , \Level4Out56[16] , \Level4Out56[15] , 
        \Level4Out56[14] , \Level4Out56[13] , \Level4Out56[12] , 
        \Level4Out56[11] , \Level4Out56[10] , \Level4Out56[9] , 
        \Level4Out56[8] , \Level4Out56[7] , \Level4Out56[6] , \Level4Out56[5] , 
        \Level4Out56[4] , \Level4Out56[3] , \Level4Out56[2] , \Level4Out56[1] , 
        \Level4Out56[0] }), .In2({\Level4Out60[31] , \Level4Out60[30] , 
        \Level4Out60[29] , \Level4Out60[28] , \Level4Out60[27] , 
        \Level4Out60[26] , \Level4Out60[25] , \Level4Out60[24] , 
        \Level4Out60[23] , \Level4Out60[22] , \Level4Out60[21] , 
        \Level4Out60[20] , \Level4Out60[19] , \Level4Out60[18] , 
        \Level4Out60[17] , \Level4Out60[16] , \Level4Out60[15] , 
        \Level4Out60[14] , \Level4Out60[13] , \Level4Out60[12] , 
        \Level4Out60[11] , \Level4Out60[10] , \Level4Out60[9] , 
        \Level4Out60[8] , \Level4Out60[7] , \Level4Out60[6] , \Level4Out60[5] , 
        \Level4Out60[4] , \Level4Out60[3] , \Level4Out60[2] , \Level4Out60[1] , 
        \Level4Out60[0] }), .Read1(\Level4Load56[0] ), .Read2(
        \Level4Load60[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load48[0] ), .Out({\Level16Out48[31] , \Level16Out48[30] , 
        \Level16Out48[29] , \Level16Out48[28] , \Level16Out48[27] , 
        \Level16Out48[26] , \Level16Out48[25] , \Level16Out48[24] , 
        \Level16Out48[23] , \Level16Out48[22] , \Level16Out48[21] , 
        \Level16Out48[20] , \Level16Out48[19] , \Level16Out48[18] , 
        \Level16Out48[17] , \Level16Out48[16] , \Level16Out48[15] , 
        \Level16Out48[14] , \Level16Out48[13] , \Level16Out48[12] , 
        \Level16Out48[11] , \Level16Out48[10] , \Level16Out48[9] , 
        \Level16Out48[8] , \Level16Out48[7] , \Level16Out48[6] , 
        \Level16Out48[5] , \Level16Out48[4] , \Level16Out48[3] , 
        \Level16Out48[2] , \Level16Out48[1] , \Level16Out48[0] }), .In1({
        \Level8Out48[31] , \Level8Out48[30] , \Level8Out48[29] , 
        \Level8Out48[28] , \Level8Out48[27] , \Level8Out48[26] , 
        \Level8Out48[25] , \Level8Out48[24] , \Level8Out48[23] , 
        \Level8Out48[22] , \Level8Out48[21] , \Level8Out48[20] , 
        \Level8Out48[19] , \Level8Out48[18] , \Level8Out48[17] , 
        \Level8Out48[16] , \Level8Out48[15] , \Level8Out48[14] , 
        \Level8Out48[13] , \Level8Out48[12] , \Level8Out48[11] , 
        \Level8Out48[10] , \Level8Out48[9] , \Level8Out48[8] , 
        \Level8Out48[7] , \Level8Out48[6] , \Level8Out48[5] , \Level8Out48[4] , 
        \Level8Out48[3] , \Level8Out48[2] , \Level8Out48[1] , \Level8Out48[0] 
        }), .In2({\Level8Out56[31] , \Level8Out56[30] , \Level8Out56[29] , 
        \Level8Out56[28] , \Level8Out56[27] , \Level8Out56[26] , 
        \Level8Out56[25] , \Level8Out56[24] , \Level8Out56[23] , 
        \Level8Out56[22] , \Level8Out56[21] , \Level8Out56[20] , 
        \Level8Out56[19] , \Level8Out56[18] , \Level8Out56[17] , 
        \Level8Out56[16] , \Level8Out56[15] , \Level8Out56[14] , 
        \Level8Out56[13] , \Level8Out56[12] , \Level8Out56[11] , 
        \Level8Out56[10] , \Level8Out56[9] , \Level8Out56[8] , 
        \Level8Out56[7] , \Level8Out56[6] , \Level8Out56[5] , \Level8Out56[4] , 
        \Level8Out56[3] , \Level8Out56[2] , \Level8Out56[1] , \Level8Out56[0] 
        }), .Read1(\Level8Load48[0] ), .Read2(\Level8Load56[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load8[0] ), .Out({\Level2Out8[31] , \Level2Out8[30] , 
        \Level2Out8[29] , \Level2Out8[28] , \Level2Out8[27] , \Level2Out8[26] , 
        \Level2Out8[25] , \Level2Out8[24] , \Level2Out8[23] , \Level2Out8[22] , 
        \Level2Out8[21] , \Level2Out8[20] , \Level2Out8[19] , \Level2Out8[18] , 
        \Level2Out8[17] , \Level2Out8[16] , \Level2Out8[15] , \Level2Out8[14] , 
        \Level2Out8[13] , \Level2Out8[12] , \Level2Out8[11] , \Level2Out8[10] , 
        \Level2Out8[9] , \Level2Out8[8] , \Level2Out8[7] , \Level2Out8[6] , 
        \Level2Out8[5] , \Level2Out8[4] , \Level2Out8[3] , \Level2Out8[2] , 
        \Level2Out8[1] , \Level2Out8[0] }), .In1({\Level1Out8[31] , 
        \Level1Out8[30] , \Level1Out8[29] , \Level1Out8[28] , \Level1Out8[27] , 
        \Level1Out8[26] , \Level1Out8[25] , \Level1Out8[24] , \Level1Out8[23] , 
        \Level1Out8[22] , \Level1Out8[21] , \Level1Out8[20] , \Level1Out8[19] , 
        \Level1Out8[18] , \Level1Out8[17] , \Level1Out8[16] , \Level1Out8[15] , 
        \Level1Out8[14] , \Level1Out8[13] , \Level1Out8[12] , \Level1Out8[11] , 
        \Level1Out8[10] , \Level1Out8[9] , \Level1Out8[8] , \Level1Out8[7] , 
        \Level1Out8[6] , \Level1Out8[5] , \Level1Out8[4] , \Level1Out8[3] , 
        \Level1Out8[2] , \Level1Out8[1] , \Level1Out8[0] }), .In2({
        \Level1Out9[31] , \Level1Out9[30] , \Level1Out9[29] , \Level1Out9[28] , 
        \Level1Out9[27] , \Level1Out9[26] , \Level1Out9[25] , \Level1Out9[24] , 
        \Level1Out9[23] , \Level1Out9[22] , \Level1Out9[21] , \Level1Out9[20] , 
        \Level1Out9[19] , \Level1Out9[18] , \Level1Out9[17] , \Level1Out9[16] , 
        \Level1Out9[15] , \Level1Out9[14] , \Level1Out9[13] , \Level1Out9[12] , 
        \Level1Out9[11] , \Level1Out9[10] , \Level1Out9[9] , \Level1Out9[8] , 
        \Level1Out9[7] , \Level1Out9[6] , \Level1Out9[5] , \Level1Out9[4] , 
        \Level1Out9[3] , \Level1Out9[2] , \Level1Out9[1] , \Level1Out9[0] }), 
        .Read1(\Level1Load8[0] ), .Read2(\Level1Load9[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_27 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink27[31] , \ScanLink27[30] , 
        \ScanLink27[29] , \ScanLink27[28] , \ScanLink27[27] , \ScanLink27[26] , 
        \ScanLink27[25] , \ScanLink27[24] , \ScanLink27[23] , \ScanLink27[22] , 
        \ScanLink27[21] , \ScanLink27[20] , \ScanLink27[19] , \ScanLink27[18] , 
        \ScanLink27[17] , \ScanLink27[16] , \ScanLink27[15] , \ScanLink27[14] , 
        \ScanLink27[13] , \ScanLink27[12] , \ScanLink27[11] , \ScanLink27[10] , 
        \ScanLink27[9] , \ScanLink27[8] , \ScanLink27[7] , \ScanLink27[6] , 
        \ScanLink27[5] , \ScanLink27[4] , \ScanLink27[3] , \ScanLink27[2] , 
        \ScanLink27[1] , \ScanLink27[0] }), .ScanOut({\ScanLink28[31] , 
        \ScanLink28[30] , \ScanLink28[29] , \ScanLink28[28] , \ScanLink28[27] , 
        \ScanLink28[26] , \ScanLink28[25] , \ScanLink28[24] , \ScanLink28[23] , 
        \ScanLink28[22] , \ScanLink28[21] , \ScanLink28[20] , \ScanLink28[19] , 
        \ScanLink28[18] , \ScanLink28[17] , \ScanLink28[16] , \ScanLink28[15] , 
        \ScanLink28[14] , \ScanLink28[13] , \ScanLink28[12] , \ScanLink28[11] , 
        \ScanLink28[10] , \ScanLink28[9] , \ScanLink28[8] , \ScanLink28[7] , 
        \ScanLink28[6] , \ScanLink28[5] , \ScanLink28[4] , \ScanLink28[3] , 
        \ScanLink28[2] , \ScanLink28[1] , \ScanLink28[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load27[0] ), .Out({
        \Level1Out27[31] , \Level1Out27[30] , \Level1Out27[29] , 
        \Level1Out27[28] , \Level1Out27[27] , \Level1Out27[26] , 
        \Level1Out27[25] , \Level1Out27[24] , \Level1Out27[23] , 
        \Level1Out27[22] , \Level1Out27[21] , \Level1Out27[20] , 
        \Level1Out27[19] , \Level1Out27[18] , \Level1Out27[17] , 
        \Level1Out27[16] , \Level1Out27[15] , \Level1Out27[14] , 
        \Level1Out27[13] , \Level1Out27[12] , \Level1Out27[11] , 
        \Level1Out27[10] , \Level1Out27[9] , \Level1Out27[8] , 
        \Level1Out27[7] , \Level1Out27[6] , \Level1Out27[5] , \Level1Out27[4] , 
        \Level1Out27[3] , \Level1Out27[2] , \Level1Out27[1] , \Level1Out27[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_50_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load50[0] ), .Out({\Level2Out50[31] , \Level2Out50[30] , 
        \Level2Out50[29] , \Level2Out50[28] , \Level2Out50[27] , 
        \Level2Out50[26] , \Level2Out50[25] , \Level2Out50[24] , 
        \Level2Out50[23] , \Level2Out50[22] , \Level2Out50[21] , 
        \Level2Out50[20] , \Level2Out50[19] , \Level2Out50[18] , 
        \Level2Out50[17] , \Level2Out50[16] , \Level2Out50[15] , 
        \Level2Out50[14] , \Level2Out50[13] , \Level2Out50[12] , 
        \Level2Out50[11] , \Level2Out50[10] , \Level2Out50[9] , 
        \Level2Out50[8] , \Level2Out50[7] , \Level2Out50[6] , \Level2Out50[5] , 
        \Level2Out50[4] , \Level2Out50[3] , \Level2Out50[2] , \Level2Out50[1] , 
        \Level2Out50[0] }), .In1({\Level1Out50[31] , \Level1Out50[30] , 
        \Level1Out50[29] , \Level1Out50[28] , \Level1Out50[27] , 
        \Level1Out50[26] , \Level1Out50[25] , \Level1Out50[24] , 
        \Level1Out50[23] , \Level1Out50[22] , \Level1Out50[21] , 
        \Level1Out50[20] , \Level1Out50[19] , \Level1Out50[18] , 
        \Level1Out50[17] , \Level1Out50[16] , \Level1Out50[15] , 
        \Level1Out50[14] , \Level1Out50[13] , \Level1Out50[12] , 
        \Level1Out50[11] , \Level1Out50[10] , \Level1Out50[9] , 
        \Level1Out50[8] , \Level1Out50[7] , \Level1Out50[6] , \Level1Out50[5] , 
        \Level1Out50[4] , \Level1Out50[3] , \Level1Out50[2] , \Level1Out50[1] , 
        \Level1Out50[0] }), .In2({\Level1Out51[31] , \Level1Out51[30] , 
        \Level1Out51[29] , \Level1Out51[28] , \Level1Out51[27] , 
        \Level1Out51[26] , \Level1Out51[25] , \Level1Out51[24] , 
        \Level1Out51[23] , \Level1Out51[22] , \Level1Out51[21] , 
        \Level1Out51[20] , \Level1Out51[19] , \Level1Out51[18] , 
        \Level1Out51[17] , \Level1Out51[16] , \Level1Out51[15] , 
        \Level1Out51[14] , \Level1Out51[13] , \Level1Out51[12] , 
        \Level1Out51[11] , \Level1Out51[10] , \Level1Out51[9] , 
        \Level1Out51[8] , \Level1Out51[7] , \Level1Out51[6] , \Level1Out51[5] , 
        \Level1Out51[4] , \Level1Out51[3] , \Level1Out51[2] , \Level1Out51[1] , 
        \Level1Out51[0] }), .Read1(\Level1Load50[0] ), .Read2(
        \Level1Load51[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_49 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink49[31] , \ScanLink49[30] , 
        \ScanLink49[29] , \ScanLink49[28] , \ScanLink49[27] , \ScanLink49[26] , 
        \ScanLink49[25] , \ScanLink49[24] , \ScanLink49[23] , \ScanLink49[22] , 
        \ScanLink49[21] , \ScanLink49[20] , \ScanLink49[19] , \ScanLink49[18] , 
        \ScanLink49[17] , \ScanLink49[16] , \ScanLink49[15] , \ScanLink49[14] , 
        \ScanLink49[13] , \ScanLink49[12] , \ScanLink49[11] , \ScanLink49[10] , 
        \ScanLink49[9] , \ScanLink49[8] , \ScanLink49[7] , \ScanLink49[6] , 
        \ScanLink49[5] , \ScanLink49[4] , \ScanLink49[3] , \ScanLink49[2] , 
        \ScanLink49[1] , \ScanLink49[0] }), .ScanOut({\ScanLink50[31] , 
        \ScanLink50[30] , \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , 
        \ScanLink50[26] , \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , 
        \ScanLink50[22] , \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , 
        \ScanLink50[18] , \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , 
        \ScanLink50[14] , \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , 
        \ScanLink50[10] , \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , 
        \ScanLink50[6] , \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , 
        \ScanLink50[2] , \ScanLink50[1] , \ScanLink50[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load49[0] ), .Out({
        \Level1Out49[31] , \Level1Out49[30] , \Level1Out49[29] , 
        \Level1Out49[28] , \Level1Out49[27] , \Level1Out49[26] , 
        \Level1Out49[25] , \Level1Out49[24] , \Level1Out49[23] , 
        \Level1Out49[22] , \Level1Out49[21] , \Level1Out49[20] , 
        \Level1Out49[19] , \Level1Out49[18] , \Level1Out49[17] , 
        \Level1Out49[16] , \Level1Out49[15] , \Level1Out49[14] , 
        \Level1Out49[13] , \Level1Out49[12] , \Level1Out49[11] , 
        \Level1Out49[10] , \Level1Out49[9] , \Level1Out49[8] , 
        \Level1Out49[7] , \Level1Out49[6] , \Level1Out49[5] , \Level1Out49[4] , 
        \Level1Out49[3] , \Level1Out49[2] , \Level1Out49[1] , \Level1Out49[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_36_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load36[0] ), .Out({\Level4Out36[31] , \Level4Out36[30] , 
        \Level4Out36[29] , \Level4Out36[28] , \Level4Out36[27] , 
        \Level4Out36[26] , \Level4Out36[25] , \Level4Out36[24] , 
        \Level4Out36[23] , \Level4Out36[22] , \Level4Out36[21] , 
        \Level4Out36[20] , \Level4Out36[19] , \Level4Out36[18] , 
        \Level4Out36[17] , \Level4Out36[16] , \Level4Out36[15] , 
        \Level4Out36[14] , \Level4Out36[13] , \Level4Out36[12] , 
        \Level4Out36[11] , \Level4Out36[10] , \Level4Out36[9] , 
        \Level4Out36[8] , \Level4Out36[7] , \Level4Out36[6] , \Level4Out36[5] , 
        \Level4Out36[4] , \Level4Out36[3] , \Level4Out36[2] , \Level4Out36[1] , 
        \Level4Out36[0] }), .In1({\Level2Out36[31] , \Level2Out36[30] , 
        \Level2Out36[29] , \Level2Out36[28] , \Level2Out36[27] , 
        \Level2Out36[26] , \Level2Out36[25] , \Level2Out36[24] , 
        \Level2Out36[23] , \Level2Out36[22] , \Level2Out36[21] , 
        \Level2Out36[20] , \Level2Out36[19] , \Level2Out36[18] , 
        \Level2Out36[17] , \Level2Out36[16] , \Level2Out36[15] , 
        \Level2Out36[14] , \Level2Out36[13] , \Level2Out36[12] , 
        \Level2Out36[11] , \Level2Out36[10] , \Level2Out36[9] , 
        \Level2Out36[8] , \Level2Out36[7] , \Level2Out36[6] , \Level2Out36[5] , 
        \Level2Out36[4] , \Level2Out36[3] , \Level2Out36[2] , \Level2Out36[1] , 
        \Level2Out36[0] }), .In2({\Level2Out38[31] , \Level2Out38[30] , 
        \Level2Out38[29] , \Level2Out38[28] , \Level2Out38[27] , 
        \Level2Out38[26] , \Level2Out38[25] , \Level2Out38[24] , 
        \Level2Out38[23] , \Level2Out38[22] , \Level2Out38[21] , 
        \Level2Out38[20] , \Level2Out38[19] , \Level2Out38[18] , 
        \Level2Out38[17] , \Level2Out38[16] , \Level2Out38[15] , 
        \Level2Out38[14] , \Level2Out38[13] , \Level2Out38[12] , 
        \Level2Out38[11] , \Level2Out38[10] , \Level2Out38[9] , 
        \Level2Out38[8] , \Level2Out38[7] , \Level2Out38[6] , \Level2Out38[5] , 
        \Level2Out38[4] , \Level2Out38[3] , \Level2Out38[2] , \Level2Out38[1] , 
        \Level2Out38[0] }), .Read1(\Level2Load36[0] ), .Read2(
        \Level2Load38[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_52 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink52[31] , \ScanLink52[30] , 
        \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , \ScanLink52[26] , 
        \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , \ScanLink52[22] , 
        \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , \ScanLink52[18] , 
        \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , \ScanLink52[14] , 
        \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , \ScanLink52[10] , 
        \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , \ScanLink52[6] , 
        \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , \ScanLink52[2] , 
        \ScanLink52[1] , \ScanLink52[0] }), .ScanOut({\ScanLink53[31] , 
        \ScanLink53[30] , \ScanLink53[29] , \ScanLink53[28] , \ScanLink53[27] , 
        \ScanLink53[26] , \ScanLink53[25] , \ScanLink53[24] , \ScanLink53[23] , 
        \ScanLink53[22] , \ScanLink53[21] , \ScanLink53[20] , \ScanLink53[19] , 
        \ScanLink53[18] , \ScanLink53[17] , \ScanLink53[16] , \ScanLink53[15] , 
        \ScanLink53[14] , \ScanLink53[13] , \ScanLink53[12] , \ScanLink53[11] , 
        \ScanLink53[10] , \ScanLink53[9] , \ScanLink53[8] , \ScanLink53[7] , 
        \ScanLink53[6] , \ScanLink53[5] , \ScanLink53[4] , \ScanLink53[3] , 
        \ScanLink53[2] , \ScanLink53[1] , \ScanLink53[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load52[0] ), .Out({
        \Level1Out52[31] , \Level1Out52[30] , \Level1Out52[29] , 
        \Level1Out52[28] , \Level1Out52[27] , \Level1Out52[26] , 
        \Level1Out52[25] , \Level1Out52[24] , \Level1Out52[23] , 
        \Level1Out52[22] , \Level1Out52[21] , \Level1Out52[20] , 
        \Level1Out52[19] , \Level1Out52[18] , \Level1Out52[17] , 
        \Level1Out52[16] , \Level1Out52[15] , \Level1Out52[14] , 
        \Level1Out52[13] , \Level1Out52[12] , \Level1Out52[11] , 
        \Level1Out52[10] , \Level1Out52[9] , \Level1Out52[8] , 
        \Level1Out52[7] , \Level1Out52[6] , \Level1Out52[5] , \Level1Out52[4] , 
        \Level1Out52[3] , \Level1Out52[2] , \Level1Out52[1] , \Level1Out52[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_18_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load18[0] ), .Out({\Level2Out18[31] , \Level2Out18[30] , 
        \Level2Out18[29] , \Level2Out18[28] , \Level2Out18[27] , 
        \Level2Out18[26] , \Level2Out18[25] , \Level2Out18[24] , 
        \Level2Out18[23] , \Level2Out18[22] , \Level2Out18[21] , 
        \Level2Out18[20] , \Level2Out18[19] , \Level2Out18[18] , 
        \Level2Out18[17] , \Level2Out18[16] , \Level2Out18[15] , 
        \Level2Out18[14] , \Level2Out18[13] , \Level2Out18[12] , 
        \Level2Out18[11] , \Level2Out18[10] , \Level2Out18[9] , 
        \Level2Out18[8] , \Level2Out18[7] , \Level2Out18[6] , \Level2Out18[5] , 
        \Level2Out18[4] , \Level2Out18[3] , \Level2Out18[2] , \Level2Out18[1] , 
        \Level2Out18[0] }), .In1({\Level1Out18[31] , \Level1Out18[30] , 
        \Level1Out18[29] , \Level1Out18[28] , \Level1Out18[27] , 
        \Level1Out18[26] , \Level1Out18[25] , \Level1Out18[24] , 
        \Level1Out18[23] , \Level1Out18[22] , \Level1Out18[21] , 
        \Level1Out18[20] , \Level1Out18[19] , \Level1Out18[18] , 
        \Level1Out18[17] , \Level1Out18[16] , \Level1Out18[15] , 
        \Level1Out18[14] , \Level1Out18[13] , \Level1Out18[12] , 
        \Level1Out18[11] , \Level1Out18[10] , \Level1Out18[9] , 
        \Level1Out18[8] , \Level1Out18[7] , \Level1Out18[6] , \Level1Out18[5] , 
        \Level1Out18[4] , \Level1Out18[3] , \Level1Out18[2] , \Level1Out18[1] , 
        \Level1Out18[0] }), .In2({\Level1Out19[31] , \Level1Out19[30] , 
        \Level1Out19[29] , \Level1Out19[28] , \Level1Out19[27] , 
        \Level1Out19[26] , \Level1Out19[25] , \Level1Out19[24] , 
        \Level1Out19[23] , \Level1Out19[22] , \Level1Out19[21] , 
        \Level1Out19[20] , \Level1Out19[19] , \Level1Out19[18] , 
        \Level1Out19[17] , \Level1Out19[16] , \Level1Out19[15] , 
        \Level1Out19[14] , \Level1Out19[13] , \Level1Out19[12] , 
        \Level1Out19[11] , \Level1Out19[10] , \Level1Out19[9] , 
        \Level1Out19[8] , \Level1Out19[7] , \Level1Out19[6] , \Level1Out19[5] , 
        \Level1Out19[4] , \Level1Out19[3] , \Level1Out19[2] , \Level1Out19[1] , 
        \Level1Out19[0] }), .Read1(\Level1Load18[0] ), .Read2(
        \Level1Load19[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load32[0] ), .Out({\Level2Out32[31] , \Level2Out32[30] , 
        \Level2Out32[29] , \Level2Out32[28] , \Level2Out32[27] , 
        \Level2Out32[26] , \Level2Out32[25] , \Level2Out32[24] , 
        \Level2Out32[23] , \Level2Out32[22] , \Level2Out32[21] , 
        \Level2Out32[20] , \Level2Out32[19] , \Level2Out32[18] , 
        \Level2Out32[17] , \Level2Out32[16] , \Level2Out32[15] , 
        \Level2Out32[14] , \Level2Out32[13] , \Level2Out32[12] , 
        \Level2Out32[11] , \Level2Out32[10] , \Level2Out32[9] , 
        \Level2Out32[8] , \Level2Out32[7] , \Level2Out32[6] , \Level2Out32[5] , 
        \Level2Out32[4] , \Level2Out32[3] , \Level2Out32[2] , \Level2Out32[1] , 
        \Level2Out32[0] }), .In1({\Level1Out32[31] , \Level1Out32[30] , 
        \Level1Out32[29] , \Level1Out32[28] , \Level1Out32[27] , 
        \Level1Out32[26] , \Level1Out32[25] , \Level1Out32[24] , 
        \Level1Out32[23] , \Level1Out32[22] , \Level1Out32[21] , 
        \Level1Out32[20] , \Level1Out32[19] , \Level1Out32[18] , 
        \Level1Out32[17] , \Level1Out32[16] , \Level1Out32[15] , 
        \Level1Out32[14] , \Level1Out32[13] , \Level1Out32[12] , 
        \Level1Out32[11] , \Level1Out32[10] , \Level1Out32[9] , 
        \Level1Out32[8] , \Level1Out32[7] , \Level1Out32[6] , \Level1Out32[5] , 
        \Level1Out32[4] , \Level1Out32[3] , \Level1Out32[2] , \Level1Out32[1] , 
        \Level1Out32[0] }), .In2({\Level1Out33[31] , \Level1Out33[30] , 
        \Level1Out33[29] , \Level1Out33[28] , \Level1Out33[27] , 
        \Level1Out33[26] , \Level1Out33[25] , \Level1Out33[24] , 
        \Level1Out33[23] , \Level1Out33[22] , \Level1Out33[21] , 
        \Level1Out33[20] , \Level1Out33[19] , \Level1Out33[18] , 
        \Level1Out33[17] , \Level1Out33[16] , \Level1Out33[15] , 
        \Level1Out33[14] , \Level1Out33[13] , \Level1Out33[12] , 
        \Level1Out33[11] , \Level1Out33[10] , \Level1Out33[9] , 
        \Level1Out33[8] , \Level1Out33[7] , \Level1Out33[6] , \Level1Out33[5] , 
        \Level1Out33[4] , \Level1Out33[3] , \Level1Out33[2] , \Level1Out33[1] , 
        \Level1Out33[0] }), .Read1(\Level1Load32[0] ), .Read2(
        \Level1Load33[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_55 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink55[31] , \ScanLink55[30] , 
        \ScanLink55[29] , \ScanLink55[28] , \ScanLink55[27] , \ScanLink55[26] , 
        \ScanLink55[25] , \ScanLink55[24] , \ScanLink55[23] , \ScanLink55[22] , 
        \ScanLink55[21] , \ScanLink55[20] , \ScanLink55[19] , \ScanLink55[18] , 
        \ScanLink55[17] , \ScanLink55[16] , \ScanLink55[15] , \ScanLink55[14] , 
        \ScanLink55[13] , \ScanLink55[12] , \ScanLink55[11] , \ScanLink55[10] , 
        \ScanLink55[9] , \ScanLink55[8] , \ScanLink55[7] , \ScanLink55[6] , 
        \ScanLink55[5] , \ScanLink55[4] , \ScanLink55[3] , \ScanLink55[2] , 
        \ScanLink55[1] , \ScanLink55[0] }), .ScanOut({\ScanLink56[31] , 
        \ScanLink56[30] , \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , 
        \ScanLink56[26] , \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , 
        \ScanLink56[22] , \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , 
        \ScanLink56[18] , \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , 
        \ScanLink56[14] , \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , 
        \ScanLink56[10] , \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , 
        \ScanLink56[6] , \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , 
        \ScanLink56[2] , \ScanLink56[1] , \ScanLink56[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load55[0] ), .Out({
        \Level1Out55[31] , \Level1Out55[30] , \Level1Out55[29] , 
        \Level1Out55[28] , \Level1Out55[27] , \Level1Out55[26] , 
        \Level1Out55[25] , \Level1Out55[24] , \Level1Out55[23] , 
        \Level1Out55[22] , \Level1Out55[21] , \Level1Out55[20] , 
        \Level1Out55[19] , \Level1Out55[18] , \Level1Out55[17] , 
        \Level1Out55[16] , \Level1Out55[15] , \Level1Out55[14] , 
        \Level1Out55[13] , \Level1Out55[12] , \Level1Out55[11] , 
        \Level1Out55[10] , \Level1Out55[9] , \Level1Out55[8] , 
        \Level1Out55[7] , \Level1Out55[6] , \Level1Out55[5] , \Level1Out55[4] , 
        \Level1Out55[3] , \Level1Out55[2] , \Level1Out55[1] , \Level1Out55[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_26_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load26[0] ), .Out({\Level2Out26[31] , \Level2Out26[30] , 
        \Level2Out26[29] , \Level2Out26[28] , \Level2Out26[27] , 
        \Level2Out26[26] , \Level2Out26[25] , \Level2Out26[24] , 
        \Level2Out26[23] , \Level2Out26[22] , \Level2Out26[21] , 
        \Level2Out26[20] , \Level2Out26[19] , \Level2Out26[18] , 
        \Level2Out26[17] , \Level2Out26[16] , \Level2Out26[15] , 
        \Level2Out26[14] , \Level2Out26[13] , \Level2Out26[12] , 
        \Level2Out26[11] , \Level2Out26[10] , \Level2Out26[9] , 
        \Level2Out26[8] , \Level2Out26[7] , \Level2Out26[6] , \Level2Out26[5] , 
        \Level2Out26[4] , \Level2Out26[3] , \Level2Out26[2] , \Level2Out26[1] , 
        \Level2Out26[0] }), .In1({\Level1Out26[31] , \Level1Out26[30] , 
        \Level1Out26[29] , \Level1Out26[28] , \Level1Out26[27] , 
        \Level1Out26[26] , \Level1Out26[25] , \Level1Out26[24] , 
        \Level1Out26[23] , \Level1Out26[22] , \Level1Out26[21] , 
        \Level1Out26[20] , \Level1Out26[19] , \Level1Out26[18] , 
        \Level1Out26[17] , \Level1Out26[16] , \Level1Out26[15] , 
        \Level1Out26[14] , \Level1Out26[13] , \Level1Out26[12] , 
        \Level1Out26[11] , \Level1Out26[10] , \Level1Out26[9] , 
        \Level1Out26[8] , \Level1Out26[7] , \Level1Out26[6] , \Level1Out26[5] , 
        \Level1Out26[4] , \Level1Out26[3] , \Level1Out26[2] , \Level1Out26[1] , 
        \Level1Out26[0] }), .In2({\Level1Out27[31] , \Level1Out27[30] , 
        \Level1Out27[29] , \Level1Out27[28] , \Level1Out27[27] , 
        \Level1Out27[26] , \Level1Out27[25] , \Level1Out27[24] , 
        \Level1Out27[23] , \Level1Out27[22] , \Level1Out27[21] , 
        \Level1Out27[20] , \Level1Out27[19] , \Level1Out27[18] , 
        \Level1Out27[17] , \Level1Out27[16] , \Level1Out27[15] , 
        \Level1Out27[14] , \Level1Out27[13] , \Level1Out27[12] , 
        \Level1Out27[11] , \Level1Out27[10] , \Level1Out27[9] , 
        \Level1Out27[8] , \Level1Out27[7] , \Level1Out27[6] , \Level1Out27[5] , 
        \Level1Out27[4] , \Level1Out27[3] , \Level1Out27[2] , \Level1Out27[1] , 
        \Level1Out27[0] }), .Read1(\Level1Load26[0] ), .Read2(
        \Level1Load27[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_9 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink9[31] , \ScanLink9[30] , 
        \ScanLink9[29] , \ScanLink9[28] , \ScanLink9[27] , \ScanLink9[26] , 
        \ScanLink9[25] , \ScanLink9[24] , \ScanLink9[23] , \ScanLink9[22] , 
        \ScanLink9[21] , \ScanLink9[20] , \ScanLink9[19] , \ScanLink9[18] , 
        \ScanLink9[17] , \ScanLink9[16] , \ScanLink9[15] , \ScanLink9[14] , 
        \ScanLink9[13] , \ScanLink9[12] , \ScanLink9[11] , \ScanLink9[10] , 
        \ScanLink9[9] , \ScanLink9[8] , \ScanLink9[7] , \ScanLink9[6] , 
        \ScanLink9[5] , \ScanLink9[4] , \ScanLink9[3] , \ScanLink9[2] , 
        \ScanLink9[1] , \ScanLink9[0] }), .ScanOut({\ScanLink10[31] , 
        \ScanLink10[30] , \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , 
        \ScanLink10[26] , \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , 
        \ScanLink10[22] , \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , 
        \ScanLink10[18] , \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , 
        \ScanLink10[14] , \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , 
        \ScanLink10[10] , \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , 
        \ScanLink10[6] , \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , 
        \ScanLink10[2] , \ScanLink10[1] , \ScanLink10[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load9[0] ), .Out({
        \Level1Out9[31] , \Level1Out9[30] , \Level1Out9[29] , \Level1Out9[28] , 
        \Level1Out9[27] , \Level1Out9[26] , \Level1Out9[25] , \Level1Out9[24] , 
        \Level1Out9[23] , \Level1Out9[22] , \Level1Out9[21] , \Level1Out9[20] , 
        \Level1Out9[19] , \Level1Out9[18] , \Level1Out9[17] , \Level1Out9[16] , 
        \Level1Out9[15] , \Level1Out9[14] , \Level1Out9[13] , \Level1Out9[12] , 
        \Level1Out9[11] , \Level1Out9[10] , \Level1Out9[9] , \Level1Out9[8] , 
        \Level1Out9[7] , \Level1Out9[6] , \Level1Out9[5] , \Level1Out9[4] , 
        \Level1Out9[3] , \Level1Out9[2] , \Level1Out9[1] , \Level1Out9[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_15 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink15[31] , \ScanLink15[30] , 
        \ScanLink15[29] , \ScanLink15[28] , \ScanLink15[27] , \ScanLink15[26] , 
        \ScanLink15[25] , \ScanLink15[24] , \ScanLink15[23] , \ScanLink15[22] , 
        \ScanLink15[21] , \ScanLink15[20] , \ScanLink15[19] , \ScanLink15[18] , 
        \ScanLink15[17] , \ScanLink15[16] , \ScanLink15[15] , \ScanLink15[14] , 
        \ScanLink15[13] , \ScanLink15[12] , \ScanLink15[11] , \ScanLink15[10] , 
        \ScanLink15[9] , \ScanLink15[8] , \ScanLink15[7] , \ScanLink15[6] , 
        \ScanLink15[5] , \ScanLink15[4] , \ScanLink15[3] , \ScanLink15[2] , 
        \ScanLink15[1] , \ScanLink15[0] }), .ScanOut({\ScanLink16[31] , 
        \ScanLink16[30] , \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , 
        \ScanLink16[26] , \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , 
        \ScanLink16[22] , \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , 
        \ScanLink16[18] , \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , 
        \ScanLink16[14] , \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , 
        \ScanLink16[10] , \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , 
        \ScanLink16[6] , \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , 
        \ScanLink16[2] , \ScanLink16[1] , \ScanLink16[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load15[0] ), .Out({
        \Level1Out15[31] , \Level1Out15[30] , \Level1Out15[29] , 
        \Level1Out15[28] , \Level1Out15[27] , \Level1Out15[26] , 
        \Level1Out15[25] , \Level1Out15[24] , \Level1Out15[23] , 
        \Level1Out15[22] , \Level1Out15[21] , \Level1Out15[20] , 
        \Level1Out15[19] , \Level1Out15[18] , \Level1Out15[17] , 
        \Level1Out15[16] , \Level1Out15[15] , \Level1Out15[14] , 
        \Level1Out15[13] , \Level1Out15[12] , \Level1Out15[11] , 
        \Level1Out15[10] , \Level1Out15[9] , \Level1Out15[8] , 
        \Level1Out15[7] , \Level1Out15[6] , \Level1Out15[5] , \Level1Out15[4] , 
        \Level1Out15[3] , \Level1Out15[2] , \Level1Out15[1] , \Level1Out15[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_20 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink20[31] , \ScanLink20[30] , 
        \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , \ScanLink20[26] , 
        \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , \ScanLink20[22] , 
        \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , \ScanLink20[18] , 
        \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , \ScanLink20[14] , 
        \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , \ScanLink20[10] , 
        \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , \ScanLink20[6] , 
        \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , \ScanLink20[2] , 
        \ScanLink20[1] , \ScanLink20[0] }), .ScanOut({\ScanLink21[31] , 
        \ScanLink21[30] , \ScanLink21[29] , \ScanLink21[28] , \ScanLink21[27] , 
        \ScanLink21[26] , \ScanLink21[25] , \ScanLink21[24] , \ScanLink21[23] , 
        \ScanLink21[22] , \ScanLink21[21] , \ScanLink21[20] , \ScanLink21[19] , 
        \ScanLink21[18] , \ScanLink21[17] , \ScanLink21[16] , \ScanLink21[15] , 
        \ScanLink21[14] , \ScanLink21[13] , \ScanLink21[12] , \ScanLink21[11] , 
        \ScanLink21[10] , \ScanLink21[9] , \ScanLink21[8] , \ScanLink21[7] , 
        \ScanLink21[6] , \ScanLink21[5] , \ScanLink21[4] , \ScanLink21[3] , 
        \ScanLink21[2] , \ScanLink21[1] , \ScanLink21[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load20[0] ), .Out({
        \Level1Out20[31] , \Level1Out20[30] , \Level1Out20[29] , 
        \Level1Out20[28] , \Level1Out20[27] , \Level1Out20[26] , 
        \Level1Out20[25] , \Level1Out20[24] , \Level1Out20[23] , 
        \Level1Out20[22] , \Level1Out20[21] , \Level1Out20[20] , 
        \Level1Out20[19] , \Level1Out20[18] , \Level1Out20[17] , 
        \Level1Out20[16] , \Level1Out20[15] , \Level1Out20[14] , 
        \Level1Out20[13] , \Level1Out20[12] , \Level1Out20[11] , 
        \Level1Out20[10] , \Level1Out20[9] , \Level1Out20[8] , 
        \Level1Out20[7] , \Level1Out20[6] , \Level1Out20[5] , \Level1Out20[4] , 
        \Level1Out20[3] , \Level1Out20[2] , \Level1Out20[1] , \Level1Out20[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_14_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load14[0] ), .Out({\Level2Out14[31] , \Level2Out14[30] , 
        \Level2Out14[29] , \Level2Out14[28] , \Level2Out14[27] , 
        \Level2Out14[26] , \Level2Out14[25] , \Level2Out14[24] , 
        \Level2Out14[23] , \Level2Out14[22] , \Level2Out14[21] , 
        \Level2Out14[20] , \Level2Out14[19] , \Level2Out14[18] , 
        \Level2Out14[17] , \Level2Out14[16] , \Level2Out14[15] , 
        \Level2Out14[14] , \Level2Out14[13] , \Level2Out14[12] , 
        \Level2Out14[11] , \Level2Out14[10] , \Level2Out14[9] , 
        \Level2Out14[8] , \Level2Out14[7] , \Level2Out14[6] , \Level2Out14[5] , 
        \Level2Out14[4] , \Level2Out14[3] , \Level2Out14[2] , \Level2Out14[1] , 
        \Level2Out14[0] }), .In1({\Level1Out14[31] , \Level1Out14[30] , 
        \Level1Out14[29] , \Level1Out14[28] , \Level1Out14[27] , 
        \Level1Out14[26] , \Level1Out14[25] , \Level1Out14[24] , 
        \Level1Out14[23] , \Level1Out14[22] , \Level1Out14[21] , 
        \Level1Out14[20] , \Level1Out14[19] , \Level1Out14[18] , 
        \Level1Out14[17] , \Level1Out14[16] , \Level1Out14[15] , 
        \Level1Out14[14] , \Level1Out14[13] , \Level1Out14[12] , 
        \Level1Out14[11] , \Level1Out14[10] , \Level1Out14[9] , 
        \Level1Out14[8] , \Level1Out14[7] , \Level1Out14[6] , \Level1Out14[5] , 
        \Level1Out14[4] , \Level1Out14[3] , \Level1Out14[2] , \Level1Out14[1] , 
        \Level1Out14[0] }), .In2({\Level1Out15[31] , \Level1Out15[30] , 
        \Level1Out15[29] , \Level1Out15[28] , \Level1Out15[27] , 
        \Level1Out15[26] , \Level1Out15[25] , \Level1Out15[24] , 
        \Level1Out15[23] , \Level1Out15[22] , \Level1Out15[21] , 
        \Level1Out15[20] , \Level1Out15[19] , \Level1Out15[18] , 
        \Level1Out15[17] , \Level1Out15[16] , \Level1Out15[15] , 
        \Level1Out15[14] , \Level1Out15[13] , \Level1Out15[12] , 
        \Level1Out15[11] , \Level1Out15[10] , \Level1Out15[9] , 
        \Level1Out15[8] , \Level1Out15[7] , \Level1Out15[6] , \Level1Out15[5] , 
        \Level1Out15[4] , \Level1Out15[3] , \Level1Out15[2] , \Level1Out15[1] , 
        \Level1Out15[0] }), .Read1(\Level1Load14[0] ), .Read2(
        \Level1Load15[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_32 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink32[31] , \ScanLink32[30] , 
        \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , \ScanLink32[26] , 
        \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , \ScanLink32[22] , 
        \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , \ScanLink32[18] , 
        \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , \ScanLink32[14] , 
        \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , \ScanLink32[10] , 
        \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , \ScanLink32[6] , 
        \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , \ScanLink32[2] , 
        \ScanLink32[1] , \ScanLink32[0] }), .ScanOut({\ScanLink33[31] , 
        \ScanLink33[30] , \ScanLink33[29] , \ScanLink33[28] , \ScanLink33[27] , 
        \ScanLink33[26] , \ScanLink33[25] , \ScanLink33[24] , \ScanLink33[23] , 
        \ScanLink33[22] , \ScanLink33[21] , \ScanLink33[20] , \ScanLink33[19] , 
        \ScanLink33[18] , \ScanLink33[17] , \ScanLink33[16] , \ScanLink33[15] , 
        \ScanLink33[14] , \ScanLink33[13] , \ScanLink33[12] , \ScanLink33[11] , 
        \ScanLink33[10] , \ScanLink33[9] , \ScanLink33[8] , \ScanLink33[7] , 
        \ScanLink33[6] , \ScanLink33[5] , \ScanLink33[4] , \ScanLink33[3] , 
        \ScanLink33[2] , \ScanLink33[1] , \ScanLink33[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load32[0] ), .Out({
        \Level1Out32[31] , \Level1Out32[30] , \Level1Out32[29] , 
        \Level1Out32[28] , \Level1Out32[27] , \Level1Out32[26] , 
        \Level1Out32[25] , \Level1Out32[24] , \Level1Out32[23] , 
        \Level1Out32[22] , \Level1Out32[21] , \Level1Out32[20] , 
        \Level1Out32[19] , \Level1Out32[18] , \Level1Out32[17] , 
        \Level1Out32[16] , \Level1Out32[15] , \Level1Out32[14] , 
        \Level1Out32[13] , \Level1Out32[12] , \Level1Out32[11] , 
        \Level1Out32[10] , \Level1Out32[9] , \Level1Out32[8] , 
        \Level1Out32[7] , \Level1Out32[6] , \Level1Out32[5] , \Level1Out32[4] , 
        \Level1Out32[3] , \Level1Out32[2] , \Level1Out32[1] , \Level1Out32[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_47 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink47[31] , \ScanLink47[30] , 
        \ScanLink47[29] , \ScanLink47[28] , \ScanLink47[27] , \ScanLink47[26] , 
        \ScanLink47[25] , \ScanLink47[24] , \ScanLink47[23] , \ScanLink47[22] , 
        \ScanLink47[21] , \ScanLink47[20] , \ScanLink47[19] , \ScanLink47[18] , 
        \ScanLink47[17] , \ScanLink47[16] , \ScanLink47[15] , \ScanLink47[14] , 
        \ScanLink47[13] , \ScanLink47[12] , \ScanLink47[11] , \ScanLink47[10] , 
        \ScanLink47[9] , \ScanLink47[8] , \ScanLink47[7] , \ScanLink47[6] , 
        \ScanLink47[5] , \ScanLink47[4] , \ScanLink47[3] , \ScanLink47[2] , 
        \ScanLink47[1] , \ScanLink47[0] }), .ScanOut({\ScanLink48[31] , 
        \ScanLink48[30] , \ScanLink48[29] , \ScanLink48[28] , \ScanLink48[27] , 
        \ScanLink48[26] , \ScanLink48[25] , \ScanLink48[24] , \ScanLink48[23] , 
        \ScanLink48[22] , \ScanLink48[21] , \ScanLink48[20] , \ScanLink48[19] , 
        \ScanLink48[18] , \ScanLink48[17] , \ScanLink48[16] , \ScanLink48[15] , 
        \ScanLink48[14] , \ScanLink48[13] , \ScanLink48[12] , \ScanLink48[11] , 
        \ScanLink48[10] , \ScanLink48[9] , \ScanLink48[8] , \ScanLink48[7] , 
        \ScanLink48[6] , \ScanLink48[5] , \ScanLink48[4] , \ScanLink48[3] , 
        \ScanLink48[2] , \ScanLink48[1] , \ScanLink48[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load47[0] ), .Out({
        \Level1Out47[31] , \Level1Out47[30] , \Level1Out47[29] , 
        \Level1Out47[28] , \Level1Out47[27] , \Level1Out47[26] , 
        \Level1Out47[25] , \Level1Out47[24] , \Level1Out47[23] , 
        \Level1Out47[22] , \Level1Out47[21] , \Level1Out47[20] , 
        \Level1Out47[19] , \Level1Out47[18] , \Level1Out47[17] , 
        \Level1Out47[16] , \Level1Out47[15] , \Level1Out47[14] , 
        \Level1Out47[13] , \Level1Out47[12] , \Level1Out47[11] , 
        \Level1Out47[10] , \Level1Out47[9] , \Level1Out47[8] , 
        \Level1Out47[7] , \Level1Out47[6] , \Level1Out47[5] , \Level1Out47[4] , 
        \Level1Out47[3] , \Level1Out47[2] , \Level1Out47[1] , \Level1Out47[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_60 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink60[31] , \ScanLink60[30] , 
        \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , \ScanLink60[26] , 
        \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , \ScanLink60[22] , 
        \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , \ScanLink60[18] , 
        \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , \ScanLink60[14] , 
        \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , \ScanLink60[10] , 
        \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , \ScanLink60[6] , 
        \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , \ScanLink60[2] , 
        \ScanLink60[1] , \ScanLink60[0] }), .ScanOut({\ScanLink61[31] , 
        \ScanLink61[30] , \ScanLink61[29] , \ScanLink61[28] , \ScanLink61[27] , 
        \ScanLink61[26] , \ScanLink61[25] , \ScanLink61[24] , \ScanLink61[23] , 
        \ScanLink61[22] , \ScanLink61[21] , \ScanLink61[20] , \ScanLink61[19] , 
        \ScanLink61[18] , \ScanLink61[17] , \ScanLink61[16] , \ScanLink61[15] , 
        \ScanLink61[14] , \ScanLink61[13] , \ScanLink61[12] , \ScanLink61[11] , 
        \ScanLink61[10] , \ScanLink61[9] , \ScanLink61[8] , \ScanLink61[7] , 
        \ScanLink61[6] , \ScanLink61[5] , \ScanLink61[4] , \ScanLink61[3] , 
        \ScanLink61[2] , \ScanLink61[1] , \ScanLink61[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load60[0] ), .Out({
        \Level1Out60[31] , \Level1Out60[30] , \Level1Out60[29] , 
        \Level1Out60[28] , \Level1Out60[27] , \Level1Out60[26] , 
        \Level1Out60[25] , \Level1Out60[24] , \Level1Out60[23] , 
        \Level1Out60[22] , \Level1Out60[21] , \Level1Out60[20] , 
        \Level1Out60[19] , \Level1Out60[18] , \Level1Out60[17] , 
        \Level1Out60[16] , \Level1Out60[15] , \Level1Out60[14] , 
        \Level1Out60[13] , \Level1Out60[12] , \Level1Out60[11] , 
        \Level1Out60[10] , \Level1Out60[9] , \Level1Out60[8] , 
        \Level1Out60[7] , \Level1Out60[6] , \Level1Out60[5] , \Level1Out60[4] , 
        \Level1Out60[3] , \Level1Out60[2] , \Level1Out60[1] , \Level1Out60[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_44_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load44[0] ), .Out({\Level2Out44[31] , \Level2Out44[30] , 
        \Level2Out44[29] , \Level2Out44[28] , \Level2Out44[27] , 
        \Level2Out44[26] , \Level2Out44[25] , \Level2Out44[24] , 
        \Level2Out44[23] , \Level2Out44[22] , \Level2Out44[21] , 
        \Level2Out44[20] , \Level2Out44[19] , \Level2Out44[18] , 
        \Level2Out44[17] , \Level2Out44[16] , \Level2Out44[15] , 
        \Level2Out44[14] , \Level2Out44[13] , \Level2Out44[12] , 
        \Level2Out44[11] , \Level2Out44[10] , \Level2Out44[9] , 
        \Level2Out44[8] , \Level2Out44[7] , \Level2Out44[6] , \Level2Out44[5] , 
        \Level2Out44[4] , \Level2Out44[3] , \Level2Out44[2] , \Level2Out44[1] , 
        \Level2Out44[0] }), .In1({\Level1Out44[31] , \Level1Out44[30] , 
        \Level1Out44[29] , \Level1Out44[28] , \Level1Out44[27] , 
        \Level1Out44[26] , \Level1Out44[25] , \Level1Out44[24] , 
        \Level1Out44[23] , \Level1Out44[22] , \Level1Out44[21] , 
        \Level1Out44[20] , \Level1Out44[19] , \Level1Out44[18] , 
        \Level1Out44[17] , \Level1Out44[16] , \Level1Out44[15] , 
        \Level1Out44[14] , \Level1Out44[13] , \Level1Out44[12] , 
        \Level1Out44[11] , \Level1Out44[10] , \Level1Out44[9] , 
        \Level1Out44[8] , \Level1Out44[7] , \Level1Out44[6] , \Level1Out44[5] , 
        \Level1Out44[4] , \Level1Out44[3] , \Level1Out44[2] , \Level1Out44[1] , 
        \Level1Out44[0] }), .In2({\Level1Out45[31] , \Level1Out45[30] , 
        \Level1Out45[29] , \Level1Out45[28] , \Level1Out45[27] , 
        \Level1Out45[26] , \Level1Out45[25] , \Level1Out45[24] , 
        \Level1Out45[23] , \Level1Out45[22] , \Level1Out45[21] , 
        \Level1Out45[20] , \Level1Out45[19] , \Level1Out45[18] , 
        \Level1Out45[17] , \Level1Out45[16] , \Level1Out45[15] , 
        \Level1Out45[14] , \Level1Out45[13] , \Level1Out45[12] , 
        \Level1Out45[11] , \Level1Out45[10] , \Level1Out45[9] , 
        \Level1Out45[8] , \Level1Out45[7] , \Level1Out45[6] , \Level1Out45[5] , 
        \Level1Out45[4] , \Level1Out45[3] , \Level1Out45[2] , \Level1Out45[1] , 
        \Level1Out45[0] }), .Read1(\Level1Load44[0] ), .Read2(
        \Level1Load45[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load0[0] ), .Out({\Level4Out0[31] , \Level4Out0[30] , 
        \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , \Level4Out0[26] , 
        \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , \Level4Out0[22] , 
        \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , \Level4Out0[18] , 
        \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , \Level4Out0[14] , 
        \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , \Level4Out0[10] , 
        \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , \Level4Out0[6] , 
        \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , \Level4Out0[2] , 
        \Level4Out0[1] , \Level4Out0[0] }), .In1({\Level2Out0[31] , 
        \Level2Out0[30] , \Level2Out0[29] , \Level2Out0[28] , \Level2Out0[27] , 
        \Level2Out0[26] , \Level2Out0[25] , \Level2Out0[24] , \Level2Out0[23] , 
        \Level2Out0[22] , \Level2Out0[21] , \Level2Out0[20] , \Level2Out0[19] , 
        \Level2Out0[18] , \Level2Out0[17] , \Level2Out0[16] , \Level2Out0[15] , 
        \Level2Out0[14] , \Level2Out0[13] , \Level2Out0[12] , \Level2Out0[11] , 
        \Level2Out0[10] , \Level2Out0[9] , \Level2Out0[8] , \Level2Out0[7] , 
        \Level2Out0[6] , \Level2Out0[5] , \Level2Out0[4] , \Level2Out0[3] , 
        \Level2Out0[2] , \Level2Out0[1] , \Level2Out0[0] }), .In2({
        \Level2Out2[31] , \Level2Out2[30] , \Level2Out2[29] , \Level2Out2[28] , 
        \Level2Out2[27] , \Level2Out2[26] , \Level2Out2[25] , \Level2Out2[24] , 
        \Level2Out2[23] , \Level2Out2[22] , \Level2Out2[21] , \Level2Out2[20] , 
        \Level2Out2[19] , \Level2Out2[18] , \Level2Out2[17] , \Level2Out2[16] , 
        \Level2Out2[15] , \Level2Out2[14] , \Level2Out2[13] , \Level2Out2[12] , 
        \Level2Out2[11] , \Level2Out2[10] , \Level2Out2[9] , \Level2Out2[8] , 
        \Level2Out2[7] , \Level2Out2[6] , \Level2Out2[5] , \Level2Out2[4] , 
        \Level2Out2[3] , \Level2Out2[2] , \Level2Out2[1] , \Level2Out2[0] }), 
        .Read1(\Level2Load0[0] ), .Read2(\Level2Load2[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load40[0] ), .Out({\Level4Out40[31] , \Level4Out40[30] , 
        \Level4Out40[29] , \Level4Out40[28] , \Level4Out40[27] , 
        \Level4Out40[26] , \Level4Out40[25] , \Level4Out40[24] , 
        \Level4Out40[23] , \Level4Out40[22] , \Level4Out40[21] , 
        \Level4Out40[20] , \Level4Out40[19] , \Level4Out40[18] , 
        \Level4Out40[17] , \Level4Out40[16] , \Level4Out40[15] , 
        \Level4Out40[14] , \Level4Out40[13] , \Level4Out40[12] , 
        \Level4Out40[11] , \Level4Out40[10] , \Level4Out40[9] , 
        \Level4Out40[8] , \Level4Out40[7] , \Level4Out40[6] , \Level4Out40[5] , 
        \Level4Out40[4] , \Level4Out40[3] , \Level4Out40[2] , \Level4Out40[1] , 
        \Level4Out40[0] }), .In1({\Level2Out40[31] , \Level2Out40[30] , 
        \Level2Out40[29] , \Level2Out40[28] , \Level2Out40[27] , 
        \Level2Out40[26] , \Level2Out40[25] , \Level2Out40[24] , 
        \Level2Out40[23] , \Level2Out40[22] , \Level2Out40[21] , 
        \Level2Out40[20] , \Level2Out40[19] , \Level2Out40[18] , 
        \Level2Out40[17] , \Level2Out40[16] , \Level2Out40[15] , 
        \Level2Out40[14] , \Level2Out40[13] , \Level2Out40[12] , 
        \Level2Out40[11] , \Level2Out40[10] , \Level2Out40[9] , 
        \Level2Out40[8] , \Level2Out40[7] , \Level2Out40[6] , \Level2Out40[5] , 
        \Level2Out40[4] , \Level2Out40[3] , \Level2Out40[2] , \Level2Out40[1] , 
        \Level2Out40[0] }), .In2({\Level2Out42[31] , \Level2Out42[30] , 
        \Level2Out42[29] , \Level2Out42[28] , \Level2Out42[27] , 
        \Level2Out42[26] , \Level2Out42[25] , \Level2Out42[24] , 
        \Level2Out42[23] , \Level2Out42[22] , \Level2Out42[21] , 
        \Level2Out42[20] , \Level2Out42[19] , \Level2Out42[18] , 
        \Level2Out42[17] , \Level2Out42[16] , \Level2Out42[15] , 
        \Level2Out42[14] , \Level2Out42[13] , \Level2Out42[12] , 
        \Level2Out42[11] , \Level2Out42[10] , \Level2Out42[9] , 
        \Level2Out42[8] , \Level2Out42[7] , \Level2Out42[6] , \Level2Out42[5] , 
        \Level2Out42[4] , \Level2Out42[3] , \Level2Out42[2] , \Level2Out42[1] , 
        \Level2Out42[0] }), .Read1(\Level2Load40[0] ), .Read2(
        \Level2Load42[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_2 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink2[31] , \ScanLink2[30] , 
        \ScanLink2[29] , \ScanLink2[28] , \ScanLink2[27] , \ScanLink2[26] , 
        \ScanLink2[25] , \ScanLink2[24] , \ScanLink2[23] , \ScanLink2[22] , 
        \ScanLink2[21] , \ScanLink2[20] , \ScanLink2[19] , \ScanLink2[18] , 
        \ScanLink2[17] , \ScanLink2[16] , \ScanLink2[15] , \ScanLink2[14] , 
        \ScanLink2[13] , \ScanLink2[12] , \ScanLink2[11] , \ScanLink2[10] , 
        \ScanLink2[9] , \ScanLink2[8] , \ScanLink2[7] , \ScanLink2[6] , 
        \ScanLink2[5] , \ScanLink2[4] , \ScanLink2[3] , \ScanLink2[2] , 
        \ScanLink2[1] , \ScanLink2[0] }), .ScanOut({\ScanLink3[31] , 
        \ScanLink3[30] , \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , 
        \ScanLink3[26] , \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , 
        \ScanLink3[22] , \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , 
        \ScanLink3[18] , \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , 
        \ScanLink3[14] , \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , 
        \ScanLink3[10] , \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , 
        \ScanLink3[6] , \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , 
        \ScanLink3[2] , \ScanLink3[1] , \ScanLink3[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load2[0] ), .Out({
        \Level1Out2[31] , \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , 
        \Level1Out2[27] , \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , 
        \Level1Out2[23] , \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , 
        \Level1Out2[19] , \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , 
        \Level1Out2[15] , \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , 
        \Level1Out2[11] , \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , 
        \Level1Out2[7] , \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , 
        \Level1Out2[3] , \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_22 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink22[31] , \ScanLink22[30] , 
        \ScanLink22[29] , \ScanLink22[28] , \ScanLink22[27] , \ScanLink22[26] , 
        \ScanLink22[25] , \ScanLink22[24] , \ScanLink22[23] , \ScanLink22[22] , 
        \ScanLink22[21] , \ScanLink22[20] , \ScanLink22[19] , \ScanLink22[18] , 
        \ScanLink22[17] , \ScanLink22[16] , \ScanLink22[15] , \ScanLink22[14] , 
        \ScanLink22[13] , \ScanLink22[12] , \ScanLink22[11] , \ScanLink22[10] , 
        \ScanLink22[9] , \ScanLink22[8] , \ScanLink22[7] , \ScanLink22[6] , 
        \ScanLink22[5] , \ScanLink22[4] , \ScanLink22[3] , \ScanLink22[2] , 
        \ScanLink22[1] , \ScanLink22[0] }), .ScanOut({\ScanLink23[31] , 
        \ScanLink23[30] , \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , 
        \ScanLink23[26] , \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , 
        \ScanLink23[22] , \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , 
        \ScanLink23[18] , \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , 
        \ScanLink23[14] , \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , 
        \ScanLink23[10] , \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , 
        \ScanLink23[6] , \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , 
        \ScanLink23[2] , \ScanLink23[1] , \ScanLink23[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load22[0] ), .Out({
        \Level1Out22[31] , \Level1Out22[30] , \Level1Out22[29] , 
        \Level1Out22[28] , \Level1Out22[27] , \Level1Out22[26] , 
        \Level1Out22[25] , \Level1Out22[24] , \Level1Out22[23] , 
        \Level1Out22[22] , \Level1Out22[21] , \Level1Out22[20] , 
        \Level1Out22[19] , \Level1Out22[18] , \Level1Out22[17] , 
        \Level1Out22[16] , \Level1Out22[15] , \Level1Out22[14] , 
        \Level1Out22[13] , \Level1Out22[12] , \Level1Out22[11] , 
        \Level1Out22[10] , \Level1Out22[9] , \Level1Out22[8] , 
        \Level1Out22[7] , \Level1Out22[6] , \Level1Out22[5] , \Level1Out22[4] , 
        \Level1Out22[3] , \Level1Out22[2] , \Level1Out22[1] , \Level1Out22[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_29 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink29[31] , \ScanLink29[30] , 
        \ScanLink29[29] , \ScanLink29[28] , \ScanLink29[27] , \ScanLink29[26] , 
        \ScanLink29[25] , \ScanLink29[24] , \ScanLink29[23] , \ScanLink29[22] , 
        \ScanLink29[21] , \ScanLink29[20] , \ScanLink29[19] , \ScanLink29[18] , 
        \ScanLink29[17] , \ScanLink29[16] , \ScanLink29[15] , \ScanLink29[14] , 
        \ScanLink29[13] , \ScanLink29[12] , \ScanLink29[11] , \ScanLink29[10] , 
        \ScanLink29[9] , \ScanLink29[8] , \ScanLink29[7] , \ScanLink29[6] , 
        \ScanLink29[5] , \ScanLink29[4] , \ScanLink29[3] , \ScanLink29[2] , 
        \ScanLink29[1] , \ScanLink29[0] }), .ScanOut({\ScanLink30[31] , 
        \ScanLink30[30] , \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , 
        \ScanLink30[26] , \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , 
        \ScanLink30[22] , \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , 
        \ScanLink30[18] , \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , 
        \ScanLink30[14] , \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , 
        \ScanLink30[10] , \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , 
        \ScanLink30[6] , \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , 
        \ScanLink30[2] , \ScanLink30[1] , \ScanLink30[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load29[0] ), .Out({
        \Level1Out29[31] , \Level1Out29[30] , \Level1Out29[29] , 
        \Level1Out29[28] , \Level1Out29[27] , \Level1Out29[26] , 
        \Level1Out29[25] , \Level1Out29[24] , \Level1Out29[23] , 
        \Level1Out29[22] , \Level1Out29[21] , \Level1Out29[20] , 
        \Level1Out29[19] , \Level1Out29[18] , \Level1Out29[17] , 
        \Level1Out29[16] , \Level1Out29[15] , \Level1Out29[14] , 
        \Level1Out29[13] , \Level1Out29[12] , \Level1Out29[11] , 
        \Level1Out29[10] , \Level1Out29[9] , \Level1Out29[8] , 
        \Level1Out29[7] , \Level1Out29[6] , \Level1Out29[5] , \Level1Out29[4] , 
        \Level1Out29[3] , \Level1Out29[2] , \Level1Out29[1] , \Level1Out29[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load4[0] ), .Out({\Level2Out4[31] , \Level2Out4[30] , 
        \Level2Out4[29] , \Level2Out4[28] , \Level2Out4[27] , \Level2Out4[26] , 
        \Level2Out4[25] , \Level2Out4[24] , \Level2Out4[23] , \Level2Out4[22] , 
        \Level2Out4[21] , \Level2Out4[20] , \Level2Out4[19] , \Level2Out4[18] , 
        \Level2Out4[17] , \Level2Out4[16] , \Level2Out4[15] , \Level2Out4[14] , 
        \Level2Out4[13] , \Level2Out4[12] , \Level2Out4[11] , \Level2Out4[10] , 
        \Level2Out4[9] , \Level2Out4[8] , \Level2Out4[7] , \Level2Out4[6] , 
        \Level2Out4[5] , \Level2Out4[4] , \Level2Out4[3] , \Level2Out4[2] , 
        \Level2Out4[1] , \Level2Out4[0] }), .In1({\Level1Out4[31] , 
        \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , \Level1Out4[27] , 
        \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , \Level1Out4[23] , 
        \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , \Level1Out4[19] , 
        \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , \Level1Out4[15] , 
        \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , \Level1Out4[11] , 
        \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , \Level1Out4[7] , 
        \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , \Level1Out4[3] , 
        \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] }), .In2({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] }), 
        .Read1(\Level1Load4[0] ), .Read2(\Level1Load5[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_60_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load60[0] ), .Out({\Level2Out60[31] , \Level2Out60[30] , 
        \Level2Out60[29] , \Level2Out60[28] , \Level2Out60[27] , 
        \Level2Out60[26] , \Level2Out60[25] , \Level2Out60[24] , 
        \Level2Out60[23] , \Level2Out60[22] , \Level2Out60[21] , 
        \Level2Out60[20] , \Level2Out60[19] , \Level2Out60[18] , 
        \Level2Out60[17] , \Level2Out60[16] , \Level2Out60[15] , 
        \Level2Out60[14] , \Level2Out60[13] , \Level2Out60[12] , 
        \Level2Out60[11] , \Level2Out60[10] , \Level2Out60[9] , 
        \Level2Out60[8] , \Level2Out60[7] , \Level2Out60[6] , \Level2Out60[5] , 
        \Level2Out60[4] , \Level2Out60[3] , \Level2Out60[2] , \Level2Out60[1] , 
        \Level2Out60[0] }), .In1({\Level1Out60[31] , \Level1Out60[30] , 
        \Level1Out60[29] , \Level1Out60[28] , \Level1Out60[27] , 
        \Level1Out60[26] , \Level1Out60[25] , \Level1Out60[24] , 
        \Level1Out60[23] , \Level1Out60[22] , \Level1Out60[21] , 
        \Level1Out60[20] , \Level1Out60[19] , \Level1Out60[18] , 
        \Level1Out60[17] , \Level1Out60[16] , \Level1Out60[15] , 
        \Level1Out60[14] , \Level1Out60[13] , \Level1Out60[12] , 
        \Level1Out60[11] , \Level1Out60[10] , \Level1Out60[9] , 
        \Level1Out60[8] , \Level1Out60[7] , \Level1Out60[6] , \Level1Out60[5] , 
        \Level1Out60[4] , \Level1Out60[3] , \Level1Out60[2] , \Level1Out60[1] , 
        \Level1Out60[0] }), .In2({\Level1Out61[31] , \Level1Out61[30] , 
        \Level1Out61[29] , \Level1Out61[28] , \Level1Out61[27] , 
        \Level1Out61[26] , \Level1Out61[25] , \Level1Out61[24] , 
        \Level1Out61[23] , \Level1Out61[22] , \Level1Out61[21] , 
        \Level1Out61[20] , \Level1Out61[19] , \Level1Out61[18] , 
        \Level1Out61[17] , \Level1Out61[16] , \Level1Out61[15] , 
        \Level1Out61[14] , \Level1Out61[13] , \Level1Out61[12] , 
        \Level1Out61[11] , \Level1Out61[10] , \Level1Out61[9] , 
        \Level1Out61[8] , \Level1Out61[7] , \Level1Out61[6] , \Level1Out61[5] , 
        \Level1Out61[4] , \Level1Out61[3] , \Level1Out61[2] , \Level1Out61[1] , 
        \Level1Out61[0] }), .Read1(\Level1Load60[0] ), .Read2(
        \Level1Load61[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load56[0] ), .Out({\Level4Out56[31] , \Level4Out56[30] , 
        \Level4Out56[29] , \Level4Out56[28] , \Level4Out56[27] , 
        \Level4Out56[26] , \Level4Out56[25] , \Level4Out56[24] , 
        \Level4Out56[23] , \Level4Out56[22] , \Level4Out56[21] , 
        \Level4Out56[20] , \Level4Out56[19] , \Level4Out56[18] , 
        \Level4Out56[17] , \Level4Out56[16] , \Level4Out56[15] , 
        \Level4Out56[14] , \Level4Out56[13] , \Level4Out56[12] , 
        \Level4Out56[11] , \Level4Out56[10] , \Level4Out56[9] , 
        \Level4Out56[8] , \Level4Out56[7] , \Level4Out56[6] , \Level4Out56[5] , 
        \Level4Out56[4] , \Level4Out56[3] , \Level4Out56[2] , \Level4Out56[1] , 
        \Level4Out56[0] }), .In1({\Level2Out56[31] , \Level2Out56[30] , 
        \Level2Out56[29] , \Level2Out56[28] , \Level2Out56[27] , 
        \Level2Out56[26] , \Level2Out56[25] , \Level2Out56[24] , 
        \Level2Out56[23] , \Level2Out56[22] , \Level2Out56[21] , 
        \Level2Out56[20] , \Level2Out56[19] , \Level2Out56[18] , 
        \Level2Out56[17] , \Level2Out56[16] , \Level2Out56[15] , 
        \Level2Out56[14] , \Level2Out56[13] , \Level2Out56[12] , 
        \Level2Out56[11] , \Level2Out56[10] , \Level2Out56[9] , 
        \Level2Out56[8] , \Level2Out56[7] , \Level2Out56[6] , \Level2Out56[5] , 
        \Level2Out56[4] , \Level2Out56[3] , \Level2Out56[2] , \Level2Out56[1] , 
        \Level2Out56[0] }), .In2({\Level2Out58[31] , \Level2Out58[30] , 
        \Level2Out58[29] , \Level2Out58[28] , \Level2Out58[27] , 
        \Level2Out58[26] , \Level2Out58[25] , \Level2Out58[24] , 
        \Level2Out58[23] , \Level2Out58[22] , \Level2Out58[21] , 
        \Level2Out58[20] , \Level2Out58[19] , \Level2Out58[18] , 
        \Level2Out58[17] , \Level2Out58[16] , \Level2Out58[15] , 
        \Level2Out58[14] , \Level2Out58[13] , \Level2Out58[12] , 
        \Level2Out58[11] , \Level2Out58[10] , \Level2Out58[9] , 
        \Level2Out58[8] , \Level2Out58[7] , \Level2Out58[6] , \Level2Out58[5] , 
        \Level2Out58[4] , \Level2Out58[3] , \Level2Out58[2] , \Level2Out58[1] , 
        \Level2Out58[0] }), .Read1(\Level2Load56[0] ), .Read2(
        \Level2Load58[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_3 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink3[31] , \ScanLink3[30] , 
        \ScanLink3[29] , \ScanLink3[28] , \ScanLink3[27] , \ScanLink3[26] , 
        \ScanLink3[25] , \ScanLink3[24] , \ScanLink3[23] , \ScanLink3[22] , 
        \ScanLink3[21] , \ScanLink3[20] , \ScanLink3[19] , \ScanLink3[18] , 
        \ScanLink3[17] , \ScanLink3[16] , \ScanLink3[15] , \ScanLink3[14] , 
        \ScanLink3[13] , \ScanLink3[12] , \ScanLink3[11] , \ScanLink3[10] , 
        \ScanLink3[9] , \ScanLink3[8] , \ScanLink3[7] , \ScanLink3[6] , 
        \ScanLink3[5] , \ScanLink3[4] , \ScanLink3[3] , \ScanLink3[2] , 
        \ScanLink3[1] , \ScanLink3[0] }), .ScanOut({\ScanLink4[31] , 
        \ScanLink4[30] , \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , 
        \ScanLink4[26] , \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , 
        \ScanLink4[22] , \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , 
        \ScanLink4[18] , \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , 
        \ScanLink4[14] , \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , 
        \ScanLink4[10] , \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , 
        \ScanLink4[6] , \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , 
        \ScanLink4[2] , \ScanLink4[1] , \ScanLink4[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load3[0] ), .Out({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_4 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink4[31] , \ScanLink4[30] , 
        \ScanLink4[29] , \ScanLink4[28] , \ScanLink4[27] , \ScanLink4[26] , 
        \ScanLink4[25] , \ScanLink4[24] , \ScanLink4[23] , \ScanLink4[22] , 
        \ScanLink4[21] , \ScanLink4[20] , \ScanLink4[19] , \ScanLink4[18] , 
        \ScanLink4[17] , \ScanLink4[16] , \ScanLink4[15] , \ScanLink4[14] , 
        \ScanLink4[13] , \ScanLink4[12] , \ScanLink4[11] , \ScanLink4[10] , 
        \ScanLink4[9] , \ScanLink4[8] , \ScanLink4[7] , \ScanLink4[6] , 
        \ScanLink4[5] , \ScanLink4[4] , \ScanLink4[3] , \ScanLink4[2] , 
        \ScanLink4[1] , \ScanLink4[0] }), .ScanOut({\ScanLink5[31] , 
        \ScanLink5[30] , \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , 
        \ScanLink5[26] , \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , 
        \ScanLink5[22] , \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , 
        \ScanLink5[18] , \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , 
        \ScanLink5[14] , \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , 
        \ScanLink5[10] , \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , 
        \ScanLink5[6] , \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , 
        \ScanLink5[2] , \ScanLink5[1] , \ScanLink5[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load4[0] ), .Out({
        \Level1Out4[31] , \Level1Out4[30] , \Level1Out4[29] , \Level1Out4[28] , 
        \Level1Out4[27] , \Level1Out4[26] , \Level1Out4[25] , \Level1Out4[24] , 
        \Level1Out4[23] , \Level1Out4[22] , \Level1Out4[21] , \Level1Out4[20] , 
        \Level1Out4[19] , \Level1Out4[18] , \Level1Out4[17] , \Level1Out4[16] , 
        \Level1Out4[15] , \Level1Out4[14] , \Level1Out4[13] , \Level1Out4[12] , 
        \Level1Out4[11] , \Level1Out4[10] , \Level1Out4[9] , \Level1Out4[8] , 
        \Level1Out4[7] , \Level1Out4[6] , \Level1Out4[5] , \Level1Out4[4] , 
        \Level1Out4[3] , \Level1Out4[2] , \Level1Out4[1] , \Level1Out4[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_5 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink5[31] , \ScanLink5[30] , 
        \ScanLink5[29] , \ScanLink5[28] , \ScanLink5[27] , \ScanLink5[26] , 
        \ScanLink5[25] , \ScanLink5[24] , \ScanLink5[23] , \ScanLink5[22] , 
        \ScanLink5[21] , \ScanLink5[20] , \ScanLink5[19] , \ScanLink5[18] , 
        \ScanLink5[17] , \ScanLink5[16] , \ScanLink5[15] , \ScanLink5[14] , 
        \ScanLink5[13] , \ScanLink5[12] , \ScanLink5[11] , \ScanLink5[10] , 
        \ScanLink5[9] , \ScanLink5[8] , \ScanLink5[7] , \ScanLink5[6] , 
        \ScanLink5[5] , \ScanLink5[4] , \ScanLink5[3] , \ScanLink5[2] , 
        \ScanLink5[1] , \ScanLink5[0] }), .ScanOut({\ScanLink6[31] , 
        \ScanLink6[30] , \ScanLink6[29] , \ScanLink6[28] , \ScanLink6[27] , 
        \ScanLink6[26] , \ScanLink6[25] , \ScanLink6[24] , \ScanLink6[23] , 
        \ScanLink6[22] , \ScanLink6[21] , \ScanLink6[20] , \ScanLink6[19] , 
        \ScanLink6[18] , \ScanLink6[17] , \ScanLink6[16] , \ScanLink6[15] , 
        \ScanLink6[14] , \ScanLink6[13] , \ScanLink6[12] , \ScanLink6[11] , 
        \ScanLink6[10] , \ScanLink6[9] , \ScanLink6[8] , \ScanLink6[7] , 
        \ScanLink6[6] , \ScanLink6[5] , \ScanLink6[4] , \ScanLink6[3] , 
        \ScanLink6[2] , \ScanLink6[1] , \ScanLink6[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load5[0] ), .Out({
        \Level1Out5[31] , \Level1Out5[30] , \Level1Out5[29] , \Level1Out5[28] , 
        \Level1Out5[27] , \Level1Out5[26] , \Level1Out5[25] , \Level1Out5[24] , 
        \Level1Out5[23] , \Level1Out5[22] , \Level1Out5[21] , \Level1Out5[20] , 
        \Level1Out5[19] , \Level1Out5[18] , \Level1Out5[17] , \Level1Out5[16] , 
        \Level1Out5[15] , \Level1Out5[14] , \Level1Out5[13] , \Level1Out5[12] , 
        \Level1Out5[11] , \Level1Out5[10] , \Level1Out5[9] , \Level1Out5[8] , 
        \Level1Out5[7] , \Level1Out5[6] , \Level1Out5[5] , \Level1Out5[4] , 
        \Level1Out5[3] , \Level1Out5[2] , \Level1Out5[1] , \Level1Out5[0] })
         );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_10 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink10[31] , \ScanLink10[30] , 
        \ScanLink10[29] , \ScanLink10[28] , \ScanLink10[27] , \ScanLink10[26] , 
        \ScanLink10[25] , \ScanLink10[24] , \ScanLink10[23] , \ScanLink10[22] , 
        \ScanLink10[21] , \ScanLink10[20] , \ScanLink10[19] , \ScanLink10[18] , 
        \ScanLink10[17] , \ScanLink10[16] , \ScanLink10[15] , \ScanLink10[14] , 
        \ScanLink10[13] , \ScanLink10[12] , \ScanLink10[11] , \ScanLink10[10] , 
        \ScanLink10[9] , \ScanLink10[8] , \ScanLink10[7] , \ScanLink10[6] , 
        \ScanLink10[5] , \ScanLink10[4] , \ScanLink10[3] , \ScanLink10[2] , 
        \ScanLink10[1] , \ScanLink10[0] }), .ScanOut({\ScanLink11[31] , 
        \ScanLink11[30] , \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , 
        \ScanLink11[26] , \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , 
        \ScanLink11[22] , \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , 
        \ScanLink11[18] , \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , 
        \ScanLink11[14] , \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , 
        \ScanLink11[10] , \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , 
        \ScanLink11[6] , \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , 
        \ScanLink11[2] , \ScanLink11[1] , \ScanLink11[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load10[0] ), .Out({
        \Level1Out10[31] , \Level1Out10[30] , \Level1Out10[29] , 
        \Level1Out10[28] , \Level1Out10[27] , \Level1Out10[26] , 
        \Level1Out10[25] , \Level1Out10[24] , \Level1Out10[23] , 
        \Level1Out10[22] , \Level1Out10[21] , \Level1Out10[20] , 
        \Level1Out10[19] , \Level1Out10[18] , \Level1Out10[17] , 
        \Level1Out10[16] , \Level1Out10[15] , \Level1Out10[14] , 
        \Level1Out10[13] , \Level1Out10[12] , \Level1Out10[11] , 
        \Level1Out10[10] , \Level1Out10[9] , \Level1Out10[8] , 
        \Level1Out10[7] , \Level1Out10[6] , \Level1Out10[5] , \Level1Out10[4] , 
        \Level1Out10[3] , \Level1Out10[2] , \Level1Out10[1] , \Level1Out10[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_17 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink17[31] , \ScanLink17[30] , 
        \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , \ScanLink17[26] , 
        \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , \ScanLink17[22] , 
        \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , \ScanLink17[18] , 
        \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , \ScanLink17[14] , 
        \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , \ScanLink17[10] , 
        \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , \ScanLink17[6] , 
        \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , \ScanLink17[2] , 
        \ScanLink17[1] , \ScanLink17[0] }), .ScanOut({\ScanLink18[31] , 
        \ScanLink18[30] , \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , 
        \ScanLink18[26] , \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , 
        \ScanLink18[22] , \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , 
        \ScanLink18[18] , \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , 
        \ScanLink18[14] , \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , 
        \ScanLink18[10] , \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , 
        \ScanLink18[6] , \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , 
        \ScanLink18[2] , \ScanLink18[1] , \ScanLink18[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load17[0] ), .Out({
        \Level1Out17[31] , \Level1Out17[30] , \Level1Out17[29] , 
        \Level1Out17[28] , \Level1Out17[27] , \Level1Out17[26] , 
        \Level1Out17[25] , \Level1Out17[24] , \Level1Out17[23] , 
        \Level1Out17[22] , \Level1Out17[21] , \Level1Out17[20] , 
        \Level1Out17[19] , \Level1Out17[18] , \Level1Out17[17] , 
        \Level1Out17[16] , \Level1Out17[15] , \Level1Out17[14] , 
        \Level1Out17[13] , \Level1Out17[12] , \Level1Out17[11] , 
        \Level1Out17[10] , \Level1Out17[9] , \Level1Out17[8] , 
        \Level1Out17[7] , \Level1Out17[6] , \Level1Out17[5] , \Level1Out17[4] , 
        \Level1Out17[3] , \Level1Out17[2] , \Level1Out17[1] , \Level1Out17[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_30 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink30[31] , \ScanLink30[30] , 
        \ScanLink30[29] , \ScanLink30[28] , \ScanLink30[27] , \ScanLink30[26] , 
        \ScanLink30[25] , \ScanLink30[24] , \ScanLink30[23] , \ScanLink30[22] , 
        \ScanLink30[21] , \ScanLink30[20] , \ScanLink30[19] , \ScanLink30[18] , 
        \ScanLink30[17] , \ScanLink30[16] , \ScanLink30[15] , \ScanLink30[14] , 
        \ScanLink30[13] , \ScanLink30[12] , \ScanLink30[11] , \ScanLink30[10] , 
        \ScanLink30[9] , \ScanLink30[8] , \ScanLink30[7] , \ScanLink30[6] , 
        \ScanLink30[5] , \ScanLink30[4] , \ScanLink30[3] , \ScanLink30[2] , 
        \ScanLink30[1] , \ScanLink30[0] }), .ScanOut({\ScanLink31[31] , 
        \ScanLink31[30] , \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , 
        \ScanLink31[26] , \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , 
        \ScanLink31[22] , \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , 
        \ScanLink31[18] , \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , 
        \ScanLink31[14] , \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , 
        \ScanLink31[10] , \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , 
        \ScanLink31[6] , \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , 
        \ScanLink31[2] , \ScanLink31[1] , \ScanLink31[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load30[0] ), .Out({
        \Level1Out30[31] , \Level1Out30[30] , \Level1Out30[29] , 
        \Level1Out30[28] , \Level1Out30[27] , \Level1Out30[26] , 
        \Level1Out30[25] , \Level1Out30[24] , \Level1Out30[23] , 
        \Level1Out30[22] , \Level1Out30[21] , \Level1Out30[20] , 
        \Level1Out30[19] , \Level1Out30[18] , \Level1Out30[17] , 
        \Level1Out30[16] , \Level1Out30[15] , \Level1Out30[14] , 
        \Level1Out30[13] , \Level1Out30[12] , \Level1Out30[11] , 
        \Level1Out30[10] , \Level1Out30[9] , \Level1Out30[8] , 
        \Level1Out30[7] , \Level1Out30[6] , \Level1Out30[5] , \Level1Out30[4] , 
        \Level1Out30[3] , \Level1Out30[2] , \Level1Out30[1] , \Level1Out30[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_39 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink39[31] , \ScanLink39[30] , 
        \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , \ScanLink39[26] , 
        \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , \ScanLink39[22] , 
        \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , \ScanLink39[18] , 
        \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , \ScanLink39[14] , 
        \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , \ScanLink39[10] , 
        \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , \ScanLink39[6] , 
        \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , \ScanLink39[2] , 
        \ScanLink39[1] , \ScanLink39[0] }), .ScanOut({\ScanLink40[31] , 
        \ScanLink40[30] , \ScanLink40[29] , \ScanLink40[28] , \ScanLink40[27] , 
        \ScanLink40[26] , \ScanLink40[25] , \ScanLink40[24] , \ScanLink40[23] , 
        \ScanLink40[22] , \ScanLink40[21] , \ScanLink40[20] , \ScanLink40[19] , 
        \ScanLink40[18] , \ScanLink40[17] , \ScanLink40[16] , \ScanLink40[15] , 
        \ScanLink40[14] , \ScanLink40[13] , \ScanLink40[12] , \ScanLink40[11] , 
        \ScanLink40[10] , \ScanLink40[9] , \ScanLink40[8] , \ScanLink40[7] , 
        \ScanLink40[6] , \ScanLink40[5] , \ScanLink40[4] , \ScanLink40[3] , 
        \ScanLink40[2] , \ScanLink40[1] , \ScanLink40[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load39[0] ), .Out({
        \Level1Out39[31] , \Level1Out39[30] , \Level1Out39[29] , 
        \Level1Out39[28] , \Level1Out39[27] , \Level1Out39[26] , 
        \Level1Out39[25] , \Level1Out39[24] , \Level1Out39[23] , 
        \Level1Out39[22] , \Level1Out39[21] , \Level1Out39[20] , 
        \Level1Out39[19] , \Level1Out39[18] , \Level1Out39[17] , 
        \Level1Out39[16] , \Level1Out39[15] , \Level1Out39[14] , 
        \Level1Out39[13] , \Level1Out39[12] , \Level1Out39[11] , 
        \Level1Out39[10] , \Level1Out39[9] , \Level1Out39[8] , 
        \Level1Out39[7] , \Level1Out39[6] , \Level1Out39[5] , \Level1Out39[4] , 
        \Level1Out39[3] , \Level1Out39[2] , \Level1Out39[1] , \Level1Out39[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_57 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink57[31] , \ScanLink57[30] , 
        \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , \ScanLink57[26] , 
        \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , \ScanLink57[22] , 
        \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , \ScanLink57[18] , 
        \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , \ScanLink57[14] , 
        \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , \ScanLink57[10] , 
        \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , \ScanLink57[6] , 
        \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , \ScanLink57[2] , 
        \ScanLink57[1] , \ScanLink57[0] }), .ScanOut({\ScanLink58[31] , 
        \ScanLink58[30] , \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , 
        \ScanLink58[26] , \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , 
        \ScanLink58[22] , \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , 
        \ScanLink58[18] , \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , 
        \ScanLink58[14] , \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , 
        \ScanLink58[10] , \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , 
        \ScanLink58[6] , \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , 
        \ScanLink58[2] , \ScanLink58[1] , \ScanLink58[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load57[0] ), .Out({
        \Level1Out57[31] , \Level1Out57[30] , \Level1Out57[29] , 
        \Level1Out57[28] , \Level1Out57[27] , \Level1Out57[26] , 
        \Level1Out57[25] , \Level1Out57[24] , \Level1Out57[23] , 
        \Level1Out57[22] , \Level1Out57[21] , \Level1Out57[20] , 
        \Level1Out57[19] , \Level1Out57[18] , \Level1Out57[17] , 
        \Level1Out57[16] , \Level1Out57[15] , \Level1Out57[14] , 
        \Level1Out57[13] , \Level1Out57[12] , \Level1Out57[11] , 
        \Level1Out57[10] , \Level1Out57[9] , \Level1Out57[8] , 
        \Level1Out57[7] , \Level1Out57[6] , \Level1Out57[5] , \Level1Out57[4] , 
        \Level1Out57[3] , \Level1Out57[2] , \Level1Out57[1] , \Level1Out57[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_45 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink45[31] , \ScanLink45[30] , 
        \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , \ScanLink45[26] , 
        \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , \ScanLink45[22] , 
        \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , \ScanLink45[18] , 
        \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , \ScanLink45[14] , 
        \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , \ScanLink45[10] , 
        \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , \ScanLink45[6] , 
        \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , \ScanLink45[2] , 
        \ScanLink45[1] , \ScanLink45[0] }), .ScanOut({\ScanLink46[31] , 
        \ScanLink46[30] , \ScanLink46[29] , \ScanLink46[28] , \ScanLink46[27] , 
        \ScanLink46[26] , \ScanLink46[25] , \ScanLink46[24] , \ScanLink46[23] , 
        \ScanLink46[22] , \ScanLink46[21] , \ScanLink46[20] , \ScanLink46[19] , 
        \ScanLink46[18] , \ScanLink46[17] , \ScanLink46[16] , \ScanLink46[15] , 
        \ScanLink46[14] , \ScanLink46[13] , \ScanLink46[12] , \ScanLink46[11] , 
        \ScanLink46[10] , \ScanLink46[9] , \ScanLink46[8] , \ScanLink46[7] , 
        \ScanLink46[6] , \ScanLink46[5] , \ScanLink46[4] , \ScanLink46[3] , 
        \ScanLink46[2] , \ScanLink46[1] , \ScanLink46[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load45[0] ), .Out({
        \Level1Out45[31] , \Level1Out45[30] , \Level1Out45[29] , 
        \Level1Out45[28] , \Level1Out45[27] , \Level1Out45[26] , 
        \Level1Out45[25] , \Level1Out45[24] , \Level1Out45[23] , 
        \Level1Out45[22] , \Level1Out45[21] , \Level1Out45[20] , 
        \Level1Out45[19] , \Level1Out45[18] , \Level1Out45[17] , 
        \Level1Out45[16] , \Level1Out45[15] , \Level1Out45[14] , 
        \Level1Out45[13] , \Level1Out45[12] , \Level1Out45[11] , 
        \Level1Out45[10] , \Level1Out45[9] , \Level1Out45[8] , 
        \Level1Out45[7] , \Level1Out45[6] , \Level1Out45[5] , \Level1Out45[4] , 
        \Level1Out45[3] , \Level1Out45[2] , \Level1Out45[1] , \Level1Out45[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_28_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load28[0] ), .Out({\Level2Out28[31] , \Level2Out28[30] , 
        \Level2Out28[29] , \Level2Out28[28] , \Level2Out28[27] , 
        \Level2Out28[26] , \Level2Out28[25] , \Level2Out28[24] , 
        \Level2Out28[23] , \Level2Out28[22] , \Level2Out28[21] , 
        \Level2Out28[20] , \Level2Out28[19] , \Level2Out28[18] , 
        \Level2Out28[17] , \Level2Out28[16] , \Level2Out28[15] , 
        \Level2Out28[14] , \Level2Out28[13] , \Level2Out28[12] , 
        \Level2Out28[11] , \Level2Out28[10] , \Level2Out28[9] , 
        \Level2Out28[8] , \Level2Out28[7] , \Level2Out28[6] , \Level2Out28[5] , 
        \Level2Out28[4] , \Level2Out28[3] , \Level2Out28[2] , \Level2Out28[1] , 
        \Level2Out28[0] }), .In1({\Level1Out28[31] , \Level1Out28[30] , 
        \Level1Out28[29] , \Level1Out28[28] , \Level1Out28[27] , 
        \Level1Out28[26] , \Level1Out28[25] , \Level1Out28[24] , 
        \Level1Out28[23] , \Level1Out28[22] , \Level1Out28[21] , 
        \Level1Out28[20] , \Level1Out28[19] , \Level1Out28[18] , 
        \Level1Out28[17] , \Level1Out28[16] , \Level1Out28[15] , 
        \Level1Out28[14] , \Level1Out28[13] , \Level1Out28[12] , 
        \Level1Out28[11] , \Level1Out28[10] , \Level1Out28[9] , 
        \Level1Out28[8] , \Level1Out28[7] , \Level1Out28[6] , \Level1Out28[5] , 
        \Level1Out28[4] , \Level1Out28[3] , \Level1Out28[2] , \Level1Out28[1] , 
        \Level1Out28[0] }), .In2({\Level1Out29[31] , \Level1Out29[30] , 
        \Level1Out29[29] , \Level1Out29[28] , \Level1Out29[27] , 
        \Level1Out29[26] , \Level1Out29[25] , \Level1Out29[24] , 
        \Level1Out29[23] , \Level1Out29[22] , \Level1Out29[21] , 
        \Level1Out29[20] , \Level1Out29[19] , \Level1Out29[18] , 
        \Level1Out29[17] , \Level1Out29[16] , \Level1Out29[15] , 
        \Level1Out29[14] , \Level1Out29[13] , \Level1Out29[12] , 
        \Level1Out29[11] , \Level1Out29[10] , \Level1Out29[9] , 
        \Level1Out29[8] , \Level1Out29[7] , \Level1Out29[6] , \Level1Out29[5] , 
        \Level1Out29[4] , \Level1Out29[3] , \Level1Out29[2] , \Level1Out29[1] , 
        \Level1Out29[0] }), .Read1(\Level1Load28[0] ), .Read2(
        \Level1Load29[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_52_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load52[0] ), .Out({\Level2Out52[31] , \Level2Out52[30] , 
        \Level2Out52[29] , \Level2Out52[28] , \Level2Out52[27] , 
        \Level2Out52[26] , \Level2Out52[25] , \Level2Out52[24] , 
        \Level2Out52[23] , \Level2Out52[22] , \Level2Out52[21] , 
        \Level2Out52[20] , \Level2Out52[19] , \Level2Out52[18] , 
        \Level2Out52[17] , \Level2Out52[16] , \Level2Out52[15] , 
        \Level2Out52[14] , \Level2Out52[13] , \Level2Out52[12] , 
        \Level2Out52[11] , \Level2Out52[10] , \Level2Out52[9] , 
        \Level2Out52[8] , \Level2Out52[7] , \Level2Out52[6] , \Level2Out52[5] , 
        \Level2Out52[4] , \Level2Out52[3] , \Level2Out52[2] , \Level2Out52[1] , 
        \Level2Out52[0] }), .In1({\Level1Out52[31] , \Level1Out52[30] , 
        \Level1Out52[29] , \Level1Out52[28] , \Level1Out52[27] , 
        \Level1Out52[26] , \Level1Out52[25] , \Level1Out52[24] , 
        \Level1Out52[23] , \Level1Out52[22] , \Level1Out52[21] , 
        \Level1Out52[20] , \Level1Out52[19] , \Level1Out52[18] , 
        \Level1Out52[17] , \Level1Out52[16] , \Level1Out52[15] , 
        \Level1Out52[14] , \Level1Out52[13] , \Level1Out52[12] , 
        \Level1Out52[11] , \Level1Out52[10] , \Level1Out52[9] , 
        \Level1Out52[8] , \Level1Out52[7] , \Level1Out52[6] , \Level1Out52[5] , 
        \Level1Out52[4] , \Level1Out52[3] , \Level1Out52[2] , \Level1Out52[1] , 
        \Level1Out52[0] }), .In2({\Level1Out53[31] , \Level1Out53[30] , 
        \Level1Out53[29] , \Level1Out53[28] , \Level1Out53[27] , 
        \Level1Out53[26] , \Level1Out53[25] , \Level1Out53[24] , 
        \Level1Out53[23] , \Level1Out53[22] , \Level1Out53[21] , 
        \Level1Out53[20] , \Level1Out53[19] , \Level1Out53[18] , 
        \Level1Out53[17] , \Level1Out53[16] , \Level1Out53[15] , 
        \Level1Out53[14] , \Level1Out53[13] , \Level1Out53[12] , 
        \Level1Out53[11] , \Level1Out53[10] , \Level1Out53[9] , 
        \Level1Out53[8] , \Level1Out53[7] , \Level1Out53[6] , \Level1Out53[5] , 
        \Level1Out53[4] , \Level1Out53[3] , \Level1Out53[2] , \Level1Out53[1] , 
        \Level1Out53[0] }), .Read1(\Level1Load52[0] ), .Read2(
        \Level1Load53[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_62 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink62[31] , \ScanLink62[30] , 
        \ScanLink62[29] , \ScanLink62[28] , \ScanLink62[27] , \ScanLink62[26] , 
        \ScanLink62[25] , \ScanLink62[24] , \ScanLink62[23] , \ScanLink62[22] , 
        \ScanLink62[21] , \ScanLink62[20] , \ScanLink62[19] , \ScanLink62[18] , 
        \ScanLink62[17] , \ScanLink62[16] , \ScanLink62[15] , \ScanLink62[14] , 
        \ScanLink62[13] , \ScanLink62[12] , \ScanLink62[11] , \ScanLink62[10] , 
        \ScanLink62[9] , \ScanLink62[8] , \ScanLink62[7] , \ScanLink62[6] , 
        \ScanLink62[5] , \ScanLink62[4] , \ScanLink62[3] , \ScanLink62[2] , 
        \ScanLink62[1] , \ScanLink62[0] }), .ScanOut({\ScanLink63[31] , 
        \ScanLink63[30] , \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , 
        \ScanLink63[26] , \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , 
        \ScanLink63[22] , \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , 
        \ScanLink63[18] , \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , 
        \ScanLink63[14] , \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , 
        \ScanLink63[10] , \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , 
        \ScanLink63[6] , \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , 
        \ScanLink63[2] , \ScanLink63[1] , \ScanLink63[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load62[0] ), .Out({
        \Level1Out62[31] , \Level1Out62[30] , \Level1Out62[29] , 
        \Level1Out62[28] , \Level1Out62[27] , \Level1Out62[26] , 
        \Level1Out62[25] , \Level1Out62[24] , \Level1Out62[23] , 
        \Level1Out62[22] , \Level1Out62[21] , \Level1Out62[20] , 
        \Level1Out62[19] , \Level1Out62[18] , \Level1Out62[17] , 
        \Level1Out62[16] , \Level1Out62[15] , \Level1Out62[14] , 
        \Level1Out62[13] , \Level1Out62[12] , \Level1Out62[11] , 
        \Level1Out62[10] , \Level1Out62[9] , \Level1Out62[8] , 
        \Level1Out62[7] , \Level1Out62[6] , \Level1Out62[5] , \Level1Out62[4] , 
        \Level1Out62[3] , \Level1Out62[2] , \Level1Out62[1] , \Level1Out62[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load16[0] ), .Out({\Level16Out16[31] , \Level16Out16[30] , 
        \Level16Out16[29] , \Level16Out16[28] , \Level16Out16[27] , 
        \Level16Out16[26] , \Level16Out16[25] , \Level16Out16[24] , 
        \Level16Out16[23] , \Level16Out16[22] , \Level16Out16[21] , 
        \Level16Out16[20] , \Level16Out16[19] , \Level16Out16[18] , 
        \Level16Out16[17] , \Level16Out16[16] , \Level16Out16[15] , 
        \Level16Out16[14] , \Level16Out16[13] , \Level16Out16[12] , 
        \Level16Out16[11] , \Level16Out16[10] , \Level16Out16[9] , 
        \Level16Out16[8] , \Level16Out16[7] , \Level16Out16[6] , 
        \Level16Out16[5] , \Level16Out16[4] , \Level16Out16[3] , 
        \Level16Out16[2] , \Level16Out16[1] , \Level16Out16[0] }), .In1({
        \Level8Out16[31] , \Level8Out16[30] , \Level8Out16[29] , 
        \Level8Out16[28] , \Level8Out16[27] , \Level8Out16[26] , 
        \Level8Out16[25] , \Level8Out16[24] , \Level8Out16[23] , 
        \Level8Out16[22] , \Level8Out16[21] , \Level8Out16[20] , 
        \Level8Out16[19] , \Level8Out16[18] , \Level8Out16[17] , 
        \Level8Out16[16] , \Level8Out16[15] , \Level8Out16[14] , 
        \Level8Out16[13] , \Level8Out16[12] , \Level8Out16[11] , 
        \Level8Out16[10] , \Level8Out16[9] , \Level8Out16[8] , 
        \Level8Out16[7] , \Level8Out16[6] , \Level8Out16[5] , \Level8Out16[4] , 
        \Level8Out16[3] , \Level8Out16[2] , \Level8Out16[1] , \Level8Out16[0] 
        }), .In2({\Level8Out24[31] , \Level8Out24[30] , \Level8Out24[29] , 
        \Level8Out24[28] , \Level8Out24[27] , \Level8Out24[26] , 
        \Level8Out24[25] , \Level8Out24[24] , \Level8Out24[23] , 
        \Level8Out24[22] , \Level8Out24[21] , \Level8Out24[20] , 
        \Level8Out24[19] , \Level8Out24[18] , \Level8Out24[17] , 
        \Level8Out24[16] , \Level8Out24[15] , \Level8Out24[14] , 
        \Level8Out24[13] , \Level8Out24[12] , \Level8Out24[11] , 
        \Level8Out24[10] , \Level8Out24[9] , \Level8Out24[8] , 
        \Level8Out24[7] , \Level8Out24[6] , \Level8Out24[5] , \Level8Out24[4] , 
        \Level8Out24[3] , \Level8Out24[2] , \Level8Out24[1] , \Level8Out24[0] 
        }), .Read1(\Level8Load16[0] ), .Read2(\Level8Load24[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_30_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load30[0] ), .Out({\Level2Out30[31] , \Level2Out30[30] , 
        \Level2Out30[29] , \Level2Out30[28] , \Level2Out30[27] , 
        \Level2Out30[26] , \Level2Out30[25] , \Level2Out30[24] , 
        \Level2Out30[23] , \Level2Out30[22] , \Level2Out30[21] , 
        \Level2Out30[20] , \Level2Out30[19] , \Level2Out30[18] , 
        \Level2Out30[17] , \Level2Out30[16] , \Level2Out30[15] , 
        \Level2Out30[14] , \Level2Out30[13] , \Level2Out30[12] , 
        \Level2Out30[11] , \Level2Out30[10] , \Level2Out30[9] , 
        \Level2Out30[8] , \Level2Out30[7] , \Level2Out30[6] , \Level2Out30[5] , 
        \Level2Out30[4] , \Level2Out30[3] , \Level2Out30[2] , \Level2Out30[1] , 
        \Level2Out30[0] }), .In1({\Level1Out30[31] , \Level1Out30[30] , 
        \Level1Out30[29] , \Level1Out30[28] , \Level1Out30[27] , 
        \Level1Out30[26] , \Level1Out30[25] , \Level1Out30[24] , 
        \Level1Out30[23] , \Level1Out30[22] , \Level1Out30[21] , 
        \Level1Out30[20] , \Level1Out30[19] , \Level1Out30[18] , 
        \Level1Out30[17] , \Level1Out30[16] , \Level1Out30[15] , 
        \Level1Out30[14] , \Level1Out30[13] , \Level1Out30[12] , 
        \Level1Out30[11] , \Level1Out30[10] , \Level1Out30[9] , 
        \Level1Out30[8] , \Level1Out30[7] , \Level1Out30[6] , \Level1Out30[5] , 
        \Level1Out30[4] , \Level1Out30[3] , \Level1Out30[2] , \Level1Out30[1] , 
        \Level1Out30[0] }), .In2({\Level1Out31[31] , \Level1Out31[30] , 
        \Level1Out31[29] , \Level1Out31[28] , \Level1Out31[27] , 
        \Level1Out31[26] , \Level1Out31[25] , \Level1Out31[24] , 
        \Level1Out31[23] , \Level1Out31[22] , \Level1Out31[21] , 
        \Level1Out31[20] , \Level1Out31[19] , \Level1Out31[18] , 
        \Level1Out31[17] , \Level1Out31[16] , \Level1Out31[15] , 
        \Level1Out31[14] , \Level1Out31[13] , \Level1Out31[12] , 
        \Level1Out31[11] , \Level1Out31[10] , \Level1Out31[9] , 
        \Level1Out31[8] , \Level1Out31[7] , \Level1Out31[6] , \Level1Out31[5] , 
        \Level1Out31[4] , \Level1Out31[3] , \Level1Out31[2] , \Level1Out31[1] , 
        \Level1Out31[0] }), .Read1(\Level1Load30[0] ), .Read2(
        \Level1Load31[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load24[0] ), .Out({\Level2Out24[31] , \Level2Out24[30] , 
        \Level2Out24[29] , \Level2Out24[28] , \Level2Out24[27] , 
        \Level2Out24[26] , \Level2Out24[25] , \Level2Out24[24] , 
        \Level2Out24[23] , \Level2Out24[22] , \Level2Out24[21] , 
        \Level2Out24[20] , \Level2Out24[19] , \Level2Out24[18] , 
        \Level2Out24[17] , \Level2Out24[16] , \Level2Out24[15] , 
        \Level2Out24[14] , \Level2Out24[13] , \Level2Out24[12] , 
        \Level2Out24[11] , \Level2Out24[10] , \Level2Out24[9] , 
        \Level2Out24[8] , \Level2Out24[7] , \Level2Out24[6] , \Level2Out24[5] , 
        \Level2Out24[4] , \Level2Out24[3] , \Level2Out24[2] , \Level2Out24[1] , 
        \Level2Out24[0] }), .In1({\Level1Out24[31] , \Level1Out24[30] , 
        \Level1Out24[29] , \Level1Out24[28] , \Level1Out24[27] , 
        \Level1Out24[26] , \Level1Out24[25] , \Level1Out24[24] , 
        \Level1Out24[23] , \Level1Out24[22] , \Level1Out24[21] , 
        \Level1Out24[20] , \Level1Out24[19] , \Level1Out24[18] , 
        \Level1Out24[17] , \Level1Out24[16] , \Level1Out24[15] , 
        \Level1Out24[14] , \Level1Out24[13] , \Level1Out24[12] , 
        \Level1Out24[11] , \Level1Out24[10] , \Level1Out24[9] , 
        \Level1Out24[8] , \Level1Out24[7] , \Level1Out24[6] , \Level1Out24[5] , 
        \Level1Out24[4] , \Level1Out24[3] , \Level1Out24[2] , \Level1Out24[1] , 
        \Level1Out24[0] }), .In2({\Level1Out25[31] , \Level1Out25[30] , 
        \Level1Out25[29] , \Level1Out25[28] , \Level1Out25[27] , 
        \Level1Out25[26] , \Level1Out25[25] , \Level1Out25[24] , 
        \Level1Out25[23] , \Level1Out25[22] , \Level1Out25[21] , 
        \Level1Out25[20] , \Level1Out25[19] , \Level1Out25[18] , 
        \Level1Out25[17] , \Level1Out25[16] , \Level1Out25[15] , 
        \Level1Out25[14] , \Level1Out25[13] , \Level1Out25[12] , 
        \Level1Out25[11] , \Level1Out25[10] , \Level1Out25[9] , 
        \Level1Out25[8] , \Level1Out25[7] , \Level1Out25[6] , \Level1Out25[5] , 
        \Level1Out25[4] , \Level1Out25[3] , \Level1Out25[2] , \Level1Out25[1] , 
        \Level1Out25[0] }), .Read1(\Level1Load24[0] ), .Read2(
        \Level1Load25[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_12_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load12[0] ), .Out({\Level4Out12[31] , \Level4Out12[30] , 
        \Level4Out12[29] , \Level4Out12[28] , \Level4Out12[27] , 
        \Level4Out12[26] , \Level4Out12[25] , \Level4Out12[24] , 
        \Level4Out12[23] , \Level4Out12[22] , \Level4Out12[21] , 
        \Level4Out12[20] , \Level4Out12[19] , \Level4Out12[18] , 
        \Level4Out12[17] , \Level4Out12[16] , \Level4Out12[15] , 
        \Level4Out12[14] , \Level4Out12[13] , \Level4Out12[12] , 
        \Level4Out12[11] , \Level4Out12[10] , \Level4Out12[9] , 
        \Level4Out12[8] , \Level4Out12[7] , \Level4Out12[6] , \Level4Out12[5] , 
        \Level4Out12[4] , \Level4Out12[3] , \Level4Out12[2] , \Level4Out12[1] , 
        \Level4Out12[0] }), .In1({\Level2Out12[31] , \Level2Out12[30] , 
        \Level2Out12[29] , \Level2Out12[28] , \Level2Out12[27] , 
        \Level2Out12[26] , \Level2Out12[25] , \Level2Out12[24] , 
        \Level2Out12[23] , \Level2Out12[22] , \Level2Out12[21] , 
        \Level2Out12[20] , \Level2Out12[19] , \Level2Out12[18] , 
        \Level2Out12[17] , \Level2Out12[16] , \Level2Out12[15] , 
        \Level2Out12[14] , \Level2Out12[13] , \Level2Out12[12] , 
        \Level2Out12[11] , \Level2Out12[10] , \Level2Out12[9] , 
        \Level2Out12[8] , \Level2Out12[7] , \Level2Out12[6] , \Level2Out12[5] , 
        \Level2Out12[4] , \Level2Out12[3] , \Level2Out12[2] , \Level2Out12[1] , 
        \Level2Out12[0] }), .In2({\Level2Out14[31] , \Level2Out14[30] , 
        \Level2Out14[29] , \Level2Out14[28] , \Level2Out14[27] , 
        \Level2Out14[26] , \Level2Out14[25] , \Level2Out14[24] , 
        \Level2Out14[23] , \Level2Out14[22] , \Level2Out14[21] , 
        \Level2Out14[20] , \Level2Out14[19] , \Level2Out14[18] , 
        \Level2Out14[17] , \Level2Out14[16] , \Level2Out14[15] , 
        \Level2Out14[14] , \Level2Out14[13] , \Level2Out14[12] , 
        \Level2Out14[11] , \Level2Out14[10] , \Level2Out14[9] , 
        \Level2Out14[8] , \Level2Out14[7] , \Level2Out14[6] , \Level2Out14[5] , 
        \Level2Out14[4] , \Level2Out14[3] , \Level2Out14[2] , \Level2Out14[1] , 
        \Level2Out14[0] }), .Read1(\Level2Load12[0] ), .Read2(
        \Level2Load14[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_19 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink19[31] , \ScanLink19[30] , 
        \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , \ScanLink19[26] , 
        \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , \ScanLink19[22] , 
        \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , \ScanLink19[18] , 
        \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , \ScanLink19[14] , 
        \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , \ScanLink19[10] , 
        \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , \ScanLink19[6] , 
        \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , \ScanLink19[2] , 
        \ScanLink19[1] , \ScanLink19[0] }), .ScanOut({\ScanLink20[31] , 
        \ScanLink20[30] , \ScanLink20[29] , \ScanLink20[28] , \ScanLink20[27] , 
        \ScanLink20[26] , \ScanLink20[25] , \ScanLink20[24] , \ScanLink20[23] , 
        \ScanLink20[22] , \ScanLink20[21] , \ScanLink20[20] , \ScanLink20[19] , 
        \ScanLink20[18] , \ScanLink20[17] , \ScanLink20[16] , \ScanLink20[15] , 
        \ScanLink20[14] , \ScanLink20[13] , \ScanLink20[12] , \ScanLink20[11] , 
        \ScanLink20[10] , \ScanLink20[9] , \ScanLink20[8] , \ScanLink20[7] , 
        \ScanLink20[6] , \ScanLink20[5] , \ScanLink20[4] , \ScanLink20[3] , 
        \ScanLink20[2] , \ScanLink20[1] , \ScanLink20[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load19[0] ), .Out({
        \Level1Out19[31] , \Level1Out19[30] , \Level1Out19[29] , 
        \Level1Out19[28] , \Level1Out19[27] , \Level1Out19[26] , 
        \Level1Out19[25] , \Level1Out19[24] , \Level1Out19[23] , 
        \Level1Out19[22] , \Level1Out19[21] , \Level1Out19[20] , 
        \Level1Out19[19] , \Level1Out19[18] , \Level1Out19[17] , 
        \Level1Out19[16] , \Level1Out19[15] , \Level1Out19[14] , 
        \Level1Out19[13] , \Level1Out19[12] , \Level1Out19[11] , 
        \Level1Out19[10] , \Level1Out19[9] , \Level1Out19[8] , 
        \Level1Out19[7] , \Level1Out19[6] , \Level1Out19[5] , \Level1Out19[4] , 
        \Level1Out19[3] , \Level1Out19[2] , \Level1Out19[1] , \Level1Out19[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_37 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink37[31] , \ScanLink37[30] , 
        \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , \ScanLink37[26] , 
        \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , \ScanLink37[22] , 
        \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , \ScanLink37[18] , 
        \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , \ScanLink37[14] , 
        \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , \ScanLink37[10] , 
        \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , \ScanLink37[6] , 
        \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , \ScanLink37[2] , 
        \ScanLink37[1] , \ScanLink37[0] }), .ScanOut({\ScanLink38[31] , 
        \ScanLink38[30] , \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , 
        \ScanLink38[26] , \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , 
        \ScanLink38[22] , \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , 
        \ScanLink38[18] , \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , 
        \ScanLink38[14] , \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , 
        \ScanLink38[10] , \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , 
        \ScanLink38[6] , \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , 
        \ScanLink38[2] , \ScanLink38[1] , \ScanLink38[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load37[0] ), .Out({
        \Level1Out37[31] , \Level1Out37[30] , \Level1Out37[29] , 
        \Level1Out37[28] , \Level1Out37[27] , \Level1Out37[26] , 
        \Level1Out37[25] , \Level1Out37[24] , \Level1Out37[23] , 
        \Level1Out37[22] , \Level1Out37[21] , \Level1Out37[20] , 
        \Level1Out37[19] , \Level1Out37[18] , \Level1Out37[17] , 
        \Level1Out37[16] , \Level1Out37[15] , \Level1Out37[14] , 
        \Level1Out37[13] , \Level1Out37[12] , \Level1Out37[11] , 
        \Level1Out37[10] , \Level1Out37[9] , \Level1Out37[8] , 
        \Level1Out37[7] , \Level1Out37[6] , \Level1Out37[5] , \Level1Out37[4] , 
        \Level1Out37[3] , \Level1Out37[2] , \Level1Out37[1] , \Level1Out37[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_42 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink42[31] , \ScanLink42[30] , 
        \ScanLink42[29] , \ScanLink42[28] , \ScanLink42[27] , \ScanLink42[26] , 
        \ScanLink42[25] , \ScanLink42[24] , \ScanLink42[23] , \ScanLink42[22] , 
        \ScanLink42[21] , \ScanLink42[20] , \ScanLink42[19] , \ScanLink42[18] , 
        \ScanLink42[17] , \ScanLink42[16] , \ScanLink42[15] , \ScanLink42[14] , 
        \ScanLink42[13] , \ScanLink42[12] , \ScanLink42[11] , \ScanLink42[10] , 
        \ScanLink42[9] , \ScanLink42[8] , \ScanLink42[7] , \ScanLink42[6] , 
        \ScanLink42[5] , \ScanLink42[4] , \ScanLink42[3] , \ScanLink42[2] , 
        \ScanLink42[1] , \ScanLink42[0] }), .ScanOut({\ScanLink43[31] , 
        \ScanLink43[30] , \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , 
        \ScanLink43[26] , \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , 
        \ScanLink43[22] , \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , 
        \ScanLink43[18] , \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , 
        \ScanLink43[14] , \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , 
        \ScanLink43[10] , \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , 
        \ScanLink43[6] , \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , 
        \ScanLink43[2] , \ScanLink43[1] , \ScanLink43[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load42[0] ), .Out({
        \Level1Out42[31] , \Level1Out42[30] , \Level1Out42[29] , 
        \Level1Out42[28] , \Level1Out42[27] , \Level1Out42[26] , 
        \Level1Out42[25] , \Level1Out42[24] , \Level1Out42[23] , 
        \Level1Out42[22] , \Level1Out42[21] , \Level1Out42[20] , 
        \Level1Out42[19] , \Level1Out42[18] , \Level1Out42[17] , 
        \Level1Out42[16] , \Level1Out42[15] , \Level1Out42[14] , 
        \Level1Out42[13] , \Level1Out42[12] , \Level1Out42[11] , 
        \Level1Out42[10] , \Level1Out42[9] , \Level1Out42[8] , 
        \Level1Out42[7] , \Level1Out42[6] , \Level1Out42[5] , \Level1Out42[4] , 
        \Level1Out42[3] , \Level1Out42[2] , \Level1Out42[1] , \Level1Out42[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_59 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink59[31] , \ScanLink59[30] , 
        \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , \ScanLink59[26] , 
        \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , \ScanLink59[22] , 
        \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , \ScanLink59[18] , 
        \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , \ScanLink59[14] , 
        \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , \ScanLink59[10] , 
        \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , \ScanLink59[6] , 
        \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , \ScanLink59[2] , 
        \ScanLink59[1] , \ScanLink59[0] }), .ScanOut({\ScanLink60[31] , 
        \ScanLink60[30] , \ScanLink60[29] , \ScanLink60[28] , \ScanLink60[27] , 
        \ScanLink60[26] , \ScanLink60[25] , \ScanLink60[24] , \ScanLink60[23] , 
        \ScanLink60[22] , \ScanLink60[21] , \ScanLink60[20] , \ScanLink60[19] , 
        \ScanLink60[18] , \ScanLink60[17] , \ScanLink60[16] , \ScanLink60[15] , 
        \ScanLink60[14] , \ScanLink60[13] , \ScanLink60[12] , \ScanLink60[11] , 
        \ScanLink60[10] , \ScanLink60[9] , \ScanLink60[8] , \ScanLink60[7] , 
        \ScanLink60[6] , \ScanLink60[5] , \ScanLink60[4] , \ScanLink60[3] , 
        \ScanLink60[2] , \ScanLink60[1] , \ScanLink60[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load59[0] ), .Out({
        \Level1Out59[31] , \Level1Out59[30] , \Level1Out59[29] , 
        \Level1Out59[28] , \Level1Out59[27] , \Level1Out59[26] , 
        \Level1Out59[25] , \Level1Out59[24] , \Level1Out59[23] , 
        \Level1Out59[22] , \Level1Out59[21] , \Level1Out59[20] , 
        \Level1Out59[19] , \Level1Out59[18] , \Level1Out59[17] , 
        \Level1Out59[16] , \Level1Out59[15] , \Level1Out59[14] , 
        \Level1Out59[13] , \Level1Out59[12] , \Level1Out59[11] , 
        \Level1Out59[10] , \Level1Out59[9] , \Level1Out59[8] , 
        \Level1Out59[7] , \Level1Out59[6] , \Level1Out59[5] , \Level1Out59[4] , 
        \Level1Out59[3] , \Level1Out59[2] , \Level1Out59[1] , \Level1Out59[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load0[0] ), .Out({\Level16Out0[31] , \Level16Out0[30] , 
        \Level16Out0[29] , \Level16Out0[28] , \Level16Out0[27] , 
        \Level16Out0[26] , \Level16Out0[25] , \Level16Out0[24] , 
        \Level16Out0[23] , \Level16Out0[22] , \Level16Out0[21] , 
        \Level16Out0[20] , \Level16Out0[19] , \Level16Out0[18] , 
        \Level16Out0[17] , \Level16Out0[16] , \Level16Out0[15] , 
        \Level16Out0[14] , \Level16Out0[13] , \Level16Out0[12] , 
        \Level16Out0[11] , \Level16Out0[10] , \Level16Out0[9] , 
        \Level16Out0[8] , \Level16Out0[7] , \Level16Out0[6] , \Level16Out0[5] , 
        \Level16Out0[4] , \Level16Out0[3] , \Level16Out0[2] , \Level16Out0[1] , 
        \Level16Out0[0] }), .In1({\Level8Out0[31] , \Level8Out0[30] , 
        \Level8Out0[29] , \Level8Out0[28] , \Level8Out0[27] , \Level8Out0[26] , 
        \Level8Out0[25] , \Level8Out0[24] , \Level8Out0[23] , \Level8Out0[22] , 
        \Level8Out0[21] , \Level8Out0[20] , \Level8Out0[19] , \Level8Out0[18] , 
        \Level8Out0[17] , \Level8Out0[16] , \Level8Out0[15] , \Level8Out0[14] , 
        \Level8Out0[13] , \Level8Out0[12] , \Level8Out0[11] , \Level8Out0[10] , 
        \Level8Out0[9] , \Level8Out0[8] , \Level8Out0[7] , \Level8Out0[6] , 
        \Level8Out0[5] , \Level8Out0[4] , \Level8Out0[3] , \Level8Out0[2] , 
        \Level8Out0[1] , \Level8Out0[0] }), .In2({\Level8Out8[31] , 
        \Level8Out8[30] , \Level8Out8[29] , \Level8Out8[28] , \Level8Out8[27] , 
        \Level8Out8[26] , \Level8Out8[25] , \Level8Out8[24] , \Level8Out8[23] , 
        \Level8Out8[22] , \Level8Out8[21] , \Level8Out8[20] , \Level8Out8[19] , 
        \Level8Out8[18] , \Level8Out8[17] , \Level8Out8[16] , \Level8Out8[15] , 
        \Level8Out8[14] , \Level8Out8[13] , \Level8Out8[12] , \Level8Out8[11] , 
        \Level8Out8[10] , \Level8Out8[9] , \Level8Out8[8] , \Level8Out8[7] , 
        \Level8Out8[6] , \Level8Out8[5] , \Level8Out8[4] , \Level8Out8[3] , 
        \Level8Out8[2] , \Level8Out8[1] , \Level8Out8[0] }), .Read1(
        \Level8Load0[0] ), .Read2(\Level8Load8[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load16[0] ), .Out({\Level2Out16[31] , \Level2Out16[30] , 
        \Level2Out16[29] , \Level2Out16[28] , \Level2Out16[27] , 
        \Level2Out16[26] , \Level2Out16[25] , \Level2Out16[24] , 
        \Level2Out16[23] , \Level2Out16[22] , \Level2Out16[21] , 
        \Level2Out16[20] , \Level2Out16[19] , \Level2Out16[18] , 
        \Level2Out16[17] , \Level2Out16[16] , \Level2Out16[15] , 
        \Level2Out16[14] , \Level2Out16[13] , \Level2Out16[12] , 
        \Level2Out16[11] , \Level2Out16[10] , \Level2Out16[9] , 
        \Level2Out16[8] , \Level2Out16[7] , \Level2Out16[6] , \Level2Out16[5] , 
        \Level2Out16[4] , \Level2Out16[3] , \Level2Out16[2] , \Level2Out16[1] , 
        \Level2Out16[0] }), .In1({\Level1Out16[31] , \Level1Out16[30] , 
        \Level1Out16[29] , \Level1Out16[28] , \Level1Out16[27] , 
        \Level1Out16[26] , \Level1Out16[25] , \Level1Out16[24] , 
        \Level1Out16[23] , \Level1Out16[22] , \Level1Out16[21] , 
        \Level1Out16[20] , \Level1Out16[19] , \Level1Out16[18] , 
        \Level1Out16[17] , \Level1Out16[16] , \Level1Out16[15] , 
        \Level1Out16[14] , \Level1Out16[13] , \Level1Out16[12] , 
        \Level1Out16[11] , \Level1Out16[10] , \Level1Out16[9] , 
        \Level1Out16[8] , \Level1Out16[7] , \Level1Out16[6] , \Level1Out16[5] , 
        \Level1Out16[4] , \Level1Out16[3] , \Level1Out16[2] , \Level1Out16[1] , 
        \Level1Out16[0] }), .In2({\Level1Out17[31] , \Level1Out17[30] , 
        \Level1Out17[29] , \Level1Out17[28] , \Level1Out17[27] , 
        \Level1Out17[26] , \Level1Out17[25] , \Level1Out17[24] , 
        \Level1Out17[23] , \Level1Out17[22] , \Level1Out17[21] , 
        \Level1Out17[20] , \Level1Out17[19] , \Level1Out17[18] , 
        \Level1Out17[17] , \Level1Out17[16] , \Level1Out17[15] , 
        \Level1Out17[14] , \Level1Out17[13] , \Level1Out17[12] , 
        \Level1Out17[11] , \Level1Out17[10] , \Level1Out17[9] , 
        \Level1Out17[8] , \Level1Out17[7] , \Level1Out17[6] , \Level1Out17[5] , 
        \Level1Out17[4] , \Level1Out17[3] , \Level1Out17[2] , \Level1Out17[1] , 
        \Level1Out17[0] }), .Read1(\Level1Load16[0] ), .Read2(
        \Level1Load17[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_20_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load20[0] ), .Out({\Level4Out20[31] , \Level4Out20[30] , 
        \Level4Out20[29] , \Level4Out20[28] , \Level4Out20[27] , 
        \Level4Out20[26] , \Level4Out20[25] , \Level4Out20[24] , 
        \Level4Out20[23] , \Level4Out20[22] , \Level4Out20[21] , 
        \Level4Out20[20] , \Level4Out20[19] , \Level4Out20[18] , 
        \Level4Out20[17] , \Level4Out20[16] , \Level4Out20[15] , 
        \Level4Out20[14] , \Level4Out20[13] , \Level4Out20[12] , 
        \Level4Out20[11] , \Level4Out20[10] , \Level4Out20[9] , 
        \Level4Out20[8] , \Level4Out20[7] , \Level4Out20[6] , \Level4Out20[5] , 
        \Level4Out20[4] , \Level4Out20[3] , \Level4Out20[2] , \Level4Out20[1] , 
        \Level4Out20[0] }), .In1({\Level2Out20[31] , \Level2Out20[30] , 
        \Level2Out20[29] , \Level2Out20[28] , \Level2Out20[27] , 
        \Level2Out20[26] , \Level2Out20[25] , \Level2Out20[24] , 
        \Level2Out20[23] , \Level2Out20[22] , \Level2Out20[21] , 
        \Level2Out20[20] , \Level2Out20[19] , \Level2Out20[18] , 
        \Level2Out20[17] , \Level2Out20[16] , \Level2Out20[15] , 
        \Level2Out20[14] , \Level2Out20[13] , \Level2Out20[12] , 
        \Level2Out20[11] , \Level2Out20[10] , \Level2Out20[9] , 
        \Level2Out20[8] , \Level2Out20[7] , \Level2Out20[6] , \Level2Out20[5] , 
        \Level2Out20[4] , \Level2Out20[3] , \Level2Out20[2] , \Level2Out20[1] , 
        \Level2Out20[0] }), .In2({\Level2Out22[31] , \Level2Out22[30] , 
        \Level2Out22[29] , \Level2Out22[28] , \Level2Out22[27] , 
        \Level2Out22[26] , \Level2Out22[25] , \Level2Out22[24] , 
        \Level2Out22[23] , \Level2Out22[22] , \Level2Out22[21] , 
        \Level2Out22[20] , \Level2Out22[19] , \Level2Out22[18] , 
        \Level2Out22[17] , \Level2Out22[16] , \Level2Out22[15] , 
        \Level2Out22[14] , \Level2Out22[13] , \Level2Out22[12] , 
        \Level2Out22[11] , \Level2Out22[10] , \Level2Out22[9] , 
        \Level2Out22[8] , \Level2Out22[7] , \Level2Out22[6] , \Level2Out22[5] , 
        \Level2Out22[4] , \Level2Out22[3] , \Level2Out22[2] , \Level2Out22[1] , 
        \Level2Out22[0] }), .Read1(\Level2Load20[0] ), .Read2(
        \Level2Load22[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_0_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load0[0] ), .Out({\Level8Out0[31] , \Level8Out0[30] , 
        \Level8Out0[29] , \Level8Out0[28] , \Level8Out0[27] , \Level8Out0[26] , 
        \Level8Out0[25] , \Level8Out0[24] , \Level8Out0[23] , \Level8Out0[22] , 
        \Level8Out0[21] , \Level8Out0[20] , \Level8Out0[19] , \Level8Out0[18] , 
        \Level8Out0[17] , \Level8Out0[16] , \Level8Out0[15] , \Level8Out0[14] , 
        \Level8Out0[13] , \Level8Out0[12] , \Level8Out0[11] , \Level8Out0[10] , 
        \Level8Out0[9] , \Level8Out0[8] , \Level8Out0[7] , \Level8Out0[6] , 
        \Level8Out0[5] , \Level8Out0[4] , \Level8Out0[3] , \Level8Out0[2] , 
        \Level8Out0[1] , \Level8Out0[0] }), .In1({\Level4Out0[31] , 
        \Level4Out0[30] , \Level4Out0[29] , \Level4Out0[28] , \Level4Out0[27] , 
        \Level4Out0[26] , \Level4Out0[25] , \Level4Out0[24] , \Level4Out0[23] , 
        \Level4Out0[22] , \Level4Out0[21] , \Level4Out0[20] , \Level4Out0[19] , 
        \Level4Out0[18] , \Level4Out0[17] , \Level4Out0[16] , \Level4Out0[15] , 
        \Level4Out0[14] , \Level4Out0[13] , \Level4Out0[12] , \Level4Out0[11] , 
        \Level4Out0[10] , \Level4Out0[9] , \Level4Out0[8] , \Level4Out0[7] , 
        \Level4Out0[6] , \Level4Out0[5] , \Level4Out0[4] , \Level4Out0[3] , 
        \Level4Out0[2] , \Level4Out0[1] , \Level4Out0[0] }), .In2({
        \Level4Out4[31] , \Level4Out4[30] , \Level4Out4[29] , \Level4Out4[28] , 
        \Level4Out4[27] , \Level4Out4[26] , \Level4Out4[25] , \Level4Out4[24] , 
        \Level4Out4[23] , \Level4Out4[22] , \Level4Out4[21] , \Level4Out4[20] , 
        \Level4Out4[19] , \Level4Out4[18] , \Level4Out4[17] , \Level4Out4[16] , 
        \Level4Out4[15] , \Level4Out4[14] , \Level4Out4[13] , \Level4Out4[12] , 
        \Level4Out4[11] , \Level4Out4[10] , \Level4Out4[9] , \Level4Out4[8] , 
        \Level4Out4[7] , \Level4Out4[6] , \Level4Out4[5] , \Level4Out4[4] , 
        \Level4Out4[3] , \Level4Out4[2] , \Level4Out4[1] , \Level4Out4[0] }), 
        .Read1(\Level4Load0[0] ), .Read2(\Level4Load4[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_50 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink50[31] , \ScanLink50[30] , 
        \ScanLink50[29] , \ScanLink50[28] , \ScanLink50[27] , \ScanLink50[26] , 
        \ScanLink50[25] , \ScanLink50[24] , \ScanLink50[23] , \ScanLink50[22] , 
        \ScanLink50[21] , \ScanLink50[20] , \ScanLink50[19] , \ScanLink50[18] , 
        \ScanLink50[17] , \ScanLink50[16] , \ScanLink50[15] , \ScanLink50[14] , 
        \ScanLink50[13] , \ScanLink50[12] , \ScanLink50[11] , \ScanLink50[10] , 
        \ScanLink50[9] , \ScanLink50[8] , \ScanLink50[7] , \ScanLink50[6] , 
        \ScanLink50[5] , \ScanLink50[4] , \ScanLink50[3] , \ScanLink50[2] , 
        \ScanLink50[1] , \ScanLink50[0] }), .ScanOut({\ScanLink51[31] , 
        \ScanLink51[30] , \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , 
        \ScanLink51[26] , \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , 
        \ScanLink51[22] , \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , 
        \ScanLink51[18] , \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , 
        \ScanLink51[14] , \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , 
        \ScanLink51[10] , \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , 
        \ScanLink51[6] , \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , 
        \ScanLink51[2] , \ScanLink51[1] , \ScanLink51[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load50[0] ), .Out({
        \Level1Out50[31] , \Level1Out50[30] , \Level1Out50[29] , 
        \Level1Out50[28] , \Level1Out50[27] , \Level1Out50[26] , 
        \Level1Out50[25] , \Level1Out50[24] , \Level1Out50[23] , 
        \Level1Out50[22] , \Level1Out50[21] , \Level1Out50[20] , 
        \Level1Out50[19] , \Level1Out50[18] , \Level1Out50[17] , 
        \Level1Out50[16] , \Level1Out50[15] , \Level1Out50[14] , 
        \Level1Out50[13] , \Level1Out50[12] , \Level1Out50[11] , 
        \Level1Out50[10] , \Level1Out50[9] , \Level1Out50[8] , 
        \Level1Out50[7] , \Level1Out50[6] , \Level1Out50[5] , \Level1Out50[4] , 
        \Level1Out50[3] , \Level1Out50[2] , \Level1Out50[1] , \Level1Out50[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_46_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load46[0] ), .Out({\Level2Out46[31] , \Level2Out46[30] , 
        \Level2Out46[29] , \Level2Out46[28] , \Level2Out46[27] , 
        \Level2Out46[26] , \Level2Out46[25] , \Level2Out46[24] , 
        \Level2Out46[23] , \Level2Out46[22] , \Level2Out46[21] , 
        \Level2Out46[20] , \Level2Out46[19] , \Level2Out46[18] , 
        \Level2Out46[17] , \Level2Out46[16] , \Level2Out46[15] , 
        \Level2Out46[14] , \Level2Out46[13] , \Level2Out46[12] , 
        \Level2Out46[11] , \Level2Out46[10] , \Level2Out46[9] , 
        \Level2Out46[8] , \Level2Out46[7] , \Level2Out46[6] , \Level2Out46[5] , 
        \Level2Out46[4] , \Level2Out46[3] , \Level2Out46[2] , \Level2Out46[1] , 
        \Level2Out46[0] }), .In1({\Level1Out46[31] , \Level1Out46[30] , 
        \Level1Out46[29] , \Level1Out46[28] , \Level1Out46[27] , 
        \Level1Out46[26] , \Level1Out46[25] , \Level1Out46[24] , 
        \Level1Out46[23] , \Level1Out46[22] , \Level1Out46[21] , 
        \Level1Out46[20] , \Level1Out46[19] , \Level1Out46[18] , 
        \Level1Out46[17] , \Level1Out46[16] , \Level1Out46[15] , 
        \Level1Out46[14] , \Level1Out46[13] , \Level1Out46[12] , 
        \Level1Out46[11] , \Level1Out46[10] , \Level1Out46[9] , 
        \Level1Out46[8] , \Level1Out46[7] , \Level1Out46[6] , \Level1Out46[5] , 
        \Level1Out46[4] , \Level1Out46[3] , \Level1Out46[2] , \Level1Out46[1] , 
        \Level1Out46[0] }), .In2({\Level1Out47[31] , \Level1Out47[30] , 
        \Level1Out47[29] , \Level1Out47[28] , \Level1Out47[27] , 
        \Level1Out47[26] , \Level1Out47[25] , \Level1Out47[24] , 
        \Level1Out47[23] , \Level1Out47[22] , \Level1Out47[21] , 
        \Level1Out47[20] , \Level1Out47[19] , \Level1Out47[18] , 
        \Level1Out47[17] , \Level1Out47[16] , \Level1Out47[15] , 
        \Level1Out47[14] , \Level1Out47[13] , \Level1Out47[12] , 
        \Level1Out47[11] , \Level1Out47[10] , \Level1Out47[9] , 
        \Level1Out47[8] , \Level1Out47[7] , \Level1Out47[6] , \Level1Out47[5] , 
        \Level1Out47[4] , \Level1Out47[3] , \Level1Out47[2] , \Level1Out47[1] , 
        \Level1Out47[0] }), .Read1(\Level1Load46[0] ), .Read2(
        \Level1Load47[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_40_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load40[0] ), .Out({\Level8Out40[31] , \Level8Out40[30] , 
        \Level8Out40[29] , \Level8Out40[28] , \Level8Out40[27] , 
        \Level8Out40[26] , \Level8Out40[25] , \Level8Out40[24] , 
        \Level8Out40[23] , \Level8Out40[22] , \Level8Out40[21] , 
        \Level8Out40[20] , \Level8Out40[19] , \Level8Out40[18] , 
        \Level8Out40[17] , \Level8Out40[16] , \Level8Out40[15] , 
        \Level8Out40[14] , \Level8Out40[13] , \Level8Out40[12] , 
        \Level8Out40[11] , \Level8Out40[10] , \Level8Out40[9] , 
        \Level8Out40[8] , \Level8Out40[7] , \Level8Out40[6] , \Level8Out40[5] , 
        \Level8Out40[4] , \Level8Out40[3] , \Level8Out40[2] , \Level8Out40[1] , 
        \Level8Out40[0] }), .In1({\Level4Out40[31] , \Level4Out40[30] , 
        \Level4Out40[29] , \Level4Out40[28] , \Level4Out40[27] , 
        \Level4Out40[26] , \Level4Out40[25] , \Level4Out40[24] , 
        \Level4Out40[23] , \Level4Out40[22] , \Level4Out40[21] , 
        \Level4Out40[20] , \Level4Out40[19] , \Level4Out40[18] , 
        \Level4Out40[17] , \Level4Out40[16] , \Level4Out40[15] , 
        \Level4Out40[14] , \Level4Out40[13] , \Level4Out40[12] , 
        \Level4Out40[11] , \Level4Out40[10] , \Level4Out40[9] , 
        \Level4Out40[8] , \Level4Out40[7] , \Level4Out40[6] , \Level4Out40[5] , 
        \Level4Out40[4] , \Level4Out40[3] , \Level4Out40[2] , \Level4Out40[1] , 
        \Level4Out40[0] }), .In2({\Level4Out44[31] , \Level4Out44[30] , 
        \Level4Out44[29] , \Level4Out44[28] , \Level4Out44[27] , 
        \Level4Out44[26] , \Level4Out44[25] , \Level4Out44[24] , 
        \Level4Out44[23] , \Level4Out44[22] , \Level4Out44[21] , 
        \Level4Out44[20] , \Level4Out44[19] , \Level4Out44[18] , 
        \Level4Out44[17] , \Level4Out44[16] , \Level4Out44[15] , 
        \Level4Out44[14] , \Level4Out44[13] , \Level4Out44[12] , 
        \Level4Out44[11] , \Level4Out44[10] , \Level4Out44[9] , 
        \Level4Out44[8] , \Level4Out44[7] , \Level4Out44[6] , \Level4Out44[5] , 
        \Level4Out44[4] , \Level4Out44[3] , \Level4Out44[2] , \Level4Out44[1] , 
        \Level4Out44[0] }), .Read1(\Level4Load40[0] ), .Read2(
        \Level4Load44[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_11 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink11[31] , \ScanLink11[30] , 
        \ScanLink11[29] , \ScanLink11[28] , \ScanLink11[27] , \ScanLink11[26] , 
        \ScanLink11[25] , \ScanLink11[24] , \ScanLink11[23] , \ScanLink11[22] , 
        \ScanLink11[21] , \ScanLink11[20] , \ScanLink11[19] , \ScanLink11[18] , 
        \ScanLink11[17] , \ScanLink11[16] , \ScanLink11[15] , \ScanLink11[14] , 
        \ScanLink11[13] , \ScanLink11[12] , \ScanLink11[11] , \ScanLink11[10] , 
        \ScanLink11[9] , \ScanLink11[8] , \ScanLink11[7] , \ScanLink11[6] , 
        \ScanLink11[5] , \ScanLink11[4] , \ScanLink11[3] , \ScanLink11[2] , 
        \ScanLink11[1] , \ScanLink11[0] }), .ScanOut({\ScanLink12[31] , 
        \ScanLink12[30] , \ScanLink12[29] , \ScanLink12[28] , \ScanLink12[27] , 
        \ScanLink12[26] , \ScanLink12[25] , \ScanLink12[24] , \ScanLink12[23] , 
        \ScanLink12[22] , \ScanLink12[21] , \ScanLink12[20] , \ScanLink12[19] , 
        \ScanLink12[18] , \ScanLink12[17] , \ScanLink12[16] , \ScanLink12[15] , 
        \ScanLink12[14] , \ScanLink12[13] , \ScanLink12[12] , \ScanLink12[11] , 
        \ScanLink12[10] , \ScanLink12[9] , \ScanLink12[8] , \ScanLink12[7] , 
        \ScanLink12[6] , \ScanLink12[5] , \ScanLink12[4] , \ScanLink12[3] , 
        \ScanLink12[2] , \ScanLink12[1] , \ScanLink12[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load11[0] ), .Out({
        \Level1Out11[31] , \Level1Out11[30] , \Level1Out11[29] , 
        \Level1Out11[28] , \Level1Out11[27] , \Level1Out11[26] , 
        \Level1Out11[25] , \Level1Out11[24] , \Level1Out11[23] , 
        \Level1Out11[22] , \Level1Out11[21] , \Level1Out11[20] , 
        \Level1Out11[19] , \Level1Out11[18] , \Level1Out11[17] , 
        \Level1Out11[16] , \Level1Out11[15] , \Level1Out11[14] , 
        \Level1Out11[13] , \Level1Out11[12] , \Level1Out11[11] , 
        \Level1Out11[10] , \Level1Out11[9] , \Level1Out11[8] , 
        \Level1Out11[7] , \Level1Out11[6] , \Level1Out11[5] , \Level1Out11[4] , 
        \Level1Out11[3] , \Level1Out11[2] , \Level1Out11[1] , \Level1Out11[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_25 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink25[31] , \ScanLink25[30] , 
        \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , \ScanLink25[26] , 
        \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , \ScanLink25[22] , 
        \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , \ScanLink25[18] , 
        \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , \ScanLink25[14] , 
        \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , \ScanLink25[10] , 
        \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , \ScanLink25[6] , 
        \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , \ScanLink25[2] , 
        \ScanLink25[1] , \ScanLink25[0] }), .ScanOut({\ScanLink26[31] , 
        \ScanLink26[30] , \ScanLink26[29] , \ScanLink26[28] , \ScanLink26[27] , 
        \ScanLink26[26] , \ScanLink26[25] , \ScanLink26[24] , \ScanLink26[23] , 
        \ScanLink26[22] , \ScanLink26[21] , \ScanLink26[20] , \ScanLink26[19] , 
        \ScanLink26[18] , \ScanLink26[17] , \ScanLink26[16] , \ScanLink26[15] , 
        \ScanLink26[14] , \ScanLink26[13] , \ScanLink26[12] , \ScanLink26[11] , 
        \ScanLink26[10] , \ScanLink26[9] , \ScanLink26[8] , \ScanLink26[7] , 
        \ScanLink26[6] , \ScanLink26[5] , \ScanLink26[4] , \ScanLink26[3] , 
        \ScanLink26[2] , \ScanLink26[1] , \ScanLink26[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load25[0] ), .Out({
        \Level1Out25[31] , \Level1Out25[30] , \Level1Out25[29] , 
        \Level1Out25[28] , \Level1Out25[27] , \Level1Out25[26] , 
        \Level1Out25[25] , \Level1Out25[24] , \Level1Out25[23] , 
        \Level1Out25[22] , \Level1Out25[21] , \Level1Out25[20] , 
        \Level1Out25[19] , \Level1Out25[18] , \Level1Out25[17] , 
        \Level1Out25[16] , \Level1Out25[15] , \Level1Out25[14] , 
        \Level1Out25[13] , \Level1Out25[12] , \Level1Out25[11] , 
        \Level1Out25[10] , \Level1Out25[9] , \Level1Out25[8] , 
        \Level1Out25[7] , \Level1Out25[6] , \Level1Out25[5] , \Level1Out25[4] , 
        \Level1Out25[3] , \Level1Out25[2] , \Level1Out25[1] , \Level1Out25[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_43 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink43[31] , \ScanLink43[30] , 
        \ScanLink43[29] , \ScanLink43[28] , \ScanLink43[27] , \ScanLink43[26] , 
        \ScanLink43[25] , \ScanLink43[24] , \ScanLink43[23] , \ScanLink43[22] , 
        \ScanLink43[21] , \ScanLink43[20] , \ScanLink43[19] , \ScanLink43[18] , 
        \ScanLink43[17] , \ScanLink43[16] , \ScanLink43[15] , \ScanLink43[14] , 
        \ScanLink43[13] , \ScanLink43[12] , \ScanLink43[11] , \ScanLink43[10] , 
        \ScanLink43[9] , \ScanLink43[8] , \ScanLink43[7] , \ScanLink43[6] , 
        \ScanLink43[5] , \ScanLink43[4] , \ScanLink43[3] , \ScanLink43[2] , 
        \ScanLink43[1] , \ScanLink43[0] }), .ScanOut({\ScanLink44[31] , 
        \ScanLink44[30] , \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , 
        \ScanLink44[26] , \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , 
        \ScanLink44[22] , \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , 
        \ScanLink44[18] , \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , 
        \ScanLink44[14] , \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , 
        \ScanLink44[10] , \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , 
        \ScanLink44[6] , \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , 
        \ScanLink44[2] , \ScanLink44[1] , \ScanLink44[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load43[0] ), .Out({
        \Level1Out43[31] , \Level1Out43[30] , \Level1Out43[29] , 
        \Level1Out43[28] , \Level1Out43[27] , \Level1Out43[26] , 
        \Level1Out43[25] , \Level1Out43[24] , \Level1Out43[23] , 
        \Level1Out43[22] , \Level1Out43[21] , \Level1Out43[20] , 
        \Level1Out43[19] , \Level1Out43[18] , \Level1Out43[17] , 
        \Level1Out43[16] , \Level1Out43[15] , \Level1Out43[14] , 
        \Level1Out43[13] , \Level1Out43[12] , \Level1Out43[11] , 
        \Level1Out43[10] , \Level1Out43[9] , \Level1Out43[8] , 
        \Level1Out43[7] , \Level1Out43[6] , \Level1Out43[5] , \Level1Out43[4] , 
        \Level1Out43[3] , \Level1Out43[2] , \Level1Out43[1] , \Level1Out43[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load6[0] ), .Out({\Level2Out6[31] , \Level2Out6[30] , 
        \Level2Out6[29] , \Level2Out6[28] , \Level2Out6[27] , \Level2Out6[26] , 
        \Level2Out6[25] , \Level2Out6[24] , \Level2Out6[23] , \Level2Out6[22] , 
        \Level2Out6[21] , \Level2Out6[20] , \Level2Out6[19] , \Level2Out6[18] , 
        \Level2Out6[17] , \Level2Out6[16] , \Level2Out6[15] , \Level2Out6[14] , 
        \Level2Out6[13] , \Level2Out6[12] , \Level2Out6[11] , \Level2Out6[10] , 
        \Level2Out6[9] , \Level2Out6[8] , \Level2Out6[7] , \Level2Out6[6] , 
        \Level2Out6[5] , \Level2Out6[4] , \Level2Out6[3] , \Level2Out6[2] , 
        \Level2Out6[1] , \Level2Out6[0] }), .In1({\Level1Out6[31] , 
        \Level1Out6[30] , \Level1Out6[29] , \Level1Out6[28] , \Level1Out6[27] , 
        \Level1Out6[26] , \Level1Out6[25] , \Level1Out6[24] , \Level1Out6[23] , 
        \Level1Out6[22] , \Level1Out6[21] , \Level1Out6[20] , \Level1Out6[19] , 
        \Level1Out6[18] , \Level1Out6[17] , \Level1Out6[16] , \Level1Out6[15] , 
        \Level1Out6[14] , \Level1Out6[13] , \Level1Out6[12] , \Level1Out6[11] , 
        \Level1Out6[10] , \Level1Out6[9] , \Level1Out6[8] , \Level1Out6[7] , 
        \Level1Out6[6] , \Level1Out6[5] , \Level1Out6[4] , \Level1Out6[3] , 
        \Level1Out6[2] , \Level1Out6[1] , \Level1Out6[0] }), .In2({
        \Level1Out7[31] , \Level1Out7[30] , \Level1Out7[29] , \Level1Out7[28] , 
        \Level1Out7[27] , \Level1Out7[26] , \Level1Out7[25] , \Level1Out7[24] , 
        \Level1Out7[23] , \Level1Out7[22] , \Level1Out7[21] , \Level1Out7[20] , 
        \Level1Out7[19] , \Level1Out7[18] , \Level1Out7[17] , \Level1Out7[16] , 
        \Level1Out7[15] , \Level1Out7[14] , \Level1Out7[13] , \Level1Out7[12] , 
        \Level1Out7[11] , \Level1Out7[10] , \Level1Out7[9] , \Level1Out7[8] , 
        \Level1Out7[7] , \Level1Out7[6] , \Level1Out7[5] , \Level1Out7[4] , 
        \Level1Out7[3] , \Level1Out7[2] , \Level1Out7[1] , \Level1Out7[0] }), 
        .Read1(\Level1Load6[0] ), .Read2(\Level1Load7[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_34_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load34[0] ), .Out({\Level2Out34[31] , \Level2Out34[30] , 
        \Level2Out34[29] , \Level2Out34[28] , \Level2Out34[27] , 
        \Level2Out34[26] , \Level2Out34[25] , \Level2Out34[24] , 
        \Level2Out34[23] , \Level2Out34[22] , \Level2Out34[21] , 
        \Level2Out34[20] , \Level2Out34[19] , \Level2Out34[18] , 
        \Level2Out34[17] , \Level2Out34[16] , \Level2Out34[15] , 
        \Level2Out34[14] , \Level2Out34[13] , \Level2Out34[12] , 
        \Level2Out34[11] , \Level2Out34[10] , \Level2Out34[9] , 
        \Level2Out34[8] , \Level2Out34[7] , \Level2Out34[6] , \Level2Out34[5] , 
        \Level2Out34[4] , \Level2Out34[3] , \Level2Out34[2] , \Level2Out34[1] , 
        \Level2Out34[0] }), .In1({\Level1Out34[31] , \Level1Out34[30] , 
        \Level1Out34[29] , \Level1Out34[28] , \Level1Out34[27] , 
        \Level1Out34[26] , \Level1Out34[25] , \Level1Out34[24] , 
        \Level1Out34[23] , \Level1Out34[22] , \Level1Out34[21] , 
        \Level1Out34[20] , \Level1Out34[19] , \Level1Out34[18] , 
        \Level1Out34[17] , \Level1Out34[16] , \Level1Out34[15] , 
        \Level1Out34[14] , \Level1Out34[13] , \Level1Out34[12] , 
        \Level1Out34[11] , \Level1Out34[10] , \Level1Out34[9] , 
        \Level1Out34[8] , \Level1Out34[7] , \Level1Out34[6] , \Level1Out34[5] , 
        \Level1Out34[4] , \Level1Out34[3] , \Level1Out34[2] , \Level1Out34[1] , 
        \Level1Out34[0] }), .In2({\Level1Out35[31] , \Level1Out35[30] , 
        \Level1Out35[29] , \Level1Out35[28] , \Level1Out35[27] , 
        \Level1Out35[26] , \Level1Out35[25] , \Level1Out35[24] , 
        \Level1Out35[23] , \Level1Out35[22] , \Level1Out35[21] , 
        \Level1Out35[20] , \Level1Out35[19] , \Level1Out35[18] , 
        \Level1Out35[17] , \Level1Out35[16] , \Level1Out35[15] , 
        \Level1Out35[14] , \Level1Out35[13] , \Level1Out35[12] , 
        \Level1Out35[11] , \Level1Out35[10] , \Level1Out35[9] , 
        \Level1Out35[8] , \Level1Out35[7] , \Level1Out35[6] , \Level1Out35[5] , 
        \Level1Out35[4] , \Level1Out35[3] , \Level1Out35[2] , \Level1Out35[1] , 
        \Level1Out35[0] }), .Read1(\Level1Load34[0] ), .Read2(
        \Level1Load35[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level16Load32[0] ), .Out({\Level16Out32[31] , \Level16Out32[30] , 
        \Level16Out32[29] , \Level16Out32[28] , \Level16Out32[27] , 
        \Level16Out32[26] , \Level16Out32[25] , \Level16Out32[24] , 
        \Level16Out32[23] , \Level16Out32[22] , \Level16Out32[21] , 
        \Level16Out32[20] , \Level16Out32[19] , \Level16Out32[18] , 
        \Level16Out32[17] , \Level16Out32[16] , \Level16Out32[15] , 
        \Level16Out32[14] , \Level16Out32[13] , \Level16Out32[12] , 
        \Level16Out32[11] , \Level16Out32[10] , \Level16Out32[9] , 
        \Level16Out32[8] , \Level16Out32[7] , \Level16Out32[6] , 
        \Level16Out32[5] , \Level16Out32[4] , \Level16Out32[3] , 
        \Level16Out32[2] , \Level16Out32[1] , \Level16Out32[0] }), .In1({
        \Level8Out32[31] , \Level8Out32[30] , \Level8Out32[29] , 
        \Level8Out32[28] , \Level8Out32[27] , \Level8Out32[26] , 
        \Level8Out32[25] , \Level8Out32[24] , \Level8Out32[23] , 
        \Level8Out32[22] , \Level8Out32[21] , \Level8Out32[20] , 
        \Level8Out32[19] , \Level8Out32[18] , \Level8Out32[17] , 
        \Level8Out32[16] , \Level8Out32[15] , \Level8Out32[14] , 
        \Level8Out32[13] , \Level8Out32[12] , \Level8Out32[11] , 
        \Level8Out32[10] , \Level8Out32[9] , \Level8Out32[8] , 
        \Level8Out32[7] , \Level8Out32[6] , \Level8Out32[5] , \Level8Out32[4] , 
        \Level8Out32[3] , \Level8Out32[2] , \Level8Out32[1] , \Level8Out32[0] 
        }), .In2({\Level8Out40[31] , \Level8Out40[30] , \Level8Out40[29] , 
        \Level8Out40[28] , \Level8Out40[27] , \Level8Out40[26] , 
        \Level8Out40[25] , \Level8Out40[24] , \Level8Out40[23] , 
        \Level8Out40[22] , \Level8Out40[21] , \Level8Out40[20] , 
        \Level8Out40[19] , \Level8Out40[18] , \Level8Out40[17] , 
        \Level8Out40[16] , \Level8Out40[15] , \Level8Out40[14] , 
        \Level8Out40[13] , \Level8Out40[12] , \Level8Out40[11] , 
        \Level8Out40[10] , \Level8Out40[9] , \Level8Out40[8] , 
        \Level8Out40[7] , \Level8Out40[6] , \Level8Out40[5] , \Level8Out40[4] , 
        \Level8Out40[3] , \Level8Out40[2] , \Level8Out40[1] , \Level8Out40[0] 
        }), .Read1(\Level8Load32[0] ), .Read2(\Level8Load40[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_28_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load28[0] ), .Out({\Level4Out28[31] , \Level4Out28[30] , 
        \Level4Out28[29] , \Level4Out28[28] , \Level4Out28[27] , 
        \Level4Out28[26] , \Level4Out28[25] , \Level4Out28[24] , 
        \Level4Out28[23] , \Level4Out28[22] , \Level4Out28[21] , 
        \Level4Out28[20] , \Level4Out28[19] , \Level4Out28[18] , 
        \Level4Out28[17] , \Level4Out28[16] , \Level4Out28[15] , 
        \Level4Out28[14] , \Level4Out28[13] , \Level4Out28[12] , 
        \Level4Out28[11] , \Level4Out28[10] , \Level4Out28[9] , 
        \Level4Out28[8] , \Level4Out28[7] , \Level4Out28[6] , \Level4Out28[5] , 
        \Level4Out28[4] , \Level4Out28[3] , \Level4Out28[2] , \Level4Out28[1] , 
        \Level4Out28[0] }), .In1({\Level2Out28[31] , \Level2Out28[30] , 
        \Level2Out28[29] , \Level2Out28[28] , \Level2Out28[27] , 
        \Level2Out28[26] , \Level2Out28[25] , \Level2Out28[24] , 
        \Level2Out28[23] , \Level2Out28[22] , \Level2Out28[21] , 
        \Level2Out28[20] , \Level2Out28[19] , \Level2Out28[18] , 
        \Level2Out28[17] , \Level2Out28[16] , \Level2Out28[15] , 
        \Level2Out28[14] , \Level2Out28[13] , \Level2Out28[12] , 
        \Level2Out28[11] , \Level2Out28[10] , \Level2Out28[9] , 
        \Level2Out28[8] , \Level2Out28[7] , \Level2Out28[6] , \Level2Out28[5] , 
        \Level2Out28[4] , \Level2Out28[3] , \Level2Out28[2] , \Level2Out28[1] , 
        \Level2Out28[0] }), .In2({\Level2Out30[31] , \Level2Out30[30] , 
        \Level2Out30[29] , \Level2Out30[28] , \Level2Out30[27] , 
        \Level2Out30[26] , \Level2Out30[25] , \Level2Out30[24] , 
        \Level2Out30[23] , \Level2Out30[22] , \Level2Out30[21] , 
        \Level2Out30[20] , \Level2Out30[19] , \Level2Out30[18] , 
        \Level2Out30[17] , \Level2Out30[16] , \Level2Out30[15] , 
        \Level2Out30[14] , \Level2Out30[13] , \Level2Out30[12] , 
        \Level2Out30[11] , \Level2Out30[10] , \Level2Out30[9] , 
        \Level2Out30[8] , \Level2Out30[7] , \Level2Out30[6] , \Level2Out30[5] , 
        \Level2Out30[4] , \Level2Out30[3] , \Level2Out30[2] , \Level2Out30[1] , 
        \Level2Out30[0] }), .Read1(\Level2Load28[0] ), .Read2(
        \Level2Load30[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_58 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink58[31] , \ScanLink58[30] , 
        \ScanLink58[29] , \ScanLink58[28] , \ScanLink58[27] , \ScanLink58[26] , 
        \ScanLink58[25] , \ScanLink58[24] , \ScanLink58[23] , \ScanLink58[22] , 
        \ScanLink58[21] , \ScanLink58[20] , \ScanLink58[19] , \ScanLink58[18] , 
        \ScanLink58[17] , \ScanLink58[16] , \ScanLink58[15] , \ScanLink58[14] , 
        \ScanLink58[13] , \ScanLink58[12] , \ScanLink58[11] , \ScanLink58[10] , 
        \ScanLink58[9] , \ScanLink58[8] , \ScanLink58[7] , \ScanLink58[6] , 
        \ScanLink58[5] , \ScanLink58[4] , \ScanLink58[3] , \ScanLink58[2] , 
        \ScanLink58[1] , \ScanLink58[0] }), .ScanOut({\ScanLink59[31] , 
        \ScanLink59[30] , \ScanLink59[29] , \ScanLink59[28] , \ScanLink59[27] , 
        \ScanLink59[26] , \ScanLink59[25] , \ScanLink59[24] , \ScanLink59[23] , 
        \ScanLink59[22] , \ScanLink59[21] , \ScanLink59[20] , \ScanLink59[19] , 
        \ScanLink59[18] , \ScanLink59[17] , \ScanLink59[16] , \ScanLink59[15] , 
        \ScanLink59[14] , \ScanLink59[13] , \ScanLink59[12] , \ScanLink59[11] , 
        \ScanLink59[10] , \ScanLink59[9] , \ScanLink59[8] , \ScanLink59[7] , 
        \ScanLink59[6] , \ScanLink59[5] , \ScanLink59[4] , \ScanLink59[3] , 
        \ScanLink59[2] , \ScanLink59[1] , \ScanLink59[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load58[0] ), .Out({
        \Level1Out58[31] , \Level1Out58[30] , \Level1Out58[29] , 
        \Level1Out58[28] , \Level1Out58[27] , \Level1Out58[26] , 
        \Level1Out58[25] , \Level1Out58[24] , \Level1Out58[23] , 
        \Level1Out58[22] , \Level1Out58[21] , \Level1Out58[20] , 
        \Level1Out58[19] , \Level1Out58[18] , \Level1Out58[17] , 
        \Level1Out58[16] , \Level1Out58[15] , \Level1Out58[14] , 
        \Level1Out58[13] , \Level1Out58[12] , \Level1Out58[11] , 
        \Level1Out58[10] , \Level1Out58[9] , \Level1Out58[8] , 
        \Level1Out58[7] , \Level1Out58[6] , \Level1Out58[5] , \Level1Out58[4] , 
        \Level1Out58[3] , \Level1Out58[2] , \Level1Out58[1] , \Level1Out58[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_32_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load32[0] ), .Out({\Level8Out32[31] , \Level8Out32[30] , 
        \Level8Out32[29] , \Level8Out32[28] , \Level8Out32[27] , 
        \Level8Out32[26] , \Level8Out32[25] , \Level8Out32[24] , 
        \Level8Out32[23] , \Level8Out32[22] , \Level8Out32[21] , 
        \Level8Out32[20] , \Level8Out32[19] , \Level8Out32[18] , 
        \Level8Out32[17] , \Level8Out32[16] , \Level8Out32[15] , 
        \Level8Out32[14] , \Level8Out32[13] , \Level8Out32[12] , 
        \Level8Out32[11] , \Level8Out32[10] , \Level8Out32[9] , 
        \Level8Out32[8] , \Level8Out32[7] , \Level8Out32[6] , \Level8Out32[5] , 
        \Level8Out32[4] , \Level8Out32[3] , \Level8Out32[2] , \Level8Out32[1] , 
        \Level8Out32[0] }), .In1({\Level4Out32[31] , \Level4Out32[30] , 
        \Level4Out32[29] , \Level4Out32[28] , \Level4Out32[27] , 
        \Level4Out32[26] , \Level4Out32[25] , \Level4Out32[24] , 
        \Level4Out32[23] , \Level4Out32[22] , \Level4Out32[21] , 
        \Level4Out32[20] , \Level4Out32[19] , \Level4Out32[18] , 
        \Level4Out32[17] , \Level4Out32[16] , \Level4Out32[15] , 
        \Level4Out32[14] , \Level4Out32[13] , \Level4Out32[12] , 
        \Level4Out32[11] , \Level4Out32[10] , \Level4Out32[9] , 
        \Level4Out32[8] , \Level4Out32[7] , \Level4Out32[6] , \Level4Out32[5] , 
        \Level4Out32[4] , \Level4Out32[3] , \Level4Out32[2] , \Level4Out32[1] , 
        \Level4Out32[0] }), .In2({\Level4Out36[31] , \Level4Out36[30] , 
        \Level4Out36[29] , \Level4Out36[28] , \Level4Out36[27] , 
        \Level4Out36[26] , \Level4Out36[25] , \Level4Out36[24] , 
        \Level4Out36[23] , \Level4Out36[22] , \Level4Out36[21] , 
        \Level4Out36[20] , \Level4Out36[19] , \Level4Out36[18] , 
        \Level4Out36[17] , \Level4Out36[16] , \Level4Out36[15] , 
        \Level4Out36[14] , \Level4Out36[13] , \Level4Out36[12] , 
        \Level4Out36[11] , \Level4Out36[10] , \Level4Out36[9] , 
        \Level4Out36[8] , \Level4Out36[7] , \Level4Out36[6] , \Level4Out36[5] , 
        \Level4Out36[4] , \Level4Out36[3] , \Level4Out36[2] , \Level4Out36[1] , 
        \Level4Out36[0] }), .Read1(\Level4Load32[0] ), .Read2(
        \Level4Load36[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_24 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink24[31] , \ScanLink24[30] , 
        \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , \ScanLink24[26] , 
        \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , \ScanLink24[22] , 
        \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , \ScanLink24[18] , 
        \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , \ScanLink24[14] , 
        \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , \ScanLink24[10] , 
        \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , \ScanLink24[6] , 
        \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , \ScanLink24[2] , 
        \ScanLink24[1] , \ScanLink24[0] }), .ScanOut({\ScanLink25[31] , 
        \ScanLink25[30] , \ScanLink25[29] , \ScanLink25[28] , \ScanLink25[27] , 
        \ScanLink25[26] , \ScanLink25[25] , \ScanLink25[24] , \ScanLink25[23] , 
        \ScanLink25[22] , \ScanLink25[21] , \ScanLink25[20] , \ScanLink25[19] , 
        \ScanLink25[18] , \ScanLink25[17] , \ScanLink25[16] , \ScanLink25[15] , 
        \ScanLink25[14] , \ScanLink25[13] , \ScanLink25[12] , \ScanLink25[11] , 
        \ScanLink25[10] , \ScanLink25[9] , \ScanLink25[8] , \ScanLink25[7] , 
        \ScanLink25[6] , \ScanLink25[5] , \ScanLink25[4] , \ScanLink25[3] , 
        \ScanLink25[2] , \ScanLink25[1] , \ScanLink25[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load24[0] ), .Out({
        \Level1Out24[31] , \Level1Out24[30] , \Level1Out24[29] , 
        \Level1Out24[28] , \Level1Out24[27] , \Level1Out24[26] , 
        \Level1Out24[25] , \Level1Out24[24] , \Level1Out24[23] , 
        \Level1Out24[22] , \Level1Out24[21] , \Level1Out24[20] , 
        \Level1Out24[19] , \Level1Out24[18] , \Level1Out24[17] , 
        \Level1Out24[16] , \Level1Out24[15] , \Level1Out24[14] , 
        \Level1Out24[13] , \Level1Out24[12] , \Level1Out24[11] , 
        \Level1Out24[10] , \Level1Out24[9] , \Level1Out24[8] , 
        \Level1Out24[7] , \Level1Out24[6] , \Level1Out24[5] , \Level1Out24[4] , 
        \Level1Out24[3] , \Level1Out24[2] , \Level1Out24[1] , \Level1Out24[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_36 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink36[31] , \ScanLink36[30] , 
        \ScanLink36[29] , \ScanLink36[28] , \ScanLink36[27] , \ScanLink36[26] , 
        \ScanLink36[25] , \ScanLink36[24] , \ScanLink36[23] , \ScanLink36[22] , 
        \ScanLink36[21] , \ScanLink36[20] , \ScanLink36[19] , \ScanLink36[18] , 
        \ScanLink36[17] , \ScanLink36[16] , \ScanLink36[15] , \ScanLink36[14] , 
        \ScanLink36[13] , \ScanLink36[12] , \ScanLink36[11] , \ScanLink36[10] , 
        \ScanLink36[9] , \ScanLink36[8] , \ScanLink36[7] , \ScanLink36[6] , 
        \ScanLink36[5] , \ScanLink36[4] , \ScanLink36[3] , \ScanLink36[2] , 
        \ScanLink36[1] , \ScanLink36[0] }), .ScanOut({\ScanLink37[31] , 
        \ScanLink37[30] , \ScanLink37[29] , \ScanLink37[28] , \ScanLink37[27] , 
        \ScanLink37[26] , \ScanLink37[25] , \ScanLink37[24] , \ScanLink37[23] , 
        \ScanLink37[22] , \ScanLink37[21] , \ScanLink37[20] , \ScanLink37[19] , 
        \ScanLink37[18] , \ScanLink37[17] , \ScanLink37[16] , \ScanLink37[15] , 
        \ScanLink37[14] , \ScanLink37[13] , \ScanLink37[12] , \ScanLink37[11] , 
        \ScanLink37[10] , \ScanLink37[9] , \ScanLink37[8] , \ScanLink37[7] , 
        \ScanLink37[6] , \ScanLink37[5] , \ScanLink37[4] , \ScanLink37[3] , 
        \ScanLink37[2] , \ScanLink37[1] , \ScanLink37[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load36[0] ), .Out({
        \Level1Out36[31] , \Level1Out36[30] , \Level1Out36[29] , 
        \Level1Out36[28] , \Level1Out36[27] , \Level1Out36[26] , 
        \Level1Out36[25] , \Level1Out36[24] , \Level1Out36[23] , 
        \Level1Out36[22] , \Level1Out36[21] , \Level1Out36[20] , 
        \Level1Out36[19] , \Level1Out36[18] , \Level1Out36[17] , 
        \Level1Out36[16] , \Level1Out36[15] , \Level1Out36[14] , 
        \Level1Out36[13] , \Level1Out36[12] , \Level1Out36[11] , 
        \Level1Out36[10] , \Level1Out36[9] , \Level1Out36[8] , 
        \Level1Out36[7] , \Level1Out36[6] , \Level1Out36[5] , \Level1Out36[4] , 
        \Level1Out36[3] , \Level1Out36[2] , \Level1Out36[1] , \Level1Out36[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_48_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load48[0] ), .Out({\Level8Out48[31] , \Level8Out48[30] , 
        \Level8Out48[29] , \Level8Out48[28] , \Level8Out48[27] , 
        \Level8Out48[26] , \Level8Out48[25] , \Level8Out48[24] , 
        \Level8Out48[23] , \Level8Out48[22] , \Level8Out48[21] , 
        \Level8Out48[20] , \Level8Out48[19] , \Level8Out48[18] , 
        \Level8Out48[17] , \Level8Out48[16] , \Level8Out48[15] , 
        \Level8Out48[14] , \Level8Out48[13] , \Level8Out48[12] , 
        \Level8Out48[11] , \Level8Out48[10] , \Level8Out48[9] , 
        \Level8Out48[8] , \Level8Out48[7] , \Level8Out48[6] , \Level8Out48[5] , 
        \Level8Out48[4] , \Level8Out48[3] , \Level8Out48[2] , \Level8Out48[1] , 
        \Level8Out48[0] }), .In1({\Level4Out48[31] , \Level4Out48[30] , 
        \Level4Out48[29] , \Level4Out48[28] , \Level4Out48[27] , 
        \Level4Out48[26] , \Level4Out48[25] , \Level4Out48[24] , 
        \Level4Out48[23] , \Level4Out48[22] , \Level4Out48[21] , 
        \Level4Out48[20] , \Level4Out48[19] , \Level4Out48[18] , 
        \Level4Out48[17] , \Level4Out48[16] , \Level4Out48[15] , 
        \Level4Out48[14] , \Level4Out48[13] , \Level4Out48[12] , 
        \Level4Out48[11] , \Level4Out48[10] , \Level4Out48[9] , 
        \Level4Out48[8] , \Level4Out48[7] , \Level4Out48[6] , \Level4Out48[5] , 
        \Level4Out48[4] , \Level4Out48[3] , \Level4Out48[2] , \Level4Out48[1] , 
        \Level4Out48[0] }), .In2({\Level4Out52[31] , \Level4Out52[30] , 
        \Level4Out52[29] , \Level4Out52[28] , \Level4Out52[27] , 
        \Level4Out52[26] , \Level4Out52[25] , \Level4Out52[24] , 
        \Level4Out52[23] , \Level4Out52[22] , \Level4Out52[21] , 
        \Level4Out52[20] , \Level4Out52[19] , \Level4Out52[18] , 
        \Level4Out52[17] , \Level4Out52[16] , \Level4Out52[15] , 
        \Level4Out52[14] , \Level4Out52[13] , \Level4Out52[12] , 
        \Level4Out52[11] , \Level4Out52[10] , \Level4Out52[9] , 
        \Level4Out52[8] , \Level4Out52[7] , \Level4Out52[6] , \Level4Out52[5] , 
        \Level4Out52[4] , \Level4Out52[3] , \Level4Out52[2] , \Level4Out52[1] , 
        \Level4Out52[0] }), .Read1(\Level4Load48[0] ), .Read2(
        \Level4Load52[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_56_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load56[0] ), .Out({\Level2Out56[31] , \Level2Out56[30] , 
        \Level2Out56[29] , \Level2Out56[28] , \Level2Out56[27] , 
        \Level2Out56[26] , \Level2Out56[25] , \Level2Out56[24] , 
        \Level2Out56[23] , \Level2Out56[22] , \Level2Out56[21] , 
        \Level2Out56[20] , \Level2Out56[19] , \Level2Out56[18] , 
        \Level2Out56[17] , \Level2Out56[16] , \Level2Out56[15] , 
        \Level2Out56[14] , \Level2Out56[13] , \Level2Out56[12] , 
        \Level2Out56[11] , \Level2Out56[10] , \Level2Out56[9] , 
        \Level2Out56[8] , \Level2Out56[7] , \Level2Out56[6] , \Level2Out56[5] , 
        \Level2Out56[4] , \Level2Out56[3] , \Level2Out56[2] , \Level2Out56[1] , 
        \Level2Out56[0] }), .In1({\Level1Out56[31] , \Level1Out56[30] , 
        \Level1Out56[29] , \Level1Out56[28] , \Level1Out56[27] , 
        \Level1Out56[26] , \Level1Out56[25] , \Level1Out56[24] , 
        \Level1Out56[23] , \Level1Out56[22] , \Level1Out56[21] , 
        \Level1Out56[20] , \Level1Out56[19] , \Level1Out56[18] , 
        \Level1Out56[17] , \Level1Out56[16] , \Level1Out56[15] , 
        \Level1Out56[14] , \Level1Out56[13] , \Level1Out56[12] , 
        \Level1Out56[11] , \Level1Out56[10] , \Level1Out56[9] , 
        \Level1Out56[8] , \Level1Out56[7] , \Level1Out56[6] , \Level1Out56[5] , 
        \Level1Out56[4] , \Level1Out56[3] , \Level1Out56[2] , \Level1Out56[1] , 
        \Level1Out56[0] }), .In2({\Level1Out57[31] , \Level1Out57[30] , 
        \Level1Out57[29] , \Level1Out57[28] , \Level1Out57[27] , 
        \Level1Out57[26] , \Level1Out57[25] , \Level1Out57[24] , 
        \Level1Out57[23] , \Level1Out57[22] , \Level1Out57[21] , 
        \Level1Out57[20] , \Level1Out57[19] , \Level1Out57[18] , 
        \Level1Out57[17] , \Level1Out57[16] , \Level1Out57[15] , 
        \Level1Out57[14] , \Level1Out57[13] , \Level1Out57[12] , 
        \Level1Out57[11] , \Level1Out57[10] , \Level1Out57[9] , 
        \Level1Out57[8] , \Level1Out57[7] , \Level1Out57[6] , \Level1Out57[5] , 
        \Level1Out57[4] , \Level1Out57[3] , \Level1Out57[2] , \Level1Out57[1] , 
        \Level1Out57[0] }), .Read1(\Level1Load56[0] ), .Read2(
        \Level1Load57[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_60_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load60[0] ), .Out({\Level4Out60[31] , \Level4Out60[30] , 
        \Level4Out60[29] , \Level4Out60[28] , \Level4Out60[27] , 
        \Level4Out60[26] , \Level4Out60[25] , \Level4Out60[24] , 
        \Level4Out60[23] , \Level4Out60[22] , \Level4Out60[21] , 
        \Level4Out60[20] , \Level4Out60[19] , \Level4Out60[18] , 
        \Level4Out60[17] , \Level4Out60[16] , \Level4Out60[15] , 
        \Level4Out60[14] , \Level4Out60[13] , \Level4Out60[12] , 
        \Level4Out60[11] , \Level4Out60[10] , \Level4Out60[9] , 
        \Level4Out60[8] , \Level4Out60[7] , \Level4Out60[6] , \Level4Out60[5] , 
        \Level4Out60[4] , \Level4Out60[3] , \Level4Out60[2] , \Level4Out60[1] , 
        \Level4Out60[0] }), .In1({\Level2Out60[31] , \Level2Out60[30] , 
        \Level2Out60[29] , \Level2Out60[28] , \Level2Out60[27] , 
        \Level2Out60[26] , \Level2Out60[25] , \Level2Out60[24] , 
        \Level2Out60[23] , \Level2Out60[22] , \Level2Out60[21] , 
        \Level2Out60[20] , \Level2Out60[19] , \Level2Out60[18] , 
        \Level2Out60[17] , \Level2Out60[16] , \Level2Out60[15] , 
        \Level2Out60[14] , \Level2Out60[13] , \Level2Out60[12] , 
        \Level2Out60[11] , \Level2Out60[10] , \Level2Out60[9] , 
        \Level2Out60[8] , \Level2Out60[7] , \Level2Out60[6] , \Level2Out60[5] , 
        \Level2Out60[4] , \Level2Out60[3] , \Level2Out60[2] , \Level2Out60[1] , 
        \Level2Out60[0] }), .In2({\Level2Out62[31] , \Level2Out62[30] , 
        \Level2Out62[29] , \Level2Out62[28] , \Level2Out62[27] , 
        \Level2Out62[26] , \Level2Out62[25] , \Level2Out62[24] , 
        \Level2Out62[23] , \Level2Out62[22] , \Level2Out62[21] , 
        \Level2Out62[20] , \Level2Out62[19] , \Level2Out62[18] , 
        \Level2Out62[17] , \Level2Out62[16] , \Level2Out62[15] , 
        \Level2Out62[14] , \Level2Out62[13] , \Level2Out62[12] , 
        \Level2Out62[11] , \Level2Out62[10] , \Level2Out62[9] , 
        \Level2Out62[8] , \Level2Out62[7] , \Level2Out62[6] , \Level2Out62[5] , 
        \Level2Out62[4] , \Level2Out62[3] , \Level2Out62[2] , \Level2Out62[1] , 
        \Level2Out62[0] }), .Read1(\Level2Load60[0] ), .Read2(
        \Level2Load62[0] ) );
    Merge_Top_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Top_Node ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink64[31] , \ScanLink64[30] , 
        \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , \ScanLink64[26] , 
        \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , \ScanLink64[22] , 
        \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , \ScanLink64[18] , 
        \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , \ScanLink64[14] , 
        \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , \ScanLink64[10] , 
        \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , \ScanLink64[6] , 
        \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , \ScanLink64[2] , 
        \ScanLink64[1] , \ScanLink64[0] }), .ScanOut({\ScanLink0[31] , 
        \ScanLink0[30] , \ScanLink0[29] , \ScanLink0[28] , \ScanLink0[27] , 
        \ScanLink0[26] , \ScanLink0[25] , \ScanLink0[24] , \ScanLink0[23] , 
        \ScanLink0[22] , \ScanLink0[21] , \ScanLink0[20] , \ScanLink0[19] , 
        \ScanLink0[18] , \ScanLink0[17] , \ScanLink0[16] , \ScanLink0[15] , 
        \ScanLink0[14] , \ScanLink0[13] , \ScanLink0[12] , \ScanLink0[11] , 
        \ScanLink0[10] , \ScanLink0[9] , \ScanLink0[8] , \ScanLink0[7] , 
        \ScanLink0[6] , \ScanLink0[5] , \ScanLink0[4] , \ScanLink0[3] , 
        \ScanLink0[2] , \ScanLink0[1] , \ScanLink0[0] }), .ScanEnable(
        \ScanEnable[0] ), .ScanId(1'b0), .Id(1'b1), .In1({\Level32Out0[31] , 
        \Level32Out0[30] , \Level32Out0[29] , \Level32Out0[28] , 
        \Level32Out0[27] , \Level32Out0[26] , \Level32Out0[25] , 
        \Level32Out0[24] , \Level32Out0[23] , \Level32Out0[22] , 
        \Level32Out0[21] , \Level32Out0[20] , \Level32Out0[19] , 
        \Level32Out0[18] , \Level32Out0[17] , \Level32Out0[16] , 
        \Level32Out0[15] , \Level32Out0[14] , \Level32Out0[13] , 
        \Level32Out0[12] , \Level32Out0[11] , \Level32Out0[10] , 
        \Level32Out0[9] , \Level32Out0[8] , \Level32Out0[7] , \Level32Out0[6] , 
        \Level32Out0[5] , \Level32Out0[4] , \Level32Out0[3] , \Level32Out0[2] , 
        \Level32Out0[1] , \Level32Out0[0] }), .In2({\Level32Out32[31] , 
        \Level32Out32[30] , \Level32Out32[29] , \Level32Out32[28] , 
        \Level32Out32[27] , \Level32Out32[26] , \Level32Out32[25] , 
        \Level32Out32[24] , \Level32Out32[23] , \Level32Out32[22] , 
        \Level32Out32[21] , \Level32Out32[20] , \Level32Out32[19] , 
        \Level32Out32[18] , \Level32Out32[17] , \Level32Out32[16] , 
        \Level32Out32[15] , \Level32Out32[14] , \Level32Out32[13] , 
        \Level32Out32[12] , \Level32Out32[11] , \Level32Out32[10] , 
        \Level32Out32[9] , \Level32Out32[8] , \Level32Out32[7] , 
        \Level32Out32[6] , \Level32Out32[5] , \Level32Out32[4] , 
        \Level32Out32[3] , \Level32Out32[2] , \Level32Out32[1] , 
        \Level32Out32[0] }), .Read1(\Level32Load0[0] ), .Read2(
        \Level32Load32[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_18 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink18[31] , \ScanLink18[30] , 
        \ScanLink18[29] , \ScanLink18[28] , \ScanLink18[27] , \ScanLink18[26] , 
        \ScanLink18[25] , \ScanLink18[24] , \ScanLink18[23] , \ScanLink18[22] , 
        \ScanLink18[21] , \ScanLink18[20] , \ScanLink18[19] , \ScanLink18[18] , 
        \ScanLink18[17] , \ScanLink18[16] , \ScanLink18[15] , \ScanLink18[14] , 
        \ScanLink18[13] , \ScanLink18[12] , \ScanLink18[11] , \ScanLink18[10] , 
        \ScanLink18[9] , \ScanLink18[8] , \ScanLink18[7] , \ScanLink18[6] , 
        \ScanLink18[5] , \ScanLink18[4] , \ScanLink18[3] , \ScanLink18[2] , 
        \ScanLink18[1] , \ScanLink18[0] }), .ScanOut({\ScanLink19[31] , 
        \ScanLink19[30] , \ScanLink19[29] , \ScanLink19[28] , \ScanLink19[27] , 
        \ScanLink19[26] , \ScanLink19[25] , \ScanLink19[24] , \ScanLink19[23] , 
        \ScanLink19[22] , \ScanLink19[21] , \ScanLink19[20] , \ScanLink19[19] , 
        \ScanLink19[18] , \ScanLink19[17] , \ScanLink19[16] , \ScanLink19[15] , 
        \ScanLink19[14] , \ScanLink19[13] , \ScanLink19[12] , \ScanLink19[11] , 
        \ScanLink19[10] , \ScanLink19[9] , \ScanLink19[8] , \ScanLink19[7] , 
        \ScanLink19[6] , \ScanLink19[5] , \ScanLink19[4] , \ScanLink19[3] , 
        \ScanLink19[2] , \ScanLink19[1] , \ScanLink19[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load18[0] ), .Out({
        \Level1Out18[31] , \Level1Out18[30] , \Level1Out18[29] , 
        \Level1Out18[28] , \Level1Out18[27] , \Level1Out18[26] , 
        \Level1Out18[25] , \Level1Out18[24] , \Level1Out18[23] , 
        \Level1Out18[22] , \Level1Out18[21] , \Level1Out18[20] , 
        \Level1Out18[19] , \Level1Out18[18] , \Level1Out18[17] , 
        \Level1Out18[16] , \Level1Out18[15] , \Level1Out18[14] , 
        \Level1Out18[13] , \Level1Out18[12] , \Level1Out18[11] , 
        \Level1Out18[10] , \Level1Out18[9] , \Level1Out18[8] , 
        \Level1Out18[7] , \Level1Out18[6] , \Level1Out18[5] , \Level1Out18[4] , 
        \Level1Out18[3] , \Level1Out18[2] , \Level1Out18[1] , \Level1Out18[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_51 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink51[31] , \ScanLink51[30] , 
        \ScanLink51[29] , \ScanLink51[28] , \ScanLink51[27] , \ScanLink51[26] , 
        \ScanLink51[25] , \ScanLink51[24] , \ScanLink51[23] , \ScanLink51[22] , 
        \ScanLink51[21] , \ScanLink51[20] , \ScanLink51[19] , \ScanLink51[18] , 
        \ScanLink51[17] , \ScanLink51[16] , \ScanLink51[15] , \ScanLink51[14] , 
        \ScanLink51[13] , \ScanLink51[12] , \ScanLink51[11] , \ScanLink51[10] , 
        \ScanLink51[9] , \ScanLink51[8] , \ScanLink51[7] , \ScanLink51[6] , 
        \ScanLink51[5] , \ScanLink51[4] , \ScanLink51[3] , \ScanLink51[2] , 
        \ScanLink51[1] , \ScanLink51[0] }), .ScanOut({\ScanLink52[31] , 
        \ScanLink52[30] , \ScanLink52[29] , \ScanLink52[28] , \ScanLink52[27] , 
        \ScanLink52[26] , \ScanLink52[25] , \ScanLink52[24] , \ScanLink52[23] , 
        \ScanLink52[22] , \ScanLink52[21] , \ScanLink52[20] , \ScanLink52[19] , 
        \ScanLink52[18] , \ScanLink52[17] , \ScanLink52[16] , \ScanLink52[15] , 
        \ScanLink52[14] , \ScanLink52[13] , \ScanLink52[12] , \ScanLink52[11] , 
        \ScanLink52[10] , \ScanLink52[9] , \ScanLink52[8] , \ScanLink52[7] , 
        \ScanLink52[6] , \ScanLink52[5] , \ScanLink52[4] , \ScanLink52[3] , 
        \ScanLink52[2] , \ScanLink52[1] , \ScanLink52[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load51[0] ), .Out({
        \Level1Out51[31] , \Level1Out51[30] , \Level1Out51[29] , 
        \Level1Out51[28] , \Level1Out51[27] , \Level1Out51[26] , 
        \Level1Out51[25] , \Level1Out51[24] , \Level1Out51[23] , 
        \Level1Out51[22] , \Level1Out51[21] , \Level1Out51[20] , 
        \Level1Out51[19] , \Level1Out51[18] , \Level1Out51[17] , 
        \Level1Out51[16] , \Level1Out51[15] , \Level1Out51[14] , 
        \Level1Out51[13] , \Level1Out51[12] , \Level1Out51[11] , 
        \Level1Out51[10] , \Level1Out51[9] , \Level1Out51[8] , 
        \Level1Out51[7] , \Level1Out51[6] , \Level1Out51[5] , \Level1Out51[4] , 
        \Level1Out51[3] , \Level1Out51[2] , \Level1Out51[1] , \Level1Out51[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_8_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level8Load8[0] ), .Out({\Level8Out8[31] , \Level8Out8[30] , 
        \Level8Out8[29] , \Level8Out8[28] , \Level8Out8[27] , \Level8Out8[26] , 
        \Level8Out8[25] , \Level8Out8[24] , \Level8Out8[23] , \Level8Out8[22] , 
        \Level8Out8[21] , \Level8Out8[20] , \Level8Out8[19] , \Level8Out8[18] , 
        \Level8Out8[17] , \Level8Out8[16] , \Level8Out8[15] , \Level8Out8[14] , 
        \Level8Out8[13] , \Level8Out8[12] , \Level8Out8[11] , \Level8Out8[10] , 
        \Level8Out8[9] , \Level8Out8[8] , \Level8Out8[7] , \Level8Out8[6] , 
        \Level8Out8[5] , \Level8Out8[4] , \Level8Out8[3] , \Level8Out8[2] , 
        \Level8Out8[1] , \Level8Out8[0] }), .In1({\Level4Out8[31] , 
        \Level4Out8[30] , \Level4Out8[29] , \Level4Out8[28] , \Level4Out8[27] , 
        \Level4Out8[26] , \Level4Out8[25] , \Level4Out8[24] , \Level4Out8[23] , 
        \Level4Out8[22] , \Level4Out8[21] , \Level4Out8[20] , \Level4Out8[19] , 
        \Level4Out8[18] , \Level4Out8[17] , \Level4Out8[16] , \Level4Out8[15] , 
        \Level4Out8[14] , \Level4Out8[13] , \Level4Out8[12] , \Level4Out8[11] , 
        \Level4Out8[10] , \Level4Out8[9] , \Level4Out8[8] , \Level4Out8[7] , 
        \Level4Out8[6] , \Level4Out8[5] , \Level4Out8[4] , \Level4Out8[3] , 
        \Level4Out8[2] , \Level4Out8[1] , \Level4Out8[0] }), .In2({
        \Level4Out12[31] , \Level4Out12[30] , \Level4Out12[29] , 
        \Level4Out12[28] , \Level4Out12[27] , \Level4Out12[26] , 
        \Level4Out12[25] , \Level4Out12[24] , \Level4Out12[23] , 
        \Level4Out12[22] , \Level4Out12[21] , \Level4Out12[20] , 
        \Level4Out12[19] , \Level4Out12[18] , \Level4Out12[17] , 
        \Level4Out12[16] , \Level4Out12[15] , \Level4Out12[14] , 
        \Level4Out12[13] , \Level4Out12[12] , \Level4Out12[11] , 
        \Level4Out12[10] , \Level4Out12[9] , \Level4Out12[8] , 
        \Level4Out12[7] , \Level4Out12[6] , \Level4Out12[5] , \Level4Out12[4] , 
        \Level4Out12[3] , \Level4Out12[2] , \Level4Out12[1] , \Level4Out12[0] 
        }), .Read1(\Level4Load8[0] ), .Read2(\Level4Load12[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_52_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load52[0] ), .Out({\Level4Out52[31] , \Level4Out52[30] , 
        \Level4Out52[29] , \Level4Out52[28] , \Level4Out52[27] , 
        \Level4Out52[26] , \Level4Out52[25] , \Level4Out52[24] , 
        \Level4Out52[23] , \Level4Out52[22] , \Level4Out52[21] , 
        \Level4Out52[20] , \Level4Out52[19] , \Level4Out52[18] , 
        \Level4Out52[17] , \Level4Out52[16] , \Level4Out52[15] , 
        \Level4Out52[14] , \Level4Out52[13] , \Level4Out52[12] , 
        \Level4Out52[11] , \Level4Out52[10] , \Level4Out52[9] , 
        \Level4Out52[8] , \Level4Out52[7] , \Level4Out52[6] , \Level4Out52[5] , 
        \Level4Out52[4] , \Level4Out52[3] , \Level4Out52[2] , \Level4Out52[1] , 
        \Level4Out52[0] }), .In1({\Level2Out52[31] , \Level2Out52[30] , 
        \Level2Out52[29] , \Level2Out52[28] , \Level2Out52[27] , 
        \Level2Out52[26] , \Level2Out52[25] , \Level2Out52[24] , 
        \Level2Out52[23] , \Level2Out52[22] , \Level2Out52[21] , 
        \Level2Out52[20] , \Level2Out52[19] , \Level2Out52[18] , 
        \Level2Out52[17] , \Level2Out52[16] , \Level2Out52[15] , 
        \Level2Out52[14] , \Level2Out52[13] , \Level2Out52[12] , 
        \Level2Out52[11] , \Level2Out52[10] , \Level2Out52[9] , 
        \Level2Out52[8] , \Level2Out52[7] , \Level2Out52[6] , \Level2Out52[5] , 
        \Level2Out52[4] , \Level2Out52[3] , \Level2Out52[2] , \Level2Out52[1] , 
        \Level2Out52[0] }), .In2({\Level2Out54[31] , \Level2Out54[30] , 
        \Level2Out54[29] , \Level2Out54[28] , \Level2Out54[27] , 
        \Level2Out54[26] , \Level2Out54[25] , \Level2Out54[24] , 
        \Level2Out54[23] , \Level2Out54[22] , \Level2Out54[21] , 
        \Level2Out54[20] , \Level2Out54[19] , \Level2Out54[18] , 
        \Level2Out54[17] , \Level2Out54[16] , \Level2Out54[15] , 
        \Level2Out54[14] , \Level2Out54[13] , \Level2Out54[12] , 
        \Level2Out54[11] , \Level2Out54[10] , \Level2Out54[9] , 
        \Level2Out54[8] , \Level2Out54[7] , \Level2Out54[6] , \Level2Out54[5] , 
        \Level2Out54[4] , \Level2Out54[3] , \Level2Out54[2] , \Level2Out54[1] , 
        \Level2Out54[0] }), .Read1(\Level2Load52[0] ), .Read2(
        \Level2Load54[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_38 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink38[31] , \ScanLink38[30] , 
        \ScanLink38[29] , \ScanLink38[28] , \ScanLink38[27] , \ScanLink38[26] , 
        \ScanLink38[25] , \ScanLink38[24] , \ScanLink38[23] , \ScanLink38[22] , 
        \ScanLink38[21] , \ScanLink38[20] , \ScanLink38[19] , \ScanLink38[18] , 
        \ScanLink38[17] , \ScanLink38[16] , \ScanLink38[15] , \ScanLink38[14] , 
        \ScanLink38[13] , \ScanLink38[12] , \ScanLink38[11] , \ScanLink38[10] , 
        \ScanLink38[9] , \ScanLink38[8] , \ScanLink38[7] , \ScanLink38[6] , 
        \ScanLink38[5] , \ScanLink38[4] , \ScanLink38[3] , \ScanLink38[2] , 
        \ScanLink38[1] , \ScanLink38[0] }), .ScanOut({\ScanLink39[31] , 
        \ScanLink39[30] , \ScanLink39[29] , \ScanLink39[28] , \ScanLink39[27] , 
        \ScanLink39[26] , \ScanLink39[25] , \ScanLink39[24] , \ScanLink39[23] , 
        \ScanLink39[22] , \ScanLink39[21] , \ScanLink39[20] , \ScanLink39[19] , 
        \ScanLink39[18] , \ScanLink39[17] , \ScanLink39[16] , \ScanLink39[15] , 
        \ScanLink39[14] , \ScanLink39[13] , \ScanLink39[12] , \ScanLink39[11] , 
        \ScanLink39[10] , \ScanLink39[9] , \ScanLink39[8] , \ScanLink39[7] , 
        \ScanLink39[6] , \ScanLink39[5] , \ScanLink39[4] , \ScanLink39[3] , 
        \ScanLink39[2] , \ScanLink39[1] , \ScanLink39[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load38[0] ), .Out({
        \Level1Out38[31] , \Level1Out38[30] , \Level1Out38[29] , 
        \Level1Out38[28] , \Level1Out38[27] , \Level1Out38[26] , 
        \Level1Out38[25] , \Level1Out38[24] , \Level1Out38[23] , 
        \Level1Out38[22] , \Level1Out38[21] , \Level1Out38[20] , 
        \Level1Out38[19] , \Level1Out38[18] , \Level1Out38[17] , 
        \Level1Out38[16] , \Level1Out38[15] , \Level1Out38[14] , 
        \Level1Out38[13] , \Level1Out38[12] , \Level1Out38[11] , 
        \Level1Out38[10] , \Level1Out38[9] , \Level1Out38[8] , 
        \Level1Out38[7] , \Level1Out38[6] , \Level1Out38[5] , \Level1Out38[4] , 
        \Level1Out38[3] , \Level1Out38[2] , \Level1Out38[1] , \Level1Out38[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_56 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink56[31] , \ScanLink56[30] , 
        \ScanLink56[29] , \ScanLink56[28] , \ScanLink56[27] , \ScanLink56[26] , 
        \ScanLink56[25] , \ScanLink56[24] , \ScanLink56[23] , \ScanLink56[22] , 
        \ScanLink56[21] , \ScanLink56[20] , \ScanLink56[19] , \ScanLink56[18] , 
        \ScanLink56[17] , \ScanLink56[16] , \ScanLink56[15] , \ScanLink56[14] , 
        \ScanLink56[13] , \ScanLink56[12] , \ScanLink56[11] , \ScanLink56[10] , 
        \ScanLink56[9] , \ScanLink56[8] , \ScanLink56[7] , \ScanLink56[6] , 
        \ScanLink56[5] , \ScanLink56[4] , \ScanLink56[3] , \ScanLink56[2] , 
        \ScanLink56[1] , \ScanLink56[0] }), .ScanOut({\ScanLink57[31] , 
        \ScanLink57[30] , \ScanLink57[29] , \ScanLink57[28] , \ScanLink57[27] , 
        \ScanLink57[26] , \ScanLink57[25] , \ScanLink57[24] , \ScanLink57[23] , 
        \ScanLink57[22] , \ScanLink57[21] , \ScanLink57[20] , \ScanLink57[19] , 
        \ScanLink57[18] , \ScanLink57[17] , \ScanLink57[16] , \ScanLink57[15] , 
        \ScanLink57[14] , \ScanLink57[13] , \ScanLink57[12] , \ScanLink57[11] , 
        \ScanLink57[10] , \ScanLink57[9] , \ScanLink57[8] , \ScanLink57[7] , 
        \ScanLink57[6] , \ScanLink57[5] , \ScanLink57[4] , \ScanLink57[3] , 
        \ScanLink57[2] , \ScanLink57[1] , \ScanLink57[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load56[0] ), .Out({
        \Level1Out56[31] , \Level1Out56[30] , \Level1Out56[29] , 
        \Level1Out56[28] , \Level1Out56[27] , \Level1Out56[26] , 
        \Level1Out56[25] , \Level1Out56[24] , \Level1Out56[23] , 
        \Level1Out56[22] , \Level1Out56[21] , \Level1Out56[20] , 
        \Level1Out56[19] , \Level1Out56[18] , \Level1Out56[17] , 
        \Level1Out56[16] , \Level1Out56[15] , \Level1Out56[14] , 
        \Level1Out56[13] , \Level1Out56[12] , \Level1Out56[11] , 
        \Level1Out56[10] , \Level1Out56[9] , \Level1Out56[8] , 
        \Level1Out56[7] , \Level1Out56[6] , \Level1Out56[5] , \Level1Out56[4] , 
        \Level1Out56[3] , \Level1Out56[2] , \Level1Out56[1] , \Level1Out56[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load2[0] ), .Out({\Level2Out2[31] , \Level2Out2[30] , 
        \Level2Out2[29] , \Level2Out2[28] , \Level2Out2[27] , \Level2Out2[26] , 
        \Level2Out2[25] , \Level2Out2[24] , \Level2Out2[23] , \Level2Out2[22] , 
        \Level2Out2[21] , \Level2Out2[20] , \Level2Out2[19] , \Level2Out2[18] , 
        \Level2Out2[17] , \Level2Out2[16] , \Level2Out2[15] , \Level2Out2[14] , 
        \Level2Out2[13] , \Level2Out2[12] , \Level2Out2[11] , \Level2Out2[10] , 
        \Level2Out2[9] , \Level2Out2[8] , \Level2Out2[7] , \Level2Out2[6] , 
        \Level2Out2[5] , \Level2Out2[4] , \Level2Out2[3] , \Level2Out2[2] , 
        \Level2Out2[1] , \Level2Out2[0] }), .In1({\Level1Out2[31] , 
        \Level1Out2[30] , \Level1Out2[29] , \Level1Out2[28] , \Level1Out2[27] , 
        \Level1Out2[26] , \Level1Out2[25] , \Level1Out2[24] , \Level1Out2[23] , 
        \Level1Out2[22] , \Level1Out2[21] , \Level1Out2[20] , \Level1Out2[19] , 
        \Level1Out2[18] , \Level1Out2[17] , \Level1Out2[16] , \Level1Out2[15] , 
        \Level1Out2[14] , \Level1Out2[13] , \Level1Out2[12] , \Level1Out2[11] , 
        \Level1Out2[10] , \Level1Out2[9] , \Level1Out2[8] , \Level1Out2[7] , 
        \Level1Out2[6] , \Level1Out2[5] , \Level1Out2[4] , \Level1Out2[3] , 
        \Level1Out2[2] , \Level1Out2[1] , \Level1Out2[0] }), .In2({
        \Level1Out3[31] , \Level1Out3[30] , \Level1Out3[29] , \Level1Out3[28] , 
        \Level1Out3[27] , \Level1Out3[26] , \Level1Out3[25] , \Level1Out3[24] , 
        \Level1Out3[23] , \Level1Out3[22] , \Level1Out3[21] , \Level1Out3[20] , 
        \Level1Out3[19] , \Level1Out3[18] , \Level1Out3[17] , \Level1Out3[16] , 
        \Level1Out3[15] , \Level1Out3[14] , \Level1Out3[13] , \Level1Out3[12] , 
        \Level1Out3[11] , \Level1Out3[10] , \Level1Out3[9] , \Level1Out3[8] , 
        \Level1Out3[7] , \Level1Out3[6] , \Level1Out3[5] , \Level1Out3[4] , 
        \Level1Out3[3] , \Level1Out3[2] , \Level1Out3[1] , \Level1Out3[0] }), 
        .Read1(\Level1Load2[0] ), .Read2(\Level1Load3[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_16 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink16[31] , \ScanLink16[30] , 
        \ScanLink16[29] , \ScanLink16[28] , \ScanLink16[27] , \ScanLink16[26] , 
        \ScanLink16[25] , \ScanLink16[24] , \ScanLink16[23] , \ScanLink16[22] , 
        \ScanLink16[21] , \ScanLink16[20] , \ScanLink16[19] , \ScanLink16[18] , 
        \ScanLink16[17] , \ScanLink16[16] , \ScanLink16[15] , \ScanLink16[14] , 
        \ScanLink16[13] , \ScanLink16[12] , \ScanLink16[11] , \ScanLink16[10] , 
        \ScanLink16[9] , \ScanLink16[8] , \ScanLink16[7] , \ScanLink16[6] , 
        \ScanLink16[5] , \ScanLink16[4] , \ScanLink16[3] , \ScanLink16[2] , 
        \ScanLink16[1] , \ScanLink16[0] }), .ScanOut({\ScanLink17[31] , 
        \ScanLink17[30] , \ScanLink17[29] , \ScanLink17[28] , \ScanLink17[27] , 
        \ScanLink17[26] , \ScanLink17[25] , \ScanLink17[24] , \ScanLink17[23] , 
        \ScanLink17[22] , \ScanLink17[21] , \ScanLink17[20] , \ScanLink17[19] , 
        \ScanLink17[18] , \ScanLink17[17] , \ScanLink17[16] , \ScanLink17[15] , 
        \ScanLink17[14] , \ScanLink17[13] , \ScanLink17[12] , \ScanLink17[11] , 
        \ScanLink17[10] , \ScanLink17[9] , \ScanLink17[8] , \ScanLink17[7] , 
        \ScanLink17[6] , \ScanLink17[5] , \ScanLink17[4] , \ScanLink17[3] , 
        \ScanLink17[2] , \ScanLink17[1] , \ScanLink17[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load16[0] ), .Out({
        \Level1Out16[31] , \Level1Out16[30] , \Level1Out16[29] , 
        \Level1Out16[28] , \Level1Out16[27] , \Level1Out16[26] , 
        \Level1Out16[25] , \Level1Out16[24] , \Level1Out16[23] , 
        \Level1Out16[22] , \Level1Out16[21] , \Level1Out16[20] , 
        \Level1Out16[19] , \Level1Out16[18] , \Level1Out16[17] , 
        \Level1Out16[16] , \Level1Out16[15] , \Level1Out16[14] , 
        \Level1Out16[13] , \Level1Out16[12] , \Level1Out16[11] , 
        \Level1Out16[10] , \Level1Out16[9] , \Level1Out16[8] , 
        \Level1Out16[7] , \Level1Out16[6] , \Level1Out16[5] , \Level1Out16[4] , 
        \Level1Out16[3] , \Level1Out16[2] , \Level1Out16[1] , \Level1Out16[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_23 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink23[31] , \ScanLink23[30] , 
        \ScanLink23[29] , \ScanLink23[28] , \ScanLink23[27] , \ScanLink23[26] , 
        \ScanLink23[25] , \ScanLink23[24] , \ScanLink23[23] , \ScanLink23[22] , 
        \ScanLink23[21] , \ScanLink23[20] , \ScanLink23[19] , \ScanLink23[18] , 
        \ScanLink23[17] , \ScanLink23[16] , \ScanLink23[15] , \ScanLink23[14] , 
        \ScanLink23[13] , \ScanLink23[12] , \ScanLink23[11] , \ScanLink23[10] , 
        \ScanLink23[9] , \ScanLink23[8] , \ScanLink23[7] , \ScanLink23[6] , 
        \ScanLink23[5] , \ScanLink23[4] , \ScanLink23[3] , \ScanLink23[2] , 
        \ScanLink23[1] , \ScanLink23[0] }), .ScanOut({\ScanLink24[31] , 
        \ScanLink24[30] , \ScanLink24[29] , \ScanLink24[28] , \ScanLink24[27] , 
        \ScanLink24[26] , \ScanLink24[25] , \ScanLink24[24] , \ScanLink24[23] , 
        \ScanLink24[22] , \ScanLink24[21] , \ScanLink24[20] , \ScanLink24[19] , 
        \ScanLink24[18] , \ScanLink24[17] , \ScanLink24[16] , \ScanLink24[15] , 
        \ScanLink24[14] , \ScanLink24[13] , \ScanLink24[12] , \ScanLink24[11] , 
        \ScanLink24[10] , \ScanLink24[9] , \ScanLink24[8] , \ScanLink24[7] , 
        \ScanLink24[6] , \ScanLink24[5] , \ScanLink24[4] , \ScanLink24[3] , 
        \ScanLink24[2] , \ScanLink24[1] , \ScanLink24[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load23[0] ), .Out({
        \Level1Out23[31] , \Level1Out23[30] , \Level1Out23[29] , 
        \Level1Out23[28] , \Level1Out23[27] , \Level1Out23[26] , 
        \Level1Out23[25] , \Level1Out23[24] , \Level1Out23[23] , 
        \Level1Out23[22] , \Level1Out23[21] , \Level1Out23[20] , 
        \Level1Out23[19] , \Level1Out23[18] , \Level1Out23[17] , 
        \Level1Out23[16] , \Level1Out23[15] , \Level1Out23[14] , 
        \Level1Out23[13] , \Level1Out23[12] , \Level1Out23[11] , 
        \Level1Out23[10] , \Level1Out23[9] , \Level1Out23[8] , 
        \Level1Out23[7] , \Level1Out23[6] , \Level1Out23[5] , \Level1Out23[4] , 
        \Level1Out23[3] , \Level1Out23[2] , \Level1Out23[1] , \Level1Out23[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_42_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load42[0] ), .Out({\Level2Out42[31] , \Level2Out42[30] , 
        \Level2Out42[29] , \Level2Out42[28] , \Level2Out42[27] , 
        \Level2Out42[26] , \Level2Out42[25] , \Level2Out42[24] , 
        \Level2Out42[23] , \Level2Out42[22] , \Level2Out42[21] , 
        \Level2Out42[20] , \Level2Out42[19] , \Level2Out42[18] , 
        \Level2Out42[17] , \Level2Out42[16] , \Level2Out42[15] , 
        \Level2Out42[14] , \Level2Out42[13] , \Level2Out42[12] , 
        \Level2Out42[11] , \Level2Out42[10] , \Level2Out42[9] , 
        \Level2Out42[8] , \Level2Out42[7] , \Level2Out42[6] , \Level2Out42[5] , 
        \Level2Out42[4] , \Level2Out42[3] , \Level2Out42[2] , \Level2Out42[1] , 
        \Level2Out42[0] }), .In1({\Level1Out42[31] , \Level1Out42[30] , 
        \Level1Out42[29] , \Level1Out42[28] , \Level1Out42[27] , 
        \Level1Out42[26] , \Level1Out42[25] , \Level1Out42[24] , 
        \Level1Out42[23] , \Level1Out42[22] , \Level1Out42[21] , 
        \Level1Out42[20] , \Level1Out42[19] , \Level1Out42[18] , 
        \Level1Out42[17] , \Level1Out42[16] , \Level1Out42[15] , 
        \Level1Out42[14] , \Level1Out42[13] , \Level1Out42[12] , 
        \Level1Out42[11] , \Level1Out42[10] , \Level1Out42[9] , 
        \Level1Out42[8] , \Level1Out42[7] , \Level1Out42[6] , \Level1Out42[5] , 
        \Level1Out42[4] , \Level1Out42[3] , \Level1Out42[2] , \Level1Out42[1] , 
        \Level1Out42[0] }), .In2({\Level1Out43[31] , \Level1Out43[30] , 
        \Level1Out43[29] , \Level1Out43[28] , \Level1Out43[27] , 
        \Level1Out43[26] , \Level1Out43[25] , \Level1Out43[24] , 
        \Level1Out43[23] , \Level1Out43[22] , \Level1Out43[21] , 
        \Level1Out43[20] , \Level1Out43[19] , \Level1Out43[18] , 
        \Level1Out43[17] , \Level1Out43[16] , \Level1Out43[15] , 
        \Level1Out43[14] , \Level1Out43[13] , \Level1Out43[12] , 
        \Level1Out43[11] , \Level1Out43[10] , \Level1Out43[9] , 
        \Level1Out43[8] , \Level1Out43[7] , \Level1Out43[6] , \Level1Out43[5] , 
        \Level1Out43[4] , \Level1Out43[3] , \Level1Out43[2] , \Level1Out43[1] , 
        \Level1Out43[0] }), .Read1(\Level1Load42[0] ), .Read2(
        \Level1Load43[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_31 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink31[31] , \ScanLink31[30] , 
        \ScanLink31[29] , \ScanLink31[28] , \ScanLink31[27] , \ScanLink31[26] , 
        \ScanLink31[25] , \ScanLink31[24] , \ScanLink31[23] , \ScanLink31[22] , 
        \ScanLink31[21] , \ScanLink31[20] , \ScanLink31[19] , \ScanLink31[18] , 
        \ScanLink31[17] , \ScanLink31[16] , \ScanLink31[15] , \ScanLink31[14] , 
        \ScanLink31[13] , \ScanLink31[12] , \ScanLink31[11] , \ScanLink31[10] , 
        \ScanLink31[9] , \ScanLink31[8] , \ScanLink31[7] , \ScanLink31[6] , 
        \ScanLink31[5] , \ScanLink31[4] , \ScanLink31[3] , \ScanLink31[2] , 
        \ScanLink31[1] , \ScanLink31[0] }), .ScanOut({\ScanLink32[31] , 
        \ScanLink32[30] , \ScanLink32[29] , \ScanLink32[28] , \ScanLink32[27] , 
        \ScanLink32[26] , \ScanLink32[25] , \ScanLink32[24] , \ScanLink32[23] , 
        \ScanLink32[22] , \ScanLink32[21] , \ScanLink32[20] , \ScanLink32[19] , 
        \ScanLink32[18] , \ScanLink32[17] , \ScanLink32[16] , \ScanLink32[15] , 
        \ScanLink32[14] , \ScanLink32[13] , \ScanLink32[12] , \ScanLink32[11] , 
        \ScanLink32[10] , \ScanLink32[9] , \ScanLink32[8] , \ScanLink32[7] , 
        \ScanLink32[6] , \ScanLink32[5] , \ScanLink32[4] , \ScanLink32[3] , 
        \ScanLink32[2] , \ScanLink32[1] , \ScanLink32[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load31[0] ), .Out({
        \Level1Out31[31] , \Level1Out31[30] , \Level1Out31[29] , 
        \Level1Out31[28] , \Level1Out31[27] , \Level1Out31[26] , 
        \Level1Out31[25] , \Level1Out31[24] , \Level1Out31[23] , 
        \Level1Out31[22] , \Level1Out31[21] , \Level1Out31[20] , 
        \Level1Out31[19] , \Level1Out31[18] , \Level1Out31[17] , 
        \Level1Out31[16] , \Level1Out31[15] , \Level1Out31[14] , 
        \Level1Out31[13] , \Level1Out31[12] , \Level1Out31[11] , 
        \Level1Out31[10] , \Level1Out31[9] , \Level1Out31[8] , 
        \Level1Out31[7] , \Level1Out31[6] , \Level1Out31[5] , \Level1Out31[4] , 
        \Level1Out31[3] , \Level1Out31[2] , \Level1Out31[1] , \Level1Out31[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_12_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load12[0] ), .Out({\Level2Out12[31] , \Level2Out12[30] , 
        \Level2Out12[29] , \Level2Out12[28] , \Level2Out12[27] , 
        \Level2Out12[26] , \Level2Out12[25] , \Level2Out12[24] , 
        \Level2Out12[23] , \Level2Out12[22] , \Level2Out12[21] , 
        \Level2Out12[20] , \Level2Out12[19] , \Level2Out12[18] , 
        \Level2Out12[17] , \Level2Out12[16] , \Level2Out12[15] , 
        \Level2Out12[14] , \Level2Out12[13] , \Level2Out12[12] , 
        \Level2Out12[11] , \Level2Out12[10] , \Level2Out12[9] , 
        \Level2Out12[8] , \Level2Out12[7] , \Level2Out12[6] , \Level2Out12[5] , 
        \Level2Out12[4] , \Level2Out12[3] , \Level2Out12[2] , \Level2Out12[1] , 
        \Level2Out12[0] }), .In1({\Level1Out12[31] , \Level1Out12[30] , 
        \Level1Out12[29] , \Level1Out12[28] , \Level1Out12[27] , 
        \Level1Out12[26] , \Level1Out12[25] , \Level1Out12[24] , 
        \Level1Out12[23] , \Level1Out12[22] , \Level1Out12[21] , 
        \Level1Out12[20] , \Level1Out12[19] , \Level1Out12[18] , 
        \Level1Out12[17] , \Level1Out12[16] , \Level1Out12[15] , 
        \Level1Out12[14] , \Level1Out12[13] , \Level1Out12[12] , 
        \Level1Out12[11] , \Level1Out12[10] , \Level1Out12[9] , 
        \Level1Out12[8] , \Level1Out12[7] , \Level1Out12[6] , \Level1Out12[5] , 
        \Level1Out12[4] , \Level1Out12[3] , \Level1Out12[2] , \Level1Out12[1] , 
        \Level1Out12[0] }), .In2({\Level1Out13[31] , \Level1Out13[30] , 
        \Level1Out13[29] , \Level1Out13[28] , \Level1Out13[27] , 
        \Level1Out13[26] , \Level1Out13[25] , \Level1Out13[24] , 
        \Level1Out13[23] , \Level1Out13[22] , \Level1Out13[21] , 
        \Level1Out13[20] , \Level1Out13[19] , \Level1Out13[18] , 
        \Level1Out13[17] , \Level1Out13[16] , \Level1Out13[15] , 
        \Level1Out13[14] , \Level1Out13[13] , \Level1Out13[12] , 
        \Level1Out13[11] , \Level1Out13[10] , \Level1Out13[9] , 
        \Level1Out13[8] , \Level1Out13[7] , \Level1Out13[6] , \Level1Out13[5] , 
        \Level1Out13[4] , \Level1Out13[3] , \Level1Out13[2] , \Level1Out13[1] , 
        \Level1Out13[0] }), .Read1(\Level1Load12[0] ), .Read2(
        \Level1Load13[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_38_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load38[0] ), .Out({\Level2Out38[31] , \Level2Out38[30] , 
        \Level2Out38[29] , \Level2Out38[28] , \Level2Out38[27] , 
        \Level2Out38[26] , \Level2Out38[25] , \Level2Out38[24] , 
        \Level2Out38[23] , \Level2Out38[22] , \Level2Out38[21] , 
        \Level2Out38[20] , \Level2Out38[19] , \Level2Out38[18] , 
        \Level2Out38[17] , \Level2Out38[16] , \Level2Out38[15] , 
        \Level2Out38[14] , \Level2Out38[13] , \Level2Out38[12] , 
        \Level2Out38[11] , \Level2Out38[10] , \Level2Out38[9] , 
        \Level2Out38[8] , \Level2Out38[7] , \Level2Out38[6] , \Level2Out38[5] , 
        \Level2Out38[4] , \Level2Out38[3] , \Level2Out38[2] , \Level2Out38[1] , 
        \Level2Out38[0] }), .In1({\Level1Out38[31] , \Level1Out38[30] , 
        \Level1Out38[29] , \Level1Out38[28] , \Level1Out38[27] , 
        \Level1Out38[26] , \Level1Out38[25] , \Level1Out38[24] , 
        \Level1Out38[23] , \Level1Out38[22] , \Level1Out38[21] , 
        \Level1Out38[20] , \Level1Out38[19] , \Level1Out38[18] , 
        \Level1Out38[17] , \Level1Out38[16] , \Level1Out38[15] , 
        \Level1Out38[14] , \Level1Out38[13] , \Level1Out38[12] , 
        \Level1Out38[11] , \Level1Out38[10] , \Level1Out38[9] , 
        \Level1Out38[8] , \Level1Out38[7] , \Level1Out38[6] , \Level1Out38[5] , 
        \Level1Out38[4] , \Level1Out38[3] , \Level1Out38[2] , \Level1Out38[1] , 
        \Level1Out38[0] }), .In2({\Level1Out39[31] , \Level1Out39[30] , 
        \Level1Out39[29] , \Level1Out39[28] , \Level1Out39[27] , 
        \Level1Out39[26] , \Level1Out39[25] , \Level1Out39[24] , 
        \Level1Out39[23] , \Level1Out39[22] , \Level1Out39[21] , 
        \Level1Out39[20] , \Level1Out39[19] , \Level1Out39[18] , 
        \Level1Out39[17] , \Level1Out39[16] , \Level1Out39[15] , 
        \Level1Out39[14] , \Level1Out39[13] , \Level1Out39[12] , 
        \Level1Out39[11] , \Level1Out39[10] , \Level1Out39[9] , 
        \Level1Out39[8] , \Level1Out39[7] , \Level1Out39[6] , \Level1Out39[5] , 
        \Level1Out39[4] , \Level1Out39[3] , \Level1Out39[2] , \Level1Out39[1] , 
        \Level1Out39[0] }), .Read1(\Level1Load38[0] ), .Read2(
        \Level1Load39[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_24_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load24[0] ), .Out({\Level4Out24[31] , \Level4Out24[30] , 
        \Level4Out24[29] , \Level4Out24[28] , \Level4Out24[27] , 
        \Level4Out24[26] , \Level4Out24[25] , \Level4Out24[24] , 
        \Level4Out24[23] , \Level4Out24[22] , \Level4Out24[21] , 
        \Level4Out24[20] , \Level4Out24[19] , \Level4Out24[18] , 
        \Level4Out24[17] , \Level4Out24[16] , \Level4Out24[15] , 
        \Level4Out24[14] , \Level4Out24[13] , \Level4Out24[12] , 
        \Level4Out24[11] , \Level4Out24[10] , \Level4Out24[9] , 
        \Level4Out24[8] , \Level4Out24[7] , \Level4Out24[6] , \Level4Out24[5] , 
        \Level4Out24[4] , \Level4Out24[3] , \Level4Out24[2] , \Level4Out24[1] , 
        \Level4Out24[0] }), .In1({\Level2Out24[31] , \Level2Out24[30] , 
        \Level2Out24[29] , \Level2Out24[28] , \Level2Out24[27] , 
        \Level2Out24[26] , \Level2Out24[25] , \Level2Out24[24] , 
        \Level2Out24[23] , \Level2Out24[22] , \Level2Out24[21] , 
        \Level2Out24[20] , \Level2Out24[19] , \Level2Out24[18] , 
        \Level2Out24[17] , \Level2Out24[16] , \Level2Out24[15] , 
        \Level2Out24[14] , \Level2Out24[13] , \Level2Out24[12] , 
        \Level2Out24[11] , \Level2Out24[10] , \Level2Out24[9] , 
        \Level2Out24[8] , \Level2Out24[7] , \Level2Out24[6] , \Level2Out24[5] , 
        \Level2Out24[4] , \Level2Out24[3] , \Level2Out24[2] , \Level2Out24[1] , 
        \Level2Out24[0] }), .In2({\Level2Out26[31] , \Level2Out26[30] , 
        \Level2Out26[29] , \Level2Out26[28] , \Level2Out26[27] , 
        \Level2Out26[26] , \Level2Out26[25] , \Level2Out26[24] , 
        \Level2Out26[23] , \Level2Out26[22] , \Level2Out26[21] , 
        \Level2Out26[20] , \Level2Out26[19] , \Level2Out26[18] , 
        \Level2Out26[17] , \Level2Out26[16] , \Level2Out26[15] , 
        \Level2Out26[14] , \Level2Out26[13] , \Level2Out26[12] , 
        \Level2Out26[11] , \Level2Out26[10] , \Level2Out26[9] , 
        \Level2Out26[8] , \Level2Out26[7] , \Level2Out26[6] , \Level2Out26[5] , 
        \Level2Out26[4] , \Level2Out26[3] , \Level2Out26[2] , \Level2Out26[1] , 
        \Level2Out26[0] }), .Read1(\Level2Load24[0] ), .Read2(
        \Level2Load26[0] ) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_44 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink44[31] , \ScanLink44[30] , 
        \ScanLink44[29] , \ScanLink44[28] , \ScanLink44[27] , \ScanLink44[26] , 
        \ScanLink44[25] , \ScanLink44[24] , \ScanLink44[23] , \ScanLink44[22] , 
        \ScanLink44[21] , \ScanLink44[20] , \ScanLink44[19] , \ScanLink44[18] , 
        \ScanLink44[17] , \ScanLink44[16] , \ScanLink44[15] , \ScanLink44[14] , 
        \ScanLink44[13] , \ScanLink44[12] , \ScanLink44[11] , \ScanLink44[10] , 
        \ScanLink44[9] , \ScanLink44[8] , \ScanLink44[7] , \ScanLink44[6] , 
        \ScanLink44[5] , \ScanLink44[4] , \ScanLink44[3] , \ScanLink44[2] , 
        \ScanLink44[1] , \ScanLink44[0] }), .ScanOut({\ScanLink45[31] , 
        \ScanLink45[30] , \ScanLink45[29] , \ScanLink45[28] , \ScanLink45[27] , 
        \ScanLink45[26] , \ScanLink45[25] , \ScanLink45[24] , \ScanLink45[23] , 
        \ScanLink45[22] , \ScanLink45[21] , \ScanLink45[20] , \ScanLink45[19] , 
        \ScanLink45[18] , \ScanLink45[17] , \ScanLink45[16] , \ScanLink45[15] , 
        \ScanLink45[14] , \ScanLink45[13] , \ScanLink45[12] , \ScanLink45[11] , 
        \ScanLink45[10] , \ScanLink45[9] , \ScanLink45[8] , \ScanLink45[7] , 
        \ScanLink45[6] , \ScanLink45[5] , \ScanLink45[4] , \ScanLink45[3] , 
        \ScanLink45[2] , \ScanLink45[1] , \ScanLink45[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b0), .Load(\Level1Load44[0] ), .Out({
        \Level1Out44[31] , \Level1Out44[30] , \Level1Out44[29] , 
        \Level1Out44[28] , \Level1Out44[27] , \Level1Out44[26] , 
        \Level1Out44[25] , \Level1Out44[24] , \Level1Out44[23] , 
        \Level1Out44[22] , \Level1Out44[21] , \Level1Out44[20] , 
        \Level1Out44[19] , \Level1Out44[18] , \Level1Out44[17] , 
        \Level1Out44[16] , \Level1Out44[15] , \Level1Out44[14] , 
        \Level1Out44[13] , \Level1Out44[12] , \Level1Out44[11] , 
        \Level1Out44[10] , \Level1Out44[9] , \Level1Out44[8] , 
        \Level1Out44[7] , \Level1Out44[6] , \Level1Out44[5] , \Level1Out44[4] , 
        \Level1Out44[3] , \Level1Out44[2] , \Level1Out44[1] , \Level1Out44[0] 
        }) );
    Merge_Low_Node_DWIDTH32_IDWIDTH1_SCAN1 U_Merge_Low_Node_63 ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\ScanLink63[31] , \ScanLink63[30] , 
        \ScanLink63[29] , \ScanLink63[28] , \ScanLink63[27] , \ScanLink63[26] , 
        \ScanLink63[25] , \ScanLink63[24] , \ScanLink63[23] , \ScanLink63[22] , 
        \ScanLink63[21] , \ScanLink63[20] , \ScanLink63[19] , \ScanLink63[18] , 
        \ScanLink63[17] , \ScanLink63[16] , \ScanLink63[15] , \ScanLink63[14] , 
        \ScanLink63[13] , \ScanLink63[12] , \ScanLink63[11] , \ScanLink63[10] , 
        \ScanLink63[9] , \ScanLink63[8] , \ScanLink63[7] , \ScanLink63[6] , 
        \ScanLink63[5] , \ScanLink63[4] , \ScanLink63[3] , \ScanLink63[2] , 
        \ScanLink63[1] , \ScanLink63[0] }), .ScanOut({\ScanLink64[31] , 
        \ScanLink64[30] , \ScanLink64[29] , \ScanLink64[28] , \ScanLink64[27] , 
        \ScanLink64[26] , \ScanLink64[25] , \ScanLink64[24] , \ScanLink64[23] , 
        \ScanLink64[22] , \ScanLink64[21] , \ScanLink64[20] , \ScanLink64[19] , 
        \ScanLink64[18] , \ScanLink64[17] , \ScanLink64[16] , \ScanLink64[15] , 
        \ScanLink64[14] , \ScanLink64[13] , \ScanLink64[12] , \ScanLink64[11] , 
        \ScanLink64[10] , \ScanLink64[9] , \ScanLink64[8] , \ScanLink64[7] , 
        \ScanLink64[6] , \ScanLink64[5] , \ScanLink64[4] , \ScanLink64[3] , 
        \ScanLink64[2] , \ScanLink64[1] , \ScanLink64[0] }), .ScanEnable(
        \ScanEnable[0] ), .Id(1'b1), .Load(\Level1Load63[0] ), .Out({
        \Level1Out63[31] , \Level1Out63[30] , \Level1Out63[29] , 
        \Level1Out63[28] , \Level1Out63[27] , \Level1Out63[26] , 
        \Level1Out63[25] , \Level1Out63[24] , \Level1Out63[23] , 
        \Level1Out63[22] , \Level1Out63[21] , \Level1Out63[20] , 
        \Level1Out63[19] , \Level1Out63[18] , \Level1Out63[17] , 
        \Level1Out63[16] , \Level1Out63[15] , \Level1Out63[14] , 
        \Level1Out63[13] , \Level1Out63[12] , \Level1Out63[11] , 
        \Level1Out63[10] , \Level1Out63[9] , \Level1Out63[8] , 
        \Level1Out63[7] , \Level1Out63[6] , \Level1Out63[5] , \Level1Out63[4] , 
        \Level1Out63[3] , \Level1Out63[2] , \Level1Out63[1] , \Level1Out63[0] 
        }) );
    Merge_Node_DWIDTH32 U_Merge_Node_20_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level2Load20[0] ), .Out({\Level2Out20[31] , \Level2Out20[30] , 
        \Level2Out20[29] , \Level2Out20[28] , \Level2Out20[27] , 
        \Level2Out20[26] , \Level2Out20[25] , \Level2Out20[24] , 
        \Level2Out20[23] , \Level2Out20[22] , \Level2Out20[21] , 
        \Level2Out20[20] , \Level2Out20[19] , \Level2Out20[18] , 
        \Level2Out20[17] , \Level2Out20[16] , \Level2Out20[15] , 
        \Level2Out20[14] , \Level2Out20[13] , \Level2Out20[12] , 
        \Level2Out20[11] , \Level2Out20[10] , \Level2Out20[9] , 
        \Level2Out20[8] , \Level2Out20[7] , \Level2Out20[6] , \Level2Out20[5] , 
        \Level2Out20[4] , \Level2Out20[3] , \Level2Out20[2] , \Level2Out20[1] , 
        \Level2Out20[0] }), .In1({\Level1Out20[31] , \Level1Out20[30] , 
        \Level1Out20[29] , \Level1Out20[28] , \Level1Out20[27] , 
        \Level1Out20[26] , \Level1Out20[25] , \Level1Out20[24] , 
        \Level1Out20[23] , \Level1Out20[22] , \Level1Out20[21] , 
        \Level1Out20[20] , \Level1Out20[19] , \Level1Out20[18] , 
        \Level1Out20[17] , \Level1Out20[16] , \Level1Out20[15] , 
        \Level1Out20[14] , \Level1Out20[13] , \Level1Out20[12] , 
        \Level1Out20[11] , \Level1Out20[10] , \Level1Out20[9] , 
        \Level1Out20[8] , \Level1Out20[7] , \Level1Out20[6] , \Level1Out20[5] , 
        \Level1Out20[4] , \Level1Out20[3] , \Level1Out20[2] , \Level1Out20[1] , 
        \Level1Out20[0] }), .In2({\Level1Out21[31] , \Level1Out21[30] , 
        \Level1Out21[29] , \Level1Out21[28] , \Level1Out21[27] , 
        \Level1Out21[26] , \Level1Out21[25] , \Level1Out21[24] , 
        \Level1Out21[23] , \Level1Out21[22] , \Level1Out21[21] , 
        \Level1Out21[20] , \Level1Out21[19] , \Level1Out21[18] , 
        \Level1Out21[17] , \Level1Out21[16] , \Level1Out21[15] , 
        \Level1Out21[14] , \Level1Out21[13] , \Level1Out21[12] , 
        \Level1Out21[11] , \Level1Out21[10] , \Level1Out21[9] , 
        \Level1Out21[8] , \Level1Out21[7] , \Level1Out21[6] , \Level1Out21[5] , 
        \Level1Out21[4] , \Level1Out21[3] , \Level1Out21[2] , \Level1Out21[1] , 
        \Level1Out21[0] }), .Read1(\Level1Load20[0] ), .Read2(
        \Level1Load21[0] ) );
    Merge_Node_DWIDTH32 U_Merge_Node_16_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), 
        .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Load(
        \Level4Load16[0] ), .Out({\Level4Out16[31] , \Level4Out16[30] , 
        \Level4Out16[29] , \Level4Out16[28] , \Level4Out16[27] , 
        \Level4Out16[26] , \Level4Out16[25] , \Level4Out16[24] , 
        \Level4Out16[23] , \Level4Out16[22] , \Level4Out16[21] , 
        \Level4Out16[20] , \Level4Out16[19] , \Level4Out16[18] , 
        \Level4Out16[17] , \Level4Out16[16] , \Level4Out16[15] , 
        \Level4Out16[14] , \Level4Out16[13] , \Level4Out16[12] , 
        \Level4Out16[11] , \Level4Out16[10] , \Level4Out16[9] , 
        \Level4Out16[8] , \Level4Out16[7] , \Level4Out16[6] , \Level4Out16[5] , 
        \Level4Out16[4] , \Level4Out16[3] , \Level4Out16[2] , \Level4Out16[1] , 
        \Level4Out16[0] }), .In1({\Level2Out16[31] , \Level2Out16[30] , 
        \Level2Out16[29] , \Level2Out16[28] , \Level2Out16[27] , 
        \Level2Out16[26] , \Level2Out16[25] , \Level2Out16[24] , 
        \Level2Out16[23] , \Level2Out16[22] , \Level2Out16[21] , 
        \Level2Out16[20] , \Level2Out16[19] , \Level2Out16[18] , 
        \Level2Out16[17] , \Level2Out16[16] , \Level2Out16[15] , 
        \Level2Out16[14] , \Level2Out16[13] , \Level2Out16[12] , 
        \Level2Out16[11] , \Level2Out16[10] , \Level2Out16[9] , 
        \Level2Out16[8] , \Level2Out16[7] , \Level2Out16[6] , \Level2Out16[5] , 
        \Level2Out16[4] , \Level2Out16[3] , \Level2Out16[2] , \Level2Out16[1] , 
        \Level2Out16[0] }), .In2({\Level2Out18[31] , \Level2Out18[30] , 
        \Level2Out18[29] , \Level2Out18[28] , \Level2Out18[27] , 
        \Level2Out18[26] , \Level2Out18[25] , \Level2Out18[24] , 
        \Level2Out18[23] , \Level2Out18[22] , \Level2Out18[21] , 
        \Level2Out18[20] , \Level2Out18[19] , \Level2Out18[18] , 
        \Level2Out18[17] , \Level2Out18[16] , \Level2Out18[15] , 
        \Level2Out18[14] , \Level2Out18[13] , \Level2Out18[12] , 
        \Level2Out18[11] , \Level2Out18[10] , \Level2Out18[9] , 
        \Level2Out18[8] , \Level2Out18[7] , \Level2Out18[6] , \Level2Out18[5] , 
        \Level2Out18[4] , \Level2Out18[3] , \Level2Out18[2] , \Level2Out18[1] , 
        \Level2Out18[0] }), .Read1(\Level2Load16[0] ), .Read2(
        \Level2Load18[0] ) );
endmodule

