
module CELL_DUMMY0_DW01_add_5_0 ( A, B, CI, SUM, CO );
input  [4:0] A;
input  [4:0] B;
output [4:0] SUM;
input  CI;
output CO;
    wire n1, \carry[2] , n2, n3, \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n1) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n2), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n2) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n1), .S(SUM[2]), .CO(SUM[3])
         );
    VMW_FADD U1_0 ( .CI(n3), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n3) );
endmodule


module CELL_DUMMY0_DW01_add_6_0 ( A, B, CI, SUM, CO );
input  [5:0] A;
input  [5:0] B;
output [5:0] SUM;
input  CI;
output CO;
    wire n4, n6, n7, \carry[2] , n5, \carry[3] , \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n4) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n6), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n5) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n5), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n7), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n6) );
    VMW_PULLDOWN U4 ( .Z(n7) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n4), .S(SUM[3]), .CO(SUM[4])
         );
endmodule


module CELL_DUMMY0_DW01_add_7_0 ( A, B, CI, SUM, CO );
input  [6:0] A;
input  [6:0] B;
output [6:0] SUM;
input  CI;
output CO;
    wire n8, n9, \carry[4] , n12, \carry[2] , n10, n11, \carry[3] , \carry[1] ;
    VMW_PULLDOWN U1 ( .Z(n8) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n11), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n9) );
    VMW_PULLDOWN U5 ( .Z(n12) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n10), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n12), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n10) );
    VMW_PULLDOWN U4 ( .Z(n11) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(n8), .S(SUM[4]), .CO(SUM[5])
         );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n9), .S(SUM[3]), .CO(
        \carry[4] ) );
endmodule


module CELL_DUMMY0_DW01_add_8_0 ( A, B, CI, SUM, CO );
input  [7:0] A;
input  [7:0] B;
output [7:0] SUM;
input  CI;
output CO;
    wire n13, n15, \carry[4] , \carry[2] , n14, n16, n17, n18, \carry[3] , 
        \carry[1] , \carry[5] ;
    VMW_PULLDOWN U1 ( .Z(n13) );
    VMW_PULLDOWN U6 ( .Z(n18) );
    VMW_FADD U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(n17), .S(SUM[1]), .CO(
        \carry[2] ) );
    VMW_PULLDOWN U2 ( .Z(n14) );
    VMW_PULLDOWN U5 ( .Z(n17) );
    VMW_FADD U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(n16), .S(SUM[2]), .CO(
        \carry[3] ) );
    VMW_FADD U1_0 ( .CI(n18), .A(A[0]), .B(B[0]), .S(SUM[0]), .CO(\carry[1] )
         );
    VMW_PULLDOWN U3 ( .Z(n15) );
    VMW_FADD U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(n13), .S(SUM[5]), .CO(SUM[6]
        ) );
    VMW_PULLDOWN U4 ( .Z(n16) );
    VMW_FADD U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(n14), .S(SUM[4]), .CO(
        \carry[5] ) );
    VMW_FADD U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(n15), .S(SUM[3]), .CO(
        \carry[4] ) );
endmodule


module CELL_DUMMY0 ( DATA_IN, cell_value, Reset, WR, Enable, Clk, NEIGHBORS );
input  [7:0] NEIGHBORS;
input  DATA_IN, Reset, WR, Enable, Clk;
output cell_value;
    wire n759, n776, \count75[6] , n758, n764, \count358[3] , \count353[1] , 
        \count75[4] , \count75[0] , \count75[2] , n771, n757, \count358[1] , 
        n763, n762, n770, \count363[2] , \count368[4] , \count368[0] , 
        \count368[2] , n773, n775, \count363[5] , \count368[6] , n765, 
        \count363[0] , n767, \count363[4] , \count368[3] , n375, \count75[5] , 
        n769, n772, \count363[3] , \count363[1] , \count368[1] , n760, 
        \count368[5] , \count353[2] , n768, \count358[0] , n774, \count358[4] , 
        n761, \count75[1] , \count75[3] , n766, \count358[2] , \count353[0] ;
    wire UNCONNECTED_1 , UNCONNECTED_2 , UNCONNECTED_3 , UNCONNECTED_4 ;
    VMW_PULLDOWN U123 ( .Z(n759) );
    VMW_PULLDOWN U125 ( .Z(n774) );
    VMW_PULLDOWN U126 ( .Z(n775) );
    VMW_AND2 U134 ( .A(NEIGHBORS[3]), .B(n758), .Z(n760) );
    VMW_XOR2 U141 ( .A(NEIGHBORS[3]), .B(n758), .Z(\count353[0] ) );
    VMW_INV U148 ( .A(\count75[1] ), .Z(n766) );
    VMW_PULLDOWN U127 ( .Z(n776) );
    VMW_PULLDOWN U128 ( .Z(n375) );
    CELL_DUMMY0_DW01_add_7_0 add_62_6 ( .A({n375, \count363[5] , \count363[4] , 
        \count363[3] , \count363[2] , \count363[1] , \count363[0] }), .B({n774, 
        n774, n774, n774, n774, n774, NEIGHBORS[6]}), .CI(n774), .SUM({
        UNCONNECTED_1, \count368[5] , \count368[4] , \count368[3] , 
        \count368[2] , \count368[1] , \count368[0] }) );
    VMW_PULLDOWN U129 ( .Z(\count358[4] ) );
    VMW_OR3 U132 ( .A(\count75[5] ), .B(\count75[4] ), .C(\count75[6] ), .Z(
        n767) );
    VMW_AND3 U133 ( .A(n757), .B(n758), .C(NEIGHBORS[3]), .Z(\count353[2] ) );
    VMW_MUX2I U146 ( .A(n768), .B(cell_value), .S(n761), .Z(n764) );
    CELL_DUMMY0_DW01_add_8_0 add_62_7 ( .A({n375, \count368[6] , \count368[5] , 
        \count368[4] , \count368[3] , \count368[2] , \count368[1] , 
        \count368[0] }), .B({n773, n773, n773, n773, n773, n773, n773, 
        NEIGHBORS[7]}), .CI(n773), .SUM({UNCONNECTED_2, \count75[6] , 
        \count75[5] , \count75[4] , \count75[3] , \count75[2] , \count75[1] , 
        \count75[0] }) );
    VMW_OR2 U147 ( .A(Reset), .B(n770), .Z(n771) );
    VMW_AND2 U135 ( .A(\count75[0] ), .B(n762), .Z(n761) );
    VMW_XOR2 U140 ( .A(n757), .B(n760), .Z(\count353[1] ) );
    VMW_XOR2 U137 ( .A(NEIGHBORS[1]), .B(NEIGHBORS[0]), .Z(n765) );
    VMW_INV U149 ( .A(cell_value), .Z(n769) );
    VMW_OR2 U142 ( .A(n762), .B(n769), .Z(n768) );
    VMW_FD cell_value_reg ( .D(n772), .CP(Clk), .Q(cell_value) );
    VMW_PULLDOWN U130 ( .Z(\count363[5] ) );
    VMW_NOR4 U139 ( .A(\count75[3] ), .B(\count75[2] ), .C(n766), .D(n767), 
        .Z(n762) );
    CELL_DUMMY0_DW01_add_6_0 add_62_5 ( .A({n375, \count358[4] , \count358[3] , 
        \count358[2] , \count358[1] , \count358[0] }), .B({n775, n775, n775, 
        n775, n775, NEIGHBORS[5]}), .CI(n775), .SUM({UNCONNECTED_3, 
        \count363[4] , \count363[3] , \count363[2] , \count363[1] , 
        \count363[0] }) );
    VMW_AO22 U145 ( .A(NEIGHBORS[1]), .B(NEIGHBORS[0]), .C(NEIGHBORS[2]), .D(
        n765), .Z(n757) );
    VMW_XOR2 U138 ( .A(NEIGHBORS[2]), .B(n765), .Z(n758) );
    VMW_PULLDOWN U124 ( .Z(n773) );
    VMW_PULLDOWN U131 ( .Z(\count368[6] ) );
    CELL_DUMMY0_DW01_add_5_0 add_62_4 ( .A({n375, n759, \count353[2] , 
        \count353[1] , \count353[0] }), .B({n776, n776, n776, n776, 
        NEIGHBORS[4]}), .CI(n776), .SUM({UNCONNECTED_4, \count358[3] , 
        \count358[2] , \count358[1] , \count358[0] }) );
    VMW_AOI211 U136 ( .A(n764), .B(Enable), .C(WR), .D(Reset), .Z(n763) );
    VMW_MUX2I U143 ( .A(n769), .B(DATA_IN), .S(WR), .Z(n770) );
    VMW_MUX2I U144 ( .A(n771), .B(n769), .S(n763), .Z(n772) );
endmodule


module Life_Block_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, DataIn, DataOut, 
    ScanIn, ScanOut, ScanEnable, Id, Enable, BLOCK_VALUE, NORTH_EDGE, 
    SOUTH_EDGE, EAST_EDGE, WEST_EDGE, NW_EDGE, SW_EDGE, NE_EDGE, SE_EDGE );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
output [31:0] BLOCK_VALUE;
input  [31:0] NORTH_EDGE;
input  [31:0] SOUTH_EDGE;
input  Clk, Reset, RD, WR, ScanEnable, Enable, EAST_EDGE, WEST_EDGE, NW_EDGE, 
    SW_EDGE, NE_EDGE, SE_EDGE;
    wire \BLOCK_VALUE[31] , \BLOCK_VALUE[5] , \BLOCK_VALUE[1] , 
        \BLOCK_VALUE[8] , \BLOCK_VALUE[7] , \BLOCK_VALUE[3] , 
        \BLOCK_VALUE[25] , \BLOCK_VALUE[16] , \BLOCK_VALUE[21] , 
        \BLOCK_VALUE[12] , \BLOCK_VALUE[28] , \BLOCK_VALUE[19] , 
        \BLOCK_VALUE[23] , \BLOCK_VALUE[10] , \BLOCK_VALUE[27] , 
        \BLOCK_VALUE[14] , \BLOCK_VALUE[26] , \BLOCK_VALUE[15] , 
        \BLOCK_VALUE[18] , \BLOCK_VALUE[22] , \BLOCK_VALUE[11] , 
        \BLOCK_VALUE[20] , \BLOCK_VALUE[13] , \BLOCK_VALUE[30] , 
        \BLOCK_VALUE[29] , \BLOCK_VALUE[24] , \BLOCK_VALUE[17] , 
        \BLOCK_VALUE[2] , \BLOCK_VALUE[6] , \BLOCK_VALUE[4] , \BLOCK_VALUE[0] , 
        \BLOCK_VALUE[9] ;
    assign ScanOut[31] = \BLOCK_VALUE[31] ;
    assign ScanOut[30] = \BLOCK_VALUE[30] ;
    assign ScanOut[29] = \BLOCK_VALUE[29] ;
    assign ScanOut[28] = \BLOCK_VALUE[28] ;
    assign ScanOut[27] = \BLOCK_VALUE[27] ;
    assign ScanOut[26] = \BLOCK_VALUE[26] ;
    assign ScanOut[25] = \BLOCK_VALUE[25] ;
    assign ScanOut[24] = \BLOCK_VALUE[24] ;
    assign ScanOut[23] = \BLOCK_VALUE[23] ;
    assign ScanOut[22] = \BLOCK_VALUE[22] ;
    assign ScanOut[21] = \BLOCK_VALUE[21] ;
    assign ScanOut[20] = \BLOCK_VALUE[20] ;
    assign ScanOut[19] = \BLOCK_VALUE[19] ;
    assign ScanOut[18] = \BLOCK_VALUE[18] ;
    assign ScanOut[17] = \BLOCK_VALUE[17] ;
    assign ScanOut[16] = \BLOCK_VALUE[16] ;
    assign ScanOut[15] = \BLOCK_VALUE[15] ;
    assign ScanOut[14] = \BLOCK_VALUE[14] ;
    assign ScanOut[13] = \BLOCK_VALUE[13] ;
    assign ScanOut[12] = \BLOCK_VALUE[12] ;
    assign ScanOut[11] = \BLOCK_VALUE[11] ;
    assign ScanOut[10] = \BLOCK_VALUE[10] ;
    assign ScanOut[9] = \BLOCK_VALUE[9] ;
    assign ScanOut[8] = \BLOCK_VALUE[8] ;
    assign ScanOut[7] = \BLOCK_VALUE[7] ;
    assign ScanOut[6] = \BLOCK_VALUE[6] ;
    assign ScanOut[5] = \BLOCK_VALUE[5] ;
    assign ScanOut[4] = \BLOCK_VALUE[4] ;
    assign ScanOut[3] = \BLOCK_VALUE[3] ;
    assign ScanOut[2] = \BLOCK_VALUE[2] ;
    assign ScanOut[1] = \BLOCK_VALUE[1] ;
    assign ScanOut[0] = \BLOCK_VALUE[0] ;
    assign BLOCK_VALUE[31] = \BLOCK_VALUE[31] ;
    assign BLOCK_VALUE[30] = \BLOCK_VALUE[30] ;
    assign BLOCK_VALUE[29] = \BLOCK_VALUE[29] ;
    assign BLOCK_VALUE[28] = \BLOCK_VALUE[28] ;
    assign BLOCK_VALUE[27] = \BLOCK_VALUE[27] ;
    assign BLOCK_VALUE[26] = \BLOCK_VALUE[26] ;
    assign BLOCK_VALUE[25] = \BLOCK_VALUE[25] ;
    assign BLOCK_VALUE[24] = \BLOCK_VALUE[24] ;
    assign BLOCK_VALUE[23] = \BLOCK_VALUE[23] ;
    assign BLOCK_VALUE[22] = \BLOCK_VALUE[22] ;
    assign BLOCK_VALUE[21] = \BLOCK_VALUE[21] ;
    assign BLOCK_VALUE[20] = \BLOCK_VALUE[20] ;
    assign BLOCK_VALUE[19] = \BLOCK_VALUE[19] ;
    assign BLOCK_VALUE[18] = \BLOCK_VALUE[18] ;
    assign BLOCK_VALUE[17] = \BLOCK_VALUE[17] ;
    assign BLOCK_VALUE[16] = \BLOCK_VALUE[16] ;
    assign BLOCK_VALUE[15] = \BLOCK_VALUE[15] ;
    assign BLOCK_VALUE[14] = \BLOCK_VALUE[14] ;
    assign BLOCK_VALUE[13] = \BLOCK_VALUE[13] ;
    assign BLOCK_VALUE[12] = \BLOCK_VALUE[12] ;
    assign BLOCK_VALUE[11] = \BLOCK_VALUE[11] ;
    assign BLOCK_VALUE[10] = \BLOCK_VALUE[10] ;
    assign BLOCK_VALUE[9] = \BLOCK_VALUE[9] ;
    assign BLOCK_VALUE[8] = \BLOCK_VALUE[8] ;
    assign BLOCK_VALUE[7] = \BLOCK_VALUE[7] ;
    assign BLOCK_VALUE[6] = \BLOCK_VALUE[6] ;
    assign BLOCK_VALUE[5] = \BLOCK_VALUE[5] ;
    assign BLOCK_VALUE[4] = \BLOCK_VALUE[4] ;
    assign BLOCK_VALUE[3] = \BLOCK_VALUE[3] ;
    assign BLOCK_VALUE[2] = \BLOCK_VALUE[2] ;
    assign BLOCK_VALUE[1] = \BLOCK_VALUE[1] ;
    assign BLOCK_VALUE[0] = \BLOCK_VALUE[0] ;
    CELL_DUMMY0 cell_4 ( .DATA_IN(ScanIn[4]), .cell_value(\BLOCK_VALUE[4] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[5], \BLOCK_VALUE[5] , SOUTH_EDGE[5], 
        SOUTH_EDGE[4], SOUTH_EDGE[3], \BLOCK_VALUE[3] , NORTH_EDGE[3], 
        NORTH_EDGE[4]}) );
    CELL_DUMMY0 cell_15 ( .DATA_IN(ScanIn[15]), .cell_value(\BLOCK_VALUE[15] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[16], \BLOCK_VALUE[16] , SOUTH_EDGE[16], 
        SOUTH_EDGE[15], SOUTH_EDGE[14], \BLOCK_VALUE[14] , NORTH_EDGE[14], 
        NORTH_EDGE[15]}) );
    CELL_DUMMY0 cell_29 ( .DATA_IN(ScanIn[29]), .cell_value(\BLOCK_VALUE[29] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[30], \BLOCK_VALUE[30] , SOUTH_EDGE[30], 
        SOUTH_EDGE[29], SOUTH_EDGE[28], \BLOCK_VALUE[28] , NORTH_EDGE[28], 
        NORTH_EDGE[29]}) );
    CELL_DUMMY0 cell_3 ( .DATA_IN(ScanIn[3]), .cell_value(\BLOCK_VALUE[3] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[4], \BLOCK_VALUE[4] , SOUTH_EDGE[4], 
        SOUTH_EDGE[3], SOUTH_EDGE[2], \BLOCK_VALUE[2] , NORTH_EDGE[2], 
        NORTH_EDGE[3]}) );
    CELL_DUMMY0 cell_20 ( .DATA_IN(ScanIn[20]), .cell_value(\BLOCK_VALUE[20] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[21], \BLOCK_VALUE[21] , SOUTH_EDGE[21], 
        SOUTH_EDGE[20], SOUTH_EDGE[19], \BLOCK_VALUE[19] , NORTH_EDGE[19], 
        NORTH_EDGE[20]}) );
    CELL_DUMMY0 cell_27 ( .DATA_IN(ScanIn[27]), .cell_value(\BLOCK_VALUE[27] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[28], \BLOCK_VALUE[28] , SOUTH_EDGE[28], 
        SOUTH_EDGE[27], SOUTH_EDGE[26], \BLOCK_VALUE[26] , NORTH_EDGE[26], 
        NORTH_EDGE[27]}) );
    CELL_DUMMY0 cell_12 ( .DATA_IN(ScanIn[12]), .cell_value(\BLOCK_VALUE[12] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[13], \BLOCK_VALUE[13] , SOUTH_EDGE[13], 
        SOUTH_EDGE[12], SOUTH_EDGE[11], \BLOCK_VALUE[11] , NORTH_EDGE[11], 
        NORTH_EDGE[12]}) );
    CELL_DUMMY0 cell_26 ( .DATA_IN(ScanIn[26]), .cell_value(\BLOCK_VALUE[26] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[27], \BLOCK_VALUE[27] , SOUTH_EDGE[27], 
        SOUTH_EDGE[26], SOUTH_EDGE[25], \BLOCK_VALUE[25] , NORTH_EDGE[25], 
        NORTH_EDGE[26]}) );
    CELL_DUMMY0 cell_2 ( .DATA_IN(ScanIn[2]), .cell_value(\BLOCK_VALUE[2] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[3], \BLOCK_VALUE[3] , SOUTH_EDGE[3], 
        SOUTH_EDGE[2], SOUTH_EDGE[1], \BLOCK_VALUE[1] , NORTH_EDGE[1], 
        NORTH_EDGE[2]}) );
    CELL_DUMMY0 cell_5 ( .DATA_IN(ScanIn[5]), .cell_value(\BLOCK_VALUE[5] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[6], \BLOCK_VALUE[6] , SOUTH_EDGE[6], 
        SOUTH_EDGE[5], SOUTH_EDGE[4], \BLOCK_VALUE[4] , NORTH_EDGE[4], 
        NORTH_EDGE[5]}) );
    CELL_DUMMY0 cell_13 ( .DATA_IN(ScanIn[13]), .cell_value(\BLOCK_VALUE[13] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[14], \BLOCK_VALUE[14] , SOUTH_EDGE[14], 
        SOUTH_EDGE[13], SOUTH_EDGE[12], \BLOCK_VALUE[12] , NORTH_EDGE[12], 
        NORTH_EDGE[13]}) );
    CELL_DUMMY0 cell_14 ( .DATA_IN(ScanIn[14]), .cell_value(\BLOCK_VALUE[14] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[15], \BLOCK_VALUE[15] , SOUTH_EDGE[15], 
        SOUTH_EDGE[14], SOUTH_EDGE[13], \BLOCK_VALUE[13] , NORTH_EDGE[13], 
        NORTH_EDGE[14]}) );
    CELL_DUMMY0 cell_21 ( .DATA_IN(ScanIn[21]), .cell_value(\BLOCK_VALUE[21] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[22], \BLOCK_VALUE[22] , SOUTH_EDGE[22], 
        SOUTH_EDGE[21], SOUTH_EDGE[20], \BLOCK_VALUE[20] , NORTH_EDGE[20], 
        NORTH_EDGE[21]}) );
    CELL_DUMMY0 cell_28 ( .DATA_IN(ScanIn[28]), .cell_value(\BLOCK_VALUE[28] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[29], \BLOCK_VALUE[29] , SOUTH_EDGE[29], 
        SOUTH_EDGE[28], SOUTH_EDGE[27], \BLOCK_VALUE[27] , NORTH_EDGE[27], 
        NORTH_EDGE[28]}) );
    CELL_DUMMY0 cell_0 ( .DATA_IN(ScanIn[0]), .cell_value(\BLOCK_VALUE[0] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[1], \BLOCK_VALUE[1] , SOUTH_EDGE[1], 
        SOUTH_EDGE[0], SE_EDGE, EAST_EDGE, NE_EDGE, NORTH_EDGE[0]}) );
    CELL_DUMMY0 cell_7 ( .DATA_IN(ScanIn[7]), .cell_value(\BLOCK_VALUE[7] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[8], \BLOCK_VALUE[8] , SOUTH_EDGE[8], 
        SOUTH_EDGE[7], SOUTH_EDGE[6], \BLOCK_VALUE[6] , NORTH_EDGE[6], 
        NORTH_EDGE[7]}) );
    CELL_DUMMY0 cell_16 ( .DATA_IN(ScanIn[16]), .cell_value(\BLOCK_VALUE[16] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[17], \BLOCK_VALUE[17] , SOUTH_EDGE[17], 
        SOUTH_EDGE[16], SOUTH_EDGE[15], \BLOCK_VALUE[15] , NORTH_EDGE[15], 
        NORTH_EDGE[16]}) );
    CELL_DUMMY0 cell_31 ( .DATA_IN(ScanIn[31]), .cell_value(\BLOCK_VALUE[31] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NW_EDGE, WEST_EDGE, SW_EDGE, SOUTH_EDGE[31], 
        SOUTH_EDGE[30], \BLOCK_VALUE[30] , NORTH_EDGE[30], NORTH_EDGE[31]}) );
    CELL_DUMMY0 cell_9 ( .DATA_IN(ScanIn[9]), .cell_value(\BLOCK_VALUE[9] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[10], \BLOCK_VALUE[10] , SOUTH_EDGE[10], 
        SOUTH_EDGE[9], SOUTH_EDGE[8], \BLOCK_VALUE[8] , NORTH_EDGE[8], 
        NORTH_EDGE[9]}) );
    CELL_DUMMY0 cell_18 ( .DATA_IN(ScanIn[18]), .cell_value(\BLOCK_VALUE[18] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[19], \BLOCK_VALUE[19] , SOUTH_EDGE[19], 
        SOUTH_EDGE[18], SOUTH_EDGE[17], \BLOCK_VALUE[17] , NORTH_EDGE[17], 
        NORTH_EDGE[18]}) );
    CELL_DUMMY0 cell_23 ( .DATA_IN(ScanIn[23]), .cell_value(\BLOCK_VALUE[23] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[24], \BLOCK_VALUE[24] , SOUTH_EDGE[24], 
        SOUTH_EDGE[23], SOUTH_EDGE[22], \BLOCK_VALUE[22] , NORTH_EDGE[22], 
        NORTH_EDGE[23]}) );
    CELL_DUMMY0 cell_24 ( .DATA_IN(ScanIn[24]), .cell_value(\BLOCK_VALUE[24] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[25], \BLOCK_VALUE[25] , SOUTH_EDGE[25], 
        SOUTH_EDGE[24], SOUTH_EDGE[23], \BLOCK_VALUE[23] , NORTH_EDGE[23], 
        NORTH_EDGE[24]}) );
    CELL_DUMMY0 cell_1 ( .DATA_IN(ScanIn[1]), .cell_value(\BLOCK_VALUE[1] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[2], \BLOCK_VALUE[2] , SOUTH_EDGE[2], 
        SOUTH_EDGE[1], SOUTH_EDGE[0], \BLOCK_VALUE[0] , NORTH_EDGE[0], 
        NORTH_EDGE[1]}) );
    CELL_DUMMY0 cell_8 ( .DATA_IN(ScanIn[8]), .cell_value(\BLOCK_VALUE[8] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[9], \BLOCK_VALUE[9] , SOUTH_EDGE[9], 
        SOUTH_EDGE[8], SOUTH_EDGE[7], \BLOCK_VALUE[7] , NORTH_EDGE[7], 
        NORTH_EDGE[8]}) );
    CELL_DUMMY0 cell_11 ( .DATA_IN(ScanIn[11]), .cell_value(\BLOCK_VALUE[11] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[12], \BLOCK_VALUE[12] , SOUTH_EDGE[12], 
        SOUTH_EDGE[11], SOUTH_EDGE[10], \BLOCK_VALUE[10] , NORTH_EDGE[10], 
        NORTH_EDGE[11]}) );
    CELL_DUMMY0 cell_19 ( .DATA_IN(ScanIn[19]), .cell_value(\BLOCK_VALUE[19] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[20], \BLOCK_VALUE[20] , SOUTH_EDGE[20], 
        SOUTH_EDGE[19], SOUTH_EDGE[18], \BLOCK_VALUE[18] , NORTH_EDGE[18], 
        NORTH_EDGE[19]}) );
    CELL_DUMMY0 cell_25 ( .DATA_IN(ScanIn[25]), .cell_value(\BLOCK_VALUE[25] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[26], \BLOCK_VALUE[26] , SOUTH_EDGE[26], 
        SOUTH_EDGE[25], SOUTH_EDGE[24], \BLOCK_VALUE[24] , NORTH_EDGE[24], 
        NORTH_EDGE[25]}) );
    CELL_DUMMY0 cell_6 ( .DATA_IN(ScanIn[6]), .cell_value(\BLOCK_VALUE[6] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[7], \BLOCK_VALUE[7] , SOUTH_EDGE[7], 
        SOUTH_EDGE[6], SOUTH_EDGE[5], \BLOCK_VALUE[5] , NORTH_EDGE[5], 
        NORTH_EDGE[6]}) );
    CELL_DUMMY0 cell_10 ( .DATA_IN(ScanIn[10]), .cell_value(\BLOCK_VALUE[10] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[11], \BLOCK_VALUE[11] , SOUTH_EDGE[11], 
        SOUTH_EDGE[10], SOUTH_EDGE[9], \BLOCK_VALUE[9] , NORTH_EDGE[9], 
        NORTH_EDGE[10]}) );
    CELL_DUMMY0 cell_17 ( .DATA_IN(ScanIn[17]), .cell_value(\BLOCK_VALUE[17] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[18], \BLOCK_VALUE[18] , SOUTH_EDGE[18], 
        SOUTH_EDGE[17], SOUTH_EDGE[16], \BLOCK_VALUE[16] , NORTH_EDGE[16], 
        NORTH_EDGE[17]}) );
    CELL_DUMMY0 cell_30 ( .DATA_IN(ScanIn[30]), .cell_value(\BLOCK_VALUE[30] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[31], \BLOCK_VALUE[31] , SOUTH_EDGE[31], 
        SOUTH_EDGE[30], SOUTH_EDGE[29], \BLOCK_VALUE[29] , NORTH_EDGE[29], 
        NORTH_EDGE[30]}) );
    CELL_DUMMY0 cell_22 ( .DATA_IN(ScanIn[22]), .cell_value(\BLOCK_VALUE[22] ), 
        .Reset(Reset), .WR(ScanEnable), .Enable(Enable), .Clk(Clk), 
        .NEIGHBORS({NORTH_EDGE[23], \BLOCK_VALUE[23] , SOUTH_EDGE[23], 
        SOUTH_EDGE[22], SOUTH_EDGE[21], \BLOCK_VALUE[21] , NORTH_EDGE[21], 
        NORTH_EDGE[22]}) );
endmodule


module Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 ( A, SUM );
input  [6:0] A;
output [6:0] SUM;
    wire n5, n9, n7, n12, n6, n13, n8, n10, n11;
    VMW_AO21 U3 ( .A(n5), .B(A[2]), .C(n6), .Z(SUM[2]) );
    VMW_AO21 U5 ( .A(A[0]), .B(A[1]), .C(n9), .Z(SUM[1]) );
    VMW_INV U6 ( .A(A[0]), .Z(SUM[0]) );
    VMW_AO22 U14 ( .A(A[5]), .B(n13), .C(n12), .D(n10), .Z(SUM[5]) );
    VMW_AO21 U7 ( .A(n8), .B(A[4]), .C(n10), .Z(SUM[4]) );
    VMW_AND2 U8 ( .A(n10), .B(n12), .Z(n11) );
    VMW_XOR2 U13 ( .A(A[6]), .B(n11), .Z(SUM[6]) );
    VMW_OR2 U9 ( .A(A[0]), .B(A[1]), .Z(n5) );
    VMW_NOR2 U12 ( .A(n8), .B(A[4]), .Z(n10) );
    VMW_INV U15 ( .A(A[5]), .Z(n12) );
    VMW_INV U17 ( .A(A[3]), .Z(n7) );
    VMW_NOR2 U10 ( .A(n5), .B(A[2]), .Z(n6) );
    VMW_NAND2 U11 ( .A(n6), .B(n7), .Z(n8) );
    VMW_OAI21 U4 ( .A(n6), .B(n7), .C(n8), .Z(SUM[3]) );
    VMW_INV U18 ( .A(n5), .Z(n9) );
    VMW_INV U16 ( .A(n10), .Z(n13) );
endmodule


module Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1 ( Clk, Reset, RD, WR, Addr, 
    DataIn, DataOut, ScanIn, ScanOut, ScanEnable, Id, ScanId, Enable );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  [0:0] Id;
input  [31:0] ScanIn;
output [31:0] ScanOut;
input  [0:0] ScanId;
input  Clk, Reset, RD, WR;
output ScanEnable, Enable;
    wire n330, n317, \count[2] , n362, n345, \count[6] , n339, n357, n322, 
        n325, n350, n319, \count[4] , n342, \count[0] , n359, n356, n337, n318, 
        n351, \ScanReg[15] , \ScanReg[26] , \ScanReg[2] , \count260[3] , n324, 
        \ScanReg[18] , n336, n358, n343, \ScanReg[22] , \ScanReg[11] , 
        \ScanReg[6] , \count260[5] , \ScanReg[20] , \ScanReg[13] , 
        \ScanReg[4] , n344, \count260[1] , n316, \ScanReg[29] , \ScanReg[30] , 
        n331, n323, \ScanReg[17] , \ScanReg[24] , \ScanReg[0] , \ScanReg[9] , 
        n338, n314, \count260[0] , n333, \ScanReg[16] , \ScanReg[25] , n361, 
        n346, \ScanReg[1] , \ScanReg[8] , \ScanReg[7] , n328, \ScanReg[5] , 
        \count260[4] , \ScanReg[21] , \ScanReg[12] , n354, \ScanReg[28] , 
        \ScanReg[31] , n321, n326, \ScanReg[19] , n348, \count260[6] , n353, 
        \ScanReg[10] , \ScanReg[23] , n341, \ScanReg[14] , \ScanReg[27] , n313, 
        \ScanReg[3] , \count260[2] , n334, \count[1] , n352, n349, n327, n335, 
        n360, n340, \count[5] , n347, n329, n332, n315, n320, \count[3] , n355;
    tri \arr[31] , \arr[22] , \arr[11] , \arr[18] , \arr[26] , \arr[15] , 
        \arr[30] , \arr[24] , \arr[17] , \arr[29] , \arr[20] , \arr[13] , 
        \arr[3] , \arr[7] , \arr[8] , \arr[5] , \arr[9] , \arr[1] , \arr[0] , 
        \arr[6] , \arr[4] , \arr[2] , \arr[28] , \arr[21] , \arr[12] , 
        \arr[27] , \arr[25] , \arr[16] , \arr[14] , \arr[23] , \arr[10] , 
        \arr[19] ;
    assign DataOut[31] = \arr[31] ;
    assign DataOut[30] = \arr[30] ;
    assign DataOut[29] = \arr[29] ;
    assign DataOut[28] = \arr[28] ;
    assign DataOut[27] = \arr[27] ;
    assign DataOut[26] = \arr[26] ;
    assign DataOut[25] = \arr[25] ;
    assign DataOut[24] = \arr[24] ;
    assign DataOut[23] = \arr[23] ;
    assign DataOut[22] = \arr[22] ;
    assign DataOut[21] = \arr[21] ;
    assign DataOut[20] = \arr[20] ;
    assign DataOut[19] = \arr[19] ;
    assign DataOut[18] = \arr[18] ;
    assign DataOut[17] = \arr[17] ;
    assign DataOut[16] = \arr[16] ;
    assign DataOut[15] = \arr[15] ;
    assign DataOut[14] = \arr[14] ;
    assign DataOut[13] = \arr[13] ;
    assign DataOut[12] = \arr[12] ;
    assign DataOut[11] = \arr[11] ;
    assign DataOut[10] = \arr[10] ;
    assign DataOut[9] = \arr[9] ;
    assign DataOut[8] = \arr[8] ;
    assign DataOut[7] = \arr[7] ;
    assign DataOut[6] = \arr[6] ;
    assign DataOut[5] = \arr[5] ;
    assign DataOut[4] = \arr[4] ;
    assign DataOut[3] = \arr[3] ;
    assign DataOut[2] = \arr[2] ;
    assign DataOut[1] = \arr[1] ;
    assign DataOut[0] = \arr[0] ;
    VMW_AND2 U54 ( .A(DataIn[29]), .B(WR), .Z(ScanOut[29]) );
    VMW_AND2 U73 ( .A(DataIn[10]), .B(WR), .Z(ScanOut[10]) );
    VMW_NOR2 U113 ( .A(n318), .B(n316), .Z(n314) );
    VMW_INV U134 ( .A(n321), .Z(ScanEnable) );
    VMW_AND2 U68 ( .A(DataIn[15]), .B(WR), .Z(ScanOut[15]) );
    VMW_AND2 U96 ( .A(\ScanReg[13] ), .B(n316), .Z(n340) );
    VMW_AO21 U108 ( .A(RD), .B(ScanEnable), .C(n317), .Z(n328) );
    VMW_BUFIZ U141 ( .A(n330), .E(n328), .Z(\arr[27] ) );
    VMW_BUFIZ U166 ( .A(n355), .E(n328), .Z(\arr[8] ) );
    VMW_FD \ScanReg_reg[5]  ( .D(ScanIn[5]), .CP(Clk), .Q(\ScanReg[5] ) );
    VMW_FD \count_reg[6]  ( .D(n356), .CP(Clk), .Q(\count[6] ) );
    VMW_AND2 U53 ( .A(DataIn[30]), .B(WR), .Z(ScanOut[30]) );
    VMW_AND2 U61 ( .A(DataIn[22]), .B(WR), .Z(ScanOut[22]) );
    VMW_AND2 U84 ( .A(\ScanReg[8] ), .B(n316), .Z(n355) );
    VMW_BUFIZ U148 ( .A(n337), .E(n328), .Z(\arr[21] ) );
    VMW_BUFIZ U153 ( .A(n342), .E(n328), .Z(\arr[29] ) );
    VMW_FD \ScanReg_reg[8]  ( .D(ScanIn[8]), .CP(Clk), .Q(\ScanReg[8] ) );
    Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1_DW01_dec_7_0 sub_281 ( .A({
        \count[6] , \count[5] , \count[4] , \count[3] , \count[2] , \count[1] , 
        \count[0] }), .SUM({\count260[6] , \count260[5] , \count260[4] , 
        \count260[3] , \count260[2] , \count260[1] , \count260[0] }) );
    VMW_FD \count_reg[2]  ( .D(n360), .CP(Clk), .Q(\count[2] ) );
    VMW_FD \ScanReg_reg[1]  ( .D(ScanIn[1]), .CP(Clk), .Q(\ScanReg[1] ) );
    VMW_AND2 U66 ( .A(DataIn[17]), .B(WR), .Z(ScanOut[17]) );
    VMW_AND2 U101 ( .A(\ScanReg[16] ), .B(n316), .Z(n333) );
    VMW_AND2 U106 ( .A(\ScanReg[10] ), .B(n316), .Z(n326) );
    VMW_OAI21 U121 ( .A(RD), .B(WR), .C(n322), .Z(n321) );
    VMW_AO22 U126 ( .A(\count[2] ), .B(n317), .C(\ScanReg[2] ), .D(n316), .Z(
        n339) );
    VMW_AO22 U83 ( .A(ScanOut[6]), .B(n314), .C(\count260[6] ), .D(n315), .Z(
        n356) );
    VMW_FD \count_reg[0]  ( .D(n362), .CP(Clk), .Q(\count[0] ) );
    VMW_AND2 U91 ( .A(\ScanReg[17] ), .B(n316), .Z(n346) );
    VMW_AND2 U98 ( .A(\ScanReg[21] ), .B(n316), .Z(n337) );
    VMW_FD \ScanReg_reg[3]  ( .D(ScanIn[3]), .CP(Clk), .Q(\ScanReg[3] ) );
    VMW_AO22 U128 ( .A(\count[0] ), .B(n317), .C(\ScanReg[0] ), .D(n316), .Z(
        n324) );
    VMW_BUFIZ U154 ( .A(n343), .E(n328), .Z(\arr[20] ) );
    VMW_FD \count_reg[4]  ( .D(n358), .CP(Clk), .Q(\count[4] ) );
    VMW_FD \ScanReg_reg[7]  ( .D(ScanIn[7]), .CP(Clk), .Q(\ScanReg[7] ) );
    VMW_BUFIZ U146 ( .A(n335), .E(n328), .Z(\arr[6] ) );
    VMW_BUFIZ U161 ( .A(n350), .E(n328), .Z(\arr[15] ) );
    VMW_AND2 U74 ( .A(DataIn[9]), .B(WR), .Z(ScanOut[9]) );
    VMW_AND2 U114 ( .A(DataIn[6]), .B(WR), .Z(ScanOut[6]) );
    VMW_INV U133 ( .A(Reset), .Z(n320) );
    VMW_AND2 U99 ( .A(\ScanReg[31] ), .B(n316), .Z(n336) );
    VMW_BUFIZ U155 ( .A(n344), .E(n328), .Z(\arr[3] ) );
    VMW_AND2 U52 ( .A(DataIn[31]), .B(WR), .Z(ScanOut[31]) );
    VMW_AND2 U67 ( .A(DataIn[16]), .B(WR), .Z(ScanOut[16]) );
    VMW_AO22 U82 ( .A(ScanOut[5]), .B(n314), .C(\count260[5] ), .D(n315), .Z(
        n357) );
    VMW_AND2 U107 ( .A(\ScanReg[23] ), .B(n316), .Z(n325) );
    VMW_AND2 U120 ( .A(DataIn[0]), .B(WR), .Z(ScanOut[0]) );
    VMW_FD \ScanReg_reg[27]  ( .D(ScanIn[27]), .CP(Clk), .Q(\ScanReg[27] ) );
    VMW_FD \ScanReg_reg[14]  ( .D(ScanIn[14]), .CP(Clk), .Q(\ScanReg[14] ) );
    VMW_AND2 U55 ( .A(DataIn[28]), .B(WR), .Z(ScanOut[28]) );
    VMW_AND2 U69 ( .A(DataIn[14]), .B(WR), .Z(ScanOut[14]) );
    VMW_AND2 U75 ( .A(DataIn[8]), .B(WR), .Z(ScanOut[8]) );
    VMW_AND2 U115 ( .A(DataIn[5]), .B(WR), .Z(ScanOut[5]) );
    VMW_XNOR2 U132 ( .A(Addr[0]), .B(ScanId), .Z(n322) );
    VMW_AND2 U90 ( .A(\ScanReg[7] ), .B(n316), .Z(n347) );
    VMW_AND2 U109 ( .A(\ScanReg[19] ), .B(n316), .Z(n323) );
    VMW_OR4 U129 ( .A(\count[3] ), .B(\count[4] ), .C(\count[5] ), .D(
        \count[6] ), .Z(n313) );
    VMW_BUFIZ U147 ( .A(n336), .E(n328), .Z(\arr[31] ) );
    VMW_FD \ScanReg_reg[19]  ( .D(ScanIn[19]), .CP(Clk), .Q(\ScanReg[19] ) );
    VMW_BUFIZ U160 ( .A(n349), .E(n328), .Z(\arr[26] ) );
    VMW_FD \ScanReg_reg[23]  ( .D(ScanIn[23]), .CP(Clk), .Q(\ScanReg[23] ) );
    VMW_FD \ScanReg_reg[10]  ( .D(ScanIn[10]), .CP(Clk), .Q(\ScanReg[10] ) );
    VMW_AND2 U72 ( .A(DataIn[11]), .B(WR), .Z(ScanOut[11]) );
    VMW_AND2 U97 ( .A(\ScanReg[28] ), .B(n316), .Z(n338) );
    VMW_BUFIZ U140 ( .A(n329), .E(n328), .Z(\arr[4] ) );
    VMW_FD \ScanReg_reg[21]  ( .D(ScanIn[21]), .CP(Clk), .Q(\ScanReg[21] ) );
    VMW_FD \ScanReg_reg[12]  ( .D(ScanIn[12]), .CP(Clk), .Q(\ScanReg[12] ) );
    VMW_FD \ScanReg_reg[31]  ( .D(ScanIn[31]), .CP(Clk), .Q(\ScanReg[31] ) );
    VMW_FD \ScanReg_reg[28]  ( .D(ScanIn[28]), .CP(Clk), .Q(\ScanReg[28] ) );
    VMW_NOR2 U112 ( .A(n318), .B(n319), .Z(n315) );
    VMW_BUFIZ U135 ( .A(n323), .E(n328), .Z(\arr[19] ) );
    VMW_AND2 U60 ( .A(DataIn[23]), .B(WR), .Z(ScanOut[23]) );
    VMW_AND2 U85 ( .A(\ScanReg[11] ), .B(n316), .Z(n353) );
    VMW_AND2 U100 ( .A(\ScanReg[12] ), .B(n316), .Z(n334) );
    VMW_AO22 U127 ( .A(\count[1] ), .B(n317), .C(\ScanReg[1] ), .D(n316), .Z(
        n354) );
    VMW_FD \ScanReg_reg[25]  ( .D(ScanIn[25]), .CP(Clk), .Q(\ScanReg[25] ) );
    VMW_BUFIZ U149 ( .A(n338), .E(n328), .Z(\arr[28] ) );
    VMW_FD \ScanReg_reg[16]  ( .D(ScanIn[16]), .CP(Clk), .Q(\ScanReg[16] ) );
    VMW_BUFIZ U152 ( .A(n341), .E(n328), .Z(\arr[30] ) );
    VMW_OR4 U51 ( .A(\count[1] ), .B(\count[2] ), .C(\count[0] ), .D(n313), 
        .Z(Enable) );
    VMW_AND2 U57 ( .A(DataIn[26]), .B(WR), .Z(ScanOut[26]) );
    VMW_BUFIZ U137 ( .A(n325), .E(n328), .Z(\arr[23] ) );
    VMW_FD \ScanReg_reg[24]  ( .D(ScanIn[24]), .CP(Clk), .Q(\ScanReg[24] ) );
    VMW_AND2 U58 ( .A(DataIn[25]), .B(WR), .Z(ScanOut[25]) );
    VMW_AND2 U59 ( .A(DataIn[24]), .B(WR), .Z(ScanOut[24]) );
    VMW_AND2 U62 ( .A(DataIn[21]), .B(WR), .Z(ScanOut[21]) );
    VMW_AND2 U70 ( .A(DataIn[13]), .B(WR), .Z(ScanOut[13]) );
    VMW_FD \ScanReg_reg[17]  ( .D(ScanIn[17]), .CP(Clk), .Q(\ScanReg[17] ) );
    VMW_AO22 U79 ( .A(ScanOut[2]), .B(n314), .C(\count260[2] ), .D(n315), .Z(
        n360) );
    VMW_AND2 U95 ( .A(\ScanReg[30] ), .B(n316), .Z(n341) );
    VMW_XOR2 U110 ( .A(Addr[0]), .B(Id), .Z(n316) );
    VMW_BUFIZ U159 ( .A(n348), .E(n328), .Z(\arr[5] ) );
    VMW_AND2 U119 ( .A(DataIn[1]), .B(WR), .Z(ScanOut[1]) );
    VMW_BUFIZ U142 ( .A(n331), .E(n328), .Z(\arr[14] ) );
    VMW_BUFIZ U165 ( .A(n354), .E(n328), .Z(\arr[1] ) );
    VMW_AND2 U87 ( .A(\ScanReg[18] ), .B(n316), .Z(n351) );
    VMW_BUFIZ U150 ( .A(n339), .E(n328), .Z(\arr[2] ) );
    VMW_FD \ScanReg_reg[20]  ( .D(ScanIn[20]), .CP(Clk), .Q(\ScanReg[20] ) );
    VMW_FD \ScanReg_reg[13]  ( .D(ScanIn[13]), .CP(Clk), .Q(\ScanReg[13] ) );
    VMW_AO22 U125 ( .A(\count[3] ), .B(n317), .C(\ScanReg[3] ), .D(n316), .Z(
        n344) );
    VMW_FD \ScanReg_reg[30]  ( .D(ScanIn[30]), .CP(Clk), .Q(\ScanReg[30] ) );
    VMW_FD \ScanReg_reg[29]  ( .D(ScanIn[29]), .CP(Clk), .Q(\ScanReg[29] ) );
    VMW_AND2 U65 ( .A(DataIn[18]), .B(WR), .Z(ScanOut[18]) );
    VMW_AND2 U102 ( .A(\ScanReg[25] ), .B(n316), .Z(n332) );
    VMW_AND2 U105 ( .A(\ScanReg[9] ), .B(n316), .Z(n327) );
    VMW_AO22 U80 ( .A(ScanOut[3]), .B(n314), .C(\count260[3] ), .D(n315), .Z(
        n359) );
    VMW_AO22 U122 ( .A(\count[6] ), .B(n317), .C(\ScanReg[6] ), .D(n316), .Z(
        n335) );
    VMW_FD \ScanReg_reg[18]  ( .D(ScanIn[18]), .CP(Clk), .Q(\ScanReg[18] ) );
    VMW_BUFIZ U139 ( .A(n327), .E(n328), .Z(\arr[9] ) );
    VMW_BUFIZ U157 ( .A(n346), .E(n328), .Z(\arr[17] ) );
    VMW_FD \ScanReg_reg[22]  ( .D(ScanIn[22]), .CP(Clk), .Q(\ScanReg[22] ) );
    VMW_FD \ScanReg_reg[11]  ( .D(ScanIn[11]), .CP(Clk), .Q(\ScanReg[11] ) );
    VMW_AO22 U77 ( .A(ScanOut[0]), .B(n314), .C(\count260[0] ), .D(n315), .Z(
        n362) );
    VMW_AND2 U89 ( .A(\ScanReg[26] ), .B(n316), .Z(n349) );
    VMW_AND2 U92 ( .A(\ScanReg[24] ), .B(n316), .Z(n345) );
    VMW_BUFIZ U145 ( .A(n334), .E(n328), .Z(\arr[12] ) );
    VMW_BUFIZ U162 ( .A(n351), .E(n328), .Z(\arr[18] ) );
    VMW_AND2 U117 ( .A(DataIn[3]), .B(WR), .Z(ScanOut[3]) );
    VMW_FD \ScanReg_reg[26]  ( .D(ScanIn[26]), .CP(Clk), .Q(\ScanReg[26] ) );
    VMW_FD \ScanReg_reg[15]  ( .D(ScanIn[15]), .CP(Clk), .Q(\ScanReg[15] ) );
    VMW_AND2 U130 ( .A(n317), .B(WR), .Z(n319) );
    VMW_BUFIZ U138 ( .A(n326), .E(n328), .Z(\arr[10] ) );
    VMW_FD \ScanReg_reg[6]  ( .D(ScanIn[6]), .CP(Clk), .Q(\ScanReg[6] ) );
    VMW_FD \count_reg[5]  ( .D(n357), .CP(Clk), .Q(\count[5] ) );
    VMW_AND2 U64 ( .A(DataIn[19]), .B(WR), .Z(ScanOut[19]) );
    VMW_AO22 U81 ( .A(ScanOut[4]), .B(n314), .C(\count260[4] ), .D(n315), .Z(
        n358) );
    VMW_BUFIZ U156 ( .A(n345), .E(n328), .Z(\arr[24] ) );
    VMW_AND2 U104 ( .A(\ScanReg[27] ), .B(n316), .Z(n330) );
    VMW_AND2 U76 ( .A(DataIn[7]), .B(WR), .Z(ScanOut[7]) );
    VMW_AND2 U116 ( .A(DataIn[4]), .B(WR), .Z(ScanOut[4]) );
    VMW_AO22 U123 ( .A(\count[5] ), .B(n317), .C(\ScanReg[5] ), .D(n316), .Z(
        n348) );
    VMW_AND2 U56 ( .A(DataIn[27]), .B(WR), .Z(ScanOut[27]) );
    VMW_AND2 U88 ( .A(\ScanReg[15] ), .B(n316), .Z(n350) );
    VMW_AND2 U93 ( .A(\ScanReg[20] ), .B(n316), .Z(n343) );
    VMW_INV U131 ( .A(n316), .Z(n317) );
    VMW_FD \count_reg[1]  ( .D(n361), .CP(Clk), .Q(\count[1] ) );
    VMW_FD \ScanReg_reg[2]  ( .D(ScanIn[2]), .CP(Clk), .Q(\ScanReg[2] ) );
    VMW_AND2 U94 ( .A(\ScanReg[29] ), .B(n316), .Z(n342) );
    VMW_BUFIZ U143 ( .A(n332), .E(n328), .Z(\arr[25] ) );
    VMW_BUFIZ U144 ( .A(n333), .E(n328), .Z(\arr[16] ) );
    VMW_BUFIZ U163 ( .A(n352), .E(n328), .Z(\arr[22] ) );
    VMW_BUFIZ U158 ( .A(n347), .E(n328), .Z(\arr[7] ) );
    VMW_BUFIZ U164 ( .A(n353), .E(n328), .Z(\arr[11] ) );
    VMW_FD \ScanReg_reg[9]  ( .D(ScanIn[9]), .CP(Clk), .Q(\ScanReg[9] ) );
    VMW_FD \count_reg[3]  ( .D(n359), .CP(Clk), .Q(\count[3] ) );
    VMW_BUFIZ U136 ( .A(n324), .E(n328), .Z(\arr[0] ) );
    VMW_FD \ScanReg_reg[0]  ( .D(ScanIn[0]), .CP(Clk), .Q(\ScanReg[0] ) );
    VMW_AND2 U63 ( .A(DataIn[20]), .B(WR), .Z(ScanOut[20]) );
    VMW_AND2 U71 ( .A(DataIn[12]), .B(WR), .Z(ScanOut[12]) );
    VMW_OAI21 U111 ( .A(n319), .B(Enable), .C(n320), .Z(n318) );
    VMW_AO22 U124 ( .A(\count[4] ), .B(n317), .C(\ScanReg[4] ), .D(n316), .Z(
        n329) );
    VMW_AO22 U78 ( .A(ScanOut[1]), .B(n314), .C(\count260[1] ), .D(n315), .Z(
        n361) );
    VMW_AND2 U86 ( .A(\ScanReg[22] ), .B(n316), .Z(n352) );
    VMW_AND2 U103 ( .A(\ScanReg[14] ), .B(n316), .Z(n331) );
    VMW_AND2 U118 ( .A(DataIn[2]), .B(WR), .Z(ScanOut[2]) );
    VMW_BUFIZ U151 ( .A(n340), .E(n328), .Z(\arr[13] ) );
    VMW_FD \ScanReg_reg[4]  ( .D(ScanIn[4]), .CP(Clk), .Q(\ScanReg[4] ) );
endmodule


module main ( Clk, Reset, RD, WR, Addr, DataIn, DataOut );
input  [14:0] Addr;
input  [31:0] DataIn;
output [31:0] DataOut;
input  Clk, Reset, RD, WR;
    wire \nScanOut2[20] , \nScanOut2[13] , \nScanOut29[23] , \nOut2_15[3] , 
        \nOut0_1[1] , \nOut0_2[2] , \nOut0_3[22] , \nScanOut11[1] , 
        \nScanOut29[10] , \nOut2_4[26] , \nOut0_3[11] , \nOut1_9[6] , 
        \nScanOut12[2] , \nScanOut14[19] , \nScanOut37[31] , \nScanOut37[28] , 
        \nScanOut42[18] , \nScanOut4[1] , \nScanOut7[2] , \nOut1_8[23] , 
        \nOut0_13[19] , \nOut2_4[15] , \nOut2_10[18] , \nOut2_14[29] , 
        \nOut2_14[30] , \nScanOut6[22] , \nOut0_7[20] , \nOut0_7[13] , 
        \nOut1_8[10] , \nOut2_0[24] , \nScanOut10[31] , \nScanOut10[28] , 
        \nScanOut46[30] , \nScanOut33[19] , \nScanOut36[4] , \nScanOut46[29] , 
        \nOut2_0[17] , \nScanOut28[8] , \nScanOut35[7] , \nScanOut38[15] , 
        \nOut1_12[27] , \nScanOut38[26] , \nOut1_12[14] , \nScanOut33[9] , 
        \nOut1_2[25] , \nOut0_6[19] , \nScanOut6[11] , \nOut0_9[9] , 
        \nOut1_11[4] , \nOut1_12[7] , \nScanOut38[2] , \nScanOut27[27] , 
        \nScanOut32[13] , \nScanOut47[23] , \nOut1_9[30] , \nScanOut9[4] , 
        \nScanOut11[22] , \nOut2_15[10] , \nScanOut32[20] , \nScanOut41[9] , 
        \nOut1_9[29] , \nScanOut11[11] , \nOut2_15[23] , \nScanOut47[10] , 
        \nOut1_14[9] , \nScanOut27[14] , \nScanOut20[0] , \nScanOut23[3] , 
        \nOut1_2[16] , \nScanOut7[31] , \nScanOut47[7] , \nScanOut7[28] , 
        \nScanOut3[19] , \nOut1_6[27] , \nScanOut44[4] , \nOut0_9[24] , 
        \nOut1_4[3] , \nOut1_6[14] , \nScanOut19[9] , \nScanOut8[26] , 
        \nOut0_9[17] , \nScanOut28[30] , \nScanOut28[29] , \nOut0_11[9] , 
        \nOut0_12[13] , \nScanOut15[20] , \nOut2_0[2] , \nScanOut36[11] , 
        \nScanOut43[21] , \nScanOut23[25] , \nOut2_11[12] , \nOut0_14[4] , 
        \nOut2_3[1] , \nScanOut23[16] , \nScanOut15[13] , \nScanOut36[22] , 
        \nScanOut43[12] , \nOut2_11[21] , \nOut0_1[8] , \nOut1_1[7] , 
        \nOut0_2[31] , \nOut0_2[28] , \nOut1_7[0] , \nOut0_2[21] , 
        \nOut0_6[23] , \nScanOut7[21] , \nScanOut8[15] , \nOut0_12[20] , 
        \nScanOut7[12] , \nOut1_13[24] , \nOut1_13[17] , \nScanOut39[16] , 
        \nOut1_14[0] , \nOut2_1[27] , \nScanOut20[9] , \nScanOut39[25] , 
        \nScanOut41[0] , \nOut0_6[10] , \nOut1_9[20] , \nScanOut11[18] , 
        \nScanOut32[29] , \nScanOut42[3] , \nScanOut47[19] , \nScanOut32[30] , 
        \nOut0_9[0] , \nOut2_1[14] , \nScanOut25[4] , \nScanOut26[7] , 
        \nOut1_9[13] , \nOut2_11[31] , \nOut2_15[19] , \nOut2_11[28] , 
        \nOut0_2[12] , \nOut1_7[9] , \nOut0_12[30] , \nOut2_5[25] , 
        \nOut0_12[29] , \nScanOut15[30] , \nScanOut36[18] , \nScanOut43[28] , 
        \nScanOut15[29] , \nScanOut43[31] , \nOut2_3[8] , \nOut2_5[16] , 
        \nOut1_2[4] , \nOut0_12[3] , \nScanOut19[0] , \nScanOut28[20] , 
        \nScanOut48[24] , \nScanOut3[23] , \nScanOut2[30] , \nScanOut2[29] , 
        \nOut0_3[18] , \nScanOut3[10] , \nOut0_11[0] , \nOut2_5[6] , 
        \nOut2_6[5] , \nScanOut48[17] , \nScanOut28[13] , \nOut1_7[24] , 
        \nOut0_8[27] , \nScanOut9[25] , \nOut0_13[10] , \nOut2_13[4] , 
        \nScanOut9[16] , \nOut0_13[23] , \nScanOut14[23] , \nScanOut22[26] , 
        \nOut2_10[11] , \nOut2_10[7] , \nScanOut37[12] , \nScanOut42[22] , 
        \nScanOut11[8] , \nScanOut14[10] , \nScanOut22[15] , \nOut2_10[22] , 
        \nScanOut37[21] , \nScanOut42[11] , \nOut2_8[3] , \nOut0_8[14] , 
        \nScanOut17[6] , \nScanOut29[19] , \nOut1_3[26] , \nOut1_7[17] , 
        \nScanOut14[5] , \nScanOut30[3] , \nScanOut33[0] , \nOut1_3[15] , 
        \nScanOut6[18] , \nScanOut1[5] , \nScanOut2[6] , \nOut0_4[5] , 
        \nScanOut4[8] , \nOut0_7[6] , \nOut1_8[19] , \nScanOut10[21] , 
        \nOut2_14[13] , \nScanOut26[24] , \nScanOut33[10] , \nScanOut46[20] , 
        \nScanOut28[1] , \nScanOut10[12] , \nScanOut26[17] , \nOut2_14[20] , 
        \nScanOut33[23] , \nScanOut46[13] , \nOut0_7[30] , \nOut0_7[29] , 
        \nOut1_7[4] , \nScanOut8[22] , \nOut0_12[17] , \nOut2_3[5] , 
        \nScanOut8[11] , \nOut0_12[24] , \nScanOut15[24] , \nScanOut23[21] , 
        \nOut2_11[16] , \nOut2_0[6] , \nScanOut36[15] , \nScanOut43[25] , 
        \nOut2_5[31] , \nOut2_5[28] , \nOut1_4[7] , \nOut0_14[0] , 
        \nScanOut15[17] , \nOut2_11[25] , \nScanOut23[12] , \nScanOut36[26] , 
        \nScanOut43[16] , \nOut0_1[5] , \nScanOut1[8] , \nOut1_2[21] , 
        \nOut1_2[9] , \nOut1_6[23] , \nOut0_9[20] , \nOut1_6[10] , 
        \nOut0_9[13] , \nOut2_6[8] , \nScanOut48[30] , \nScanOut39[31] , 
        \nScanOut48[29] , \nOut1_2[12] , \nScanOut20[4] , \nScanOut39[28] , 
        \nScanOut23[7] , \nScanOut44[0] , \nOut1_3[18] , \nScanOut6[26] , 
        \nScanOut9[0] , \nOut1_11[0] , \nScanOut11[26] , \nOut1_13[30] , 
        \nOut1_13[29] , \nScanOut47[3] , \nOut2_15[14] , \nScanOut11[15] , 
        \nOut1_12[3] , \nScanOut27[23] , \nScanOut32[17] , \nScanOut47[27] , 
        \nOut2_1[19] , \nScanOut25[9] , \nScanOut27[10] , \nScanOut38[6] , 
        \nOut2_15[27] , \nScanOut32[24] , \nScanOut47[14] , \nOut1_12[23] , 
        \nScanOut38[11] , \nOut0_2[6] , \nScanOut6[15] , \nOut1_12[10] , 
        \nScanOut2[24] , \nOut0_3[26] , \nOut0_4[8] , \nScanOut4[5] , 
        \nOut0_7[24] , \nOut2_0[20] , \nScanOut38[22] , \nOut0_7[17] , 
        \nScanOut7[6] , \nOut1_8[27] , \nOut1_8[14] , \nOut2_0[13] , 
        \nScanOut35[3] , \nScanOut36[0] , \nScanOut26[30] , \nScanOut26[29] , 
        \nOut1_9[2] , \nScanOut12[6] , \nScanOut22[18] , \nOut0_3[15] , 
        \nScanOut9[31] , \nScanOut11[5] , \nOut2_4[22] , \nScanOut9[28] , 
        \nOut2_4[11] , \nOut2_13[9] , \nScanOut14[8] , \nScanOut29[27] , 
        \nOut1_7[30] , \nOut0_8[19] , \nOut1_7[29] , \nScanOut29[14] , 
        \nScanOut1[1] , \nScanOut2[17] , \nOut2_15[7] , \nScanOut2[2] , 
        \nOut1_3[22] , \nOut0_4[1] , \nOut0_7[2] , \nScanOut10[25] , 
        \nScanOut26[20] , \nScanOut28[5] , \nScanOut33[14] , \nScanOut36[9] , 
        \nScanOut46[24] , \nOut2_14[17] , \nScanOut10[16] , \nOut2_0[30] , 
        \nOut2_0[29] , \nScanOut33[27] , \nScanOut46[17] , \nOut1_12[19] , 
        \nScanOut26[13] , \nOut2_14[24] , \nScanOut30[7] , \nScanOut33[4] , 
        \nOut1_3[11] , \nScanOut38[18] , \nOut1_7[20] , \nOut1_1[3] , 
        \nOut1_7[13] , \nOut0_8[23] , \nScanOut14[1] , \nOut2_8[7] , 
        \nOut0_8[10] , \nScanOut9[21] , \nOut0_13[14] , \nScanOut14[27] , 
        \nScanOut17[2] , \nOut2_10[15] , \nOut2_10[3] , \nScanOut37[16] , 
        \nScanOut42[26] , \nOut2_4[18] , \nScanOut22[22] , \nScanOut9[12] , 
        \nOut0_13[27] , \nScanOut14[14] , \nScanOut22[11] , \nOut2_13[0] , 
        \nOut2_10[26] , \nScanOut37[25] , \nScanOut42[15] , \nOut0_11[4] , 
        \nOut0_2[25] , \nOut1_2[0] , \nScanOut3[27] , \nOut1_6[19] , 
        \nScanOut3[14] , \nOut0_12[7] , \nScanOut19[4] , \nScanOut48[20] , 
        \nScanOut28[24] , \nScanOut8[18] , \nOut0_9[30] , \nOut2_5[2] , 
        \nOut0_9[29] , \nOut2_6[1] , \nScanOut28[17] , \nScanOut48[13] , 
        \nOut2_5[21] , \nOut1_1[1] , \nOut0_2[16] , \nOut0_14[9] , 
        \nOut1_2[31] , \nOut1_2[28] , \nOut0_6[27] , \nOut1_9[24] , 
        \nOut2_5[12] , \nScanOut23[31] , \nScanOut23[28] , \nScanOut27[19] , 
        \nScanOut42[7] , \nOut0_6[14] , \nOut0_9[4] , \nScanOut9[9] , 
        \nOut2_1[23] , \nScanOut41[4] , \nOut1_9[17] , \nOut1_11[9] , 
        \nOut2_1[10] , \nScanOut26[3] , \nScanOut25[0] , \nScanOut7[25] , 
        \nScanOut39[12] , \nScanOut44[9] , \nOut1_13[20] , \nScanOut39[21] , 
        \nOut1_2[2] , \nScanOut7[16] , \nOut1_13[13] , \nOut1_14[4] , 
        \nOut0_12[5] , \nScanOut28[26] , \nScanOut3[25] , \nScanOut19[6] , 
        \nScanOut48[22] , \nScanOut1[3] , \nOut0_2[27] , \nScanOut3[16] , 
        \nOut1_6[31] , \nOut1_6[28] , \nOut0_9[18] , \nOut0_11[6] , 
        \nOut2_6[3] , \nOut2_5[0] , \nScanOut28[15] , \nScanOut48[11] , 
        \nScanOut23[19] , \nOut0_2[14] , \nScanOut8[30] , \nScanOut8[29] , 
        \nOut2_5[23] , \nOut2_5[10] , \nOut1_2[19] , \nOut0_6[25] , 
        \nOut2_1[21] , \nScanOut41[6] , \nOut0_6[16] , \nOut1_9[26] , 
        \nScanOut42[5] , \nScanOut7[27] , \nOut0_9[6] , \nOut1_12[8] , 
        \nOut2_1[12] , \nScanOut25[2] , \nOut1_9[15] , \nOut1_13[22] , 
        \nScanOut26[1] , \nScanOut27[31] , \nScanOut27[28] , \nScanOut47[8] , 
        \nOut1_3[20] , \nOut0_4[3] , \nScanOut7[14] , \nScanOut39[10] , 
        \nOut1_13[11] , \nOut1_14[6] , \nScanOut39[23] , \nOut0_7[0] , 
        \nScanOut10[27] , \nOut2_14[15] , \nScanOut33[16] , \nScanOut46[26] , 
        \nOut2_0[18] , \nScanOut26[22] , \nScanOut35[8] , \nScanOut10[14] , 
        \nScanOut26[11] , \nScanOut28[7] , \nOut2_14[26] , \nScanOut33[25] , 
        \nScanOut46[15] , \nScanOut38[29] , \nOut1_3[13] , \nScanOut30[5] , 
        \nScanOut38[30] , \nScanOut33[6] , \nScanOut2[0] , \nOut1_12[31] , 
        \nOut1_7[22] , \nOut0_8[21] , \nOut1_12[28] , \nOut2_8[5] , 
        \nOut0_1[7] , \nScanEnable[0] , \nScanOut2[9] , \nOut1_7[11] , 
        \nOut0_8[12] , \nScanOut17[0] , \nOut1_9[9] , \nScanOut9[23] , 
        \nOut0_13[16] , \nScanOut14[3] , \nOut2_13[2] , \nScanOut9[10] , 
        \nOut0_13[25] , \nScanOut14[25] , \nScanOut22[20] , \nScanOut37[14] , 
        \nScanOut42[24] , \nOut2_4[30] , \nOut2_10[17] , \nOut2_10[1] , 
        \nOut2_4[29] , \nScanOut14[16] , \nScanOut37[27] , \nScanOut42[17] , 
        \nOut2_10[24] , \nScanOut22[13] , \nScanOut38[13] , \nScanOut6[24] , 
        \nOut1_12[21] , \nOut0_2[4] , \nOut1_3[30] , \nOut1_3[29] , 
        \nScanOut38[20] , \nScanOut6[17] , \nOut1_12[12] , \nOut0_3[24] , 
        \nScanOut4[7] , \nOut0_7[26] , \nScanOut7[4] , \nOut1_8[25] , 
        \nScanOut26[18] , \nOut0_7[15] , \nOut0_7[9] , \nOut1_8[16] , 
        \nOut2_0[22] , \nScanOut36[2] , \nOut2_0[11] , \nScanOut35[1] , 
        \nScanOut9[19] , \nScanOut11[7] , \nOut2_4[20] , \nOut0_3[17] , 
        \nOut1_9[0] , \nScanOut12[4] , \nScanOut17[9] , \nOut2_4[13] , 
        \nScanOut22[30] , \nScanOut22[29] , \nOut2_10[8] , \nScanOut2[26] , 
        \nScanOut2[15] , \nOut1_7[18] , \nScanOut29[25] , \nOut2_15[5] , 
        \nOut0_8[31] , \nOut0_8[28] , \nScanOut8[20] , \nOut0_12[15] , 
        \nScanOut15[26] , \nOut2_0[4] , \nScanOut29[16] , \nOut2_5[19] , 
        \nScanOut23[23] , \nOut2_11[14] , \nScanOut36[17] , \nScanOut43[27] , 
        \nOut0_14[2] , \nOut2_3[7] , \nScanOut23[10] , \nScanOut15[15] , 
        \nOut2_11[27] , \nScanOut36[24] , \nScanOut43[14] , \nOut1_1[8] , 
        \nOut1_4[5] , \nOut1_6[21] , \nOut1_7[6] , \nScanOut8[13] , 
        \nOut0_12[26] , \nOut1_6[12] , \nOut0_9[22] , \nScanOut48[18] , 
        \nOut2_5[9] , \nScanOut1[7] , \nOut0_2[9] , \nOut1_2[23] , 
        \nOut0_9[11] , \nOut1_13[18] , \nScanOut20[6] , \nScanOut23[5] , 
        \nOut1_2[10] , \nScanOut47[1] , \nScanOut2[18] , \nOut0_3[30] , 
        \nScanOut9[27] , \nScanOut9[2] , \nOut1_11[2] , \nScanOut11[24] , 
        \nOut1_12[1] , \nScanOut38[4] , \nScanOut39[19] , \nScanOut44[2] , 
        \nScanOut27[21] , \nOut2_15[16] , \nScanOut26[8] , \nScanOut32[15] , 
        \nOut2_1[28] , \nScanOut47[25] , \nScanOut11[17] , \nOut2_1[31] , 
        \nOut2_15[25] , \nOut0_13[12] , \nScanOut14[21] , \nOut2_10[13] , 
        \nOut2_10[5] , \nScanOut27[12] , \nScanOut32[26] , \nScanOut47[16] , 
        \nScanOut22[24] , \nScanOut37[10] , \nScanOut42[20] , \nScanOut12[9] , 
        \nOut2_13[6] , \nScanOut14[12] , \nScanOut22[17] , \nOut2_10[20] , 
        \nScanOut37[23] , \nScanOut42[13] , \nOut0_3[29] , \nOut1_7[26] , 
        \nScanOut9[14] , \nOut0_13[21] , \nOut0_8[25] , \nOut2_8[1] , 
        \nOut1_3[24] , \nOut1_7[15] , \nScanOut14[7] , \nOut2_15[8] , 
        \nOut0_8[16] , \nScanOut17[4] , \nScanOut29[31] , \nScanOut29[28] , 
        \nScanOut30[1] , \nScanOut33[2] , \nScanOut2[4] , \nScanOut6[29] , 
        \nScanOut6[30] , \nOut1_1[5] , \nOut0_2[23] , \nOut1_3[17] , 
        \nOut0_4[7] , \nOut0_7[18] , \nOut0_7[4] , \nScanOut28[3] , 
        \nScanOut10[23] , \nScanOut26[26] , \nOut2_14[11] , \nScanOut33[12] , 
        \nScanOut46[22] , \nOut0_6[21] , \nScanOut7[23] , \nScanOut7[9] , 
        \nOut1_8[31] , \nOut1_8[28] , \nScanOut10[10] , \nOut2_14[22] , 
        \nScanOut46[11] , \nOut1_13[26] , \nScanOut26[15] , \nScanOut33[21] , 
        \nScanOut39[14] , \nScanOut7[10] , \nOut1_14[2] , \nScanOut23[8] , 
        \nScanOut39[27] , \nOut1_9[22] , \nOut1_13[15] , \nOut2_15[31] , 
        \nOut2_15[28] , \nScanOut42[1] , \nOut0_6[12] , \nOut0_9[2] , 
        \nScanOut11[30] , \nOut2_1[25] , \nScanOut26[5] , \nScanOut41[2] , 
        \nScanOut11[29] , \nScanOut32[18] , \nScanOut47[28] , \nOut1_9[11] , 
        \nScanOut47[31] , \nOut2_1[16] , \nScanOut25[6] , \nOut2_5[27] , 
        \nScanOut38[9] , \nOut0_2[10] , \nOut1_4[8] , \nScanOut15[18] , 
        \nScanOut36[30] , \nScanOut36[29] , \nScanOut43[19] , \nOut0_11[2] , 
        \nOut0_12[18] , \nOut2_5[14] , \nOut2_0[9] , \nOut2_11[19] , 
        \nOut0_2[19] , \nOut1_2[27] , \nOut1_2[6] , \nScanOut3[21] , 
        \nScanOut19[2] , \nScanOut48[26] , \nScanOut3[12] , \nOut0_12[1] , 
        \nScanOut28[22] , \nOut0_6[31] , \nOut0_6[28] , \nOut1_9[18] , 
        \nOut1_11[6] , \nOut2_5[4] , \nOut2_6[7] , \nScanOut28[11] , 
        \nScanOut32[11] , \nScanOut48[15] , \nScanOut11[20] , \nScanOut47[21] , 
        \nOut2_15[12] , \nScanOut11[13] , \nOut1_12[5] , \nScanOut27[25] , 
        \nScanOut27[16] , \nScanOut38[0] , \nScanOut42[8] , \nScanOut32[22] , 
        \nScanOut47[12] , \nOut2_15[21] , \nScanOut9[6] , \nOut1_2[14] , 
        \nScanOut7[19] , \nScanOut20[2] , \nScanOut23[1] , \nScanOut44[6] , 
        \nScanOut3[31] , \nOut1_6[25] , \nOut0_9[26] , \nScanOut47[5] , 
        \nOut0_9[15] , \nScanOut28[18] , \nScanOut3[28] , \nOut1_6[16] , 
        \nOut0_12[8] , \nOut2_3[3] , \nOut1_4[1] , \nOut1_7[2] , 
        \nScanOut8[24] , \nOut0_12[11] , \nScanOut8[17] , \nOut0_12[22] , 
        \nScanOut15[22] , \nScanOut23[27] , \nOut2_11[10] , \nScanOut36[13] , 
        \nScanOut43[23] , \nOut2_0[0] , \nScanOut2[22] , \nOut0_14[6] , 
        \nScanOut15[11] , \nOut2_11[23] , \nScanOut36[20] , \nScanOut43[10] , 
        \nScanOut23[14] , \nScanOut29[21] , \nOut2_8[8] , \nScanOut29[12] , 
        \nOut0_1[26] , \nOut0_1[15] , \nOut0_1[3] , \nScanOut2[11] , 
        \nOut0_3[20] , \nOut1_9[4] , \nScanOut12[0] , \nOut2_10[30] , 
        \nOut2_10[29] , \nOut2_15[1] , \nOut0_3[13] , \nScanOut11[3] , 
        \nOut0_13[31] , \nOut0_13[28] , \nOut2_4[24] , \nScanOut14[31] , 
        \nScanOut14[28] , \nScanOut42[30] , \nOut2_4[17] , \nScanOut37[19] , 
        \nScanOut42[29] , \nScanOut4[3] , \nOut2_0[26] , \nScanOut6[20] , 
        \nOut0_7[22] , \nOut0_7[11] , \nScanOut7[0] , \nOut1_8[21] , 
        \nScanOut10[19] , \nScanOut33[31] , \nScanOut33[28] , \nScanOut46[18] , 
        \nOut1_8[12] , \nOut2_0[15] , \nScanOut35[5] , \nOut2_14[18] , 
        \nOut1_12[25] , \nScanOut36[6] , \nScanOut6[13] , \nScanOut38[17] , 
        \nScanOut0[24] , \nScanOut0[17] , \nOut0_2[0] , \nOut1_12[16] , 
        \nScanOut30[8] , \nOut1_5[30] , \nOut1_5[29] , \nScanOut38[24] , 
        \nOut0_5[3] , \nOut0_6[0] , \nOut1_14[12] , \nScanOut34[8] , 
        \nScanOut29[7] , \nOut1_14[21] , \nScanOut3[0] , \nOut2_6[11] , 
        \nScanOut0[3] , \nScanOut20[18] , \nScanOut32[6] , \nScanOut4[26] , 
        \nScanOut4[15] , \nOut0_5[24] , \nOut0_5[17] , \nOut2_6[22] , 
        \nScanOut31[5] , \nScanOut15[3] , \nScanOut16[0] , \nOut2_2[13] , 
        \nScanOut24[30] , \nScanOut24[29] , \nOut2_2[20] , \nOut2_9[5] , 
        \nOut1_8[9] , \nOut1_10[10] , \nOut1_10[23] , \nScanOut19[13] , 
        \nOut1_0[21] , \nOut1_0[12] , \nOut1_0[1] , \nOut1_1[18] , 
        \nScanOut19[20] , \nOut2_11[1] , \nScanOut13[15] , \nOut2_12[2] , 
        \nScanOut30[24] , \nScanOut45[14] , \nOut0_14[26] , \nOut2_4[0] , 
        \nScanOut25[10] , \nOut2_7[3] , \nOut1_3[2] , \nOut0_10[6] , 
        \nScanOut25[23] , \nScanOut30[17] , \nScanOut45[27] , \nOut0_13[5] , 
        \nScanOut13[26] , \nOut0_14[15] , \nOut2_3[19] , \nScanOut18[6] , 
        \nOut1_11[30] , \nOut1_11[29] , \nOut2_8[15] , \nScanOut18[19] , 
        \nOut0_8[6] , \nOut2_8[26] , \nScanOut27[1] , \nOut1_4[10] , 
        \nOut1_13[8] , \nScanOut24[2] , \nOut1_15[18] , \nScanOut43[5] , 
        \nOut0_0[25] , \nOut0_0[16] , \nOut1_0[31] , \nOut1_4[23] , 
        \nScanOut40[6] , \nOut1_6[6] , \nOut0_10[24] , \nOut0_10[17] , 
        \nOut1_15[6] , \nOut2_7[31] , \nOut2_7[28] , \nScanOut17[17] , 
        \nScanOut21[12] , \nOut2_13[25] , \nScanOut34[26] , \nScanOut41[16] , 
        \nScanOut17[24] , \nOut2_13[16] , \nScanOut34[15] , \nScanOut41[25] , 
        \nScanOut46[8] , \nScanOut21[21] , \nOut1_0[28] , \nOut1_0[8] , 
        \nOut1_5[5] , \nScanOut5[16] , \nOut0_15[2] , \nScanOut18[10] , 
        \nScanOut5[25] , \nOut1_11[20] , \nOut1_11[13] , \nOut2_1[4] , 
        \nOut2_2[7] , \nScanOut18[23] , \nOut0_4[27] , \nOut0_4[14] , 
        \nOut2_3[10] , \nOut2_4[9] , \nScanOut25[19] , \nOut2_3[23] , 
        \nScanOut21[31] , \nOut2_7[12] , \nScanOut45[2] , \nScanOut21[28] , 
        \nScanOut21[6] , \nOut2_7[21] , \nScanOut46[1] , \nScanOut1[14] , 
        \nScanOut22[5] , \nOut1_15[11] , \nScanOut1[27] , \nScanOut8[2] , 
        \nOut1_10[2] , \nScanOut27[8] , \nOut1_15[22] , \nOut0_0[31] , 
        \nOut0_0[7] , \nOut1_4[19] , \nScanOut39[4] , \nOut1_13[1] , 
        \nScanOut16[14] , \nOut2_12[26] , \nScanOut20[11] , \nScanOut35[25] , 
        \nScanOut40[15] , \nOut1_1[22] , \nOut1_1[11] , \nOut0_3[4] , 
        \nScanOut3[9] , \nOut0_11[27] , \nOut1_5[20] , \nOut1_5[13] , 
        \nOut0_6[9] , \nOut0_11[14] , \nScanOut16[27] , \nScanOut20[22] , 
        \nOut2_12[15] , \nScanOut35[16] , \nScanOut40[26] , \nOut2_6[18] , 
        \nScanOut34[1] , \nScanOut48[7] , \nOut1_14[31] , \nOut1_14[28] , 
        \nScanOut37[2] , \nScanOut5[7] , \nScanOut6[4] , \nScanOut19[29] , 
        \nOut2_9[16] , \nOut2_11[8] , \nOut1_8[0] , \nOut1_10[19] , 
        \nScanOut19[30] , \nOut2_9[25] , \nScanOut10[7] , \nScanOut13[4] , 
        \nScanOut12[25] , \nScanOut12[16] , \nOut0_15[25] , \nOut2_2[30] , 
        \nOut2_2[29] , \nScanOut24[13] , \nOut2_14[5] , \nOut0_15[16] , 
        \nScanOut31[27] , \nScanOut44[17] , \nOut1_15[2] , \nScanOut16[9] , 
        \nScanOut31[14] , \nScanOut17[13] , \nScanOut24[20] , \nScanOut44[24] , 
        \nScanOut22[8] , \nOut2_13[21] , \nScanOut34[22] , \nScanOut41[12] , 
        \nScanOut21[16] , \nOut0_0[28] , \nOut1_4[14] , \nOut0_10[20] , 
        \nOut0_10[13] , \nScanOut17[20] , \nScanOut21[25] , \nOut2_13[12] , 
        \nScanOut34[11] , \nScanOut41[21] , \nScanOut24[6] , \nScanOut39[9] , 
        \nOut1_4[27] , \nOut0_8[2] , \nScanOut27[5] , \nScanOut40[2] , 
        \nOut1_0[25] , \nOut1_0[16] , \nScanOut1[19] , \nScanOut43[1] , 
        \nScanOut5[31] , \nScanOut5[28] , \nOut2_8[11] , \nOut2_1[9] , 
        \nOut1_5[8] , \nOut2_8[22] , \nOut1_0[5] , \nOut1_3[6] , 
        \nScanOut13[11] , \nOut0_14[22] , \nOut2_4[4] , \nOut2_7[7] , 
        \nScanOut25[14] , \nScanOut18[2] , \nScanOut30[20] , \nScanOut45[10] , 
        \nOut0_4[19] , \nOut0_10[2] , \nOut0_13[1] , \nScanOut13[22] , 
        \nOut0_14[11] , \nScanOut30[13] , \nScanOut45[23] , \nScanOut25[27] , 
        \nScanOut4[11] , \nScanOut13[9] , \nScanOut19[17] , \nOut1_10[14] , 
        \nScanOut19[24] , \nOut2_9[31] , \nOut2_9[28] , \nOut2_12[6] , 
        \nOut0_0[3] , \nOut0_1[22] , \nOut0_1[11] , \nScanOut0[7] , 
        \nScanOut4[22] , \nOut1_10[27] , \nOut2_11[5] , \nOut0_5[20] , 
        \nOut0_5[13] , \nScanOut12[31] , \nScanOut31[19] , \nScanOut12[28] , 
        \nScanOut16[4] , \nScanOut44[29] , \nScanOut15[7] , \nScanOut44[30] , 
        \nOut2_2[17] , \nOut2_9[1] , \nOut2_14[8] , \nOut0_15[31] , 
        \nOut0_15[28] , \nOut2_2[24] , \nScanOut3[4] , \nOut0_11[19] , 
        \nOut2_6[15] , \nOut2_12[18] , \nOut2_6[26] , \nScanOut31[1] , 
        \nOut1_1[26] , \nOut1_1[15] , \nScanOut0[20] , \nScanOut0[13] , 
        \nOut0_3[9] , \nScanOut6[9] , \nScanOut16[19] , \nScanOut35[28] , 
        \nScanOut40[18] , \nScanOut32[2] , \nScanOut35[31] , \nOut1_14[25] , 
        \nOut1_14[16] , \nOut0_5[30] , \nOut0_5[29] , \nOut0_5[7] , 
        \nOut0_6[4] , \nScanOut29[3] , \nScanOut12[12] , \nOut2_9[8] , 
        \nScanOut44[13] , \nScanOut31[23] , \nScanOut24[17] , \nOut2_14[1] , 
        \nScanOut12[21] , \nOut0_15[21] , \nScanOut24[24] , \nScanOut31[10] , 
        \nScanOut44[20] , \nOut0_15[12] , \nOut2_9[12] , \nScanOut0[30] , 
        \nScanOut4[18] , \nOut1_8[4] , \nScanOut10[3] , \nScanOut13[0] , 
        \nOut2_9[21] , \nScanOut37[6] , \nScanOut0[29] , \nOut0_3[0] , 
        \nOut1_5[24] , \nOut1_5[17] , \nScanOut5[3] , \nScanOut6[0] , 
        \nScanOut34[5] , \nOut0_11[23] , \nScanOut31[8] , \nOut0_1[18] , 
        \nScanOut16[10] , \nScanOut20[15] , \nScanOut35[21] , \nScanOut40[11] , 
        \nOut2_12[22] , \nScanOut1[10] , \nScanOut8[6] , \nOut0_11[10] , 
        \nScanOut48[3] , \nScanOut16[23] , \nScanOut35[12] , \nScanOut40[22] , 
        \nScanOut20[26] , \nOut2_12[11] , \nScanOut43[8] , \nOut1_13[5] , 
        \nOut1_15[15] , \nScanOut39[0] , \nOut0_0[21] , \nOut0_0[12] , 
        \nScanOut1[23] , \nOut1_15[26] , \nOut1_10[6] , \nScanOut17[30] , 
        \nScanOut17[29] , \nScanOut34[18] , \nScanOut41[31] , \nOut2_7[16] , 
        \nScanOut41[28] , \nScanOut46[5] , \nScanOut45[6] , \nScanOut22[1] , 
        \nOut2_13[31] , \nOut2_13[28] , \nOut0_4[10] , \nOut0_10[30] , 
        \nOut0_10[29] , \nScanOut21[2] , \nOut2_7[25] , \nOut0_14[18] , 
        \nScanOut1[21] , \nScanOut1[12] , \nOut0_4[23] , \nOut0_13[8] , 
        \nOut2_3[14] , \nOut2_3[27] , \nOut1_5[1] , \nScanOut5[12] , 
        \nScanOut13[18] , \nScanOut30[30] , \nScanOut30[29] , \nScanOut45[19] , 
        \nScanOut5[21] , \nOut1_6[2] , \nOut1_11[17] , \nOut0_15[6] , 
        \nScanOut18[14] , \nOut1_11[24] , \nOut1_15[17] , \nOut2_1[0] , 
        \nOut2_2[3] , \nOut2_8[18] , \nScanOut18[27] , \nOut0_8[9] , 
        \nScanOut8[4] , \nOut1_10[4] , \nScanOut40[9] , \nOut1_15[24] , 
        \nOut0_0[23] , \nOut0_0[10] , \nOut1_13[7] , \nScanOut39[2] , 
        \nOut0_10[18] , \nScanOut21[0] , \nOut2_7[27] , \nOut2_7[14] , 
        \nOut2_13[19] , \nScanOut45[4] , \nScanOut46[7] , \nOut0_4[21] , 
        \nOut0_4[12] , \nOut0_10[9] , \nScanOut13[29] , \nOut1_15[9] , 
        \nScanOut17[18] , \nScanOut34[30] , \nScanOut34[29] , \nScanOut41[19] , 
        \nScanOut22[3] , \nScanOut45[31] , \nScanOut45[28] , \nScanOut13[30] , 
        \nScanOut18[9] , \nOut2_3[16] , \nScanOut30[18] , \nOut0_5[18] , 
        \nOut1_5[3] , \nOut1_6[0] , \nOut0_14[30] , \nOut0_14[29] , 
        \nOut2_3[25] , \nOut1_11[15] , \nOut0_15[4] , \nScanOut18[16] , 
        \nScanOut5[23] , \nScanOut5[10] , \nOut2_2[1] , \nScanOut18[25] , 
        \nOut2_8[30] , \nOut2_8[29] , \nOut1_11[26] , \nScanOut12[10] , 
        \nOut0_15[23] , \nOut2_1[2] , \nScanOut24[15] , \nOut2_14[3] , 
        \nScanOut31[21] , \nScanOut44[11] , \nScanOut12[23] , \nOut0_15[10] , 
        \nScanOut31[12] , \nScanOut44[22] , \nScanOut24[26] , \nOut0_0[1] , 
        \nOut1_1[24] , \nOut1_1[17] , \nScanOut4[30] , \nOut2_9[10] , 
        \nScanOut4[29] , \nOut1_8[6] , \nScanOut13[2] , \nOut2_9[23] , 
        \nScanOut10[1] , \nScanOut0[18] , \nOut1_5[26] , \nOut1_5[15] , 
        \nScanOut29[8] , \nScanOut34[7] , \nScanOut5[1] , \nScanOut37[4] , 
        \nScanOut6[2] , \nScanOut16[12] , \nOut2_12[20] , \nScanOut35[23] , 
        \nScanOut40[13] , \nScanOut20[17] , \nScanOut32[9] , \nOut0_1[30] , 
        \nOut0_1[29] , \nOut0_3[2] , \nScanOut4[20] , \nScanOut4[13] , 
        \nOut1_10[16] , \nOut0_11[21] , \nOut0_11[12] , \nScanOut16[21] , 
        \nScanOut20[24] , \nOut2_12[13] , \nScanOut35[10] , \nScanOut40[20] , 
        \nScanOut48[1] , \nScanOut10[8] , \nScanOut19[15] , \nOut1_10[25] , 
        \nOut0_5[11] , \nScanOut19[26] , \nOut2_9[19] , \nOut2_11[7] , 
        \nOut2_12[4] , \nOut0_15[19] , \nScanOut15[5] , \nOut2_2[15] , 
        \nScanOut16[6] , \nOut2_2[26] , \nOut0_0[19] , \nOut0_0[8] , 
        \nOut0_1[13] , \nScanOut3[6] , \nOut0_5[22] , \nScanOut12[19] , 
        \nOut2_9[3] , \nScanOut31[28] , \nScanOut44[18] , \nScanOut31[31] , 
        \nScanOut16[31] , \nScanOut40[29] , \nScanOut16[28] , \nScanOut35[19] , 
        \nScanOut40[30] , \nOut2_6[17] , \nScanOut0[5] , \nScanOut48[8] , 
        \nOut2_12[30] , \nScanOut32[0] , \nOut2_12[29] , \nOut0_1[20] , 
        \nScanOut0[22] , \nScanOut0[11] , \nScanOut5[8] , \nOut0_11[31] , 
        \nOut0_11[28] , \nScanOut31[3] , \nOut2_6[24] , \nOut1_14[14] , 
        \nOut0_5[5] , \nOut0_6[6] , \nScanOut29[1] , \nOut0_10[22] , 
        \nOut1_14[27] , \nOut1_15[0] , \nScanOut21[9] , \nScanOut17[11] , 
        \nScanOut21[14] , \nOut2_13[23] , \nScanOut34[20] , \nScanOut41[10] , 
        \nOut0_8[0] , \nOut0_10[11] , \nScanOut17[22] , \nOut2_13[10] , 
        \nScanOut21[27] , \nScanOut34[13] , \nScanOut41[23] , \nScanOut27[7] , 
        \nScanOut1[31] , \nScanOut1[28] , \nOut1_4[16] , \nScanOut24[4] , 
        \nOut0_0[27] , \nOut0_0[14] , \nOut0_0[5] , \nOut1_0[27] , 
        \nOut1_0[14] , \nOut1_4[25] , \nScanOut40[0] , \nScanOut43[3] , 
        \nOut2_2[8] , \nOut2_8[13] , \nOut1_0[7] , \nOut0_4[31] , 
        \nScanOut5[19] , \nOut1_6[9] , \nOut2_8[20] , \nScanOut13[13] , 
        \nOut2_4[6] , \nScanOut25[16] , \nScanOut30[22] , \nScanOut45[12] , 
        \nOut0_4[28] , \nOut2_7[5] , \nOut0_14[20] , \nOut0_3[6] , 
        \nOut1_3[4] , \nOut0_10[0] , \nScanOut13[20] , \nScanOut25[25] , 
        \nScanOut45[21] , \nOut0_13[3] , \nOut0_14[13] , \nScanOut30[11] , 
        \nScanOut18[0] , \nOut0_11[25] , \nOut2_6[30] , \nOut2_6[29] , 
        \nOut1_0[19] , \nOut1_1[20] , \nOut1_1[13] , \nScanOut0[8] , 
        \nScanOut16[16] , \nScanOut20[13] , \nOut2_12[24] , \nScanOut35[27] , 
        \nScanOut40[17] , \nScanOut48[5] , \nOut0_5[8] , \nOut0_11[16] , 
        \nScanOut16[25] , \nScanOut20[20] , \nOut2_12[17] , \nScanOut35[14] , 
        \nScanOut40[24] , \nScanOut37[0] , \nOut1_5[22] , \nOut1_5[11] , 
        \nScanOut6[6] , \nOut1_14[19] , \nScanOut34[3] , \nScanOut5[5] , 
        \nOut2_12[9] , \nOut1_10[31] , \nOut1_10[28] , \nScanOut19[18] , 
        \nOut2_9[14] , \nOut1_5[7] , \nOut1_8[2] , \nScanOut10[5] , 
        \nOut1_11[11] , \nScanOut12[27] , \nScanOut12[14] , \nScanOut13[6] , 
        \nOut2_9[27] , \nOut0_15[27] , \nScanOut24[11] , \nScanOut31[25] , 
        \nScanOut44[15] , \nOut2_14[7] , \nScanOut24[22] , \nOut0_15[14] , 
        \nScanOut31[16] , \nScanOut44[26] , \nScanOut15[8] , \nOut2_2[18] , 
        \nScanOut5[27] , \nScanOut5[14] , \nOut1_6[4] , \nOut0_15[0] , 
        \nScanOut18[12] , \nOut2_1[6] , \nOut1_11[22] , \nOut2_2[5] , 
        \nOut1_3[9] , \nOut0_4[16] , \nScanOut18[21] , \nOut0_4[25] , 
        \nOut2_3[21] , \nOut2_3[12] , \nScanOut25[31] , \nScanOut25[28] , 
        \nOut2_7[10] , \nOut2_7[8] , \nScanOut46[3] , \nScanOut45[0] , 
        \nScanOut21[19] , \nScanOut22[7] , \nScanOut1[16] , \nOut1_4[31] , 
        \nScanOut21[4] , \nOut2_7[23] , \nOut1_4[28] , \nScanOut8[0] , 
        \nOut1_15[13] , \nOut1_13[3] , \nScanOut24[9] , \nScanOut39[6] , 
        \nScanOut1[25] , \nOut1_10[0] , \nOut1_15[20] , \nOut1_0[23] , 
        \nOut1_0[10] , \nOut1_0[3] , \nOut1_3[0] , \nScanOut13[17] , 
        \nOut0_14[24] , \nOut2_3[31] , \nOut2_3[28] , \nOut2_4[2] , 
        \nOut2_7[1] , \nScanOut25[12] , \nScanOut30[26] , \nScanOut45[16] , 
        \nOut0_10[4] , \nOut0_13[7] , \nScanOut18[4] , \nOut0_14[17] , 
        \nScanOut45[25] , \nScanOut13[24] , \nScanOut30[15] , \nScanOut25[21] , 
        \nScanOut18[31] , \nOut2_8[17] , \nOut1_11[18] , \nScanOut18[28] , 
        \nOut0_15[9] , \nOut2_8[24] , \nScanOut24[0] , \nOut1_4[12] , 
        \nOut1_15[30] , \nOut1_15[29] , \nOut1_4[21] , \nOut0_8[4] , 
        \nOut1_10[9] , \nScanOut27[3] , \nScanOut8[9] , \nScanOut40[4] , 
        \nScanOut43[7] , \nOut0_1[24] , \nOut0_1[17] , \nScanOut0[26] , 
        \nScanOut0[15] , \nOut0_10[26] , \nOut1_15[4] , \nScanOut17[15] , 
        \nScanOut34[24] , \nScanOut41[14] , \nOut2_13[27] , \nScanOut21[10] , 
        \nOut0_10[15] , \nScanOut17[26] , \nScanOut21[23] , \nScanOut34[17] , 
        \nScanOut41[27] , \nOut2_13[14] , \nOut1_14[10] , \nOut2_7[19] , 
        \nScanOut45[9] , \nScanOut37[9] , \nScanOut0[1] , \nOut0_5[1] , 
        \nOut1_14[23] , \nOut1_5[18] , \nOut0_6[2] , \nScanOut29[5] , 
        \nScanOut3[2] , \nScanOut20[30] , \nScanOut20[29] , \nOut2_6[13] , 
        \nOut2_6[20] , \nScanOut31[7] , \nOut1_1[30] , \nOut1_1[29] , 
        \nOut0_5[26] , \nOut0_5[15] , \nScanOut15[1] , \nScanOut16[2] , 
        \nScanOut32[4] , \nOut2_2[11] , \nScanOut24[18] , \nOut2_9[7] , 
        \nOut2_2[22] , \nScanOut19[11] , \nScanOut4[17] , \nOut1_10[12] , 
        \nScanOut19[22] , \nOut2_12[0] , \nOut0_0[4] , \nScanOut4[24] , 
        \nOut2_11[3] , \nOut0_5[9] , \nOut1_5[10] , \nOut1_10[21] , 
        \nScanOut34[2] , \nScanOut37[1] , \nOut1_5[23] , \nScanOut5[4] , 
        \nScanOut6[7] , \nOut1_14[18] , \nOut1_0[18] , \nOut1_1[21] , 
        \nOut1_1[12] , \nScanOut0[9] , \nOut0_3[7] , \nOut0_11[24] , 
        \nScanOut16[17] , \nOut2_12[25] , \nScanOut35[26] , \nScanOut40[16] , 
        \nScanOut20[12] , \nOut2_6[31] , \nOut2_6[28] , \nScanOut16[24] , 
        \nScanOut20[21] , \nOut2_12[16] , \nScanOut35[15] , \nScanOut40[25] , 
        \nOut1_10[30] , \nOut0_11[17] , \nScanOut48[4] , \nScanOut12[26] , 
        \nScanOut12[15] , \nOut0_15[26] , \nScanOut24[10] , \nScanOut31[24] , 
        \nScanOut44[14] , \nOut0_15[15] , \nScanOut15[9] , \nOut2_2[19] , 
        \nOut2_14[6] , \nScanOut31[17] , \nScanOut44[27] , \nScanOut24[23] , 
        \nOut2_9[15] , \nOut1_10[29] , \nOut1_8[3] , \nScanOut13[7] , 
        \nOut2_12[8] , \nScanOut19[19] , \nOut2_9[26] , \nOut1_3[8] , 
        \nOut0_4[17] , \nScanOut10[4] , \nScanOut25[30] , \nScanOut25[29] , 
        \nOut0_4[24] , \nOut2_3[20] , \nOut2_3[13] , \nOut2_7[9] , 
        \nOut1_5[6] , \nScanOut5[15] , \nOut1_6[5] , \nOut1_11[10] , 
        \nScanOut18[13] , \nOut0_15[1] , \nScanOut1[24] , \nScanOut1[17] , 
        \nScanOut5[26] , \nOut2_2[4] , \nScanOut18[20] , \nOut1_11[23] , 
        \nOut1_15[12] , \nOut2_1[7] , \nOut1_4[30] , \nOut1_4[29] , 
        \nScanOut8[1] , \nOut1_15[21] , \nOut1_10[1] , \nOut1_13[2] , 
        \nScanOut24[8] , \nOut0_0[26] , \nOut0_0[15] , \nOut2_7[11] , 
        \nScanOut39[7] , \nScanOut45[1] , \nScanOut46[2] , \nOut1_0[22] , 
        \nOut1_0[11] , \nScanOut21[18] , \nScanOut21[5] , \nOut2_7[22] , 
        \nScanOut22[6] , \nScanOut18[30] , \nScanOut18[29] , \nOut2_8[16] , 
        \nOut1_0[2] , \nOut0_10[5] , \nOut1_11[19] , \nOut2_8[25] , 
        \nScanOut13[25] , \nScanOut13[16] , \nOut0_15[8] , \nOut2_4[3] , 
        \nOut0_14[25] , \nOut2_3[30] , \nOut2_3[29] , \nScanOut25[13] , 
        \nScanOut30[27] , \nScanOut45[17] , \nOut2_7[0] , \nScanOut25[20] , 
        \nScanOut30[14] , \nScanOut45[24] , \nOut1_3[1] , \nScanOut18[5] , 
        \nOut0_8[5] , \nOut0_10[27] , \nOut0_13[6] , \nOut0_14[16] , 
        \nOut0_10[14] , \nOut1_15[5] , \nScanOut21[11] , \nScanOut17[14] , 
        \nOut2_13[26] , \nOut2_7[18] , \nScanOut34[25] , \nScanOut41[15] , 
        \nScanOut45[8] , \nOut1_10[8] , \nOut1_15[31] , \nOut1_15[28] , 
        \nScanOut17[27] , \nOut2_13[15] , \nScanOut21[22] , \nScanOut34[16] , 
        \nScanOut41[26] , \nScanOut27[2] , \nOut1_4[13] , \nScanOut24[1] , 
        \nOut0_1[25] , \nOut0_1[16] , \nScanOut3[3] , \nOut1_4[20] , 
        \nScanOut43[6] , \nScanOut8[8] , \nScanOut40[5] , \nScanOut20[31] , 
        \nScanOut20[28] , \nScanOut0[0] , \nOut2_6[21] , \nOut2_6[12] , 
        \nScanOut31[6] , \nScanOut32[5] , \nOut1_1[31] , \nScanOut0[27] , 
        \nScanOut0[14] , \nOut1_14[11] , \nOut0_5[0] , \nOut1_5[19] , 
        \nOut0_6[3] , \nScanOut29[4] , \nScanOut37[8] , \nScanOut4[16] , 
        \nOut1_10[13] , \nOut1_14[22] , \nOut1_1[28] , \nScanOut19[10] , 
        \nScanOut4[25] , \nOut1_10[20] , \nOut2_11[2] , \nOut0_0[22] , 
        \nOut0_0[11] , \nOut0_5[27] , \nOut0_5[14] , \nScanOut15[0] , 
        \nOut2_2[10] , \nScanOut19[23] , \nOut2_12[1] , \nScanOut16[3] , 
        \nOut2_2[23] , \nScanOut24[19] , \nOut2_9[6] , \nOut2_13[18] , 
        \nScanOut46[6] , \nOut0_10[19] , \nOut2_7[15] , \nScanOut45[5] , 
        \nOut1_15[8] , \nScanOut17[19] , \nScanOut22[2] , \nScanOut34[31] , 
        \nScanOut34[28] , \nScanOut41[18] , \nScanOut21[1] , \nOut2_7[26] , 
        \nScanOut1[13] , \nScanOut8[5] , \nScanOut40[8] , \nOut1_15[16] , 
        \nScanOut39[3] , \nOut1_1[16] , \nScanOut1[20] , \nOut0_8[8] , 
        \nOut1_13[6] , \nOut1_10[5] , \nOut0_4[20] , \nOut0_4[13] , 
        \nOut1_5[2] , \nScanOut5[11] , \nOut1_11[14] , \nOut0_15[5] , 
        \nOut1_15[25] , \nOut2_8[31] , \nOut2_8[28] , \nScanOut5[22] , 
        \nOut1_6[1] , \nScanOut18[17] , \nOut2_1[3] , \nOut1_11[27] , 
        \nOut2_2[0] , \nScanOut18[24] , \nOut2_3[17] , \nOut0_10[8] , 
        \nScanOut18[8] , \nScanOut13[31] , \nScanOut45[29] , \nScanOut13[28] , 
        \nScanOut30[19] , \nScanOut45[30] , \nOut0_14[31] , \nOut2_3[24] , 
        \nOut0_14[28] , \nScanOut4[31] , \nScanOut4[28] , \nOut2_9[11] , 
        \nOut0_0[0] , \nOut0_1[31] , \nOut1_1[25] , \nScanOut10[0] , 
        \nOut0_3[3] , \nOut0_5[19] , \nOut1_8[7] , \nOut2_9[22] , 
        \nScanOut12[22] , \nScanOut12[11] , \nScanOut13[3] , \nOut2_14[2] , 
        \nOut0_15[22] , \nScanOut24[14] , \nScanOut31[20] , \nScanOut44[10] , 
        \nScanOut24[27] , \nScanOut31[13] , \nScanOut44[23] , \nOut0_15[11] , 
        \nOut0_1[28] , \nOut0_11[20] , \nScanOut16[13] , \nScanOut20[16] , 
        \nScanOut32[8] , \nOut2_12[21] , \nScanOut35[22] , \nScanOut40[12] , 
        \nScanOut0[19] , \nOut1_5[14] , \nOut0_11[13] , \nScanOut16[20] , 
        \nScanOut48[0] , \nScanOut20[25] , \nOut2_12[12] , \nScanOut35[11] , 
        \nScanOut40[21] , \nScanOut34[6] , \nScanOut37[5] , \nScanOut29[9] , 
        \nScanOut4[12] , \nOut0_5[23] , \nOut0_5[10] , \nOut1_5[27] , 
        \nScanOut6[3] , \nScanOut5[0] , \nScanOut16[7] , \nScanOut12[18] , 
        \nOut0_15[18] , \nScanOut15[4] , \nOut2_2[14] , \nScanOut31[30] , 
        \nOut2_2[27] , \nOut2_9[2] , \nScanOut31[29] , \nScanOut44[19] , 
        \nOut1_10[17] , \nScanOut10[9] , \nScanOut19[14] , \nScanOut19[27] , 
        \nOut2_12[5] , \nOut2_9[18] , \nOut2_11[6] , \nOut0_0[9] , 
        \nOut0_1[21] , \nOut0_1[12] , \nScanOut0[23] , \nScanOut0[10] , 
        \nScanOut4[21] , \nOut1_10[24] , \nOut1_14[15] , \nScanOut5[9] , 
        \nScanOut0[4] , \nOut0_5[4] , \nOut1_14[26] , \nOut0_6[7] , 
        \nOut2_6[16] , \nScanOut29[0] , \nScanOut48[9] , \nScanOut3[7] , 
        \nScanOut16[30] , \nScanOut16[29] , \nScanOut40[31] , \nScanOut40[28] , 
        \nScanOut35[18] , \nOut0_11[30] , \nOut0_11[29] , \nOut2_6[25] , 
        \nScanOut31[2] , \nOut2_12[31] , \nOut2_12[28] , \nScanOut32[1] , 
        \nOut1_4[17] , \nScanOut24[5] , \nScanOut1[30] , \nOut0_8[1] , 
        \nScanOut27[6] , \nScanOut1[29] , \nOut1_4[24] , \nScanOut40[1] , 
        \nScanOut43[2] , \nOut0_0[18] , \nOut0_10[23] , \nOut1_15[1] , 
        \nScanOut17[10] , \nScanOut34[21] , \nScanOut41[11] , \nScanOut21[15] , 
        \nOut2_13[22] , \nScanOut21[8] , \nScanOut17[23] , \nScanOut21[26] , 
        \nScanOut34[12] , \nScanOut41[22] , \nOut2_13[11] , \nOut1_0[26] , 
        \nOut1_0[15] , \nOut1_0[6] , \nOut1_3[5] , \nOut0_4[30] , 
        \nOut0_4[29] , \nOut0_10[10] , \nOut0_13[2] , \nScanOut13[12] , 
        \nOut0_14[21] , \nOut2_7[4] , \nScanOut25[17] , \nScanOut30[23] , 
        \nScanOut45[13] , \nOut2_4[7] , \nOut0_14[12] , \nScanOut18[1] , 
        \nOut0_10[1] , \nScanOut13[21] , \nScanOut30[10] , \nScanOut45[20] , 
        \nOut2_8[12] , \nScanOut25[24] , \nScanOut5[18] , \nOut2_2[9] , 
        \nOut1_6[8] , \nOut2_8[21] , \nOut0_8[3] , \nScanOut27[4] , 
        \nOut1_4[15] , \nScanOut24[7] , \nScanOut39[8] , \nScanOut43[0] , 
        \nOut0_0[30] , \nOut0_0[29] , \nScanOut1[18] , \nOut1_4[26] , 
        \nScanOut40[3] , \nOut1_0[24] , \nOut1_0[17] , \nOut1_0[4] , 
        \nOut0_10[21] , \nOut0_10[12] , \nOut1_15[3] , \nScanOut21[17] , 
        \nScanOut22[9] , \nScanOut17[12] , \nOut2_13[20] , \nScanOut34[23] , 
        \nScanOut41[13] , \nOut0_10[3] , \nScanOut13[10] , \nScanOut17[21] , 
        \nOut2_13[13] , \nScanOut34[10] , \nScanOut41[20] , \nOut2_4[5] , 
        \nScanOut21[24] , \nScanOut30[21] , \nScanOut45[11] , \nOut0_14[23] , 
        \nScanOut25[15] , \nOut2_7[6] , \nScanOut25[26] , \nScanOut30[12] , 
        \nScanOut13[23] , \nScanOut45[22] , \nOut1_3[7] , \nOut0_4[18] , 
        \nOut0_13[0] , \nOut0_14[10] , \nScanOut18[3] , \nScanOut5[30] , 
        \nOut2_1[8] , \nScanOut5[29] , \nOut2_8[10] , \nScanOut4[23] , 
        \nScanOut4[10] , \nOut0_5[21] , \nOut0_5[12] , \nOut1_5[9] , 
        \nOut2_8[23] , \nScanOut15[6] , \nOut2_2[16] , \nScanOut12[30] , 
        \nScanOut12[29] , \nScanOut16[5] , \nScanOut44[31] , \nScanOut31[18] , 
        \nScanOut44[28] , \nScanOut13[8] , \nOut0_15[30] , \nOut0_15[29] , 
        \nOut2_2[25] , \nOut2_9[0] , \nOut2_14[9] , \nOut2_9[30] , 
        \nOut2_9[29] , \nOut1_10[26] , \nOut1_10[15] , \nScanOut19[16] , 
        \nOut2_11[4] , \nOut0_0[13] , \nOut0_0[2] , \nOut0_1[23] , 
        \nOut0_1[10] , \nScanOut0[21] , \nScanOut0[12] , \nScanOut19[25] , 
        \nOut2_12[7] , \nOut0_5[6] , \nOut0_6[5] , \nScanOut6[8] , 
        \nOut1_14[17] , \nScanOut29[2] , \nOut1_14[24] , \nScanOut3[5] , 
        \nOut2_12[19] , \nScanOut0[6] , \nOut0_3[8] , \nOut0_11[18] , 
        \nOut2_6[14] , \nScanOut16[18] , \nScanOut32[3] , \nOut2_6[27] , 
        \nScanOut31[0] , \nScanOut35[30] , \nScanOut35[29] , \nScanOut40[19] , 
        \nOut1_1[27] , \nOut1_1[14] , \nOut2_9[13] , \nScanOut4[19] , 
        \nOut1_8[5] , \nScanOut13[1] , \nOut2_9[20] , \nOut0_5[31] , 
        \nScanOut10[2] , \nOut0_5[28] , \nScanOut12[20] , \nScanOut12[13] , 
        \nOut0_15[20] , \nScanOut24[16] , \nOut0_15[13] , \nOut2_9[9] , 
        \nOut2_14[0] , \nScanOut31[22] , \nScanOut44[12] , \nScanOut24[25] , 
        \nScanOut31[11] , \nScanOut44[21] , \nOut0_1[19] , \nOut0_3[1] , 
        \nOut0_11[22] , \nScanOut16[11] , \nOut2_12[23] , \nScanOut20[14] , 
        \nScanOut35[20] , \nScanOut40[10] , \nScanOut31[9] , \nScanOut16[22] , 
        \nScanOut20[27] , \nOut2_12[10] , \nScanOut35[13] , \nScanOut40[23] , 
        \nScanOut48[2] , \nScanOut0[31] , \nScanOut0[28] , \nOut1_5[16] , 
        \nOut0_11[11] , \nScanOut34[4] , \nScanOut37[7] , \nOut1_5[25] , 
        \nScanOut5[2] , \nScanOut6[1] , \nOut2_7[17] , \nScanOut45[7] , 
        \nOut0_0[20] , \nScanOut17[31] , \nScanOut34[19] , \nScanOut46[4] , 
        \nScanOut17[28] , \nScanOut41[29] , \nScanOut41[30] , \nScanOut1[22] , 
        \nScanOut1[11] , \nOut0_10[31] , \nOut2_7[24] , \nOut0_10[28] , 
        \nScanOut21[3] , \nScanOut22[0] , \nOut2_13[30] , \nOut2_13[29] , 
        \nScanOut43[9] , \nScanOut8[7] , \nOut1_15[14] , \nOut1_15[27] , 
        \nOut1_10[7] , \nOut1_13[4] , \nOut0_1[27] , \nOut0_1[14] , 
        \nScanOut0[2] , \nOut0_4[22] , \nOut0_4[11] , \nOut1_5[0] , 
        \nOut1_6[3] , \nScanOut39[1] , \nScanOut18[15] , \nScanOut5[20] , 
        \nScanOut5[13] , \nOut1_11[25] , \nOut1_11[16] , \nOut0_15[7] , 
        \nOut2_1[1] , \nOut2_2[2] , \nScanOut18[26] , \nOut2_8[19] , 
        \nOut0_13[9] , \nOut2_3[15] , \nScanOut13[19] , \nOut0_14[19] , 
        \nScanOut30[28] , \nScanOut45[18] , \nOut2_3[26] , \nScanOut30[31] , 
        \nOut2_6[10] , \nScanOut3[1] , \nOut1_1[19] , \nScanOut0[25] , 
        \nScanOut0[16] , \nScanOut20[19] , \nOut2_6[23] , \nScanOut31[4] , 
        \nScanOut32[7] , \nOut1_5[31] , \nOut1_14[13] , \nOut1_5[28] , 
        \nOut1_14[20] , \nScanOut4[14] , \nOut0_5[2] , \nOut0_6[1] , 
        \nScanOut29[6] , \nScanOut34[9] , \nScanOut19[12] , \nOut1_8[8] , 
        \nOut1_10[11] , \nScanOut19[21] , \nOut2_12[3] , \nOut2_11[0] , 
        \nOut1_0[20] , \nOut1_0[13] , \nScanOut4[27] , \nOut1_10[22] , 
        \nOut0_5[25] , \nOut0_5[16] , \nScanOut16[1] , \nScanOut24[31] , 
        \nScanOut24[28] , \nScanOut15[2] , \nOut2_2[21] , \nOut2_2[12] , 
        \nOut2_9[4] , \nOut1_11[31] , \nOut1_11[28] , \nOut2_8[14] , 
        \nOut2_8[27] , \nOut1_0[0] , \nOut1_3[3] , \nOut0_13[4] , 
        \nScanOut13[14] , \nOut0_14[27] , \nScanOut18[18] , \nOut2_7[2] , 
        \nScanOut25[11] , \nOut2_4[1] , \nScanOut30[25] , \nScanOut45[15] , 
        \nOut0_14[14] , \nOut2_3[18] , \nScanOut18[7] , \nOut1_4[11] , 
        \nOut0_10[25] , \nOut0_10[7] , \nScanOut13[27] , \nScanOut30[16] , 
        \nOut1_15[7] , \nScanOut17[16] , \nScanOut25[22] , \nScanOut45[26] , 
        \nScanOut21[13] , \nOut2_13[24] , \nScanOut34[27] , \nScanOut41[17] , 
        \nOut2_7[30] , \nOut2_7[29] , \nOut0_10[16] , \nScanOut17[25] , 
        \nScanOut21[20] , \nOut2_13[17] , \nScanOut34[14] , \nScanOut46[9] , 
        \nScanOut41[24] , \nOut1_13[9] , \nScanOut24[3] , \nOut1_4[22] , 
        \nOut0_8[7] , \nScanOut27[0] , \nScanOut40[7] , \nOut1_15[19] , 
        \nOut1_0[30] , \nOut1_0[29] , \nOut1_0[9] , \nOut0_4[15] , 
        \nOut2_3[11] , \nScanOut43[4] , \nOut0_4[26] , \nOut1_5[4] , 
        \nOut0_15[3] , \nOut2_3[22] , \nOut2_4[8] , \nScanOut25[18] , 
        \nScanOut5[17] , \nOut1_11[12] , \nScanOut18[11] , \nScanOut1[15] , 
        \nScanOut5[24] , \nOut1_6[7] , \nOut1_11[21] , \nScanOut8[3] , 
        \nOut2_1[5] , \nOut2_2[6] , \nScanOut18[22] , \nOut1_15[10] , 
        \nOut1_4[18] , \nScanOut39[5] , \nOut0_0[24] , \nOut0_0[17] , 
        \nScanOut1[26] , \nOut1_10[3] , \nOut1_13[0] , \nScanOut27[9] , 
        \nOut1_15[23] , \nScanOut21[30] , \nScanOut21[29] , \nScanOut46[0] , 
        \nScanOut21[7] , \nScanOut22[4] , \nOut2_7[13] , \nScanOut45[3] , 
        \nOut2_7[20] , \nOut0_0[6] , \nOut0_3[5] , \nOut1_5[21] , 
        \nOut1_5[12] , \nOut0_6[8] , \nOut1_14[30] , \nOut1_14[29] , 
        \nScanOut34[0] , \nScanOut37[3] , \nScanOut5[6] , \nScanOut6[5] , 
        \nOut0_11[26] , \nScanOut16[15] , \nScanOut20[10] , \nScanOut35[24] , 
        \nScanOut40[14] , \nOut2_12[27] , \nOut1_1[23] , \nOut1_1[10] , 
        \nScanOut3[8] , \nOut0_11[15] , \nOut2_6[19] , \nScanOut48[6] , 
        \nScanOut12[24] , \nScanOut12[17] , \nScanOut16[26] , \nScanOut35[17] , 
        \nScanOut40[27] , \nScanOut20[23] , \nOut2_12[14] , \nOut2_14[4] , 
        \nScanOut31[26] , \nScanOut44[16] , \nOut0_15[24] , \nOut2_2[31] , 
        \nScanOut24[12] , \nOut2_2[28] , \nScanOut16[8] , \nScanOut24[21] , 
        \nScanOut31[15] , \nScanOut44[25] , \nOut0_15[17] , \nScanOut19[31] , 
        \nScanOut19[28] , \nScanOut10[6] , \nOut2_9[17] , \nOut2_11[9] , 
        \nOut0_2[8] , \nScanOut2[19] , \nOut0_8[24] , \nOut1_8[1] , 
        \nOut1_10[18] , \nOut2_9[24] , \nScanOut13[5] , \nOut2_8[0] , 
        \nOut0_3[31] , \nOut0_3[28] , \nOut1_7[27] , \nOut2_15[9] , 
        \nOut1_7[14] , \nOut0_8[17] , \nScanOut14[6] , \nScanOut17[5] , 
        \nScanOut29[30] , \nScanOut29[29] , \nScanOut9[26] , \nOut0_13[13] , 
        \nScanOut14[20] , \nScanOut22[25] , \nOut2_10[4] , \nOut2_13[7] , 
        \nScanOut37[11] , \nScanOut42[21] , \nOut2_10[12] , \nOut0_4[6] , 
        \nScanOut9[15] , \nScanOut10[22] , \nScanOut12[8] , \nOut0_13[20] , 
        \nScanOut14[13] , \nScanOut37[22] , \nScanOut42[12] , \nOut2_10[21] , 
        \nScanOut22[16] , \nOut2_14[10] , \nScanOut33[13] , \nScanOut46[23] , 
        \nScanOut26[27] , \nOut0_7[19] , \nOut0_7[5] , \nScanOut7[8] , 
        \nScanOut28[2] , \nOut1_8[30] , \nScanOut26[14] , \nScanOut46[10] , 
        \nOut1_8[29] , \nScanOut33[20] , \nScanOut10[11] , \nOut2_14[23] , 
        \nScanOut30[0] , \nOut1_3[25] , \nScanOut33[3] , \nOut1_1[4] , 
        \nScanOut1[6] , \nOut1_3[16] , \nOut1_2[7] , \nScanOut2[5] , 
        \nScanOut6[31] , \nOut0_6[20] , \nScanOut6[28] , \nOut0_6[13] , 
        \nOut1_9[23] , \nOut2_1[24] , \nScanOut41[3] , \nScanOut42[0] , 
        \nOut2_1[17] , \nScanOut25[7] , \nOut2_15[30] , \nOut2_15[29] , 
        \nScanOut38[8] , \nScanOut7[22] , \nOut0_9[3] , \nOut1_9[10] , 
        \nScanOut11[28] , \nScanOut47[30] , \nScanOut11[31] , \nOut1_13[27] , 
        \nScanOut26[4] , \nScanOut32[19] , \nScanOut47[29] , \nScanOut7[11] , 
        \nOut1_14[3] , \nScanOut23[9] , \nScanOut39[15] , \nOut1_13[14] , 
        \nScanOut28[23] , \nScanOut39[26] , \nScanOut3[20] , \nOut0_11[3] , 
        \nOut0_12[0] , \nScanOut19[3] , \nScanOut48[27] , \nOut0_2[22] , 
        \nScanOut3[13] , \nOut2_5[5] , \nOut2_6[6] , \nScanOut28[10] , 
        \nScanOut48[14] , \nOut1_4[9] , \nScanOut15[19] , \nScanOut36[31] , 
        \nOut2_5[26] , \nScanOut36[28] , \nScanOut43[18] , \nOut0_2[18] , 
        \nOut0_2[11] , \nOut2_0[8] , \nOut2_11[18] , \nOut1_2[26] , 
        \nScanOut7[18] , \nOut0_12[19] , \nOut2_5[15] , \nScanOut23[0] , 
        \nOut1_2[15] , \nScanOut20[3] , \nScanOut44[7] , \nScanOut47[4] , 
        \nOut0_6[30] , \nOut1_9[19] , \nScanOut11[21] , \nOut1_12[4] , 
        \nScanOut27[24] , \nScanOut38[1] , \nOut2_15[13] , \nOut1_11[7] , 
        \nScanOut32[10] , \nScanOut47[20] , \nOut0_6[29] , \nScanOut9[7] , 
        \nScanOut11[12] , \nOut2_15[20] , \nScanOut15[23] , \nScanOut27[17] , 
        \nScanOut32[23] , \nScanOut47[13] , \nScanOut42[9] , \nOut2_0[1] , 
        \nScanOut23[26] , \nOut2_11[11] , \nScanOut36[12] , \nScanOut43[22] , 
        \nScanOut8[25] , \nOut2_3[2] , \nOut0_12[10] , \nScanOut2[23] , 
        \nOut0_3[21] , \nScanOut3[30] , \nScanOut3[29] , \nOut1_4[0] , 
        \nOut1_6[24] , \nOut1_7[3] , \nScanOut8[16] , \nOut0_14[7] , 
        \nScanOut15[10] , \nScanOut23[15] , \nOut2_11[22] , \nScanOut36[21] , 
        \nScanOut43[11] , \nOut0_12[23] , \nScanOut28[19] , \nOut1_6[17] , 
        \nOut0_9[27] , \nOut0_9[14] , \nOut0_12[9] , \nOut0_3[12] , 
        \nOut1_9[5] , \nScanOut11[2] , \nOut0_13[30] , \nOut0_13[29] , 
        \nOut2_4[25] , \nScanOut12[1] , \nOut2_4[16] , \nOut2_10[31] , 
        \nOut2_10[28] , \nScanOut14[30] , \nScanOut14[29] , \nScanOut37[18] , 
        \nScanOut42[28] , \nScanOut42[31] , \nScanOut29[20] , \nOut0_1[2] , 
        \nOut0_2[1] , \nScanOut2[10] , \nOut2_8[9] , \nScanOut6[21] , 
        \nOut1_12[24] , \nScanOut29[13] , \nOut2_15[0] , \nScanOut38[16] , 
        \nScanOut30[9] , \nScanOut38[25] , \nScanOut6[12] , \nOut1_12[17] , 
        \nOut1_1[0] , \nOut0_2[26] , \nScanOut4[2] , \nOut0_7[23] , 
        \nScanOut7[1] , \nOut1_8[20] , \nScanOut33[29] , \nScanOut46[19] , 
        \nScanOut10[18] , \nScanOut33[30] , \nOut2_0[27] , \nOut0_7[10] , 
        \nOut1_8[13] , \nOut2_14[19] , \nScanOut36[7] , \nOut2_0[14] , 
        \nScanOut35[4] , \nOut0_2[15] , \nScanOut8[31] , \nOut2_5[22] , 
        \nOut2_5[11] , \nScanOut23[18] , \nScanOut8[28] , \nScanOut1[2] , 
        \nOut1_2[18] , \nOut1_2[3] , \nScanOut3[24] , \nOut0_9[19] , 
        \nOut0_11[7] , \nOut0_12[4] , \nScanOut19[7] , \nScanOut48[23] , 
        \nScanOut3[17] , \nScanOut28[27] , \nOut1_6[30] , \nOut2_5[1] , 
        \nScanOut28[14] , \nOut1_6[29] , \nOut2_6[2] , \nScanOut48[10] , 
        \nScanOut39[11] , \nScanOut2[1] , \nOut1_3[21] , \nOut0_6[24] , 
        \nScanOut7[26] , \nOut1_13[23] , \nScanOut47[9] , \nScanOut7[15] , 
        \nScanOut39[22] , \nOut1_9[27] , \nOut1_13[10] , \nOut1_14[7] , 
        \nOut2_1[20] , \nScanOut42[4] , \nScanOut41[7] , \nOut0_6[17] , 
        \nOut0_9[7] , \nOut1_9[14] , \nScanOut26[0] , \nScanOut27[30] , 
        \nScanOut27[29] , \nOut1_12[9] , \nScanOut25[3] , \nOut2_1[13] , 
        \nScanOut33[7] , \nOut1_12[30] , \nOut1_12[29] , \nScanOut30[4] , 
        \nScanOut38[31] , \nScanOut38[28] , \nOut1_3[12] , \nOut0_4[2] , 
        \nOut0_7[1] , \nOut2_0[19] , \nScanOut35[9] , \nScanOut28[6] , 
        \nOut1_7[23] , \nOut1_9[8] , \nScanOut9[22] , \nScanOut10[26] , 
        \nScanOut26[23] , \nScanOut10[15] , \nOut2_14[14] , \nScanOut33[17] , 
        \nScanOut46[27] , \nScanOut14[24] , \nOut2_10[16] , \nScanOut26[10] , 
        \nOut2_14[27] , \nScanOut33[24] , \nScanOut46[14] , \nScanOut22[21] , 
        \nScanOut37[15] , \nScanOut42[25] , \nOut2_10[0] , \nOut2_13[3] , 
        \nOut0_13[17] , \nScanOut22[12] , \nScanOut9[11] , \nScanOut14[17] , 
        \nOut2_10[25] , \nScanOut37[26] , \nScanOut42[16] , \nOut0_13[24] , 
        \nOut2_4[31] , \nOut2_4[28] , \nOut1_7[10] , \nOut0_8[20] , 
        \nOut2_8[4] , \nOut0_8[13] , \nScanOut14[2] , \nScanOut17[1] , 
        \nOut0_1[6] , \nScanOut2[8] , \nScanOut4[6] , \nScanOut6[25] , 
        \nOut0_7[27] , \nOut0_7[14] , \nScanOut7[5] , \nOut1_8[24] , 
        \nOut2_0[23] , \nScanOut26[19] , \nOut2_0[10] , \nScanOut35[0] , 
        \nOut0_7[8] , \nOut1_8[17] , \nOut1_12[20] , \nScanOut36[3] , 
        \nScanOut6[16] , \nScanOut38[12] , \nOut0_2[5] , \nOut1_12[13] , 
        \nOut1_3[31] , \nOut1_3[28] , \nOut1_7[19] , \nScanOut29[24] , 
        \nScanOut38[21] , \nScanOut2[27] , \nScanOut17[8] , \nScanOut2[14] , 
        \nScanOut29[17] , \nOut0_8[30] , \nOut2_15[4] , \nOut0_8[29] , 
        \nOut1_1[9] , \nOut0_3[25] , \nOut1_9[1] , \nScanOut12[5] , 
        \nScanOut9[18] , \nOut2_4[21] , \nScanOut11[6] , \nOut0_3[16] , 
        \nScanOut22[31] , \nScanOut22[28] , \nOut2_10[9] , \nOut1_6[20] , 
        \nOut0_9[23] , \nOut2_4[12] , \nOut2_5[8] , \nScanOut48[19] , 
        \nOut1_4[4] , \nOut1_6[13] , \nOut0_9[10] , \nOut1_7[7] , 
        \nScanOut8[21] , \nOut0_12[14] , \nScanOut15[27] , \nOut2_0[5] , 
        \nOut2_3[6] , \nOut2_5[18] , \nScanOut23[22] , \nOut2_11[15] , 
        \nScanOut36[16] , \nScanOut43[26] , \nScanOut8[12] , \nOut0_12[27] , 
        \nOut0_14[3] , \nScanOut15[14] , \nOut2_11[26] , \nScanOut36[25] , 
        \nScanOut43[15] , \nScanOut23[11] , \nOut1_2[22] , \nScanOut9[3] , 
        \nOut1_11[3] , \nScanOut26[9] , \nScanOut32[14] , \nScanOut47[24] , 
        \nScanOut11[25] , \nScanOut11[16] , \nOut1_12[0] , \nScanOut27[20] , 
        \nOut2_15[17] , \nScanOut38[5] , \nScanOut27[13] , \nScanOut32[27] , 
        \nScanOut47[17] , \nOut2_1[30] , \nOut2_15[24] , \nOut2_1[29] , 
        \nScanOut20[7] , \nOut1_2[11] , \nOut1_13[19] , \nScanOut23[4] , 
        \nScanOut39[18] , \nOut1_2[8] , \nOut1_6[22] , \nOut2_6[9] , 
        \nScanOut44[3] , \nScanOut47[0] , \nOut1_6[11] , \nOut0_9[21] , 
        \nScanOut48[31] , \nScanOut48[28] , \nOut1_4[6] , \nScanOut8[23] , 
        \nOut0_9[12] , \nScanOut15[25] , \nScanOut36[14] , \nScanOut43[24] , 
        \nOut2_0[7] , \nScanOut23[20] , \nOut2_11[17] , \nOut2_3[4] , 
        \nOut0_12[16] , \nOut0_1[4] , \nScanOut1[9] , \nOut1_2[20] , 
        \nOut1_7[5] , \nScanOut8[10] , \nOut0_14[1] , \nScanOut15[16] , 
        \nScanOut23[13] , \nScanOut36[27] , \nScanOut43[17] , \nOut2_11[24] , 
        \nOut0_12[25] , \nOut2_5[30] , \nOut2_5[29] , \nScanOut9[1] , 
        \nOut1_11[1] , \nOut1_12[2] , \nOut2_1[18] , \nScanOut25[8] , 
        \nScanOut27[22] , \nScanOut38[7] , \nScanOut47[26] , \nScanOut11[27] , 
        \nOut2_15[15] , \nScanOut32[16] , \nScanOut11[14] , \nOut2_15[26] , 
        \nScanOut32[25] , \nScanOut47[15] , \nScanOut23[6] , \nScanOut27[11] , 
        \nScanOut39[30] , \nScanOut39[29] , \nOut1_2[13] , \nOut1_13[31] , 
        \nScanOut20[5] , \nOut1_13[28] , \nScanOut44[1] , \nScanOut47[2] , 
        \nOut0_4[9] , \nScanOut4[4] , \nScanOut7[7] , \nOut1_8[26] , 
        \nOut2_0[21] , \nOut0_7[25] , \nOut1_8[15] , \nScanOut26[31] , 
        \nScanOut26[28] , \nScanOut36[1] , \nOut0_7[16] , \nOut2_0[12] , 
        \nScanOut35[2] , \nOut0_2[7] , \nOut1_3[19] , \nScanOut6[27] , 
        \nScanOut38[10] , \nOut1_12[22] , \nScanOut38[23] , \nOut1_12[11] , 
        \nScanOut2[25] , \nScanOut6[14] , \nOut0_8[18] , \nScanOut14[9] , 
        \nScanOut29[26] , \nScanOut1[0] , \nScanOut2[16] , \nOut2_15[6] , 
        \nOut0_3[27] , \nOut1_7[31] , \nOut1_7[28] , \nScanOut29[15] , 
        \nOut0_3[14] , \nOut1_9[3] , \nScanOut11[4] , \nScanOut12[7] , 
        \nOut2_4[23] , \nScanOut22[19] , \nScanOut9[30] , \nScanOut9[29] , 
        \nOut2_4[10] , \nOut2_13[8] , \nOut1_3[23] , \nScanOut30[6] , 
        \nOut1_3[10] , \nOut1_12[18] , \nScanOut33[5] , \nScanOut38[19] , 
        \nScanOut2[3] , \nOut0_4[0] , \nScanOut10[24] , \nOut2_14[16] , 
        \nScanOut26[21] , \nScanOut33[15] , \nScanOut46[25] , \nScanOut36[8] , 
        \nOut0_7[3] , \nScanOut28[4] , \nOut0_8[22] , \nScanOut9[20] , 
        \nScanOut10[17] , \nScanOut26[12] , \nOut2_14[25] , \nOut2_0[31] , 
        \nOut2_0[28] , \nScanOut33[26] , \nScanOut46[16] , \nScanOut9[13] , 
        \nOut0_13[15] , \nScanOut14[26] , \nOut2_4[19] , \nScanOut22[23] , 
        \nOut2_10[2] , \nOut2_13[1] , \nOut2_10[14] , \nScanOut37[17] , 
        \nScanOut42[27] , \nOut0_13[26] , \nScanOut14[15] , \nScanOut22[10] , 
        \nOut2_10[27] , \nScanOut37[24] , \nScanOut42[14] , \nOut2_8[6] , 
        \nOut1_7[21] , \nOut1_7[12] , \nOut0_8[11] , \nScanOut17[3] , 
        \nScanOut14[0] , \nEnable[0] , \nOut1_1[2] , \nOut0_2[24] , 
        \nScanOut8[19] , \nOut0_14[8] , \nOut2_5[20] , \nOut0_2[17] , 
        \nScanOut23[30] , \nScanOut23[29] , \nOut1_2[1] , \nOut1_6[18] , 
        \nScanOut19[5] , \nOut2_5[13] , \nScanOut28[25] , \nScanOut48[21] , 
        \nScanOut3[26] , \nOut0_11[5] , \nOut0_12[6] , \nScanOut3[15] , 
        \nOut2_5[3] , \nOut2_6[0] , \nScanOut48[12] , \nScanOut28[16] , 
        \nOut0_9[31] , \nOut0_9[28] , \nOut1_2[30] , \nScanOut7[24] , 
        \nScanOut7[17] , \nOut1_13[21] , \nOut1_13[12] , \nOut1_14[5] , 
        \nScanOut39[13] , \nScanOut44[8] , \nScanOut39[20] , \nOut1_2[29] , 
        \nOut0_3[23] , \nOut0_6[26] , \nOut0_6[15] , \nOut1_9[25] , 
        \nScanOut9[8] , \nScanOut41[5] , \nOut2_1[22] , \nScanOut27[18] , 
        \nScanOut42[6] , \nOut2_1[11] , \nScanOut25[1] , \nOut0_9[5] , 
        \nOut1_9[16] , \nOut1_11[8] , \nScanOut26[2] , \nOut1_9[7] , 
        \nScanOut14[18] , \nScanOut37[29] , \nScanOut42[19] , \nScanOut37[30] , 
        \nScanOut11[0] , \nScanOut12[3] , \nOut2_4[27] , \nOut0_3[10] , 
        \nOut2_10[19] , \nOut0_13[18] , \nOut2_4[14] , \nScanOut29[22] , 
        \nScanOut2[21] , \nScanOut2[12] , \nScanOut29[11] , \nOut2_15[2] , 
        \nOut0_1[0] , \nScanOut6[23] , \nOut1_12[26] , \nScanOut33[8] , 
        \nScanOut38[14] , \nOut0_2[30] , \nOut0_2[3] , \nScanOut6[10] , 
        \nOut1_12[15] , \nOut1_2[24] , \nScanOut4[0] , \nOut0_7[21] , 
        \nScanOut38[27] , \nOut0_7[12] , \nScanOut7[3] , \nOut1_8[22] , 
        \nOut2_0[25] , \nOut2_14[31] , \nOut2_14[28] , \nOut2_0[16] , 
        \nScanOut35[6] , \nOut1_8[11] , \nScanOut10[30] , \nScanOut28[9] , 
        \nScanOut33[18] , \nScanOut46[28] , \nScanOut36[5] , \nScanOut10[29] , 
        \nScanOut46[31] , \nScanOut20[1] , \nOut1_2[17] , \nOut1_14[8] , 
        \nScanOut23[2] , \nOut0_6[18] , \nScanOut7[30] , \nScanOut7[29] , 
        \nScanOut44[5] , \nScanOut47[6] , \nOut0_9[8] , \nOut1_11[5] , 
        \nScanOut11[23] , \nOut2_15[11] , \nScanOut47[22] , \nScanOut27[26] , 
        \nScanOut32[12] , \nScanOut38[3] , \nScanOut8[27] , \nOut1_9[31] , 
        \nOut1_9[28] , \nScanOut11[10] , \nOut1_12[6] , \nScanOut27[15] , 
        \nOut2_15[22] , \nScanOut32[21] , \nScanOut9[5] , \nScanOut41[8] , 
        \nScanOut47[11] , \nOut0_12[12] , \nScanOut15[21] , \nOut2_0[3] , 
        \nOut2_3[0] , \nScanOut23[24] , \nOut2_11[13] , \nScanOut36[10] , 
        \nScanOut43[20] , \nOut0_2[29] , \nOut1_7[1] , \nScanOut8[14] , 
        \nOut0_12[21] , \nOut0_14[5] , \nScanOut15[12] , \nOut2_11[20] , 
        \nScanOut36[23] , \nScanOut43[13] , \nScanOut23[17] , \nOut0_1[9] , 
        \nOut1_1[6] , \nScanOut3[18] , \nOut1_4[2] , \nOut0_9[25] , 
        \nOut0_6[22] , \nOut1_6[26] , \nOut1_6[15] , \nOut0_9[16] , 
        \nOut0_11[8] , \nScanOut28[31] , \nScanOut28[28] , \nOut1_9[21] , 
        \nScanOut11[19] , \nScanOut19[8] , \nScanOut32[31] , \nOut2_1[26] , 
        \nScanOut32[28] , \nScanOut42[2] , \nScanOut47[18] , \nScanOut41[1] , 
        \nOut0_6[11] , \nOut0_9[1] , \nOut1_9[12] , \nScanOut26[6] , 
        \nOut2_15[18] , \nScanOut7[20] , \nOut2_1[15] , \nScanOut25[5] , 
        \nScanOut39[17] , \nScanOut7[13] , \nOut1_13[25] , \nOut1_13[16] , 
        \nScanOut20[8] , \nScanOut39[24] , \nOut1_14[1] , \nOut0_2[20] , 
        \nOut1_2[5] , \nScanOut3[22] , \nOut0_11[1] , \nOut0_12[2] , 
        \nScanOut3[11] , \nScanOut19[1] , \nScanOut48[25] , \nScanOut28[21] , 
        \nOut1_7[8] , \nOut2_5[7] , \nOut2_6[4] , \nScanOut28[12] , 
        \nScanOut48[16] , \nOut0_2[13] , \nOut0_12[31] , \nOut0_12[28] , 
        \nOut2_5[24] , \nOut2_5[17] , \nOut2_11[30] , \nOut2_11[29] , 
        \nScanOut2[31] , \nOut1_7[25] , \nScanOut15[31] , \nScanOut15[28] , 
        \nOut2_3[9] , \nScanOut43[30] , \nScanOut36[19] , \nScanOut43[29] , 
        \nScanOut29[18] , \nOut1_7[16] , \nOut0_8[26] , \nOut2_8[2] , 
        \nOut0_8[15] , \nScanOut14[4] , \nScanOut17[7] , \nScanOut2[28] , 
        \nOut0_3[19] , \nScanOut14[22] , \nOut2_10[10] , \nScanOut37[13] , 
        \nScanOut42[23] , \nScanOut22[27] , \nOut2_10[6] , \nOut0_4[4] , 
        \nOut0_7[7] , \nScanOut9[24] , \nOut2_13[5] , \nScanOut9[17] , 
        \nScanOut11[9] , \nOut0_13[11] , \nScanOut14[11] , \nScanOut22[14] , 
        \nOut2_10[23] , \nScanOut37[20] , \nScanOut42[10] , \nOut0_13[22] , 
        \nScanOut28[0] , \nScanOut4[9] , \nOut0_7[28] , \nOut1_8[18] , 
        \nScanOut26[25] , \nScanOut33[11] , \nScanOut46[21] , \nScanOut10[20] , 
        \nOut2_14[12] , \nOut0_7[31] , \nScanOut10[13] , \nScanOut33[22] , 
        \nScanOut46[12] , \nScanOut26[16] , \nOut2_14[21] , \nScanOut33[1] , 
        \nScanOut1[4] , \nScanOut2[7] , \nOut1_3[27] , \nScanOut6[19] , 
        \nScanOut30[2] , \nOut1_3[14] ;
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_3 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut4[31] , \nScanOut4[30] , \nScanOut4[29] , 
        \nScanOut4[28] , \nScanOut4[27] , \nScanOut4[26] , \nScanOut4[25] , 
        \nScanOut4[24] , \nScanOut4[23] , \nScanOut4[22] , \nScanOut4[21] , 
        \nScanOut4[20] , \nScanOut4[19] , \nScanOut4[18] , \nScanOut4[17] , 
        \nScanOut4[16] , \nScanOut4[15] , \nScanOut4[14] , \nScanOut4[13] , 
        \nScanOut4[12] , \nScanOut4[11] , \nScanOut4[10] , \nScanOut4[9] , 
        \nScanOut4[8] , \nScanOut4[7] , \nScanOut4[6] , \nScanOut4[5] , 
        \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , \nScanOut4[1] , 
        \nScanOut4[0] }), .ScanOut({\nScanOut3[31] , \nScanOut3[30] , 
        \nScanOut3[29] , \nScanOut3[28] , \nScanOut3[27] , \nScanOut3[26] , 
        \nScanOut3[25] , \nScanOut3[24] , \nScanOut3[23] , \nScanOut3[22] , 
        \nScanOut3[21] , \nScanOut3[20] , \nScanOut3[19] , \nScanOut3[18] , 
        \nScanOut3[17] , \nScanOut3[16] , \nScanOut3[15] , \nScanOut3[14] , 
        \nScanOut3[13] , \nScanOut3[12] , \nScanOut3[11] , \nScanOut3[10] , 
        \nScanOut3[9] , \nScanOut3[8] , \nScanOut3[7] , \nScanOut3[6] , 
        \nScanOut3[5] , \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , 
        \nScanOut3[1] , \nScanOut3[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_3[31] , 
        \nOut0_3[30] , \nOut0_3[29] , \nOut0_3[28] , \nOut0_3[27] , 
        \nOut0_3[26] , \nOut0_3[25] , \nOut0_3[24] , \nOut0_3[23] , 
        \nOut0_3[22] , \nOut0_3[21] , \nOut0_3[20] , \nOut0_3[19] , 
        \nOut0_3[18] , \nOut0_3[17] , \nOut0_3[16] , \nOut0_3[15] , 
        \nOut0_3[14] , \nOut0_3[13] , \nOut0_3[12] , \nOut0_3[11] , 
        \nOut0_3[10] , \nOut0_3[9] , \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , 
        \nOut0_3[5] , \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , 
        \nOut0_3[0] }), .NORTH_EDGE({\nOut0_2[31] , \nOut0_2[30] , 
        \nOut0_2[29] , \nOut0_2[28] , \nOut0_2[27] , \nOut0_2[26] , 
        \nOut0_2[25] , \nOut0_2[24] , \nOut0_2[23] , \nOut0_2[22] , 
        \nOut0_2[21] , \nOut0_2[20] , \nOut0_2[19] , \nOut0_2[18] , 
        \nOut0_2[17] , \nOut0_2[16] , \nOut0_2[15] , \nOut0_2[14] , 
        \nOut0_2[13] , \nOut0_2[12] , \nOut0_2[11] , \nOut0_2[10] , 
        \nOut0_2[9] , \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , 
        \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), 
        .SOUTH_EDGE({\nOut0_4[31] , \nOut0_4[30] , \nOut0_4[29] , 
        \nOut0_4[28] , \nOut0_4[27] , \nOut0_4[26] , \nOut0_4[25] , 
        \nOut0_4[24] , \nOut0_4[23] , \nOut0_4[22] , \nOut0_4[21] , 
        \nOut0_4[20] , \nOut0_4[19] , \nOut0_4[18] , \nOut0_4[17] , 
        \nOut0_4[16] , \nOut0_4[15] , \nOut0_4[14] , \nOut0_4[13] , 
        \nOut0_4[12] , \nOut0_4[11] , \nOut0_4[10] , \nOut0_4[9] , 
        \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , \nOut0_4[4] , 
        \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), .EAST_EDGE(
        \nOut1_3[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_2[31] ), .SE_EDGE(\nOut1_4[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_21 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut22[31] , \nScanOut22[30] , \nScanOut22[29] , 
        \nScanOut22[28] , \nScanOut22[27] , \nScanOut22[26] , \nScanOut22[25] , 
        \nScanOut22[24] , \nScanOut22[23] , \nScanOut22[22] , \nScanOut22[21] , 
        \nScanOut22[20] , \nScanOut22[19] , \nScanOut22[18] , \nScanOut22[17] , 
        \nScanOut22[16] , \nScanOut22[15] , \nScanOut22[14] , \nScanOut22[13] , 
        \nScanOut22[12] , \nScanOut22[11] , \nScanOut22[10] , \nScanOut22[9] , 
        \nScanOut22[8] , \nScanOut22[7] , \nScanOut22[6] , \nScanOut22[5] , 
        \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , \nScanOut22[1] , 
        \nScanOut22[0] }), .ScanOut({\nScanOut21[31] , \nScanOut21[30] , 
        \nScanOut21[29] , \nScanOut21[28] , \nScanOut21[27] , \nScanOut21[26] , 
        \nScanOut21[25] , \nScanOut21[24] , \nScanOut21[23] , \nScanOut21[22] , 
        \nScanOut21[21] , \nScanOut21[20] , \nScanOut21[19] , \nScanOut21[18] , 
        \nScanOut21[17] , \nScanOut21[16] , \nScanOut21[15] , \nScanOut21[14] , 
        \nScanOut21[13] , \nScanOut21[12] , \nScanOut21[11] , \nScanOut21[10] , 
        \nScanOut21[9] , \nScanOut21[8] , \nScanOut21[7] , \nScanOut21[6] , 
        \nScanOut21[5] , \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , 
        \nScanOut21[1] , \nScanOut21[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_5[31] , 
        \nOut1_5[30] , \nOut1_5[29] , \nOut1_5[28] , \nOut1_5[27] , 
        \nOut1_5[26] , \nOut1_5[25] , \nOut1_5[24] , \nOut1_5[23] , 
        \nOut1_5[22] , \nOut1_5[21] , \nOut1_5[20] , \nOut1_5[19] , 
        \nOut1_5[18] , \nOut1_5[17] , \nOut1_5[16] , \nOut1_5[15] , 
        \nOut1_5[14] , \nOut1_5[13] , \nOut1_5[12] , \nOut1_5[11] , 
        \nOut1_5[10] , \nOut1_5[9] , \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , 
        \nOut1_5[5] , \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , 
        \nOut1_5[0] }), .NORTH_EDGE({\nOut1_4[31] , \nOut1_4[30] , 
        \nOut1_4[29] , \nOut1_4[28] , \nOut1_4[27] , \nOut1_4[26] , 
        \nOut1_4[25] , \nOut1_4[24] , \nOut1_4[23] , \nOut1_4[22] , 
        \nOut1_4[21] , \nOut1_4[20] , \nOut1_4[19] , \nOut1_4[18] , 
        \nOut1_4[17] , \nOut1_4[16] , \nOut1_4[15] , \nOut1_4[14] , 
        \nOut1_4[13] , \nOut1_4[12] , \nOut1_4[11] , \nOut1_4[10] , 
        \nOut1_4[9] , \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , 
        \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), 
        .SOUTH_EDGE({\nOut1_6[31] , \nOut1_6[30] , \nOut1_6[29] , 
        \nOut1_6[28] , \nOut1_6[27] , \nOut1_6[26] , \nOut1_6[25] , 
        \nOut1_6[24] , \nOut1_6[23] , \nOut1_6[22] , \nOut1_6[21] , 
        \nOut1_6[20] , \nOut1_6[19] , \nOut1_6[18] , \nOut1_6[17] , 
        \nOut1_6[16] , \nOut1_6[15] , \nOut1_6[14] , \nOut1_6[13] , 
        \nOut1_6[12] , \nOut1_6[11] , \nOut1_6[10] , \nOut1_6[9] , 
        \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , \nOut1_6[4] , 
        \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), .EAST_EDGE(
        \nOut2_5[31] ), .WEST_EDGE(\nOut0_5[0] ), .NW_EDGE(\nOut0_4[0] ), 
        .SW_EDGE(\nOut0_6[0] ), .NE_EDGE(\nOut2_4[31] ), .SE_EDGE(
        \nOut2_6[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_0 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut1[31] , \nScanOut1[30] , \nScanOut1[29] , 
        \nScanOut1[28] , \nScanOut1[27] , \nScanOut1[26] , \nScanOut1[25] , 
        \nScanOut1[24] , \nScanOut1[23] , \nScanOut1[22] , \nScanOut1[21] , 
        \nScanOut1[20] , \nScanOut1[19] , \nScanOut1[18] , \nScanOut1[17] , 
        \nScanOut1[16] , \nScanOut1[15] , \nScanOut1[14] , \nScanOut1[13] , 
        \nScanOut1[12] , \nScanOut1[11] , \nScanOut1[10] , \nScanOut1[9] , 
        \nScanOut1[8] , \nScanOut1[7] , \nScanOut1[6] , \nScanOut1[5] , 
        \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , \nScanOut1[1] , 
        \nScanOut1[0] }), .ScanOut({\nScanOut0[31] , \nScanOut0[30] , 
        \nScanOut0[29] , \nScanOut0[28] , \nScanOut0[27] , \nScanOut0[26] , 
        \nScanOut0[25] , \nScanOut0[24] , \nScanOut0[23] , \nScanOut0[22] , 
        \nScanOut0[21] , \nScanOut0[20] , \nScanOut0[19] , \nScanOut0[18] , 
        \nScanOut0[17] , \nScanOut0[16] , \nScanOut0[15] , \nScanOut0[14] , 
        \nScanOut0[13] , \nScanOut0[12] , \nScanOut0[11] , \nScanOut0[10] , 
        \nScanOut0[9] , \nScanOut0[8] , \nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_0[31] , 
        \nOut0_0[30] , \nOut0_0[29] , \nOut0_0[28] , \nOut0_0[27] , 
        \nOut0_0[26] , \nOut0_0[25] , \nOut0_0[24] , \nOut0_0[23] , 
        \nOut0_0[22] , \nOut0_0[21] , \nOut0_0[20] , \nOut0_0[19] , 
        \nOut0_0[18] , \nOut0_0[17] , \nOut0_0[16] , \nOut0_0[15] , 
        \nOut0_0[14] , \nOut0_0[13] , \nOut0_0[12] , \nOut0_0[11] , 
        \nOut0_0[10] , \nOut0_0[9] , \nOut0_0[8] , \nOut0_0[7] , \nOut0_0[6] , 
        \nOut0_0[5] , \nOut0_0[4] , \nOut0_0[3] , \nOut0_0[2] , \nOut0_0[1] , 
        \nOut0_0[0] }), .NORTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SOUTH_EDGE({\nOut0_1[31] , \nOut0_1[30] , \nOut0_1[29] , 
        \nOut0_1[28] , \nOut0_1[27] , \nOut0_1[26] , \nOut0_1[25] , 
        \nOut0_1[24] , \nOut0_1[23] , \nOut0_1[22] , \nOut0_1[21] , 
        \nOut0_1[20] , \nOut0_1[19] , \nOut0_1[18] , \nOut0_1[17] , 
        \nOut0_1[16] , \nOut0_1[15] , \nOut0_1[14] , \nOut0_1[13] , 
        \nOut0_1[12] , \nOut0_1[11] , \nOut0_1[10] , \nOut0_1[9] , 
        \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , \nOut0_1[4] , 
        \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), .EAST_EDGE(
        \nOut1_0[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(1'b0), .SE_EDGE(\nOut1_1[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_2 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut3[31] , \nScanOut3[30] , \nScanOut3[29] , 
        \nScanOut3[28] , \nScanOut3[27] , \nScanOut3[26] , \nScanOut3[25] , 
        \nScanOut3[24] , \nScanOut3[23] , \nScanOut3[22] , \nScanOut3[21] , 
        \nScanOut3[20] , \nScanOut3[19] , \nScanOut3[18] , \nScanOut3[17] , 
        \nScanOut3[16] , \nScanOut3[15] , \nScanOut3[14] , \nScanOut3[13] , 
        \nScanOut3[12] , \nScanOut3[11] , \nScanOut3[10] , \nScanOut3[9] , 
        \nScanOut3[8] , \nScanOut3[7] , \nScanOut3[6] , \nScanOut3[5] , 
        \nScanOut3[4] , \nScanOut3[3] , \nScanOut3[2] , \nScanOut3[1] , 
        \nScanOut3[0] }), .ScanOut({\nScanOut2[31] , \nScanOut2[30] , 
        \nScanOut2[29] , \nScanOut2[28] , \nScanOut2[27] , \nScanOut2[26] , 
        \nScanOut2[25] , \nScanOut2[24] , \nScanOut2[23] , \nScanOut2[22] , 
        \nScanOut2[21] , \nScanOut2[20] , \nScanOut2[19] , \nScanOut2[18] , 
        \nScanOut2[17] , \nScanOut2[16] , \nScanOut2[15] , \nScanOut2[14] , 
        \nScanOut2[13] , \nScanOut2[12] , \nScanOut2[11] , \nScanOut2[10] , 
        \nScanOut2[9] , \nScanOut2[8] , \nScanOut2[7] , \nScanOut2[6] , 
        \nScanOut2[5] , \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , 
        \nScanOut2[1] , \nScanOut2[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_2[31] , 
        \nOut0_2[30] , \nOut0_2[29] , \nOut0_2[28] , \nOut0_2[27] , 
        \nOut0_2[26] , \nOut0_2[25] , \nOut0_2[24] , \nOut0_2[23] , 
        \nOut0_2[22] , \nOut0_2[21] , \nOut0_2[20] , \nOut0_2[19] , 
        \nOut0_2[18] , \nOut0_2[17] , \nOut0_2[16] , \nOut0_2[15] , 
        \nOut0_2[14] , \nOut0_2[13] , \nOut0_2[12] , \nOut0_2[11] , 
        \nOut0_2[10] , \nOut0_2[9] , \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , 
        \nOut0_2[5] , \nOut0_2[4] , \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , 
        \nOut0_2[0] }), .NORTH_EDGE({\nOut0_1[31] , \nOut0_1[30] , 
        \nOut0_1[29] , \nOut0_1[28] , \nOut0_1[27] , \nOut0_1[26] , 
        \nOut0_1[25] , \nOut0_1[24] , \nOut0_1[23] , \nOut0_1[22] , 
        \nOut0_1[21] , \nOut0_1[20] , \nOut0_1[19] , \nOut0_1[18] , 
        \nOut0_1[17] , \nOut0_1[16] , \nOut0_1[15] , \nOut0_1[14] , 
        \nOut0_1[13] , \nOut0_1[12] , \nOut0_1[11] , \nOut0_1[10] , 
        \nOut0_1[9] , \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , \nOut0_1[5] , 
        \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , \nOut0_1[0] }), 
        .SOUTH_EDGE({\nOut0_3[31] , \nOut0_3[30] , \nOut0_3[29] , 
        \nOut0_3[28] , \nOut0_3[27] , \nOut0_3[26] , \nOut0_3[25] , 
        \nOut0_3[24] , \nOut0_3[23] , \nOut0_3[22] , \nOut0_3[21] , 
        \nOut0_3[20] , \nOut0_3[19] , \nOut0_3[18] , \nOut0_3[17] , 
        \nOut0_3[16] , \nOut0_3[15] , \nOut0_3[14] , \nOut0_3[13] , 
        \nOut0_3[12] , \nOut0_3[11] , \nOut0_3[10] , \nOut0_3[9] , 
        \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , \nOut0_3[4] , 
        \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), .EAST_EDGE(
        \nOut1_2[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_1[31] ), .SE_EDGE(\nOut1_3[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_4 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut5[31] , \nScanOut5[30] , \nScanOut5[29] , 
        \nScanOut5[28] , \nScanOut5[27] , \nScanOut5[26] , \nScanOut5[25] , 
        \nScanOut5[24] , \nScanOut5[23] , \nScanOut5[22] , \nScanOut5[21] , 
        \nScanOut5[20] , \nScanOut5[19] , \nScanOut5[18] , \nScanOut5[17] , 
        \nScanOut5[16] , \nScanOut5[15] , \nScanOut5[14] , \nScanOut5[13] , 
        \nScanOut5[12] , \nScanOut5[11] , \nScanOut5[10] , \nScanOut5[9] , 
        \nScanOut5[8] , \nScanOut5[7] , \nScanOut5[6] , \nScanOut5[5] , 
        \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , \nScanOut5[1] , 
        \nScanOut5[0] }), .ScanOut({\nScanOut4[31] , \nScanOut4[30] , 
        \nScanOut4[29] , \nScanOut4[28] , \nScanOut4[27] , \nScanOut4[26] , 
        \nScanOut4[25] , \nScanOut4[24] , \nScanOut4[23] , \nScanOut4[22] , 
        \nScanOut4[21] , \nScanOut4[20] , \nScanOut4[19] , \nScanOut4[18] , 
        \nScanOut4[17] , \nScanOut4[16] , \nScanOut4[15] , \nScanOut4[14] , 
        \nScanOut4[13] , \nScanOut4[12] , \nScanOut4[11] , \nScanOut4[10] , 
        \nScanOut4[9] , \nScanOut4[8] , \nScanOut4[7] , \nScanOut4[6] , 
        \nScanOut4[5] , \nScanOut4[4] , \nScanOut4[3] , \nScanOut4[2] , 
        \nScanOut4[1] , \nScanOut4[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_4[31] , 
        \nOut0_4[30] , \nOut0_4[29] , \nOut0_4[28] , \nOut0_4[27] , 
        \nOut0_4[26] , \nOut0_4[25] , \nOut0_4[24] , \nOut0_4[23] , 
        \nOut0_4[22] , \nOut0_4[21] , \nOut0_4[20] , \nOut0_4[19] , 
        \nOut0_4[18] , \nOut0_4[17] , \nOut0_4[16] , \nOut0_4[15] , 
        \nOut0_4[14] , \nOut0_4[13] , \nOut0_4[12] , \nOut0_4[11] , 
        \nOut0_4[10] , \nOut0_4[9] , \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , 
        \nOut0_4[5] , \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , 
        \nOut0_4[0] }), .NORTH_EDGE({\nOut0_3[31] , \nOut0_3[30] , 
        \nOut0_3[29] , \nOut0_3[28] , \nOut0_3[27] , \nOut0_3[26] , 
        \nOut0_3[25] , \nOut0_3[24] , \nOut0_3[23] , \nOut0_3[22] , 
        \nOut0_3[21] , \nOut0_3[20] , \nOut0_3[19] , \nOut0_3[18] , 
        \nOut0_3[17] , \nOut0_3[16] , \nOut0_3[15] , \nOut0_3[14] , 
        \nOut0_3[13] , \nOut0_3[12] , \nOut0_3[11] , \nOut0_3[10] , 
        \nOut0_3[9] , \nOut0_3[8] , \nOut0_3[7] , \nOut0_3[6] , \nOut0_3[5] , 
        \nOut0_3[4] , \nOut0_3[3] , \nOut0_3[2] , \nOut0_3[1] , \nOut0_3[0] }), 
        .SOUTH_EDGE({\nOut0_5[31] , \nOut0_5[30] , \nOut0_5[29] , 
        \nOut0_5[28] , \nOut0_5[27] , \nOut0_5[26] , \nOut0_5[25] , 
        \nOut0_5[24] , \nOut0_5[23] , \nOut0_5[22] , \nOut0_5[21] , 
        \nOut0_5[20] , \nOut0_5[19] , \nOut0_5[18] , \nOut0_5[17] , 
        \nOut0_5[16] , \nOut0_5[15] , \nOut0_5[14] , \nOut0_5[13] , 
        \nOut0_5[12] , \nOut0_5[11] , \nOut0_5[10] , \nOut0_5[9] , 
        \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , \nOut0_5[4] , 
        \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), .EAST_EDGE(
        \nOut1_4[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_3[31] ), .SE_EDGE(\nOut1_5[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_13 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut14[31] , \nScanOut14[30] , \nScanOut14[29] , 
        \nScanOut14[28] , \nScanOut14[27] , \nScanOut14[26] , \nScanOut14[25] , 
        \nScanOut14[24] , \nScanOut14[23] , \nScanOut14[22] , \nScanOut14[21] , 
        \nScanOut14[20] , \nScanOut14[19] , \nScanOut14[18] , \nScanOut14[17] , 
        \nScanOut14[16] , \nScanOut14[15] , \nScanOut14[14] , \nScanOut14[13] , 
        \nScanOut14[12] , \nScanOut14[11] , \nScanOut14[10] , \nScanOut14[9] , 
        \nScanOut14[8] , \nScanOut14[7] , \nScanOut14[6] , \nScanOut14[5] , 
        \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , \nScanOut14[1] , 
        \nScanOut14[0] }), .ScanOut({\nScanOut13[31] , \nScanOut13[30] , 
        \nScanOut13[29] , \nScanOut13[28] , \nScanOut13[27] , \nScanOut13[26] , 
        \nScanOut13[25] , \nScanOut13[24] , \nScanOut13[23] , \nScanOut13[22] , 
        \nScanOut13[21] , \nScanOut13[20] , \nScanOut13[19] , \nScanOut13[18] , 
        \nScanOut13[17] , \nScanOut13[16] , \nScanOut13[15] , \nScanOut13[14] , 
        \nScanOut13[13] , \nScanOut13[12] , \nScanOut13[11] , \nScanOut13[10] , 
        \nScanOut13[9] , \nScanOut13[8] , \nScanOut13[7] , \nScanOut13[6] , 
        \nScanOut13[5] , \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , 
        \nScanOut13[1] , \nScanOut13[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_13[31] , 
        \nOut0_13[30] , \nOut0_13[29] , \nOut0_13[28] , \nOut0_13[27] , 
        \nOut0_13[26] , \nOut0_13[25] , \nOut0_13[24] , \nOut0_13[23] , 
        \nOut0_13[22] , \nOut0_13[21] , \nOut0_13[20] , \nOut0_13[19] , 
        \nOut0_13[18] , \nOut0_13[17] , \nOut0_13[16] , \nOut0_13[15] , 
        \nOut0_13[14] , \nOut0_13[13] , \nOut0_13[12] , \nOut0_13[11] , 
        \nOut0_13[10] , \nOut0_13[9] , \nOut0_13[8] , \nOut0_13[7] , 
        \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , \nOut0_13[3] , 
        \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), .NORTH_EDGE({
        \nOut0_12[31] , \nOut0_12[30] , \nOut0_12[29] , \nOut0_12[28] , 
        \nOut0_12[27] , \nOut0_12[26] , \nOut0_12[25] , \nOut0_12[24] , 
        \nOut0_12[23] , \nOut0_12[22] , \nOut0_12[21] , \nOut0_12[20] , 
        \nOut0_12[19] , \nOut0_12[18] , \nOut0_12[17] , \nOut0_12[16] , 
        \nOut0_12[15] , \nOut0_12[14] , \nOut0_12[13] , \nOut0_12[12] , 
        \nOut0_12[11] , \nOut0_12[10] , \nOut0_12[9] , \nOut0_12[8] , 
        \nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , 
        \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), 
        .SOUTH_EDGE({\nOut0_14[31] , \nOut0_14[30] , \nOut0_14[29] , 
        \nOut0_14[28] , \nOut0_14[27] , \nOut0_14[26] , \nOut0_14[25] , 
        \nOut0_14[24] , \nOut0_14[23] , \nOut0_14[22] , \nOut0_14[21] , 
        \nOut0_14[20] , \nOut0_14[19] , \nOut0_14[18] , \nOut0_14[17] , 
        \nOut0_14[16] , \nOut0_14[15] , \nOut0_14[14] , \nOut0_14[13] , 
        \nOut0_14[12] , \nOut0_14[11] , \nOut0_14[10] , \nOut0_14[9] , 
        \nOut0_14[8] , \nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , 
        \nOut0_14[4] , \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , 
        \nOut0_14[0] }), .EAST_EDGE(\nOut1_13[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_12[31] ), .SE_EDGE(
        \nOut1_14[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_14 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut15[31] , \nScanOut15[30] , \nScanOut15[29] , 
        \nScanOut15[28] , \nScanOut15[27] , \nScanOut15[26] , \nScanOut15[25] , 
        \nScanOut15[24] , \nScanOut15[23] , \nScanOut15[22] , \nScanOut15[21] , 
        \nScanOut15[20] , \nScanOut15[19] , \nScanOut15[18] , \nScanOut15[17] , 
        \nScanOut15[16] , \nScanOut15[15] , \nScanOut15[14] , \nScanOut15[13] , 
        \nScanOut15[12] , \nScanOut15[11] , \nScanOut15[10] , \nScanOut15[9] , 
        \nScanOut15[8] , \nScanOut15[7] , \nScanOut15[6] , \nScanOut15[5] , 
        \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , \nScanOut15[1] , 
        \nScanOut15[0] }), .ScanOut({\nScanOut14[31] , \nScanOut14[30] , 
        \nScanOut14[29] , \nScanOut14[28] , \nScanOut14[27] , \nScanOut14[26] , 
        \nScanOut14[25] , \nScanOut14[24] , \nScanOut14[23] , \nScanOut14[22] , 
        \nScanOut14[21] , \nScanOut14[20] , \nScanOut14[19] , \nScanOut14[18] , 
        \nScanOut14[17] , \nScanOut14[16] , \nScanOut14[15] , \nScanOut14[14] , 
        \nScanOut14[13] , \nScanOut14[12] , \nScanOut14[11] , \nScanOut14[10] , 
        \nScanOut14[9] , \nScanOut14[8] , \nScanOut14[7] , \nScanOut14[6] , 
        \nScanOut14[5] , \nScanOut14[4] , \nScanOut14[3] , \nScanOut14[2] , 
        \nScanOut14[1] , \nScanOut14[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_14[31] , 
        \nOut0_14[30] , \nOut0_14[29] , \nOut0_14[28] , \nOut0_14[27] , 
        \nOut0_14[26] , \nOut0_14[25] , \nOut0_14[24] , \nOut0_14[23] , 
        \nOut0_14[22] , \nOut0_14[21] , \nOut0_14[20] , \nOut0_14[19] , 
        \nOut0_14[18] , \nOut0_14[17] , \nOut0_14[16] , \nOut0_14[15] , 
        \nOut0_14[14] , \nOut0_14[13] , \nOut0_14[12] , \nOut0_14[11] , 
        \nOut0_14[10] , \nOut0_14[9] , \nOut0_14[8] , \nOut0_14[7] , 
        \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , \nOut0_14[3] , 
        \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), .NORTH_EDGE({
        \nOut0_13[31] , \nOut0_13[30] , \nOut0_13[29] , \nOut0_13[28] , 
        \nOut0_13[27] , \nOut0_13[26] , \nOut0_13[25] , \nOut0_13[24] , 
        \nOut0_13[23] , \nOut0_13[22] , \nOut0_13[21] , \nOut0_13[20] , 
        \nOut0_13[19] , \nOut0_13[18] , \nOut0_13[17] , \nOut0_13[16] , 
        \nOut0_13[15] , \nOut0_13[14] , \nOut0_13[13] , \nOut0_13[12] , 
        \nOut0_13[11] , \nOut0_13[10] , \nOut0_13[9] , \nOut0_13[8] , 
        \nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , \nOut0_13[4] , 
        \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , \nOut0_13[0] }), 
        .SOUTH_EDGE({\nOut0_15[31] , \nOut0_15[30] , \nOut0_15[29] , 
        \nOut0_15[28] , \nOut0_15[27] , \nOut0_15[26] , \nOut0_15[25] , 
        \nOut0_15[24] , \nOut0_15[23] , \nOut0_15[22] , \nOut0_15[21] , 
        \nOut0_15[20] , \nOut0_15[19] , \nOut0_15[18] , \nOut0_15[17] , 
        \nOut0_15[16] , \nOut0_15[15] , \nOut0_15[14] , \nOut0_15[13] , 
        \nOut0_15[12] , \nOut0_15[11] , \nOut0_15[10] , \nOut0_15[9] , 
        \nOut0_15[8] , \nOut0_15[7] , \nOut0_15[6] , \nOut0_15[5] , 
        \nOut0_15[4] , \nOut0_15[3] , \nOut0_15[2] , \nOut0_15[1] , 
        \nOut0_15[0] }), .EAST_EDGE(\nOut1_14[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_13[31] ), .SE_EDGE(
        \nOut1_15[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_33 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut34[31] , \nScanOut34[30] , \nScanOut34[29] , 
        \nScanOut34[28] , \nScanOut34[27] , \nScanOut34[26] , \nScanOut34[25] , 
        \nScanOut34[24] , \nScanOut34[23] , \nScanOut34[22] , \nScanOut34[21] , 
        \nScanOut34[20] , \nScanOut34[19] , \nScanOut34[18] , \nScanOut34[17] , 
        \nScanOut34[16] , \nScanOut34[15] , \nScanOut34[14] , \nScanOut34[13] , 
        \nScanOut34[12] , \nScanOut34[11] , \nScanOut34[10] , \nScanOut34[9] , 
        \nScanOut34[8] , \nScanOut34[7] , \nScanOut34[6] , \nScanOut34[5] , 
        \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , \nScanOut34[1] , 
        \nScanOut34[0] }), .ScanOut({\nScanOut33[31] , \nScanOut33[30] , 
        \nScanOut33[29] , \nScanOut33[28] , \nScanOut33[27] , \nScanOut33[26] , 
        \nScanOut33[25] , \nScanOut33[24] , \nScanOut33[23] , \nScanOut33[22] , 
        \nScanOut33[21] , \nScanOut33[20] , \nScanOut33[19] , \nScanOut33[18] , 
        \nScanOut33[17] , \nScanOut33[16] , \nScanOut33[15] , \nScanOut33[14] , 
        \nScanOut33[13] , \nScanOut33[12] , \nScanOut33[11] , \nScanOut33[10] , 
        \nScanOut33[9] , \nScanOut33[8] , \nScanOut33[7] , \nScanOut33[6] , 
        \nScanOut33[5] , \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , 
        \nScanOut33[1] , \nScanOut33[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_1[31] , 
        \nOut2_1[30] , \nOut2_1[29] , \nOut2_1[28] , \nOut2_1[27] , 
        \nOut2_1[26] , \nOut2_1[25] , \nOut2_1[24] , \nOut2_1[23] , 
        \nOut2_1[22] , \nOut2_1[21] , \nOut2_1[20] , \nOut2_1[19] , 
        \nOut2_1[18] , \nOut2_1[17] , \nOut2_1[16] , \nOut2_1[15] , 
        \nOut2_1[14] , \nOut2_1[13] , \nOut2_1[12] , \nOut2_1[11] , 
        \nOut2_1[10] , \nOut2_1[9] , \nOut2_1[8] , \nOut2_1[7] , \nOut2_1[6] , 
        \nOut2_1[5] , \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , 
        \nOut2_1[0] }), .NORTH_EDGE({\nOut2_0[31] , \nOut2_0[30] , 
        \nOut2_0[29] , \nOut2_0[28] , \nOut2_0[27] , \nOut2_0[26] , 
        \nOut2_0[25] , \nOut2_0[24] , \nOut2_0[23] , \nOut2_0[22] , 
        \nOut2_0[21] , \nOut2_0[20] , \nOut2_0[19] , \nOut2_0[18] , 
        \nOut2_0[17] , \nOut2_0[16] , \nOut2_0[15] , \nOut2_0[14] , 
        \nOut2_0[13] , \nOut2_0[12] , \nOut2_0[11] , \nOut2_0[10] , 
        \nOut2_0[9] , \nOut2_0[8] , \nOut2_0[7] , \nOut2_0[6] , \nOut2_0[5] , 
        \nOut2_0[4] , \nOut2_0[3] , \nOut2_0[2] , \nOut2_0[1] , \nOut2_0[0] }), 
        .SOUTH_EDGE({\nOut2_2[31] , \nOut2_2[30] , \nOut2_2[29] , 
        \nOut2_2[28] , \nOut2_2[27] , \nOut2_2[26] , \nOut2_2[25] , 
        \nOut2_2[24] , \nOut2_2[23] , \nOut2_2[22] , \nOut2_2[21] , 
        \nOut2_2[20] , \nOut2_2[19] , \nOut2_2[18] , \nOut2_2[17] , 
        \nOut2_2[16] , \nOut2_2[15] , \nOut2_2[14] , \nOut2_2[13] , 
        \nOut2_2[12] , \nOut2_2[11] , \nOut2_2[10] , \nOut2_2[9] , 
        \nOut2_2[8] , \nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , \nOut2_2[4] , 
        \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_1[0] ), .NW_EDGE(\nOut1_0[0] ), .SW_EDGE(
        \nOut1_2[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_28 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut29[31] , \nScanOut29[30] , \nScanOut29[29] , 
        \nScanOut29[28] , \nScanOut29[27] , \nScanOut29[26] , \nScanOut29[25] , 
        \nScanOut29[24] , \nScanOut29[23] , \nScanOut29[22] , \nScanOut29[21] , 
        \nScanOut29[20] , \nScanOut29[19] , \nScanOut29[18] , \nScanOut29[17] , 
        \nScanOut29[16] , \nScanOut29[15] , \nScanOut29[14] , \nScanOut29[13] , 
        \nScanOut29[12] , \nScanOut29[11] , \nScanOut29[10] , \nScanOut29[9] , 
        \nScanOut29[8] , \nScanOut29[7] , \nScanOut29[6] , \nScanOut29[5] , 
        \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , \nScanOut29[1] , 
        \nScanOut29[0] }), .ScanOut({\nScanOut28[31] , \nScanOut28[30] , 
        \nScanOut28[29] , \nScanOut28[28] , \nScanOut28[27] , \nScanOut28[26] , 
        \nScanOut28[25] , \nScanOut28[24] , \nScanOut28[23] , \nScanOut28[22] , 
        \nScanOut28[21] , \nScanOut28[20] , \nScanOut28[19] , \nScanOut28[18] , 
        \nScanOut28[17] , \nScanOut28[16] , \nScanOut28[15] , \nScanOut28[14] , 
        \nScanOut28[13] , \nScanOut28[12] , \nScanOut28[11] , \nScanOut28[10] , 
        \nScanOut28[9] , \nScanOut28[8] , \nScanOut28[7] , \nScanOut28[6] , 
        \nScanOut28[5] , \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , 
        \nScanOut28[1] , \nScanOut28[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_12[31] , 
        \nOut1_12[30] , \nOut1_12[29] , \nOut1_12[28] , \nOut1_12[27] , 
        \nOut1_12[26] , \nOut1_12[25] , \nOut1_12[24] , \nOut1_12[23] , 
        \nOut1_12[22] , \nOut1_12[21] , \nOut1_12[20] , \nOut1_12[19] , 
        \nOut1_12[18] , \nOut1_12[17] , \nOut1_12[16] , \nOut1_12[15] , 
        \nOut1_12[14] , \nOut1_12[13] , \nOut1_12[12] , \nOut1_12[11] , 
        \nOut1_12[10] , \nOut1_12[9] , \nOut1_12[8] , \nOut1_12[7] , 
        \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , \nOut1_12[3] , 
        \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), .NORTH_EDGE({
        \nOut1_11[31] , \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , 
        \nOut1_11[27] , \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , 
        \nOut1_11[23] , \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , 
        \nOut1_11[19] , \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , 
        \nOut1_11[15] , \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , 
        \nOut1_11[11] , \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , 
        \nOut1_11[7] , \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , 
        \nOut1_11[3] , \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), 
        .SOUTH_EDGE({\nOut1_13[31] , \nOut1_13[30] , \nOut1_13[29] , 
        \nOut1_13[28] , \nOut1_13[27] , \nOut1_13[26] , \nOut1_13[25] , 
        \nOut1_13[24] , \nOut1_13[23] , \nOut1_13[22] , \nOut1_13[21] , 
        \nOut1_13[20] , \nOut1_13[19] , \nOut1_13[18] , \nOut1_13[17] , 
        \nOut1_13[16] , \nOut1_13[15] , \nOut1_13[14] , \nOut1_13[13] , 
        \nOut1_13[12] , \nOut1_13[11] , \nOut1_13[10] , \nOut1_13[9] , 
        \nOut1_13[8] , \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , 
        \nOut1_13[4] , \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , 
        \nOut1_13[0] }), .EAST_EDGE(\nOut2_12[31] ), .WEST_EDGE(\nOut0_12[0] ), 
        .NW_EDGE(\nOut0_11[0] ), .SW_EDGE(\nOut0_13[0] ), .NE_EDGE(
        \nOut2_11[31] ), .SE_EDGE(\nOut2_13[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_46 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut47[31] , \nScanOut47[30] , \nScanOut47[29] , 
        \nScanOut47[28] , \nScanOut47[27] , \nScanOut47[26] , \nScanOut47[25] , 
        \nScanOut47[24] , \nScanOut47[23] , \nScanOut47[22] , \nScanOut47[21] , 
        \nScanOut47[20] , \nScanOut47[19] , \nScanOut47[18] , \nScanOut47[17] , 
        \nScanOut47[16] , \nScanOut47[15] , \nScanOut47[14] , \nScanOut47[13] , 
        \nScanOut47[12] , \nScanOut47[11] , \nScanOut47[10] , \nScanOut47[9] , 
        \nScanOut47[8] , \nScanOut47[7] , \nScanOut47[6] , \nScanOut47[5] , 
        \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , \nScanOut47[1] , 
        \nScanOut47[0] }), .ScanOut({\nScanOut46[31] , \nScanOut46[30] , 
        \nScanOut46[29] , \nScanOut46[28] , \nScanOut46[27] , \nScanOut46[26] , 
        \nScanOut46[25] , \nScanOut46[24] , \nScanOut46[23] , \nScanOut46[22] , 
        \nScanOut46[21] , \nScanOut46[20] , \nScanOut46[19] , \nScanOut46[18] , 
        \nScanOut46[17] , \nScanOut46[16] , \nScanOut46[15] , \nScanOut46[14] , 
        \nScanOut46[13] , \nScanOut46[12] , \nScanOut46[11] , \nScanOut46[10] , 
        \nScanOut46[9] , \nScanOut46[8] , \nScanOut46[7] , \nScanOut46[6] , 
        \nScanOut46[5] , \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , 
        \nScanOut46[1] , \nScanOut46[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_14[31] , 
        \nOut2_14[30] , \nOut2_14[29] , \nOut2_14[28] , \nOut2_14[27] , 
        \nOut2_14[26] , \nOut2_14[25] , \nOut2_14[24] , \nOut2_14[23] , 
        \nOut2_14[22] , \nOut2_14[21] , \nOut2_14[20] , \nOut2_14[19] , 
        \nOut2_14[18] , \nOut2_14[17] , \nOut2_14[16] , \nOut2_14[15] , 
        \nOut2_14[14] , \nOut2_14[13] , \nOut2_14[12] , \nOut2_14[11] , 
        \nOut2_14[10] , \nOut2_14[9] , \nOut2_14[8] , \nOut2_14[7] , 
        \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , \nOut2_14[3] , 
        \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), .NORTH_EDGE({
        \nOut2_13[31] , \nOut2_13[30] , \nOut2_13[29] , \nOut2_13[28] , 
        \nOut2_13[27] , \nOut2_13[26] , \nOut2_13[25] , \nOut2_13[24] , 
        \nOut2_13[23] , \nOut2_13[22] , \nOut2_13[21] , \nOut2_13[20] , 
        \nOut2_13[19] , \nOut2_13[18] , \nOut2_13[17] , \nOut2_13[16] , 
        \nOut2_13[15] , \nOut2_13[14] , \nOut2_13[13] , \nOut2_13[12] , 
        \nOut2_13[11] , \nOut2_13[10] , \nOut2_13[9] , \nOut2_13[8] , 
        \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , 
        \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), 
        .SOUTH_EDGE({\nOut2_15[31] , \nOut2_15[30] , \nOut2_15[29] , 
        \nOut2_15[28] , \nOut2_15[27] , \nOut2_15[26] , \nOut2_15[25] , 
        \nOut2_15[24] , \nOut2_15[23] , \nOut2_15[22] , \nOut2_15[21] , 
        \nOut2_15[20] , \nOut2_15[19] , \nOut2_15[18] , \nOut2_15[17] , 
        \nOut2_15[16] , \nOut2_15[15] , \nOut2_15[14] , \nOut2_15[13] , 
        \nOut2_15[12] , \nOut2_15[11] , \nOut2_15[10] , \nOut2_15[9] , 
        \nOut2_15[8] , \nOut2_15[7] , \nOut2_15[6] , \nOut2_15[5] , 
        \nOut2_15[4] , \nOut2_15[3] , \nOut2_15[2] , \nOut2_15[1] , 
        \nOut2_15[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_14[0] ), 
        .NW_EDGE(\nOut1_13[0] ), .SW_EDGE(\nOut1_15[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_41 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut42[31] , \nScanOut42[30] , \nScanOut42[29] , 
        \nScanOut42[28] , \nScanOut42[27] , \nScanOut42[26] , \nScanOut42[25] , 
        \nScanOut42[24] , \nScanOut42[23] , \nScanOut42[22] , \nScanOut42[21] , 
        \nScanOut42[20] , \nScanOut42[19] , \nScanOut42[18] , \nScanOut42[17] , 
        \nScanOut42[16] , \nScanOut42[15] , \nScanOut42[14] , \nScanOut42[13] , 
        \nScanOut42[12] , \nScanOut42[11] , \nScanOut42[10] , \nScanOut42[9] , 
        \nScanOut42[8] , \nScanOut42[7] , \nScanOut42[6] , \nScanOut42[5] , 
        \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , \nScanOut42[1] , 
        \nScanOut42[0] }), .ScanOut({\nScanOut41[31] , \nScanOut41[30] , 
        \nScanOut41[29] , \nScanOut41[28] , \nScanOut41[27] , \nScanOut41[26] , 
        \nScanOut41[25] , \nScanOut41[24] , \nScanOut41[23] , \nScanOut41[22] , 
        \nScanOut41[21] , \nScanOut41[20] , \nScanOut41[19] , \nScanOut41[18] , 
        \nScanOut41[17] , \nScanOut41[16] , \nScanOut41[15] , \nScanOut41[14] , 
        \nScanOut41[13] , \nScanOut41[12] , \nScanOut41[11] , \nScanOut41[10] , 
        \nScanOut41[9] , \nScanOut41[8] , \nScanOut41[7] , \nScanOut41[6] , 
        \nScanOut41[5] , \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , 
        \nScanOut41[1] , \nScanOut41[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_9[31] , 
        \nOut2_9[30] , \nOut2_9[29] , \nOut2_9[28] , \nOut2_9[27] , 
        \nOut2_9[26] , \nOut2_9[25] , \nOut2_9[24] , \nOut2_9[23] , 
        \nOut2_9[22] , \nOut2_9[21] , \nOut2_9[20] , \nOut2_9[19] , 
        \nOut2_9[18] , \nOut2_9[17] , \nOut2_9[16] , \nOut2_9[15] , 
        \nOut2_9[14] , \nOut2_9[13] , \nOut2_9[12] , \nOut2_9[11] , 
        \nOut2_9[10] , \nOut2_9[9] , \nOut2_9[8] , \nOut2_9[7] , \nOut2_9[6] , 
        \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , 
        \nOut2_9[0] }), .NORTH_EDGE({\nOut2_8[31] , \nOut2_8[30] , 
        \nOut2_8[29] , \nOut2_8[28] , \nOut2_8[27] , \nOut2_8[26] , 
        \nOut2_8[25] , \nOut2_8[24] , \nOut2_8[23] , \nOut2_8[22] , 
        \nOut2_8[21] , \nOut2_8[20] , \nOut2_8[19] , \nOut2_8[18] , 
        \nOut2_8[17] , \nOut2_8[16] , \nOut2_8[15] , \nOut2_8[14] , 
        \nOut2_8[13] , \nOut2_8[12] , \nOut2_8[11] , \nOut2_8[10] , 
        \nOut2_8[9] , \nOut2_8[8] , \nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , 
        \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), 
        .SOUTH_EDGE({\nOut2_10[31] , \nOut2_10[30] , \nOut2_10[29] , 
        \nOut2_10[28] , \nOut2_10[27] , \nOut2_10[26] , \nOut2_10[25] , 
        \nOut2_10[24] , \nOut2_10[23] , \nOut2_10[22] , \nOut2_10[21] , 
        \nOut2_10[20] , \nOut2_10[19] , \nOut2_10[18] , \nOut2_10[17] , 
        \nOut2_10[16] , \nOut2_10[15] , \nOut2_10[14] , \nOut2_10[13] , 
        \nOut2_10[12] , \nOut2_10[11] , \nOut2_10[10] , \nOut2_10[9] , 
        \nOut2_10[8] , \nOut2_10[7] , \nOut2_10[6] , \nOut2_10[5] , 
        \nOut2_10[4] , \nOut2_10[3] , \nOut2_10[2] , \nOut2_10[1] , 
        \nOut2_10[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_9[0] ), .NW_EDGE(
        \nOut1_8[0] ), .SW_EDGE(\nOut1_10[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0)
         );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_26 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut27[31] , \nScanOut27[30] , \nScanOut27[29] , 
        \nScanOut27[28] , \nScanOut27[27] , \nScanOut27[26] , \nScanOut27[25] , 
        \nScanOut27[24] , \nScanOut27[23] , \nScanOut27[22] , \nScanOut27[21] , 
        \nScanOut27[20] , \nScanOut27[19] , \nScanOut27[18] , \nScanOut27[17] , 
        \nScanOut27[16] , \nScanOut27[15] , \nScanOut27[14] , \nScanOut27[13] , 
        \nScanOut27[12] , \nScanOut27[11] , \nScanOut27[10] , \nScanOut27[9] , 
        \nScanOut27[8] , \nScanOut27[7] , \nScanOut27[6] , \nScanOut27[5] , 
        \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , \nScanOut27[1] , 
        \nScanOut27[0] }), .ScanOut({\nScanOut26[31] , \nScanOut26[30] , 
        \nScanOut26[29] , \nScanOut26[28] , \nScanOut26[27] , \nScanOut26[26] , 
        \nScanOut26[25] , \nScanOut26[24] , \nScanOut26[23] , \nScanOut26[22] , 
        \nScanOut26[21] , \nScanOut26[20] , \nScanOut26[19] , \nScanOut26[18] , 
        \nScanOut26[17] , \nScanOut26[16] , \nScanOut26[15] , \nScanOut26[14] , 
        \nScanOut26[13] , \nScanOut26[12] , \nScanOut26[11] , \nScanOut26[10] , 
        \nScanOut26[9] , \nScanOut26[8] , \nScanOut26[7] , \nScanOut26[6] , 
        \nScanOut26[5] , \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , 
        \nScanOut26[1] , \nScanOut26[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_10[31] , 
        \nOut1_10[30] , \nOut1_10[29] , \nOut1_10[28] , \nOut1_10[27] , 
        \nOut1_10[26] , \nOut1_10[25] , \nOut1_10[24] , \nOut1_10[23] , 
        \nOut1_10[22] , \nOut1_10[21] , \nOut1_10[20] , \nOut1_10[19] , 
        \nOut1_10[18] , \nOut1_10[17] , \nOut1_10[16] , \nOut1_10[15] , 
        \nOut1_10[14] , \nOut1_10[13] , \nOut1_10[12] , \nOut1_10[11] , 
        \nOut1_10[10] , \nOut1_10[9] , \nOut1_10[8] , \nOut1_10[7] , 
        \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , \nOut1_10[3] , 
        \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), .NORTH_EDGE({
        \nOut1_9[31] , \nOut1_9[30] , \nOut1_9[29] , \nOut1_9[28] , 
        \nOut1_9[27] , \nOut1_9[26] , \nOut1_9[25] , \nOut1_9[24] , 
        \nOut1_9[23] , \nOut1_9[22] , \nOut1_9[21] , \nOut1_9[20] , 
        \nOut1_9[19] , \nOut1_9[18] , \nOut1_9[17] , \nOut1_9[16] , 
        \nOut1_9[15] , \nOut1_9[14] , \nOut1_9[13] , \nOut1_9[12] , 
        \nOut1_9[11] , \nOut1_9[10] , \nOut1_9[9] , \nOut1_9[8] , \nOut1_9[7] , 
        \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , 
        \nOut1_9[1] , \nOut1_9[0] }), .SOUTH_EDGE({\nOut1_11[31] , 
        \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , \nOut1_11[27] , 
        \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , \nOut1_11[23] , 
        \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , \nOut1_11[19] , 
        \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , \nOut1_11[15] , 
        \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , \nOut1_11[11] , 
        \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , \nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .EAST_EDGE(
        \nOut2_10[31] ), .WEST_EDGE(\nOut0_10[0] ), .NW_EDGE(\nOut0_9[0] ), 
        .SW_EDGE(\nOut0_11[0] ), .NE_EDGE(\nOut2_9[31] ), .SE_EDGE(
        \nOut2_11[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_34 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut35[31] , \nScanOut35[30] , \nScanOut35[29] , 
        \nScanOut35[28] , \nScanOut35[27] , \nScanOut35[26] , \nScanOut35[25] , 
        \nScanOut35[24] , \nScanOut35[23] , \nScanOut35[22] , \nScanOut35[21] , 
        \nScanOut35[20] , \nScanOut35[19] , \nScanOut35[18] , \nScanOut35[17] , 
        \nScanOut35[16] , \nScanOut35[15] , \nScanOut35[14] , \nScanOut35[13] , 
        \nScanOut35[12] , \nScanOut35[11] , \nScanOut35[10] , \nScanOut35[9] , 
        \nScanOut35[8] , \nScanOut35[7] , \nScanOut35[6] , \nScanOut35[5] , 
        \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , \nScanOut35[1] , 
        \nScanOut35[0] }), .ScanOut({\nScanOut34[31] , \nScanOut34[30] , 
        \nScanOut34[29] , \nScanOut34[28] , \nScanOut34[27] , \nScanOut34[26] , 
        \nScanOut34[25] , \nScanOut34[24] , \nScanOut34[23] , \nScanOut34[22] , 
        \nScanOut34[21] , \nScanOut34[20] , \nScanOut34[19] , \nScanOut34[18] , 
        \nScanOut34[17] , \nScanOut34[16] , \nScanOut34[15] , \nScanOut34[14] , 
        \nScanOut34[13] , \nScanOut34[12] , \nScanOut34[11] , \nScanOut34[10] , 
        \nScanOut34[9] , \nScanOut34[8] , \nScanOut34[7] , \nScanOut34[6] , 
        \nScanOut34[5] , \nScanOut34[4] , \nScanOut34[3] , \nScanOut34[2] , 
        \nScanOut34[1] , \nScanOut34[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_2[31] , 
        \nOut2_2[30] , \nOut2_2[29] , \nOut2_2[28] , \nOut2_2[27] , 
        \nOut2_2[26] , \nOut2_2[25] , \nOut2_2[24] , \nOut2_2[23] , 
        \nOut2_2[22] , \nOut2_2[21] , \nOut2_2[20] , \nOut2_2[19] , 
        \nOut2_2[18] , \nOut2_2[17] , \nOut2_2[16] , \nOut2_2[15] , 
        \nOut2_2[14] , \nOut2_2[13] , \nOut2_2[12] , \nOut2_2[11] , 
        \nOut2_2[10] , \nOut2_2[9] , \nOut2_2[8] , \nOut2_2[7] , \nOut2_2[6] , 
        \nOut2_2[5] , \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , 
        \nOut2_2[0] }), .NORTH_EDGE({\nOut2_1[31] , \nOut2_1[30] , 
        \nOut2_1[29] , \nOut2_1[28] , \nOut2_1[27] , \nOut2_1[26] , 
        \nOut2_1[25] , \nOut2_1[24] , \nOut2_1[23] , \nOut2_1[22] , 
        \nOut2_1[21] , \nOut2_1[20] , \nOut2_1[19] , \nOut2_1[18] , 
        \nOut2_1[17] , \nOut2_1[16] , \nOut2_1[15] , \nOut2_1[14] , 
        \nOut2_1[13] , \nOut2_1[12] , \nOut2_1[11] , \nOut2_1[10] , 
        \nOut2_1[9] , \nOut2_1[8] , \nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , 
        \nOut2_1[4] , \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), 
        .SOUTH_EDGE({\nOut2_3[31] , \nOut2_3[30] , \nOut2_3[29] , 
        \nOut2_3[28] , \nOut2_3[27] , \nOut2_3[26] , \nOut2_3[25] , 
        \nOut2_3[24] , \nOut2_3[23] , \nOut2_3[22] , \nOut2_3[21] , 
        \nOut2_3[20] , \nOut2_3[19] , \nOut2_3[18] , \nOut2_3[17] , 
        \nOut2_3[16] , \nOut2_3[15] , \nOut2_3[14] , \nOut2_3[13] , 
        \nOut2_3[12] , \nOut2_3[11] , \nOut2_3[10] , \nOut2_3[9] , 
        \nOut2_3[8] , \nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , \nOut2_3[4] , 
        \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_2[0] ), .NW_EDGE(\nOut1_1[0] ), .SW_EDGE(
        \nOut1_3[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_5 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut6[31] , \nScanOut6[30] , \nScanOut6[29] , 
        \nScanOut6[28] , \nScanOut6[27] , \nScanOut6[26] , \nScanOut6[25] , 
        \nScanOut6[24] , \nScanOut6[23] , \nScanOut6[22] , \nScanOut6[21] , 
        \nScanOut6[20] , \nScanOut6[19] , \nScanOut6[18] , \nScanOut6[17] , 
        \nScanOut6[16] , \nScanOut6[15] , \nScanOut6[14] , \nScanOut6[13] , 
        \nScanOut6[12] , \nScanOut6[11] , \nScanOut6[10] , \nScanOut6[9] , 
        \nScanOut6[8] , \nScanOut6[7] , \nScanOut6[6] , \nScanOut6[5] , 
        \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , \nScanOut6[1] , 
        \nScanOut6[0] }), .ScanOut({\nScanOut5[31] , \nScanOut5[30] , 
        \nScanOut5[29] , \nScanOut5[28] , \nScanOut5[27] , \nScanOut5[26] , 
        \nScanOut5[25] , \nScanOut5[24] , \nScanOut5[23] , \nScanOut5[22] , 
        \nScanOut5[21] , \nScanOut5[20] , \nScanOut5[19] , \nScanOut5[18] , 
        \nScanOut5[17] , \nScanOut5[16] , \nScanOut5[15] , \nScanOut5[14] , 
        \nScanOut5[13] , \nScanOut5[12] , \nScanOut5[11] , \nScanOut5[10] , 
        \nScanOut5[9] , \nScanOut5[8] , \nScanOut5[7] , \nScanOut5[6] , 
        \nScanOut5[5] , \nScanOut5[4] , \nScanOut5[3] , \nScanOut5[2] , 
        \nScanOut5[1] , \nScanOut5[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_5[31] , 
        \nOut0_5[30] , \nOut0_5[29] , \nOut0_5[28] , \nOut0_5[27] , 
        \nOut0_5[26] , \nOut0_5[25] , \nOut0_5[24] , \nOut0_5[23] , 
        \nOut0_5[22] , \nOut0_5[21] , \nOut0_5[20] , \nOut0_5[19] , 
        \nOut0_5[18] , \nOut0_5[17] , \nOut0_5[16] , \nOut0_5[15] , 
        \nOut0_5[14] , \nOut0_5[13] , \nOut0_5[12] , \nOut0_5[11] , 
        \nOut0_5[10] , \nOut0_5[9] , \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , 
        \nOut0_5[5] , \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , 
        \nOut0_5[0] }), .NORTH_EDGE({\nOut0_4[31] , \nOut0_4[30] , 
        \nOut0_4[29] , \nOut0_4[28] , \nOut0_4[27] , \nOut0_4[26] , 
        \nOut0_4[25] , \nOut0_4[24] , \nOut0_4[23] , \nOut0_4[22] , 
        \nOut0_4[21] , \nOut0_4[20] , \nOut0_4[19] , \nOut0_4[18] , 
        \nOut0_4[17] , \nOut0_4[16] , \nOut0_4[15] , \nOut0_4[14] , 
        \nOut0_4[13] , \nOut0_4[12] , \nOut0_4[11] , \nOut0_4[10] , 
        \nOut0_4[9] , \nOut0_4[8] , \nOut0_4[7] , \nOut0_4[6] , \nOut0_4[5] , 
        \nOut0_4[4] , \nOut0_4[3] , \nOut0_4[2] , \nOut0_4[1] , \nOut0_4[0] }), 
        .SOUTH_EDGE({\nOut0_6[31] , \nOut0_6[30] , \nOut0_6[29] , 
        \nOut0_6[28] , \nOut0_6[27] , \nOut0_6[26] , \nOut0_6[25] , 
        \nOut0_6[24] , \nOut0_6[23] , \nOut0_6[22] , \nOut0_6[21] , 
        \nOut0_6[20] , \nOut0_6[19] , \nOut0_6[18] , \nOut0_6[17] , 
        \nOut0_6[16] , \nOut0_6[15] , \nOut0_6[14] , \nOut0_6[13] , 
        \nOut0_6[12] , \nOut0_6[11] , \nOut0_6[10] , \nOut0_6[9] , 
        \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , \nOut0_6[4] , 
        \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), .EAST_EDGE(
        \nOut1_5[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_4[31] ), .SE_EDGE(\nOut1_6[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_12 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut13[31] , \nScanOut13[30] , \nScanOut13[29] , 
        \nScanOut13[28] , \nScanOut13[27] , \nScanOut13[26] , \nScanOut13[25] , 
        \nScanOut13[24] , \nScanOut13[23] , \nScanOut13[22] , \nScanOut13[21] , 
        \nScanOut13[20] , \nScanOut13[19] , \nScanOut13[18] , \nScanOut13[17] , 
        \nScanOut13[16] , \nScanOut13[15] , \nScanOut13[14] , \nScanOut13[13] , 
        \nScanOut13[12] , \nScanOut13[11] , \nScanOut13[10] , \nScanOut13[9] , 
        \nScanOut13[8] , \nScanOut13[7] , \nScanOut13[6] , \nScanOut13[5] , 
        \nScanOut13[4] , \nScanOut13[3] , \nScanOut13[2] , \nScanOut13[1] , 
        \nScanOut13[0] }), .ScanOut({\nScanOut12[31] , \nScanOut12[30] , 
        \nScanOut12[29] , \nScanOut12[28] , \nScanOut12[27] , \nScanOut12[26] , 
        \nScanOut12[25] , \nScanOut12[24] , \nScanOut12[23] , \nScanOut12[22] , 
        \nScanOut12[21] , \nScanOut12[20] , \nScanOut12[19] , \nScanOut12[18] , 
        \nScanOut12[17] , \nScanOut12[16] , \nScanOut12[15] , \nScanOut12[14] , 
        \nScanOut12[13] , \nScanOut12[12] , \nScanOut12[11] , \nScanOut12[10] , 
        \nScanOut12[9] , \nScanOut12[8] , \nScanOut12[7] , \nScanOut12[6] , 
        \nScanOut12[5] , \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , 
        \nScanOut12[1] , \nScanOut12[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_12[31] , 
        \nOut0_12[30] , \nOut0_12[29] , \nOut0_12[28] , \nOut0_12[27] , 
        \nOut0_12[26] , \nOut0_12[25] , \nOut0_12[24] , \nOut0_12[23] , 
        \nOut0_12[22] , \nOut0_12[21] , \nOut0_12[20] , \nOut0_12[19] , 
        \nOut0_12[18] , \nOut0_12[17] , \nOut0_12[16] , \nOut0_12[15] , 
        \nOut0_12[14] , \nOut0_12[13] , \nOut0_12[12] , \nOut0_12[11] , 
        \nOut0_12[10] , \nOut0_12[9] , \nOut0_12[8] , \nOut0_12[7] , 
        \nOut0_12[6] , \nOut0_12[5] , \nOut0_12[4] , \nOut0_12[3] , 
        \nOut0_12[2] , \nOut0_12[1] , \nOut0_12[0] }), .NORTH_EDGE({
        \nOut0_11[31] , \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , 
        \nOut0_11[27] , \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , 
        \nOut0_11[23] , \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , 
        \nOut0_11[19] , \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , 
        \nOut0_11[15] , \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , 
        \nOut0_11[11] , \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , 
        \nOut0_11[7] , \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , 
        \nOut0_11[3] , \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), 
        .SOUTH_EDGE({\nOut0_13[31] , \nOut0_13[30] , \nOut0_13[29] , 
        \nOut0_13[28] , \nOut0_13[27] , \nOut0_13[26] , \nOut0_13[25] , 
        \nOut0_13[24] , \nOut0_13[23] , \nOut0_13[22] , \nOut0_13[21] , 
        \nOut0_13[20] , \nOut0_13[19] , \nOut0_13[18] , \nOut0_13[17] , 
        \nOut0_13[16] , \nOut0_13[15] , \nOut0_13[14] , \nOut0_13[13] , 
        \nOut0_13[12] , \nOut0_13[11] , \nOut0_13[10] , \nOut0_13[9] , 
        \nOut0_13[8] , \nOut0_13[7] , \nOut0_13[6] , \nOut0_13[5] , 
        \nOut0_13[4] , \nOut0_13[3] , \nOut0_13[2] , \nOut0_13[1] , 
        \nOut0_13[0] }), .EAST_EDGE(\nOut1_12[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_11[31] ), .SE_EDGE(
        \nOut1_13[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_35 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut36[31] , \nScanOut36[30] , \nScanOut36[29] , 
        \nScanOut36[28] , \nScanOut36[27] , \nScanOut36[26] , \nScanOut36[25] , 
        \nScanOut36[24] , \nScanOut36[23] , \nScanOut36[22] , \nScanOut36[21] , 
        \nScanOut36[20] , \nScanOut36[19] , \nScanOut36[18] , \nScanOut36[17] , 
        \nScanOut36[16] , \nScanOut36[15] , \nScanOut36[14] , \nScanOut36[13] , 
        \nScanOut36[12] , \nScanOut36[11] , \nScanOut36[10] , \nScanOut36[9] , 
        \nScanOut36[8] , \nScanOut36[7] , \nScanOut36[6] , \nScanOut36[5] , 
        \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , \nScanOut36[1] , 
        \nScanOut36[0] }), .ScanOut({\nScanOut35[31] , \nScanOut35[30] , 
        \nScanOut35[29] , \nScanOut35[28] , \nScanOut35[27] , \nScanOut35[26] , 
        \nScanOut35[25] , \nScanOut35[24] , \nScanOut35[23] , \nScanOut35[22] , 
        \nScanOut35[21] , \nScanOut35[20] , \nScanOut35[19] , \nScanOut35[18] , 
        \nScanOut35[17] , \nScanOut35[16] , \nScanOut35[15] , \nScanOut35[14] , 
        \nScanOut35[13] , \nScanOut35[12] , \nScanOut35[11] , \nScanOut35[10] , 
        \nScanOut35[9] , \nScanOut35[8] , \nScanOut35[7] , \nScanOut35[6] , 
        \nScanOut35[5] , \nScanOut35[4] , \nScanOut35[3] , \nScanOut35[2] , 
        \nScanOut35[1] , \nScanOut35[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_3[31] , 
        \nOut2_3[30] , \nOut2_3[29] , \nOut2_3[28] , \nOut2_3[27] , 
        \nOut2_3[26] , \nOut2_3[25] , \nOut2_3[24] , \nOut2_3[23] , 
        \nOut2_3[22] , \nOut2_3[21] , \nOut2_3[20] , \nOut2_3[19] , 
        \nOut2_3[18] , \nOut2_3[17] , \nOut2_3[16] , \nOut2_3[15] , 
        \nOut2_3[14] , \nOut2_3[13] , \nOut2_3[12] , \nOut2_3[11] , 
        \nOut2_3[10] , \nOut2_3[9] , \nOut2_3[8] , \nOut2_3[7] , \nOut2_3[6] , 
        \nOut2_3[5] , \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , 
        \nOut2_3[0] }), .NORTH_EDGE({\nOut2_2[31] , \nOut2_2[30] , 
        \nOut2_2[29] , \nOut2_2[28] , \nOut2_2[27] , \nOut2_2[26] , 
        \nOut2_2[25] , \nOut2_2[24] , \nOut2_2[23] , \nOut2_2[22] , 
        \nOut2_2[21] , \nOut2_2[20] , \nOut2_2[19] , \nOut2_2[18] , 
        \nOut2_2[17] , \nOut2_2[16] , \nOut2_2[15] , \nOut2_2[14] , 
        \nOut2_2[13] , \nOut2_2[12] , \nOut2_2[11] , \nOut2_2[10] , 
        \nOut2_2[9] , \nOut2_2[8] , \nOut2_2[7] , \nOut2_2[6] , \nOut2_2[5] , 
        \nOut2_2[4] , \nOut2_2[3] , \nOut2_2[2] , \nOut2_2[1] , \nOut2_2[0] }), 
        .SOUTH_EDGE({\nOut2_4[31] , \nOut2_4[30] , \nOut2_4[29] , 
        \nOut2_4[28] , \nOut2_4[27] , \nOut2_4[26] , \nOut2_4[25] , 
        \nOut2_4[24] , \nOut2_4[23] , \nOut2_4[22] , \nOut2_4[21] , 
        \nOut2_4[20] , \nOut2_4[19] , \nOut2_4[18] , \nOut2_4[17] , 
        \nOut2_4[16] , \nOut2_4[15] , \nOut2_4[14] , \nOut2_4[13] , 
        \nOut2_4[12] , \nOut2_4[11] , \nOut2_4[10] , \nOut2_4[9] , 
        \nOut2_4[8] , \nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , \nOut2_4[4] , 
        \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_3[0] ), .NW_EDGE(\nOut1_2[0] ), .SW_EDGE(
        \nOut1_4[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_40 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut41[31] , \nScanOut41[30] , \nScanOut41[29] , 
        \nScanOut41[28] , \nScanOut41[27] , \nScanOut41[26] , \nScanOut41[25] , 
        \nScanOut41[24] , \nScanOut41[23] , \nScanOut41[22] , \nScanOut41[21] , 
        \nScanOut41[20] , \nScanOut41[19] , \nScanOut41[18] , \nScanOut41[17] , 
        \nScanOut41[16] , \nScanOut41[15] , \nScanOut41[14] , \nScanOut41[13] , 
        \nScanOut41[12] , \nScanOut41[11] , \nScanOut41[10] , \nScanOut41[9] , 
        \nScanOut41[8] , \nScanOut41[7] , \nScanOut41[6] , \nScanOut41[5] , 
        \nScanOut41[4] , \nScanOut41[3] , \nScanOut41[2] , \nScanOut41[1] , 
        \nScanOut41[0] }), .ScanOut({\nScanOut40[31] , \nScanOut40[30] , 
        \nScanOut40[29] , \nScanOut40[28] , \nScanOut40[27] , \nScanOut40[26] , 
        \nScanOut40[25] , \nScanOut40[24] , \nScanOut40[23] , \nScanOut40[22] , 
        \nScanOut40[21] , \nScanOut40[20] , \nScanOut40[19] , \nScanOut40[18] , 
        \nScanOut40[17] , \nScanOut40[16] , \nScanOut40[15] , \nScanOut40[14] , 
        \nScanOut40[13] , \nScanOut40[12] , \nScanOut40[11] , \nScanOut40[10] , 
        \nScanOut40[9] , \nScanOut40[8] , \nScanOut40[7] , \nScanOut40[6] , 
        \nScanOut40[5] , \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , 
        \nScanOut40[1] , \nScanOut40[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_8[31] , 
        \nOut2_8[30] , \nOut2_8[29] , \nOut2_8[28] , \nOut2_8[27] , 
        \nOut2_8[26] , \nOut2_8[25] , \nOut2_8[24] , \nOut2_8[23] , 
        \nOut2_8[22] , \nOut2_8[21] , \nOut2_8[20] , \nOut2_8[19] , 
        \nOut2_8[18] , \nOut2_8[17] , \nOut2_8[16] , \nOut2_8[15] , 
        \nOut2_8[14] , \nOut2_8[13] , \nOut2_8[12] , \nOut2_8[11] , 
        \nOut2_8[10] , \nOut2_8[9] , \nOut2_8[8] , \nOut2_8[7] , \nOut2_8[6] , 
        \nOut2_8[5] , \nOut2_8[4] , \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , 
        \nOut2_8[0] }), .NORTH_EDGE({\nOut2_7[31] , \nOut2_7[30] , 
        \nOut2_7[29] , \nOut2_7[28] , \nOut2_7[27] , \nOut2_7[26] , 
        \nOut2_7[25] , \nOut2_7[24] , \nOut2_7[23] , \nOut2_7[22] , 
        \nOut2_7[21] , \nOut2_7[20] , \nOut2_7[19] , \nOut2_7[18] , 
        \nOut2_7[17] , \nOut2_7[16] , \nOut2_7[15] , \nOut2_7[14] , 
        \nOut2_7[13] , \nOut2_7[12] , \nOut2_7[11] , \nOut2_7[10] , 
        \nOut2_7[9] , \nOut2_7[8] , \nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , 
        \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), 
        .SOUTH_EDGE({\nOut2_9[31] , \nOut2_9[30] , \nOut2_9[29] , 
        \nOut2_9[28] , \nOut2_9[27] , \nOut2_9[26] , \nOut2_9[25] , 
        \nOut2_9[24] , \nOut2_9[23] , \nOut2_9[22] , \nOut2_9[21] , 
        \nOut2_9[20] , \nOut2_9[19] , \nOut2_9[18] , \nOut2_9[17] , 
        \nOut2_9[16] , \nOut2_9[15] , \nOut2_9[14] , \nOut2_9[13] , 
        \nOut2_9[12] , \nOut2_9[11] , \nOut2_9[10] , \nOut2_9[9] , 
        \nOut2_9[8] , \nOut2_9[7] , \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , 
        \nOut2_9[3] , \nOut2_9[2] , \nOut2_9[1] , \nOut2_9[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_8[0] ), .NW_EDGE(\nOut1_7[0] ), .SW_EDGE(
        \nOut1_9[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_20 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut21[31] , \nScanOut21[30] , \nScanOut21[29] , 
        \nScanOut21[28] , \nScanOut21[27] , \nScanOut21[26] , \nScanOut21[25] , 
        \nScanOut21[24] , \nScanOut21[23] , \nScanOut21[22] , \nScanOut21[21] , 
        \nScanOut21[20] , \nScanOut21[19] , \nScanOut21[18] , \nScanOut21[17] , 
        \nScanOut21[16] , \nScanOut21[15] , \nScanOut21[14] , \nScanOut21[13] , 
        \nScanOut21[12] , \nScanOut21[11] , \nScanOut21[10] , \nScanOut21[9] , 
        \nScanOut21[8] , \nScanOut21[7] , \nScanOut21[6] , \nScanOut21[5] , 
        \nScanOut21[4] , \nScanOut21[3] , \nScanOut21[2] , \nScanOut21[1] , 
        \nScanOut21[0] }), .ScanOut({\nScanOut20[31] , \nScanOut20[30] , 
        \nScanOut20[29] , \nScanOut20[28] , \nScanOut20[27] , \nScanOut20[26] , 
        \nScanOut20[25] , \nScanOut20[24] , \nScanOut20[23] , \nScanOut20[22] , 
        \nScanOut20[21] , \nScanOut20[20] , \nScanOut20[19] , \nScanOut20[18] , 
        \nScanOut20[17] , \nScanOut20[16] , \nScanOut20[15] , \nScanOut20[14] , 
        \nScanOut20[13] , \nScanOut20[12] , \nScanOut20[11] , \nScanOut20[10] , 
        \nScanOut20[9] , \nScanOut20[8] , \nScanOut20[7] , \nScanOut20[6] , 
        \nScanOut20[5] , \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , 
        \nScanOut20[1] , \nScanOut20[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_4[31] , 
        \nOut1_4[30] , \nOut1_4[29] , \nOut1_4[28] , \nOut1_4[27] , 
        \nOut1_4[26] , \nOut1_4[25] , \nOut1_4[24] , \nOut1_4[23] , 
        \nOut1_4[22] , \nOut1_4[21] , \nOut1_4[20] , \nOut1_4[19] , 
        \nOut1_4[18] , \nOut1_4[17] , \nOut1_4[16] , \nOut1_4[15] , 
        \nOut1_4[14] , \nOut1_4[13] , \nOut1_4[12] , \nOut1_4[11] , 
        \nOut1_4[10] , \nOut1_4[9] , \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , 
        \nOut1_4[5] , \nOut1_4[4] , \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , 
        \nOut1_4[0] }), .NORTH_EDGE({\nOut1_3[31] , \nOut1_3[30] , 
        \nOut1_3[29] , \nOut1_3[28] , \nOut1_3[27] , \nOut1_3[26] , 
        \nOut1_3[25] , \nOut1_3[24] , \nOut1_3[23] , \nOut1_3[22] , 
        \nOut1_3[21] , \nOut1_3[20] , \nOut1_3[19] , \nOut1_3[18] , 
        \nOut1_3[17] , \nOut1_3[16] , \nOut1_3[15] , \nOut1_3[14] , 
        \nOut1_3[13] , \nOut1_3[12] , \nOut1_3[11] , \nOut1_3[10] , 
        \nOut1_3[9] , \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , 
        \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), 
        .SOUTH_EDGE({\nOut1_5[31] , \nOut1_5[30] , \nOut1_5[29] , 
        \nOut1_5[28] , \nOut1_5[27] , \nOut1_5[26] , \nOut1_5[25] , 
        \nOut1_5[24] , \nOut1_5[23] , \nOut1_5[22] , \nOut1_5[21] , 
        \nOut1_5[20] , \nOut1_5[19] , \nOut1_5[18] , \nOut1_5[17] , 
        \nOut1_5[16] , \nOut1_5[15] , \nOut1_5[14] , \nOut1_5[13] , 
        \nOut1_5[12] , \nOut1_5[11] , \nOut1_5[10] , \nOut1_5[9] , 
        \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , \nOut1_5[4] , 
        \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), .EAST_EDGE(
        \nOut2_4[31] ), .WEST_EDGE(\nOut0_4[0] ), .NW_EDGE(\nOut0_3[0] ), 
        .SW_EDGE(\nOut0_5[0] ), .NE_EDGE(\nOut2_3[31] ), .SE_EDGE(
        \nOut2_5[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_27 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut28[31] , \nScanOut28[30] , \nScanOut28[29] , 
        \nScanOut28[28] , \nScanOut28[27] , \nScanOut28[26] , \nScanOut28[25] , 
        \nScanOut28[24] , \nScanOut28[23] , \nScanOut28[22] , \nScanOut28[21] , 
        \nScanOut28[20] , \nScanOut28[19] , \nScanOut28[18] , \nScanOut28[17] , 
        \nScanOut28[16] , \nScanOut28[15] , \nScanOut28[14] , \nScanOut28[13] , 
        \nScanOut28[12] , \nScanOut28[11] , \nScanOut28[10] , \nScanOut28[9] , 
        \nScanOut28[8] , \nScanOut28[7] , \nScanOut28[6] , \nScanOut28[5] , 
        \nScanOut28[4] , \nScanOut28[3] , \nScanOut28[2] , \nScanOut28[1] , 
        \nScanOut28[0] }), .ScanOut({\nScanOut27[31] , \nScanOut27[30] , 
        \nScanOut27[29] , \nScanOut27[28] , \nScanOut27[27] , \nScanOut27[26] , 
        \nScanOut27[25] , \nScanOut27[24] , \nScanOut27[23] , \nScanOut27[22] , 
        \nScanOut27[21] , \nScanOut27[20] , \nScanOut27[19] , \nScanOut27[18] , 
        \nScanOut27[17] , \nScanOut27[16] , \nScanOut27[15] , \nScanOut27[14] , 
        \nScanOut27[13] , \nScanOut27[12] , \nScanOut27[11] , \nScanOut27[10] , 
        \nScanOut27[9] , \nScanOut27[8] , \nScanOut27[7] , \nScanOut27[6] , 
        \nScanOut27[5] , \nScanOut27[4] , \nScanOut27[3] , \nScanOut27[2] , 
        \nScanOut27[1] , \nScanOut27[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_11[31] , 
        \nOut1_11[30] , \nOut1_11[29] , \nOut1_11[28] , \nOut1_11[27] , 
        \nOut1_11[26] , \nOut1_11[25] , \nOut1_11[24] , \nOut1_11[23] , 
        \nOut1_11[22] , \nOut1_11[21] , \nOut1_11[20] , \nOut1_11[19] , 
        \nOut1_11[18] , \nOut1_11[17] , \nOut1_11[16] , \nOut1_11[15] , 
        \nOut1_11[14] , \nOut1_11[13] , \nOut1_11[12] , \nOut1_11[11] , 
        \nOut1_11[10] , \nOut1_11[9] , \nOut1_11[8] , \nOut1_11[7] , 
        \nOut1_11[6] , \nOut1_11[5] , \nOut1_11[4] , \nOut1_11[3] , 
        \nOut1_11[2] , \nOut1_11[1] , \nOut1_11[0] }), .NORTH_EDGE({
        \nOut1_10[31] , \nOut1_10[30] , \nOut1_10[29] , \nOut1_10[28] , 
        \nOut1_10[27] , \nOut1_10[26] , \nOut1_10[25] , \nOut1_10[24] , 
        \nOut1_10[23] , \nOut1_10[22] , \nOut1_10[21] , \nOut1_10[20] , 
        \nOut1_10[19] , \nOut1_10[18] , \nOut1_10[17] , \nOut1_10[16] , 
        \nOut1_10[15] , \nOut1_10[14] , \nOut1_10[13] , \nOut1_10[12] , 
        \nOut1_10[11] , \nOut1_10[10] , \nOut1_10[9] , \nOut1_10[8] , 
        \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , \nOut1_10[4] , 
        \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , \nOut1_10[0] }), 
        .SOUTH_EDGE({\nOut1_12[31] , \nOut1_12[30] , \nOut1_12[29] , 
        \nOut1_12[28] , \nOut1_12[27] , \nOut1_12[26] , \nOut1_12[25] , 
        \nOut1_12[24] , \nOut1_12[23] , \nOut1_12[22] , \nOut1_12[21] , 
        \nOut1_12[20] , \nOut1_12[19] , \nOut1_12[18] , \nOut1_12[17] , 
        \nOut1_12[16] , \nOut1_12[15] , \nOut1_12[14] , \nOut1_12[13] , 
        \nOut1_12[12] , \nOut1_12[11] , \nOut1_12[10] , \nOut1_12[9] , 
        \nOut1_12[8] , \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , 
        \nOut1_12[4] , \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , 
        \nOut1_12[0] }), .EAST_EDGE(\nOut2_11[31] ), .WEST_EDGE(\nOut0_11[0] ), 
        .NW_EDGE(\nOut0_10[0] ), .SW_EDGE(\nOut0_12[0] ), .NE_EDGE(
        \nOut2_10[31] ), .SE_EDGE(\nOut2_12[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_15 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut16[31] , \nScanOut16[30] , \nScanOut16[29] , 
        \nScanOut16[28] , \nScanOut16[27] , \nScanOut16[26] , \nScanOut16[25] , 
        \nScanOut16[24] , \nScanOut16[23] , \nScanOut16[22] , \nScanOut16[21] , 
        \nScanOut16[20] , \nScanOut16[19] , \nScanOut16[18] , \nScanOut16[17] , 
        \nScanOut16[16] , \nScanOut16[15] , \nScanOut16[14] , \nScanOut16[13] , 
        \nScanOut16[12] , \nScanOut16[11] , \nScanOut16[10] , \nScanOut16[9] , 
        \nScanOut16[8] , \nScanOut16[7] , \nScanOut16[6] , \nScanOut16[5] , 
        \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , \nScanOut16[1] , 
        \nScanOut16[0] }), .ScanOut({\nScanOut15[31] , \nScanOut15[30] , 
        \nScanOut15[29] , \nScanOut15[28] , \nScanOut15[27] , \nScanOut15[26] , 
        \nScanOut15[25] , \nScanOut15[24] , \nScanOut15[23] , \nScanOut15[22] , 
        \nScanOut15[21] , \nScanOut15[20] , \nScanOut15[19] , \nScanOut15[18] , 
        \nScanOut15[17] , \nScanOut15[16] , \nScanOut15[15] , \nScanOut15[14] , 
        \nScanOut15[13] , \nScanOut15[12] , \nScanOut15[11] , \nScanOut15[10] , 
        \nScanOut15[9] , \nScanOut15[8] , \nScanOut15[7] , \nScanOut15[6] , 
        \nScanOut15[5] , \nScanOut15[4] , \nScanOut15[3] , \nScanOut15[2] , 
        \nScanOut15[1] , \nScanOut15[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_15[31] , 
        \nOut0_15[30] , \nOut0_15[29] , \nOut0_15[28] , \nOut0_15[27] , 
        \nOut0_15[26] , \nOut0_15[25] , \nOut0_15[24] , \nOut0_15[23] , 
        \nOut0_15[22] , \nOut0_15[21] , \nOut0_15[20] , \nOut0_15[19] , 
        \nOut0_15[18] , \nOut0_15[17] , \nOut0_15[16] , \nOut0_15[15] , 
        \nOut0_15[14] , \nOut0_15[13] , \nOut0_15[12] , \nOut0_15[11] , 
        \nOut0_15[10] , \nOut0_15[9] , \nOut0_15[8] , \nOut0_15[7] , 
        \nOut0_15[6] , \nOut0_15[5] , \nOut0_15[4] , \nOut0_15[3] , 
        \nOut0_15[2] , \nOut0_15[1] , \nOut0_15[0] }), .NORTH_EDGE({
        \nOut0_14[31] , \nOut0_14[30] , \nOut0_14[29] , \nOut0_14[28] , 
        \nOut0_14[27] , \nOut0_14[26] , \nOut0_14[25] , \nOut0_14[24] , 
        \nOut0_14[23] , \nOut0_14[22] , \nOut0_14[21] , \nOut0_14[20] , 
        \nOut0_14[19] , \nOut0_14[18] , \nOut0_14[17] , \nOut0_14[16] , 
        \nOut0_14[15] , \nOut0_14[14] , \nOut0_14[13] , \nOut0_14[12] , 
        \nOut0_14[11] , \nOut0_14[10] , \nOut0_14[9] , \nOut0_14[8] , 
        \nOut0_14[7] , \nOut0_14[6] , \nOut0_14[5] , \nOut0_14[4] , 
        \nOut0_14[3] , \nOut0_14[2] , \nOut0_14[1] , \nOut0_14[0] }), 
        .SOUTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .EAST_EDGE(\nOut1_15[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), 
        .SW_EDGE(1'b0), .NE_EDGE(\nOut1_14[31] ), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_29 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut30[31] , \nScanOut30[30] , \nScanOut30[29] , 
        \nScanOut30[28] , \nScanOut30[27] , \nScanOut30[26] , \nScanOut30[25] , 
        \nScanOut30[24] , \nScanOut30[23] , \nScanOut30[22] , \nScanOut30[21] , 
        \nScanOut30[20] , \nScanOut30[19] , \nScanOut30[18] , \nScanOut30[17] , 
        \nScanOut30[16] , \nScanOut30[15] , \nScanOut30[14] , \nScanOut30[13] , 
        \nScanOut30[12] , \nScanOut30[11] , \nScanOut30[10] , \nScanOut30[9] , 
        \nScanOut30[8] , \nScanOut30[7] , \nScanOut30[6] , \nScanOut30[5] , 
        \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , \nScanOut30[1] , 
        \nScanOut30[0] }), .ScanOut({\nScanOut29[31] , \nScanOut29[30] , 
        \nScanOut29[29] , \nScanOut29[28] , \nScanOut29[27] , \nScanOut29[26] , 
        \nScanOut29[25] , \nScanOut29[24] , \nScanOut29[23] , \nScanOut29[22] , 
        \nScanOut29[21] , \nScanOut29[20] , \nScanOut29[19] , \nScanOut29[18] , 
        \nScanOut29[17] , \nScanOut29[16] , \nScanOut29[15] , \nScanOut29[14] , 
        \nScanOut29[13] , \nScanOut29[12] , \nScanOut29[11] , \nScanOut29[10] , 
        \nScanOut29[9] , \nScanOut29[8] , \nScanOut29[7] , \nScanOut29[6] , 
        \nScanOut29[5] , \nScanOut29[4] , \nScanOut29[3] , \nScanOut29[2] , 
        \nScanOut29[1] , \nScanOut29[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_13[31] , 
        \nOut1_13[30] , \nOut1_13[29] , \nOut1_13[28] , \nOut1_13[27] , 
        \nOut1_13[26] , \nOut1_13[25] , \nOut1_13[24] , \nOut1_13[23] , 
        \nOut1_13[22] , \nOut1_13[21] , \nOut1_13[20] , \nOut1_13[19] , 
        \nOut1_13[18] , \nOut1_13[17] , \nOut1_13[16] , \nOut1_13[15] , 
        \nOut1_13[14] , \nOut1_13[13] , \nOut1_13[12] , \nOut1_13[11] , 
        \nOut1_13[10] , \nOut1_13[9] , \nOut1_13[8] , \nOut1_13[7] , 
        \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , \nOut1_13[3] , 
        \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), .NORTH_EDGE({
        \nOut1_12[31] , \nOut1_12[30] , \nOut1_12[29] , \nOut1_12[28] , 
        \nOut1_12[27] , \nOut1_12[26] , \nOut1_12[25] , \nOut1_12[24] , 
        \nOut1_12[23] , \nOut1_12[22] , \nOut1_12[21] , \nOut1_12[20] , 
        \nOut1_12[19] , \nOut1_12[18] , \nOut1_12[17] , \nOut1_12[16] , 
        \nOut1_12[15] , \nOut1_12[14] , \nOut1_12[13] , \nOut1_12[12] , 
        \nOut1_12[11] , \nOut1_12[10] , \nOut1_12[9] , \nOut1_12[8] , 
        \nOut1_12[7] , \nOut1_12[6] , \nOut1_12[5] , \nOut1_12[4] , 
        \nOut1_12[3] , \nOut1_12[2] , \nOut1_12[1] , \nOut1_12[0] }), 
        .SOUTH_EDGE({\nOut1_14[31] , \nOut1_14[30] , \nOut1_14[29] , 
        \nOut1_14[28] , \nOut1_14[27] , \nOut1_14[26] , \nOut1_14[25] , 
        \nOut1_14[24] , \nOut1_14[23] , \nOut1_14[22] , \nOut1_14[21] , 
        \nOut1_14[20] , \nOut1_14[19] , \nOut1_14[18] , \nOut1_14[17] , 
        \nOut1_14[16] , \nOut1_14[15] , \nOut1_14[14] , \nOut1_14[13] , 
        \nOut1_14[12] , \nOut1_14[11] , \nOut1_14[10] , \nOut1_14[9] , 
        \nOut1_14[8] , \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , 
        \nOut1_14[4] , \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , 
        \nOut1_14[0] }), .EAST_EDGE(\nOut2_13[31] ), .WEST_EDGE(\nOut0_13[0] ), 
        .NW_EDGE(\nOut0_12[0] ), .SW_EDGE(\nOut0_14[0] ), .NE_EDGE(
        \nOut2_12[31] ), .SE_EDGE(\nOut2_14[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_32 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut33[31] , \nScanOut33[30] , \nScanOut33[29] , 
        \nScanOut33[28] , \nScanOut33[27] , \nScanOut33[26] , \nScanOut33[25] , 
        \nScanOut33[24] , \nScanOut33[23] , \nScanOut33[22] , \nScanOut33[21] , 
        \nScanOut33[20] , \nScanOut33[19] , \nScanOut33[18] , \nScanOut33[17] , 
        \nScanOut33[16] , \nScanOut33[15] , \nScanOut33[14] , \nScanOut33[13] , 
        \nScanOut33[12] , \nScanOut33[11] , \nScanOut33[10] , \nScanOut33[9] , 
        \nScanOut33[8] , \nScanOut33[7] , \nScanOut33[6] , \nScanOut33[5] , 
        \nScanOut33[4] , \nScanOut33[3] , \nScanOut33[2] , \nScanOut33[1] , 
        \nScanOut33[0] }), .ScanOut({\nScanOut32[31] , \nScanOut32[30] , 
        \nScanOut32[29] , \nScanOut32[28] , \nScanOut32[27] , \nScanOut32[26] , 
        \nScanOut32[25] , \nScanOut32[24] , \nScanOut32[23] , \nScanOut32[22] , 
        \nScanOut32[21] , \nScanOut32[20] , \nScanOut32[19] , \nScanOut32[18] , 
        \nScanOut32[17] , \nScanOut32[16] , \nScanOut32[15] , \nScanOut32[14] , 
        \nScanOut32[13] , \nScanOut32[12] , \nScanOut32[11] , \nScanOut32[10] , 
        \nScanOut32[9] , \nScanOut32[8] , \nScanOut32[7] , \nScanOut32[6] , 
        \nScanOut32[5] , \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , 
        \nScanOut32[1] , \nScanOut32[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_0[31] , 
        \nOut2_0[30] , \nOut2_0[29] , \nOut2_0[28] , \nOut2_0[27] , 
        \nOut2_0[26] , \nOut2_0[25] , \nOut2_0[24] , \nOut2_0[23] , 
        \nOut2_0[22] , \nOut2_0[21] , \nOut2_0[20] , \nOut2_0[19] , 
        \nOut2_0[18] , \nOut2_0[17] , \nOut2_0[16] , \nOut2_0[15] , 
        \nOut2_0[14] , \nOut2_0[13] , \nOut2_0[12] , \nOut2_0[11] , 
        \nOut2_0[10] , \nOut2_0[9] , \nOut2_0[8] , \nOut2_0[7] , \nOut2_0[6] , 
        \nOut2_0[5] , \nOut2_0[4] , \nOut2_0[3] , \nOut2_0[2] , \nOut2_0[1] , 
        \nOut2_0[0] }), .NORTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SOUTH_EDGE({\nOut2_1[31] , \nOut2_1[30] , \nOut2_1[29] , 
        \nOut2_1[28] , \nOut2_1[27] , \nOut2_1[26] , \nOut2_1[25] , 
        \nOut2_1[24] , \nOut2_1[23] , \nOut2_1[22] , \nOut2_1[21] , 
        \nOut2_1[20] , \nOut2_1[19] , \nOut2_1[18] , \nOut2_1[17] , 
        \nOut2_1[16] , \nOut2_1[15] , \nOut2_1[14] , \nOut2_1[13] , 
        \nOut2_1[12] , \nOut2_1[11] , \nOut2_1[10] , \nOut2_1[9] , 
        \nOut2_1[8] , \nOut2_1[7] , \nOut2_1[6] , \nOut2_1[5] , \nOut2_1[4] , 
        \nOut2_1[3] , \nOut2_1[2] , \nOut2_1[1] , \nOut2_1[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_0[0] ), .NW_EDGE(1'b0), .SW_EDGE(\nOut1_1[0] 
        ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_47 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut48[31] , \nScanOut48[30] , \nScanOut48[29] , 
        \nScanOut48[28] , \nScanOut48[27] , \nScanOut48[26] , \nScanOut48[25] , 
        \nScanOut48[24] , \nScanOut48[23] , \nScanOut48[22] , \nScanOut48[21] , 
        \nScanOut48[20] , \nScanOut48[19] , \nScanOut48[18] , \nScanOut48[17] , 
        \nScanOut48[16] , \nScanOut48[15] , \nScanOut48[14] , \nScanOut48[13] , 
        \nScanOut48[12] , \nScanOut48[11] , \nScanOut48[10] , \nScanOut48[9] , 
        \nScanOut48[8] , \nScanOut48[7] , \nScanOut48[6] , \nScanOut48[5] , 
        \nScanOut48[4] , \nScanOut48[3] , \nScanOut48[2] , \nScanOut48[1] , 
        \nScanOut48[0] }), .ScanOut({\nScanOut47[31] , \nScanOut47[30] , 
        \nScanOut47[29] , \nScanOut47[28] , \nScanOut47[27] , \nScanOut47[26] , 
        \nScanOut47[25] , \nScanOut47[24] , \nScanOut47[23] , \nScanOut47[22] , 
        \nScanOut47[21] , \nScanOut47[20] , \nScanOut47[19] , \nScanOut47[18] , 
        \nScanOut47[17] , \nScanOut47[16] , \nScanOut47[15] , \nScanOut47[14] , 
        \nScanOut47[13] , \nScanOut47[12] , \nScanOut47[11] , \nScanOut47[10] , 
        \nScanOut47[9] , \nScanOut47[8] , \nScanOut47[7] , \nScanOut47[6] , 
        \nScanOut47[5] , \nScanOut47[4] , \nScanOut47[3] , \nScanOut47[2] , 
        \nScanOut47[1] , \nScanOut47[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_15[31] , 
        \nOut2_15[30] , \nOut2_15[29] , \nOut2_15[28] , \nOut2_15[27] , 
        \nOut2_15[26] , \nOut2_15[25] , \nOut2_15[24] , \nOut2_15[23] , 
        \nOut2_15[22] , \nOut2_15[21] , \nOut2_15[20] , \nOut2_15[19] , 
        \nOut2_15[18] , \nOut2_15[17] , \nOut2_15[16] , \nOut2_15[15] , 
        \nOut2_15[14] , \nOut2_15[13] , \nOut2_15[12] , \nOut2_15[11] , 
        \nOut2_15[10] , \nOut2_15[9] , \nOut2_15[8] , \nOut2_15[7] , 
        \nOut2_15[6] , \nOut2_15[5] , \nOut2_15[4] , \nOut2_15[3] , 
        \nOut2_15[2] , \nOut2_15[1] , \nOut2_15[0] }), .NORTH_EDGE({
        \nOut2_14[31] , \nOut2_14[30] , \nOut2_14[29] , \nOut2_14[28] , 
        \nOut2_14[27] , \nOut2_14[26] , \nOut2_14[25] , \nOut2_14[24] , 
        \nOut2_14[23] , \nOut2_14[22] , \nOut2_14[21] , \nOut2_14[20] , 
        \nOut2_14[19] , \nOut2_14[18] , \nOut2_14[17] , \nOut2_14[16] , 
        \nOut2_14[15] , \nOut2_14[14] , \nOut2_14[13] , \nOut2_14[12] , 
        \nOut2_14[11] , \nOut2_14[10] , \nOut2_14[9] , \nOut2_14[8] , 
        \nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , \nOut2_14[4] , 
        \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , \nOut2_14[0] }), 
        .SOUTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_15[0] ), .NW_EDGE(\nOut1_14[0] ), 
        .SW_EDGE(1'b0), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_39 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut40[31] , \nScanOut40[30] , \nScanOut40[29] , 
        \nScanOut40[28] , \nScanOut40[27] , \nScanOut40[26] , \nScanOut40[25] , 
        \nScanOut40[24] , \nScanOut40[23] , \nScanOut40[22] , \nScanOut40[21] , 
        \nScanOut40[20] , \nScanOut40[19] , \nScanOut40[18] , \nScanOut40[17] , 
        \nScanOut40[16] , \nScanOut40[15] , \nScanOut40[14] , \nScanOut40[13] , 
        \nScanOut40[12] , \nScanOut40[11] , \nScanOut40[10] , \nScanOut40[9] , 
        \nScanOut40[8] , \nScanOut40[7] , \nScanOut40[6] , \nScanOut40[5] , 
        \nScanOut40[4] , \nScanOut40[3] , \nScanOut40[2] , \nScanOut40[1] , 
        \nScanOut40[0] }), .ScanOut({\nScanOut39[31] , \nScanOut39[30] , 
        \nScanOut39[29] , \nScanOut39[28] , \nScanOut39[27] , \nScanOut39[26] , 
        \nScanOut39[25] , \nScanOut39[24] , \nScanOut39[23] , \nScanOut39[22] , 
        \nScanOut39[21] , \nScanOut39[20] , \nScanOut39[19] , \nScanOut39[18] , 
        \nScanOut39[17] , \nScanOut39[16] , \nScanOut39[15] , \nScanOut39[14] , 
        \nScanOut39[13] , \nScanOut39[12] , \nScanOut39[11] , \nScanOut39[10] , 
        \nScanOut39[9] , \nScanOut39[8] , \nScanOut39[7] , \nScanOut39[6] , 
        \nScanOut39[5] , \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , 
        \nScanOut39[1] , \nScanOut39[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_7[31] , 
        \nOut2_7[30] , \nOut2_7[29] , \nOut2_7[28] , \nOut2_7[27] , 
        \nOut2_7[26] , \nOut2_7[25] , \nOut2_7[24] , \nOut2_7[23] , 
        \nOut2_7[22] , \nOut2_7[21] , \nOut2_7[20] , \nOut2_7[19] , 
        \nOut2_7[18] , \nOut2_7[17] , \nOut2_7[16] , \nOut2_7[15] , 
        \nOut2_7[14] , \nOut2_7[13] , \nOut2_7[12] , \nOut2_7[11] , 
        \nOut2_7[10] , \nOut2_7[9] , \nOut2_7[8] , \nOut2_7[7] , \nOut2_7[6] , 
        \nOut2_7[5] , \nOut2_7[4] , \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , 
        \nOut2_7[0] }), .NORTH_EDGE({\nOut2_6[31] , \nOut2_6[30] , 
        \nOut2_6[29] , \nOut2_6[28] , \nOut2_6[27] , \nOut2_6[26] , 
        \nOut2_6[25] , \nOut2_6[24] , \nOut2_6[23] , \nOut2_6[22] , 
        \nOut2_6[21] , \nOut2_6[20] , \nOut2_6[19] , \nOut2_6[18] , 
        \nOut2_6[17] , \nOut2_6[16] , \nOut2_6[15] , \nOut2_6[14] , 
        \nOut2_6[13] , \nOut2_6[12] , \nOut2_6[11] , \nOut2_6[10] , 
        \nOut2_6[9] , \nOut2_6[8] , \nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , 
        \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), 
        .SOUTH_EDGE({\nOut2_8[31] , \nOut2_8[30] , \nOut2_8[29] , 
        \nOut2_8[28] , \nOut2_8[27] , \nOut2_8[26] , \nOut2_8[25] , 
        \nOut2_8[24] , \nOut2_8[23] , \nOut2_8[22] , \nOut2_8[21] , 
        \nOut2_8[20] , \nOut2_8[19] , \nOut2_8[18] , \nOut2_8[17] , 
        \nOut2_8[16] , \nOut2_8[15] , \nOut2_8[14] , \nOut2_8[13] , 
        \nOut2_8[12] , \nOut2_8[11] , \nOut2_8[10] , \nOut2_8[9] , 
        \nOut2_8[8] , \nOut2_8[7] , \nOut2_8[6] , \nOut2_8[5] , \nOut2_8[4] , 
        \nOut2_8[3] , \nOut2_8[2] , \nOut2_8[1] , \nOut2_8[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_7[0] ), .NW_EDGE(\nOut1_6[0] ), .SW_EDGE(
        \nOut1_8[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_1 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut2[31] , \nScanOut2[30] , \nScanOut2[29] , 
        \nScanOut2[28] , \nScanOut2[27] , \nScanOut2[26] , \nScanOut2[25] , 
        \nScanOut2[24] , \nScanOut2[23] , \nScanOut2[22] , \nScanOut2[21] , 
        \nScanOut2[20] , \nScanOut2[19] , \nScanOut2[18] , \nScanOut2[17] , 
        \nScanOut2[16] , \nScanOut2[15] , \nScanOut2[14] , \nScanOut2[13] , 
        \nScanOut2[12] , \nScanOut2[11] , \nScanOut2[10] , \nScanOut2[9] , 
        \nScanOut2[8] , \nScanOut2[7] , \nScanOut2[6] , \nScanOut2[5] , 
        \nScanOut2[4] , \nScanOut2[3] , \nScanOut2[2] , \nScanOut2[1] , 
        \nScanOut2[0] }), .ScanOut({\nScanOut1[31] , \nScanOut1[30] , 
        \nScanOut1[29] , \nScanOut1[28] , \nScanOut1[27] , \nScanOut1[26] , 
        \nScanOut1[25] , \nScanOut1[24] , \nScanOut1[23] , \nScanOut1[22] , 
        \nScanOut1[21] , \nScanOut1[20] , \nScanOut1[19] , \nScanOut1[18] , 
        \nScanOut1[17] , \nScanOut1[16] , \nScanOut1[15] , \nScanOut1[14] , 
        \nScanOut1[13] , \nScanOut1[12] , \nScanOut1[11] , \nScanOut1[10] , 
        \nScanOut1[9] , \nScanOut1[8] , \nScanOut1[7] , \nScanOut1[6] , 
        \nScanOut1[5] , \nScanOut1[4] , \nScanOut1[3] , \nScanOut1[2] , 
        \nScanOut1[1] , \nScanOut1[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_1[31] , 
        \nOut0_1[30] , \nOut0_1[29] , \nOut0_1[28] , \nOut0_1[27] , 
        \nOut0_1[26] , \nOut0_1[25] , \nOut0_1[24] , \nOut0_1[23] , 
        \nOut0_1[22] , \nOut0_1[21] , \nOut0_1[20] , \nOut0_1[19] , 
        \nOut0_1[18] , \nOut0_1[17] , \nOut0_1[16] , \nOut0_1[15] , 
        \nOut0_1[14] , \nOut0_1[13] , \nOut0_1[12] , \nOut0_1[11] , 
        \nOut0_1[10] , \nOut0_1[9] , \nOut0_1[8] , \nOut0_1[7] , \nOut0_1[6] , 
        \nOut0_1[5] , \nOut0_1[4] , \nOut0_1[3] , \nOut0_1[2] , \nOut0_1[1] , 
        \nOut0_1[0] }), .NORTH_EDGE({\nOut0_0[31] , \nOut0_0[30] , 
        \nOut0_0[29] , \nOut0_0[28] , \nOut0_0[27] , \nOut0_0[26] , 
        \nOut0_0[25] , \nOut0_0[24] , \nOut0_0[23] , \nOut0_0[22] , 
        \nOut0_0[21] , \nOut0_0[20] , \nOut0_0[19] , \nOut0_0[18] , 
        \nOut0_0[17] , \nOut0_0[16] , \nOut0_0[15] , \nOut0_0[14] , 
        \nOut0_0[13] , \nOut0_0[12] , \nOut0_0[11] , \nOut0_0[10] , 
        \nOut0_0[9] , \nOut0_0[8] , \nOut0_0[7] , \nOut0_0[6] , \nOut0_0[5] , 
        \nOut0_0[4] , \nOut0_0[3] , \nOut0_0[2] , \nOut0_0[1] , \nOut0_0[0] }), 
        .SOUTH_EDGE({\nOut0_2[31] , \nOut0_2[30] , \nOut0_2[29] , 
        \nOut0_2[28] , \nOut0_2[27] , \nOut0_2[26] , \nOut0_2[25] , 
        \nOut0_2[24] , \nOut0_2[23] , \nOut0_2[22] , \nOut0_2[21] , 
        \nOut0_2[20] , \nOut0_2[19] , \nOut0_2[18] , \nOut0_2[17] , 
        \nOut0_2[16] , \nOut0_2[15] , \nOut0_2[14] , \nOut0_2[13] , 
        \nOut0_2[12] , \nOut0_2[11] , \nOut0_2[10] , \nOut0_2[9] , 
        \nOut0_2[8] , \nOut0_2[7] , \nOut0_2[6] , \nOut0_2[5] , \nOut0_2[4] , 
        \nOut0_2[3] , \nOut0_2[2] , \nOut0_2[1] , \nOut0_2[0] }), .EAST_EDGE(
        \nOut1_1[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_0[31] ), .SE_EDGE(\nOut1_2[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_6 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut7[31] , \nScanOut7[30] , \nScanOut7[29] , 
        \nScanOut7[28] , \nScanOut7[27] , \nScanOut7[26] , \nScanOut7[25] , 
        \nScanOut7[24] , \nScanOut7[23] , \nScanOut7[22] , \nScanOut7[21] , 
        \nScanOut7[20] , \nScanOut7[19] , \nScanOut7[18] , \nScanOut7[17] , 
        \nScanOut7[16] , \nScanOut7[15] , \nScanOut7[14] , \nScanOut7[13] , 
        \nScanOut7[12] , \nScanOut7[11] , \nScanOut7[10] , \nScanOut7[9] , 
        \nScanOut7[8] , \nScanOut7[7] , \nScanOut7[6] , \nScanOut7[5] , 
        \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , \nScanOut7[1] , 
        \nScanOut7[0] }), .ScanOut({\nScanOut6[31] , \nScanOut6[30] , 
        \nScanOut6[29] , \nScanOut6[28] , \nScanOut6[27] , \nScanOut6[26] , 
        \nScanOut6[25] , \nScanOut6[24] , \nScanOut6[23] , \nScanOut6[22] , 
        \nScanOut6[21] , \nScanOut6[20] , \nScanOut6[19] , \nScanOut6[18] , 
        \nScanOut6[17] , \nScanOut6[16] , \nScanOut6[15] , \nScanOut6[14] , 
        \nScanOut6[13] , \nScanOut6[12] , \nScanOut6[11] , \nScanOut6[10] , 
        \nScanOut6[9] , \nScanOut6[8] , \nScanOut6[7] , \nScanOut6[6] , 
        \nScanOut6[5] , \nScanOut6[4] , \nScanOut6[3] , \nScanOut6[2] , 
        \nScanOut6[1] , \nScanOut6[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_6[31] , 
        \nOut0_6[30] , \nOut0_6[29] , \nOut0_6[28] , \nOut0_6[27] , 
        \nOut0_6[26] , \nOut0_6[25] , \nOut0_6[24] , \nOut0_6[23] , 
        \nOut0_6[22] , \nOut0_6[21] , \nOut0_6[20] , \nOut0_6[19] , 
        \nOut0_6[18] , \nOut0_6[17] , \nOut0_6[16] , \nOut0_6[15] , 
        \nOut0_6[14] , \nOut0_6[13] , \nOut0_6[12] , \nOut0_6[11] , 
        \nOut0_6[10] , \nOut0_6[9] , \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , 
        \nOut0_6[5] , \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , 
        \nOut0_6[0] }), .NORTH_EDGE({\nOut0_5[31] , \nOut0_5[30] , 
        \nOut0_5[29] , \nOut0_5[28] , \nOut0_5[27] , \nOut0_5[26] , 
        \nOut0_5[25] , \nOut0_5[24] , \nOut0_5[23] , \nOut0_5[22] , 
        \nOut0_5[21] , \nOut0_5[20] , \nOut0_5[19] , \nOut0_5[18] , 
        \nOut0_5[17] , \nOut0_5[16] , \nOut0_5[15] , \nOut0_5[14] , 
        \nOut0_5[13] , \nOut0_5[12] , \nOut0_5[11] , \nOut0_5[10] , 
        \nOut0_5[9] , \nOut0_5[8] , \nOut0_5[7] , \nOut0_5[6] , \nOut0_5[5] , 
        \nOut0_5[4] , \nOut0_5[3] , \nOut0_5[2] , \nOut0_5[1] , \nOut0_5[0] }), 
        .SOUTH_EDGE({\nOut0_7[31] , \nOut0_7[30] , \nOut0_7[29] , 
        \nOut0_7[28] , \nOut0_7[27] , \nOut0_7[26] , \nOut0_7[25] , 
        \nOut0_7[24] , \nOut0_7[23] , \nOut0_7[22] , \nOut0_7[21] , 
        \nOut0_7[20] , \nOut0_7[19] , \nOut0_7[18] , \nOut0_7[17] , 
        \nOut0_7[16] , \nOut0_7[15] , \nOut0_7[14] , \nOut0_7[13] , 
        \nOut0_7[12] , \nOut0_7[11] , \nOut0_7[10] , \nOut0_7[9] , 
        \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , \nOut0_7[4] , 
        \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), .EAST_EDGE(
        \nOut1_6[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_5[31] ), .SE_EDGE(\nOut1_7[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_7 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut8[31] , \nScanOut8[30] , \nScanOut8[29] , 
        \nScanOut8[28] , \nScanOut8[27] , \nScanOut8[26] , \nScanOut8[25] , 
        \nScanOut8[24] , \nScanOut8[23] , \nScanOut8[22] , \nScanOut8[21] , 
        \nScanOut8[20] , \nScanOut8[19] , \nScanOut8[18] , \nScanOut8[17] , 
        \nScanOut8[16] , \nScanOut8[15] , \nScanOut8[14] , \nScanOut8[13] , 
        \nScanOut8[12] , \nScanOut8[11] , \nScanOut8[10] , \nScanOut8[9] , 
        \nScanOut8[8] , \nScanOut8[7] , \nScanOut8[6] , \nScanOut8[5] , 
        \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , \nScanOut8[1] , 
        \nScanOut8[0] }), .ScanOut({\nScanOut7[31] , \nScanOut7[30] , 
        \nScanOut7[29] , \nScanOut7[28] , \nScanOut7[27] , \nScanOut7[26] , 
        \nScanOut7[25] , \nScanOut7[24] , \nScanOut7[23] , \nScanOut7[22] , 
        \nScanOut7[21] , \nScanOut7[20] , \nScanOut7[19] , \nScanOut7[18] , 
        \nScanOut7[17] , \nScanOut7[16] , \nScanOut7[15] , \nScanOut7[14] , 
        \nScanOut7[13] , \nScanOut7[12] , \nScanOut7[11] , \nScanOut7[10] , 
        \nScanOut7[9] , \nScanOut7[8] , \nScanOut7[7] , \nScanOut7[6] , 
        \nScanOut7[5] , \nScanOut7[4] , \nScanOut7[3] , \nScanOut7[2] , 
        \nScanOut7[1] , \nScanOut7[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_7[31] , 
        \nOut0_7[30] , \nOut0_7[29] , \nOut0_7[28] , \nOut0_7[27] , 
        \nOut0_7[26] , \nOut0_7[25] , \nOut0_7[24] , \nOut0_7[23] , 
        \nOut0_7[22] , \nOut0_7[21] , \nOut0_7[20] , \nOut0_7[19] , 
        \nOut0_7[18] , \nOut0_7[17] , \nOut0_7[16] , \nOut0_7[15] , 
        \nOut0_7[14] , \nOut0_7[13] , \nOut0_7[12] , \nOut0_7[11] , 
        \nOut0_7[10] , \nOut0_7[9] , \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , 
        \nOut0_7[5] , \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , 
        \nOut0_7[0] }), .NORTH_EDGE({\nOut0_6[31] , \nOut0_6[30] , 
        \nOut0_6[29] , \nOut0_6[28] , \nOut0_6[27] , \nOut0_6[26] , 
        \nOut0_6[25] , \nOut0_6[24] , \nOut0_6[23] , \nOut0_6[22] , 
        \nOut0_6[21] , \nOut0_6[20] , \nOut0_6[19] , \nOut0_6[18] , 
        \nOut0_6[17] , \nOut0_6[16] , \nOut0_6[15] , \nOut0_6[14] , 
        \nOut0_6[13] , \nOut0_6[12] , \nOut0_6[11] , \nOut0_6[10] , 
        \nOut0_6[9] , \nOut0_6[8] , \nOut0_6[7] , \nOut0_6[6] , \nOut0_6[5] , 
        \nOut0_6[4] , \nOut0_6[3] , \nOut0_6[2] , \nOut0_6[1] , \nOut0_6[0] }), 
        .SOUTH_EDGE({\nOut0_8[31] , \nOut0_8[30] , \nOut0_8[29] , 
        \nOut0_8[28] , \nOut0_8[27] , \nOut0_8[26] , \nOut0_8[25] , 
        \nOut0_8[24] , \nOut0_8[23] , \nOut0_8[22] , \nOut0_8[21] , 
        \nOut0_8[20] , \nOut0_8[19] , \nOut0_8[18] , \nOut0_8[17] , 
        \nOut0_8[16] , \nOut0_8[15] , \nOut0_8[14] , \nOut0_8[13] , 
        \nOut0_8[12] , \nOut0_8[11] , \nOut0_8[10] , \nOut0_8[9] , 
        \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , \nOut0_8[4] , 
        \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), .EAST_EDGE(
        \nOut1_7[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_6[31] ), .SE_EDGE(\nOut1_8[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_9 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut10[31] , \nScanOut10[30] , \nScanOut10[29] , 
        \nScanOut10[28] , \nScanOut10[27] , \nScanOut10[26] , \nScanOut10[25] , 
        \nScanOut10[24] , \nScanOut10[23] , \nScanOut10[22] , \nScanOut10[21] , 
        \nScanOut10[20] , \nScanOut10[19] , \nScanOut10[18] , \nScanOut10[17] , 
        \nScanOut10[16] , \nScanOut10[15] , \nScanOut10[14] , \nScanOut10[13] , 
        \nScanOut10[12] , \nScanOut10[11] , \nScanOut10[10] , \nScanOut10[9] , 
        \nScanOut10[8] , \nScanOut10[7] , \nScanOut10[6] , \nScanOut10[5] , 
        \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , \nScanOut10[1] , 
        \nScanOut10[0] }), .ScanOut({\nScanOut9[31] , \nScanOut9[30] , 
        \nScanOut9[29] , \nScanOut9[28] , \nScanOut9[27] , \nScanOut9[26] , 
        \nScanOut9[25] , \nScanOut9[24] , \nScanOut9[23] , \nScanOut9[22] , 
        \nScanOut9[21] , \nScanOut9[20] , \nScanOut9[19] , \nScanOut9[18] , 
        \nScanOut9[17] , \nScanOut9[16] , \nScanOut9[15] , \nScanOut9[14] , 
        \nScanOut9[13] , \nScanOut9[12] , \nScanOut9[11] , \nScanOut9[10] , 
        \nScanOut9[9] , \nScanOut9[8] , \nScanOut9[7] , \nScanOut9[6] , 
        \nScanOut9[5] , \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , 
        \nScanOut9[1] , \nScanOut9[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_9[31] , 
        \nOut0_9[30] , \nOut0_9[29] , \nOut0_9[28] , \nOut0_9[27] , 
        \nOut0_9[26] , \nOut0_9[25] , \nOut0_9[24] , \nOut0_9[23] , 
        \nOut0_9[22] , \nOut0_9[21] , \nOut0_9[20] , \nOut0_9[19] , 
        \nOut0_9[18] , \nOut0_9[17] , \nOut0_9[16] , \nOut0_9[15] , 
        \nOut0_9[14] , \nOut0_9[13] , \nOut0_9[12] , \nOut0_9[11] , 
        \nOut0_9[10] , \nOut0_9[9] , \nOut0_9[8] , \nOut0_9[7] , \nOut0_9[6] , 
        \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , 
        \nOut0_9[0] }), .NORTH_EDGE({\nOut0_8[31] , \nOut0_8[30] , 
        \nOut0_8[29] , \nOut0_8[28] , \nOut0_8[27] , \nOut0_8[26] , 
        \nOut0_8[25] , \nOut0_8[24] , \nOut0_8[23] , \nOut0_8[22] , 
        \nOut0_8[21] , \nOut0_8[20] , \nOut0_8[19] , \nOut0_8[18] , 
        \nOut0_8[17] , \nOut0_8[16] , \nOut0_8[15] , \nOut0_8[14] , 
        \nOut0_8[13] , \nOut0_8[12] , \nOut0_8[11] , \nOut0_8[10] , 
        \nOut0_8[9] , \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , \nOut0_8[5] , 
        \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , \nOut0_8[0] }), 
        .SOUTH_EDGE({\nOut0_10[31] , \nOut0_10[30] , \nOut0_10[29] , 
        \nOut0_10[28] , \nOut0_10[27] , \nOut0_10[26] , \nOut0_10[25] , 
        \nOut0_10[24] , \nOut0_10[23] , \nOut0_10[22] , \nOut0_10[21] , 
        \nOut0_10[20] , \nOut0_10[19] , \nOut0_10[18] , \nOut0_10[17] , 
        \nOut0_10[16] , \nOut0_10[15] , \nOut0_10[14] , \nOut0_10[13] , 
        \nOut0_10[12] , \nOut0_10[11] , \nOut0_10[10] , \nOut0_10[9] , 
        \nOut0_10[8] , \nOut0_10[7] , \nOut0_10[6] , \nOut0_10[5] , 
        \nOut0_10[4] , \nOut0_10[3] , \nOut0_10[2] , \nOut0_10[1] , 
        \nOut0_10[0] }), .EAST_EDGE(\nOut1_9[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_8[31] ), .SE_EDGE(
        \nOut1_10[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_17 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut18[31] , \nScanOut18[30] , \nScanOut18[29] , 
        \nScanOut18[28] , \nScanOut18[27] , \nScanOut18[26] , \nScanOut18[25] , 
        \nScanOut18[24] , \nScanOut18[23] , \nScanOut18[22] , \nScanOut18[21] , 
        \nScanOut18[20] , \nScanOut18[19] , \nScanOut18[18] , \nScanOut18[17] , 
        \nScanOut18[16] , \nScanOut18[15] , \nScanOut18[14] , \nScanOut18[13] , 
        \nScanOut18[12] , \nScanOut18[11] , \nScanOut18[10] , \nScanOut18[9] , 
        \nScanOut18[8] , \nScanOut18[7] , \nScanOut18[6] , \nScanOut18[5] , 
        \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , \nScanOut18[1] , 
        \nScanOut18[0] }), .ScanOut({\nScanOut17[31] , \nScanOut17[30] , 
        \nScanOut17[29] , \nScanOut17[28] , \nScanOut17[27] , \nScanOut17[26] , 
        \nScanOut17[25] , \nScanOut17[24] , \nScanOut17[23] , \nScanOut17[22] , 
        \nScanOut17[21] , \nScanOut17[20] , \nScanOut17[19] , \nScanOut17[18] , 
        \nScanOut17[17] , \nScanOut17[16] , \nScanOut17[15] , \nScanOut17[14] , 
        \nScanOut17[13] , \nScanOut17[12] , \nScanOut17[11] , \nScanOut17[10] , 
        \nScanOut17[9] , \nScanOut17[8] , \nScanOut17[7] , \nScanOut17[6] , 
        \nScanOut17[5] , \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , 
        \nScanOut17[1] , \nScanOut17[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_1[31] , 
        \nOut1_1[30] , \nOut1_1[29] , \nOut1_1[28] , \nOut1_1[27] , 
        \nOut1_1[26] , \nOut1_1[25] , \nOut1_1[24] , \nOut1_1[23] , 
        \nOut1_1[22] , \nOut1_1[21] , \nOut1_1[20] , \nOut1_1[19] , 
        \nOut1_1[18] , \nOut1_1[17] , \nOut1_1[16] , \nOut1_1[15] , 
        \nOut1_1[14] , \nOut1_1[13] , \nOut1_1[12] , \nOut1_1[11] , 
        \nOut1_1[10] , \nOut1_1[9] , \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , 
        \nOut1_1[5] , \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , 
        \nOut1_1[0] }), .NORTH_EDGE({\nOut1_0[31] , \nOut1_0[30] , 
        \nOut1_0[29] , \nOut1_0[28] , \nOut1_0[27] , \nOut1_0[26] , 
        \nOut1_0[25] , \nOut1_0[24] , \nOut1_0[23] , \nOut1_0[22] , 
        \nOut1_0[21] , \nOut1_0[20] , \nOut1_0[19] , \nOut1_0[18] , 
        \nOut1_0[17] , \nOut1_0[16] , \nOut1_0[15] , \nOut1_0[14] , 
        \nOut1_0[13] , \nOut1_0[12] , \nOut1_0[11] , \nOut1_0[10] , 
        \nOut1_0[9] , \nOut1_0[8] , \nOut1_0[7] , \nOut1_0[6] , \nOut1_0[5] , 
        \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , \nOut1_0[0] }), 
        .SOUTH_EDGE({\nOut1_2[31] , \nOut1_2[30] , \nOut1_2[29] , 
        \nOut1_2[28] , \nOut1_2[27] , \nOut1_2[26] , \nOut1_2[25] , 
        \nOut1_2[24] , \nOut1_2[23] , \nOut1_2[22] , \nOut1_2[21] , 
        \nOut1_2[20] , \nOut1_2[19] , \nOut1_2[18] , \nOut1_2[17] , 
        \nOut1_2[16] , \nOut1_2[15] , \nOut1_2[14] , \nOut1_2[13] , 
        \nOut1_2[12] , \nOut1_2[11] , \nOut1_2[10] , \nOut1_2[9] , 
        \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , \nOut1_2[4] , 
        \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), .EAST_EDGE(
        \nOut2_1[31] ), .WEST_EDGE(\nOut0_1[0] ), .NW_EDGE(\nOut0_0[0] ), 
        .SW_EDGE(\nOut0_2[0] ), .NE_EDGE(\nOut2_0[31] ), .SE_EDGE(
        \nOut2_2[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_22 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut23[31] , \nScanOut23[30] , \nScanOut23[29] , 
        \nScanOut23[28] , \nScanOut23[27] , \nScanOut23[26] , \nScanOut23[25] , 
        \nScanOut23[24] , \nScanOut23[23] , \nScanOut23[22] , \nScanOut23[21] , 
        \nScanOut23[20] , \nScanOut23[19] , \nScanOut23[18] , \nScanOut23[17] , 
        \nScanOut23[16] , \nScanOut23[15] , \nScanOut23[14] , \nScanOut23[13] , 
        \nScanOut23[12] , \nScanOut23[11] , \nScanOut23[10] , \nScanOut23[9] , 
        \nScanOut23[8] , \nScanOut23[7] , \nScanOut23[6] , \nScanOut23[5] , 
        \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , \nScanOut23[1] , 
        \nScanOut23[0] }), .ScanOut({\nScanOut22[31] , \nScanOut22[30] , 
        \nScanOut22[29] , \nScanOut22[28] , \nScanOut22[27] , \nScanOut22[26] , 
        \nScanOut22[25] , \nScanOut22[24] , \nScanOut22[23] , \nScanOut22[22] , 
        \nScanOut22[21] , \nScanOut22[20] , \nScanOut22[19] , \nScanOut22[18] , 
        \nScanOut22[17] , \nScanOut22[16] , \nScanOut22[15] , \nScanOut22[14] , 
        \nScanOut22[13] , \nScanOut22[12] , \nScanOut22[11] , \nScanOut22[10] , 
        \nScanOut22[9] , \nScanOut22[8] , \nScanOut22[7] , \nScanOut22[6] , 
        \nScanOut22[5] , \nScanOut22[4] , \nScanOut22[3] , \nScanOut22[2] , 
        \nScanOut22[1] , \nScanOut22[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_6[31] , 
        \nOut1_6[30] , \nOut1_6[29] , \nOut1_6[28] , \nOut1_6[27] , 
        \nOut1_6[26] , \nOut1_6[25] , \nOut1_6[24] , \nOut1_6[23] , 
        \nOut1_6[22] , \nOut1_6[21] , \nOut1_6[20] , \nOut1_6[19] , 
        \nOut1_6[18] , \nOut1_6[17] , \nOut1_6[16] , \nOut1_6[15] , 
        \nOut1_6[14] , \nOut1_6[13] , \nOut1_6[12] , \nOut1_6[11] , 
        \nOut1_6[10] , \nOut1_6[9] , \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , 
        \nOut1_6[5] , \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , 
        \nOut1_6[0] }), .NORTH_EDGE({\nOut1_5[31] , \nOut1_5[30] , 
        \nOut1_5[29] , \nOut1_5[28] , \nOut1_5[27] , \nOut1_5[26] , 
        \nOut1_5[25] , \nOut1_5[24] , \nOut1_5[23] , \nOut1_5[22] , 
        \nOut1_5[21] , \nOut1_5[20] , \nOut1_5[19] , \nOut1_5[18] , 
        \nOut1_5[17] , \nOut1_5[16] , \nOut1_5[15] , \nOut1_5[14] , 
        \nOut1_5[13] , \nOut1_5[12] , \nOut1_5[11] , \nOut1_5[10] , 
        \nOut1_5[9] , \nOut1_5[8] , \nOut1_5[7] , \nOut1_5[6] , \nOut1_5[5] , 
        \nOut1_5[4] , \nOut1_5[3] , \nOut1_5[2] , \nOut1_5[1] , \nOut1_5[0] }), 
        .SOUTH_EDGE({\nOut1_7[31] , \nOut1_7[30] , \nOut1_7[29] , 
        \nOut1_7[28] , \nOut1_7[27] , \nOut1_7[26] , \nOut1_7[25] , 
        \nOut1_7[24] , \nOut1_7[23] , \nOut1_7[22] , \nOut1_7[21] , 
        \nOut1_7[20] , \nOut1_7[19] , \nOut1_7[18] , \nOut1_7[17] , 
        \nOut1_7[16] , \nOut1_7[15] , \nOut1_7[14] , \nOut1_7[13] , 
        \nOut1_7[12] , \nOut1_7[11] , \nOut1_7[10] , \nOut1_7[9] , 
        \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , \nOut1_7[4] , 
        \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), .EAST_EDGE(
        \nOut2_6[31] ), .WEST_EDGE(\nOut0_6[0] ), .NW_EDGE(\nOut0_5[0] ), 
        .SW_EDGE(\nOut0_7[0] ), .NE_EDGE(\nOut2_5[31] ), .SE_EDGE(
        \nOut2_7[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_30 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut31[31] , \nScanOut31[30] , \nScanOut31[29] , 
        \nScanOut31[28] , \nScanOut31[27] , \nScanOut31[26] , \nScanOut31[25] , 
        \nScanOut31[24] , \nScanOut31[23] , \nScanOut31[22] , \nScanOut31[21] , 
        \nScanOut31[20] , \nScanOut31[19] , \nScanOut31[18] , \nScanOut31[17] , 
        \nScanOut31[16] , \nScanOut31[15] , \nScanOut31[14] , \nScanOut31[13] , 
        \nScanOut31[12] , \nScanOut31[11] , \nScanOut31[10] , \nScanOut31[9] , 
        \nScanOut31[8] , \nScanOut31[7] , \nScanOut31[6] , \nScanOut31[5] , 
        \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , \nScanOut31[1] , 
        \nScanOut31[0] }), .ScanOut({\nScanOut30[31] , \nScanOut30[30] , 
        \nScanOut30[29] , \nScanOut30[28] , \nScanOut30[27] , \nScanOut30[26] , 
        \nScanOut30[25] , \nScanOut30[24] , \nScanOut30[23] , \nScanOut30[22] , 
        \nScanOut30[21] , \nScanOut30[20] , \nScanOut30[19] , \nScanOut30[18] , 
        \nScanOut30[17] , \nScanOut30[16] , \nScanOut30[15] , \nScanOut30[14] , 
        \nScanOut30[13] , \nScanOut30[12] , \nScanOut30[11] , \nScanOut30[10] , 
        \nScanOut30[9] , \nScanOut30[8] , \nScanOut30[7] , \nScanOut30[6] , 
        \nScanOut30[5] , \nScanOut30[4] , \nScanOut30[3] , \nScanOut30[2] , 
        \nScanOut30[1] , \nScanOut30[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_14[31] , 
        \nOut1_14[30] , \nOut1_14[29] , \nOut1_14[28] , \nOut1_14[27] , 
        \nOut1_14[26] , \nOut1_14[25] , \nOut1_14[24] , \nOut1_14[23] , 
        \nOut1_14[22] , \nOut1_14[21] , \nOut1_14[20] , \nOut1_14[19] , 
        \nOut1_14[18] , \nOut1_14[17] , \nOut1_14[16] , \nOut1_14[15] , 
        \nOut1_14[14] , \nOut1_14[13] , \nOut1_14[12] , \nOut1_14[11] , 
        \nOut1_14[10] , \nOut1_14[9] , \nOut1_14[8] , \nOut1_14[7] , 
        \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , \nOut1_14[3] , 
        \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), .NORTH_EDGE({
        \nOut1_13[31] , \nOut1_13[30] , \nOut1_13[29] , \nOut1_13[28] , 
        \nOut1_13[27] , \nOut1_13[26] , \nOut1_13[25] , \nOut1_13[24] , 
        \nOut1_13[23] , \nOut1_13[22] , \nOut1_13[21] , \nOut1_13[20] , 
        \nOut1_13[19] , \nOut1_13[18] , \nOut1_13[17] , \nOut1_13[16] , 
        \nOut1_13[15] , \nOut1_13[14] , \nOut1_13[13] , \nOut1_13[12] , 
        \nOut1_13[11] , \nOut1_13[10] , \nOut1_13[9] , \nOut1_13[8] , 
        \nOut1_13[7] , \nOut1_13[6] , \nOut1_13[5] , \nOut1_13[4] , 
        \nOut1_13[3] , \nOut1_13[2] , \nOut1_13[1] , \nOut1_13[0] }), 
        .SOUTH_EDGE({\nOut1_15[31] , \nOut1_15[30] , \nOut1_15[29] , 
        \nOut1_15[28] , \nOut1_15[27] , \nOut1_15[26] , \nOut1_15[25] , 
        \nOut1_15[24] , \nOut1_15[23] , \nOut1_15[22] , \nOut1_15[21] , 
        \nOut1_15[20] , \nOut1_15[19] , \nOut1_15[18] , \nOut1_15[17] , 
        \nOut1_15[16] , \nOut1_15[15] , \nOut1_15[14] , \nOut1_15[13] , 
        \nOut1_15[12] , \nOut1_15[11] , \nOut1_15[10] , \nOut1_15[9] , 
        \nOut1_15[8] , \nOut1_15[7] , \nOut1_15[6] , \nOut1_15[5] , 
        \nOut1_15[4] , \nOut1_15[3] , \nOut1_15[2] , \nOut1_15[1] , 
        \nOut1_15[0] }), .EAST_EDGE(\nOut2_14[31] ), .WEST_EDGE(\nOut0_14[0] ), 
        .NW_EDGE(\nOut0_13[0] ), .SW_EDGE(\nOut0_15[0] ), .NE_EDGE(
        \nOut2_13[31] ), .SE_EDGE(\nOut2_15[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_10 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut11[31] , \nScanOut11[30] , \nScanOut11[29] , 
        \nScanOut11[28] , \nScanOut11[27] , \nScanOut11[26] , \nScanOut11[25] , 
        \nScanOut11[24] , \nScanOut11[23] , \nScanOut11[22] , \nScanOut11[21] , 
        \nScanOut11[20] , \nScanOut11[19] , \nScanOut11[18] , \nScanOut11[17] , 
        \nScanOut11[16] , \nScanOut11[15] , \nScanOut11[14] , \nScanOut11[13] , 
        \nScanOut11[12] , \nScanOut11[11] , \nScanOut11[10] , \nScanOut11[9] , 
        \nScanOut11[8] , \nScanOut11[7] , \nScanOut11[6] , \nScanOut11[5] , 
        \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , \nScanOut11[1] , 
        \nScanOut11[0] }), .ScanOut({\nScanOut10[31] , \nScanOut10[30] , 
        \nScanOut10[29] , \nScanOut10[28] , \nScanOut10[27] , \nScanOut10[26] , 
        \nScanOut10[25] , \nScanOut10[24] , \nScanOut10[23] , \nScanOut10[22] , 
        \nScanOut10[21] , \nScanOut10[20] , \nScanOut10[19] , \nScanOut10[18] , 
        \nScanOut10[17] , \nScanOut10[16] , \nScanOut10[15] , \nScanOut10[14] , 
        \nScanOut10[13] , \nScanOut10[12] , \nScanOut10[11] , \nScanOut10[10] , 
        \nScanOut10[9] , \nScanOut10[8] , \nScanOut10[7] , \nScanOut10[6] , 
        \nScanOut10[5] , \nScanOut10[4] , \nScanOut10[3] , \nScanOut10[2] , 
        \nScanOut10[1] , \nScanOut10[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_10[31] , 
        \nOut0_10[30] , \nOut0_10[29] , \nOut0_10[28] , \nOut0_10[27] , 
        \nOut0_10[26] , \nOut0_10[25] , \nOut0_10[24] , \nOut0_10[23] , 
        \nOut0_10[22] , \nOut0_10[21] , \nOut0_10[20] , \nOut0_10[19] , 
        \nOut0_10[18] , \nOut0_10[17] , \nOut0_10[16] , \nOut0_10[15] , 
        \nOut0_10[14] , \nOut0_10[13] , \nOut0_10[12] , \nOut0_10[11] , 
        \nOut0_10[10] , \nOut0_10[9] , \nOut0_10[8] , \nOut0_10[7] , 
        \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , \nOut0_10[3] , 
        \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), .NORTH_EDGE({
        \nOut0_9[31] , \nOut0_9[30] , \nOut0_9[29] , \nOut0_9[28] , 
        \nOut0_9[27] , \nOut0_9[26] , \nOut0_9[25] , \nOut0_9[24] , 
        \nOut0_9[23] , \nOut0_9[22] , \nOut0_9[21] , \nOut0_9[20] , 
        \nOut0_9[19] , \nOut0_9[18] , \nOut0_9[17] , \nOut0_9[16] , 
        \nOut0_9[15] , \nOut0_9[14] , \nOut0_9[13] , \nOut0_9[12] , 
        \nOut0_9[11] , \nOut0_9[10] , \nOut0_9[9] , \nOut0_9[8] , \nOut0_9[7] , 
        \nOut0_9[6] , \nOut0_9[5] , \nOut0_9[4] , \nOut0_9[3] , \nOut0_9[2] , 
        \nOut0_9[1] , \nOut0_9[0] }), .SOUTH_EDGE({\nOut0_11[31] , 
        \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , \nOut0_11[27] , 
        \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , \nOut0_11[23] , 
        \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , \nOut0_11[19] , 
        \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , \nOut0_11[15] , 
        \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , \nOut0_11[11] , 
        \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , \nOut0_11[7] , 
        \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , 
        \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .EAST_EDGE(
        \nOut1_10[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_9[31] ), .SE_EDGE(\nOut1_11[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_37 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut38[31] , \nScanOut38[30] , \nScanOut38[29] , 
        \nScanOut38[28] , \nScanOut38[27] , \nScanOut38[26] , \nScanOut38[25] , 
        \nScanOut38[24] , \nScanOut38[23] , \nScanOut38[22] , \nScanOut38[21] , 
        \nScanOut38[20] , \nScanOut38[19] , \nScanOut38[18] , \nScanOut38[17] , 
        \nScanOut38[16] , \nScanOut38[15] , \nScanOut38[14] , \nScanOut38[13] , 
        \nScanOut38[12] , \nScanOut38[11] , \nScanOut38[10] , \nScanOut38[9] , 
        \nScanOut38[8] , \nScanOut38[7] , \nScanOut38[6] , \nScanOut38[5] , 
        \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , \nScanOut38[1] , 
        \nScanOut38[0] }), .ScanOut({\nScanOut37[31] , \nScanOut37[30] , 
        \nScanOut37[29] , \nScanOut37[28] , \nScanOut37[27] , \nScanOut37[26] , 
        \nScanOut37[25] , \nScanOut37[24] , \nScanOut37[23] , \nScanOut37[22] , 
        \nScanOut37[21] , \nScanOut37[20] , \nScanOut37[19] , \nScanOut37[18] , 
        \nScanOut37[17] , \nScanOut37[16] , \nScanOut37[15] , \nScanOut37[14] , 
        \nScanOut37[13] , \nScanOut37[12] , \nScanOut37[11] , \nScanOut37[10] , 
        \nScanOut37[9] , \nScanOut37[8] , \nScanOut37[7] , \nScanOut37[6] , 
        \nScanOut37[5] , \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , 
        \nScanOut37[1] , \nScanOut37[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_5[31] , 
        \nOut2_5[30] , \nOut2_5[29] , \nOut2_5[28] , \nOut2_5[27] , 
        \nOut2_5[26] , \nOut2_5[25] , \nOut2_5[24] , \nOut2_5[23] , 
        \nOut2_5[22] , \nOut2_5[21] , \nOut2_5[20] , \nOut2_5[19] , 
        \nOut2_5[18] , \nOut2_5[17] , \nOut2_5[16] , \nOut2_5[15] , 
        \nOut2_5[14] , \nOut2_5[13] , \nOut2_5[12] , \nOut2_5[11] , 
        \nOut2_5[10] , \nOut2_5[9] , \nOut2_5[8] , \nOut2_5[7] , \nOut2_5[6] , 
        \nOut2_5[5] , \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , 
        \nOut2_5[0] }), .NORTH_EDGE({\nOut2_4[31] , \nOut2_4[30] , 
        \nOut2_4[29] , \nOut2_4[28] , \nOut2_4[27] , \nOut2_4[26] , 
        \nOut2_4[25] , \nOut2_4[24] , \nOut2_4[23] , \nOut2_4[22] , 
        \nOut2_4[21] , \nOut2_4[20] , \nOut2_4[19] , \nOut2_4[18] , 
        \nOut2_4[17] , \nOut2_4[16] , \nOut2_4[15] , \nOut2_4[14] , 
        \nOut2_4[13] , \nOut2_4[12] , \nOut2_4[11] , \nOut2_4[10] , 
        \nOut2_4[9] , \nOut2_4[8] , \nOut2_4[7] , \nOut2_4[6] , \nOut2_4[5] , 
        \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , \nOut2_4[0] }), 
        .SOUTH_EDGE({\nOut2_6[31] , \nOut2_6[30] , \nOut2_6[29] , 
        \nOut2_6[28] , \nOut2_6[27] , \nOut2_6[26] , \nOut2_6[25] , 
        \nOut2_6[24] , \nOut2_6[23] , \nOut2_6[22] , \nOut2_6[21] , 
        \nOut2_6[20] , \nOut2_6[19] , \nOut2_6[18] , \nOut2_6[17] , 
        \nOut2_6[16] , \nOut2_6[15] , \nOut2_6[14] , \nOut2_6[13] , 
        \nOut2_6[12] , \nOut2_6[11] , \nOut2_6[10] , \nOut2_6[9] , 
        \nOut2_6[8] , \nOut2_6[7] , \nOut2_6[6] , \nOut2_6[5] , \nOut2_6[4] , 
        \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , \nOut2_6[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_5[0] ), .NW_EDGE(\nOut1_4[0] ), .SW_EDGE(
        \nOut1_6[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_42 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut43[31] , \nScanOut43[30] , \nScanOut43[29] , 
        \nScanOut43[28] , \nScanOut43[27] , \nScanOut43[26] , \nScanOut43[25] , 
        \nScanOut43[24] , \nScanOut43[23] , \nScanOut43[22] , \nScanOut43[21] , 
        \nScanOut43[20] , \nScanOut43[19] , \nScanOut43[18] , \nScanOut43[17] , 
        \nScanOut43[16] , \nScanOut43[15] , \nScanOut43[14] , \nScanOut43[13] , 
        \nScanOut43[12] , \nScanOut43[11] , \nScanOut43[10] , \nScanOut43[9] , 
        \nScanOut43[8] , \nScanOut43[7] , \nScanOut43[6] , \nScanOut43[5] , 
        \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , \nScanOut43[1] , 
        \nScanOut43[0] }), .ScanOut({\nScanOut42[31] , \nScanOut42[30] , 
        \nScanOut42[29] , \nScanOut42[28] , \nScanOut42[27] , \nScanOut42[26] , 
        \nScanOut42[25] , \nScanOut42[24] , \nScanOut42[23] , \nScanOut42[22] , 
        \nScanOut42[21] , \nScanOut42[20] , \nScanOut42[19] , \nScanOut42[18] , 
        \nScanOut42[17] , \nScanOut42[16] , \nScanOut42[15] , \nScanOut42[14] , 
        \nScanOut42[13] , \nScanOut42[12] , \nScanOut42[11] , \nScanOut42[10] , 
        \nScanOut42[9] , \nScanOut42[8] , \nScanOut42[7] , \nScanOut42[6] , 
        \nScanOut42[5] , \nScanOut42[4] , \nScanOut42[3] , \nScanOut42[2] , 
        \nScanOut42[1] , \nScanOut42[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_10[31] , 
        \nOut2_10[30] , \nOut2_10[29] , \nOut2_10[28] , \nOut2_10[27] , 
        \nOut2_10[26] , \nOut2_10[25] , \nOut2_10[24] , \nOut2_10[23] , 
        \nOut2_10[22] , \nOut2_10[21] , \nOut2_10[20] , \nOut2_10[19] , 
        \nOut2_10[18] , \nOut2_10[17] , \nOut2_10[16] , \nOut2_10[15] , 
        \nOut2_10[14] , \nOut2_10[13] , \nOut2_10[12] , \nOut2_10[11] , 
        \nOut2_10[10] , \nOut2_10[9] , \nOut2_10[8] , \nOut2_10[7] , 
        \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , \nOut2_10[3] , 
        \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), .NORTH_EDGE({
        \nOut2_9[31] , \nOut2_9[30] , \nOut2_9[29] , \nOut2_9[28] , 
        \nOut2_9[27] , \nOut2_9[26] , \nOut2_9[25] , \nOut2_9[24] , 
        \nOut2_9[23] , \nOut2_9[22] , \nOut2_9[21] , \nOut2_9[20] , 
        \nOut2_9[19] , \nOut2_9[18] , \nOut2_9[17] , \nOut2_9[16] , 
        \nOut2_9[15] , \nOut2_9[14] , \nOut2_9[13] , \nOut2_9[12] , 
        \nOut2_9[11] , \nOut2_9[10] , \nOut2_9[9] , \nOut2_9[8] , \nOut2_9[7] , 
        \nOut2_9[6] , \nOut2_9[5] , \nOut2_9[4] , \nOut2_9[3] , \nOut2_9[2] , 
        \nOut2_9[1] , \nOut2_9[0] }), .SOUTH_EDGE({\nOut2_11[31] , 
        \nOut2_11[30] , \nOut2_11[29] , \nOut2_11[28] , \nOut2_11[27] , 
        \nOut2_11[26] , \nOut2_11[25] , \nOut2_11[24] , \nOut2_11[23] , 
        \nOut2_11[22] , \nOut2_11[21] , \nOut2_11[20] , \nOut2_11[19] , 
        \nOut2_11[18] , \nOut2_11[17] , \nOut2_11[16] , \nOut2_11[15] , 
        \nOut2_11[14] , \nOut2_11[13] , \nOut2_11[12] , \nOut2_11[11] , 
        \nOut2_11[10] , \nOut2_11[9] , \nOut2_11[8] , \nOut2_11[7] , 
        \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , \nOut2_11[3] , 
        \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .EAST_EDGE(1'b0), 
        .WEST_EDGE(\nOut1_10[0] ), .NW_EDGE(\nOut1_9[0] ), .SW_EDGE(
        \nOut1_11[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_45 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut46[31] , \nScanOut46[30] , \nScanOut46[29] , 
        \nScanOut46[28] , \nScanOut46[27] , \nScanOut46[26] , \nScanOut46[25] , 
        \nScanOut46[24] , \nScanOut46[23] , \nScanOut46[22] , \nScanOut46[21] , 
        \nScanOut46[20] , \nScanOut46[19] , \nScanOut46[18] , \nScanOut46[17] , 
        \nScanOut46[16] , \nScanOut46[15] , \nScanOut46[14] , \nScanOut46[13] , 
        \nScanOut46[12] , \nScanOut46[11] , \nScanOut46[10] , \nScanOut46[9] , 
        \nScanOut46[8] , \nScanOut46[7] , \nScanOut46[6] , \nScanOut46[5] , 
        \nScanOut46[4] , \nScanOut46[3] , \nScanOut46[2] , \nScanOut46[1] , 
        \nScanOut46[0] }), .ScanOut({\nScanOut45[31] , \nScanOut45[30] , 
        \nScanOut45[29] , \nScanOut45[28] , \nScanOut45[27] , \nScanOut45[26] , 
        \nScanOut45[25] , \nScanOut45[24] , \nScanOut45[23] , \nScanOut45[22] , 
        \nScanOut45[21] , \nScanOut45[20] , \nScanOut45[19] , \nScanOut45[18] , 
        \nScanOut45[17] , \nScanOut45[16] , \nScanOut45[15] , \nScanOut45[14] , 
        \nScanOut45[13] , \nScanOut45[12] , \nScanOut45[11] , \nScanOut45[10] , 
        \nScanOut45[9] , \nScanOut45[8] , \nScanOut45[7] , \nScanOut45[6] , 
        \nScanOut45[5] , \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , 
        \nScanOut45[1] , \nScanOut45[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_13[31] , 
        \nOut2_13[30] , \nOut2_13[29] , \nOut2_13[28] , \nOut2_13[27] , 
        \nOut2_13[26] , \nOut2_13[25] , \nOut2_13[24] , \nOut2_13[23] , 
        \nOut2_13[22] , \nOut2_13[21] , \nOut2_13[20] , \nOut2_13[19] , 
        \nOut2_13[18] , \nOut2_13[17] , \nOut2_13[16] , \nOut2_13[15] , 
        \nOut2_13[14] , \nOut2_13[13] , \nOut2_13[12] , \nOut2_13[11] , 
        \nOut2_13[10] , \nOut2_13[9] , \nOut2_13[8] , \nOut2_13[7] , 
        \nOut2_13[6] , \nOut2_13[5] , \nOut2_13[4] , \nOut2_13[3] , 
        \nOut2_13[2] , \nOut2_13[1] , \nOut2_13[0] }), .NORTH_EDGE({
        \nOut2_12[31] , \nOut2_12[30] , \nOut2_12[29] , \nOut2_12[28] , 
        \nOut2_12[27] , \nOut2_12[26] , \nOut2_12[25] , \nOut2_12[24] , 
        \nOut2_12[23] , \nOut2_12[22] , \nOut2_12[21] , \nOut2_12[20] , 
        \nOut2_12[19] , \nOut2_12[18] , \nOut2_12[17] , \nOut2_12[16] , 
        \nOut2_12[15] , \nOut2_12[14] , \nOut2_12[13] , \nOut2_12[12] , 
        \nOut2_12[11] , \nOut2_12[10] , \nOut2_12[9] , \nOut2_12[8] , 
        \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , 
        \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), 
        .SOUTH_EDGE({\nOut2_14[31] , \nOut2_14[30] , \nOut2_14[29] , 
        \nOut2_14[28] , \nOut2_14[27] , \nOut2_14[26] , \nOut2_14[25] , 
        \nOut2_14[24] , \nOut2_14[23] , \nOut2_14[22] , \nOut2_14[21] , 
        \nOut2_14[20] , \nOut2_14[19] , \nOut2_14[18] , \nOut2_14[17] , 
        \nOut2_14[16] , \nOut2_14[15] , \nOut2_14[14] , \nOut2_14[13] , 
        \nOut2_14[12] , \nOut2_14[11] , \nOut2_14[10] , \nOut2_14[9] , 
        \nOut2_14[8] , \nOut2_14[7] , \nOut2_14[6] , \nOut2_14[5] , 
        \nOut2_14[4] , \nOut2_14[3] , \nOut2_14[2] , \nOut2_14[1] , 
        \nOut2_14[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_13[0] ), 
        .NW_EDGE(\nOut1_12[0] ), .SW_EDGE(\nOut1_14[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_25 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut26[31] , \nScanOut26[30] , \nScanOut26[29] , 
        \nScanOut26[28] , \nScanOut26[27] , \nScanOut26[26] , \nScanOut26[25] , 
        \nScanOut26[24] , \nScanOut26[23] , \nScanOut26[22] , \nScanOut26[21] , 
        \nScanOut26[20] , \nScanOut26[19] , \nScanOut26[18] , \nScanOut26[17] , 
        \nScanOut26[16] , \nScanOut26[15] , \nScanOut26[14] , \nScanOut26[13] , 
        \nScanOut26[12] , \nScanOut26[11] , \nScanOut26[10] , \nScanOut26[9] , 
        \nScanOut26[8] , \nScanOut26[7] , \nScanOut26[6] , \nScanOut26[5] , 
        \nScanOut26[4] , \nScanOut26[3] , \nScanOut26[2] , \nScanOut26[1] , 
        \nScanOut26[0] }), .ScanOut({\nScanOut25[31] , \nScanOut25[30] , 
        \nScanOut25[29] , \nScanOut25[28] , \nScanOut25[27] , \nScanOut25[26] , 
        \nScanOut25[25] , \nScanOut25[24] , \nScanOut25[23] , \nScanOut25[22] , 
        \nScanOut25[21] , \nScanOut25[20] , \nScanOut25[19] , \nScanOut25[18] , 
        \nScanOut25[17] , \nScanOut25[16] , \nScanOut25[15] , \nScanOut25[14] , 
        \nScanOut25[13] , \nScanOut25[12] , \nScanOut25[11] , \nScanOut25[10] , 
        \nScanOut25[9] , \nScanOut25[8] , \nScanOut25[7] , \nScanOut25[6] , 
        \nScanOut25[5] , \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , 
        \nScanOut25[1] , \nScanOut25[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_9[31] , 
        \nOut1_9[30] , \nOut1_9[29] , \nOut1_9[28] , \nOut1_9[27] , 
        \nOut1_9[26] , \nOut1_9[25] , \nOut1_9[24] , \nOut1_9[23] , 
        \nOut1_9[22] , \nOut1_9[21] , \nOut1_9[20] , \nOut1_9[19] , 
        \nOut1_9[18] , \nOut1_9[17] , \nOut1_9[16] , \nOut1_9[15] , 
        \nOut1_9[14] , \nOut1_9[13] , \nOut1_9[12] , \nOut1_9[11] , 
        \nOut1_9[10] , \nOut1_9[9] , \nOut1_9[8] , \nOut1_9[7] , \nOut1_9[6] , 
        \nOut1_9[5] , \nOut1_9[4] , \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , 
        \nOut1_9[0] }), .NORTH_EDGE({\nOut1_8[31] , \nOut1_8[30] , 
        \nOut1_8[29] , \nOut1_8[28] , \nOut1_8[27] , \nOut1_8[26] , 
        \nOut1_8[25] , \nOut1_8[24] , \nOut1_8[23] , \nOut1_8[22] , 
        \nOut1_8[21] , \nOut1_8[20] , \nOut1_8[19] , \nOut1_8[18] , 
        \nOut1_8[17] , \nOut1_8[16] , \nOut1_8[15] , \nOut1_8[14] , 
        \nOut1_8[13] , \nOut1_8[12] , \nOut1_8[11] , \nOut1_8[10] , 
        \nOut1_8[9] , \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , 
        \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), 
        .SOUTH_EDGE({\nOut1_10[31] , \nOut1_10[30] , \nOut1_10[29] , 
        \nOut1_10[28] , \nOut1_10[27] , \nOut1_10[26] , \nOut1_10[25] , 
        \nOut1_10[24] , \nOut1_10[23] , \nOut1_10[22] , \nOut1_10[21] , 
        \nOut1_10[20] , \nOut1_10[19] , \nOut1_10[18] , \nOut1_10[17] , 
        \nOut1_10[16] , \nOut1_10[15] , \nOut1_10[14] , \nOut1_10[13] , 
        \nOut1_10[12] , \nOut1_10[11] , \nOut1_10[10] , \nOut1_10[9] , 
        \nOut1_10[8] , \nOut1_10[7] , \nOut1_10[6] , \nOut1_10[5] , 
        \nOut1_10[4] , \nOut1_10[3] , \nOut1_10[2] , \nOut1_10[1] , 
        \nOut1_10[0] }), .EAST_EDGE(\nOut2_9[31] ), .WEST_EDGE(\nOut0_9[0] ), 
        .NW_EDGE(\nOut0_8[0] ), .SW_EDGE(\nOut0_10[0] ), .NE_EDGE(
        \nOut2_8[31] ), .SE_EDGE(\nOut2_10[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_11 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut12[31] , \nScanOut12[30] , \nScanOut12[29] , 
        \nScanOut12[28] , \nScanOut12[27] , \nScanOut12[26] , \nScanOut12[25] , 
        \nScanOut12[24] , \nScanOut12[23] , \nScanOut12[22] , \nScanOut12[21] , 
        \nScanOut12[20] , \nScanOut12[19] , \nScanOut12[18] , \nScanOut12[17] , 
        \nScanOut12[16] , \nScanOut12[15] , \nScanOut12[14] , \nScanOut12[13] , 
        \nScanOut12[12] , \nScanOut12[11] , \nScanOut12[10] , \nScanOut12[9] , 
        \nScanOut12[8] , \nScanOut12[7] , \nScanOut12[6] , \nScanOut12[5] , 
        \nScanOut12[4] , \nScanOut12[3] , \nScanOut12[2] , \nScanOut12[1] , 
        \nScanOut12[0] }), .ScanOut({\nScanOut11[31] , \nScanOut11[30] , 
        \nScanOut11[29] , \nScanOut11[28] , \nScanOut11[27] , \nScanOut11[26] , 
        \nScanOut11[25] , \nScanOut11[24] , \nScanOut11[23] , \nScanOut11[22] , 
        \nScanOut11[21] , \nScanOut11[20] , \nScanOut11[19] , \nScanOut11[18] , 
        \nScanOut11[17] , \nScanOut11[16] , \nScanOut11[15] , \nScanOut11[14] , 
        \nScanOut11[13] , \nScanOut11[12] , \nScanOut11[11] , \nScanOut11[10] , 
        \nScanOut11[9] , \nScanOut11[8] , \nScanOut11[7] , \nScanOut11[6] , 
        \nScanOut11[5] , \nScanOut11[4] , \nScanOut11[3] , \nScanOut11[2] , 
        \nScanOut11[1] , \nScanOut11[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_11[31] , 
        \nOut0_11[30] , \nOut0_11[29] , \nOut0_11[28] , \nOut0_11[27] , 
        \nOut0_11[26] , \nOut0_11[25] , \nOut0_11[24] , \nOut0_11[23] , 
        \nOut0_11[22] , \nOut0_11[21] , \nOut0_11[20] , \nOut0_11[19] , 
        \nOut0_11[18] , \nOut0_11[17] , \nOut0_11[16] , \nOut0_11[15] , 
        \nOut0_11[14] , \nOut0_11[13] , \nOut0_11[12] , \nOut0_11[11] , 
        \nOut0_11[10] , \nOut0_11[9] , \nOut0_11[8] , \nOut0_11[7] , 
        \nOut0_11[6] , \nOut0_11[5] , \nOut0_11[4] , \nOut0_11[3] , 
        \nOut0_11[2] , \nOut0_11[1] , \nOut0_11[0] }), .NORTH_EDGE({
        \nOut0_10[31] , \nOut0_10[30] , \nOut0_10[29] , \nOut0_10[28] , 
        \nOut0_10[27] , \nOut0_10[26] , \nOut0_10[25] , \nOut0_10[24] , 
        \nOut0_10[23] , \nOut0_10[22] , \nOut0_10[21] , \nOut0_10[20] , 
        \nOut0_10[19] , \nOut0_10[18] , \nOut0_10[17] , \nOut0_10[16] , 
        \nOut0_10[15] , \nOut0_10[14] , \nOut0_10[13] , \nOut0_10[12] , 
        \nOut0_10[11] , \nOut0_10[10] , \nOut0_10[9] , \nOut0_10[8] , 
        \nOut0_10[7] , \nOut0_10[6] , \nOut0_10[5] , \nOut0_10[4] , 
        \nOut0_10[3] , \nOut0_10[2] , \nOut0_10[1] , \nOut0_10[0] }), 
        .SOUTH_EDGE({\nOut0_12[31] , \nOut0_12[30] , \nOut0_12[29] , 
        \nOut0_12[28] , \nOut0_12[27] , \nOut0_12[26] , \nOut0_12[25] , 
        \nOut0_12[24] , \nOut0_12[23] , \nOut0_12[22] , \nOut0_12[21] , 
        \nOut0_12[20] , \nOut0_12[19] , \nOut0_12[18] , \nOut0_12[17] , 
        \nOut0_12[16] , \nOut0_12[15] , \nOut0_12[14] , \nOut0_12[13] , 
        \nOut0_12[12] , \nOut0_12[11] , \nOut0_12[10] , \nOut0_12[9] , 
        \nOut0_12[8] , \nOut0_12[7] , \nOut0_12[6] , \nOut0_12[5] , 
        \nOut0_12[4] , \nOut0_12[3] , \nOut0_12[2] , \nOut0_12[1] , 
        \nOut0_12[0] }), .EAST_EDGE(\nOut1_11[31] ), .WEST_EDGE(1'b0), 
        .NW_EDGE(1'b0), .SW_EDGE(1'b0), .NE_EDGE(\nOut1_10[31] ), .SE_EDGE(
        \nOut1_12[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_19 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut20[31] , \nScanOut20[30] , \nScanOut20[29] , 
        \nScanOut20[28] , \nScanOut20[27] , \nScanOut20[26] , \nScanOut20[25] , 
        \nScanOut20[24] , \nScanOut20[23] , \nScanOut20[22] , \nScanOut20[21] , 
        \nScanOut20[20] , \nScanOut20[19] , \nScanOut20[18] , \nScanOut20[17] , 
        \nScanOut20[16] , \nScanOut20[15] , \nScanOut20[14] , \nScanOut20[13] , 
        \nScanOut20[12] , \nScanOut20[11] , \nScanOut20[10] , \nScanOut20[9] , 
        \nScanOut20[8] , \nScanOut20[7] , \nScanOut20[6] , \nScanOut20[5] , 
        \nScanOut20[4] , \nScanOut20[3] , \nScanOut20[2] , \nScanOut20[1] , 
        \nScanOut20[0] }), .ScanOut({\nScanOut19[31] , \nScanOut19[30] , 
        \nScanOut19[29] , \nScanOut19[28] , \nScanOut19[27] , \nScanOut19[26] , 
        \nScanOut19[25] , \nScanOut19[24] , \nScanOut19[23] , \nScanOut19[22] , 
        \nScanOut19[21] , \nScanOut19[20] , \nScanOut19[19] , \nScanOut19[18] , 
        \nScanOut19[17] , \nScanOut19[16] , \nScanOut19[15] , \nScanOut19[14] , 
        \nScanOut19[13] , \nScanOut19[12] , \nScanOut19[11] , \nScanOut19[10] , 
        \nScanOut19[9] , \nScanOut19[8] , \nScanOut19[7] , \nScanOut19[6] , 
        \nScanOut19[5] , \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , 
        \nScanOut19[1] , \nScanOut19[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_3[31] , 
        \nOut1_3[30] , \nOut1_3[29] , \nOut1_3[28] , \nOut1_3[27] , 
        \nOut1_3[26] , \nOut1_3[25] , \nOut1_3[24] , \nOut1_3[23] , 
        \nOut1_3[22] , \nOut1_3[21] , \nOut1_3[20] , \nOut1_3[19] , 
        \nOut1_3[18] , \nOut1_3[17] , \nOut1_3[16] , \nOut1_3[15] , 
        \nOut1_3[14] , \nOut1_3[13] , \nOut1_3[12] , \nOut1_3[11] , 
        \nOut1_3[10] , \nOut1_3[9] , \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , 
        \nOut1_3[5] , \nOut1_3[4] , \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , 
        \nOut1_3[0] }), .NORTH_EDGE({\nOut1_2[31] , \nOut1_2[30] , 
        \nOut1_2[29] , \nOut1_2[28] , \nOut1_2[27] , \nOut1_2[26] , 
        \nOut1_2[25] , \nOut1_2[24] , \nOut1_2[23] , \nOut1_2[22] , 
        \nOut1_2[21] , \nOut1_2[20] , \nOut1_2[19] , \nOut1_2[18] , 
        \nOut1_2[17] , \nOut1_2[16] , \nOut1_2[15] , \nOut1_2[14] , 
        \nOut1_2[13] , \nOut1_2[12] , \nOut1_2[11] , \nOut1_2[10] , 
        \nOut1_2[9] , \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , \nOut1_2[5] , 
        \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , \nOut1_2[0] }), 
        .SOUTH_EDGE({\nOut1_4[31] , \nOut1_4[30] , \nOut1_4[29] , 
        \nOut1_4[28] , \nOut1_4[27] , \nOut1_4[26] , \nOut1_4[25] , 
        \nOut1_4[24] , \nOut1_4[23] , \nOut1_4[22] , \nOut1_4[21] , 
        \nOut1_4[20] , \nOut1_4[19] , \nOut1_4[18] , \nOut1_4[17] , 
        \nOut1_4[16] , \nOut1_4[15] , \nOut1_4[14] , \nOut1_4[13] , 
        \nOut1_4[12] , \nOut1_4[11] , \nOut1_4[10] , \nOut1_4[9] , 
        \nOut1_4[8] , \nOut1_4[7] , \nOut1_4[6] , \nOut1_4[5] , \nOut1_4[4] , 
        \nOut1_4[3] , \nOut1_4[2] , \nOut1_4[1] , \nOut1_4[0] }), .EAST_EDGE(
        \nOut2_3[31] ), .WEST_EDGE(\nOut0_3[0] ), .NW_EDGE(\nOut0_2[0] ), 
        .SW_EDGE(\nOut0_4[0] ), .NE_EDGE(\nOut2_2[31] ), .SE_EDGE(
        \nOut2_4[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_36 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut37[31] , \nScanOut37[30] , \nScanOut37[29] , 
        \nScanOut37[28] , \nScanOut37[27] , \nScanOut37[26] , \nScanOut37[25] , 
        \nScanOut37[24] , \nScanOut37[23] , \nScanOut37[22] , \nScanOut37[21] , 
        \nScanOut37[20] , \nScanOut37[19] , \nScanOut37[18] , \nScanOut37[17] , 
        \nScanOut37[16] , \nScanOut37[15] , \nScanOut37[14] , \nScanOut37[13] , 
        \nScanOut37[12] , \nScanOut37[11] , \nScanOut37[10] , \nScanOut37[9] , 
        \nScanOut37[8] , \nScanOut37[7] , \nScanOut37[6] , \nScanOut37[5] , 
        \nScanOut37[4] , \nScanOut37[3] , \nScanOut37[2] , \nScanOut37[1] , 
        \nScanOut37[0] }), .ScanOut({\nScanOut36[31] , \nScanOut36[30] , 
        \nScanOut36[29] , \nScanOut36[28] , \nScanOut36[27] , \nScanOut36[26] , 
        \nScanOut36[25] , \nScanOut36[24] , \nScanOut36[23] , \nScanOut36[22] , 
        \nScanOut36[21] , \nScanOut36[20] , \nScanOut36[19] , \nScanOut36[18] , 
        \nScanOut36[17] , \nScanOut36[16] , \nScanOut36[15] , \nScanOut36[14] , 
        \nScanOut36[13] , \nScanOut36[12] , \nScanOut36[11] , \nScanOut36[10] , 
        \nScanOut36[9] , \nScanOut36[8] , \nScanOut36[7] , \nScanOut36[6] , 
        \nScanOut36[5] , \nScanOut36[4] , \nScanOut36[3] , \nScanOut36[2] , 
        \nScanOut36[1] , \nScanOut36[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_4[31] , 
        \nOut2_4[30] , \nOut2_4[29] , \nOut2_4[28] , \nOut2_4[27] , 
        \nOut2_4[26] , \nOut2_4[25] , \nOut2_4[24] , \nOut2_4[23] , 
        \nOut2_4[22] , \nOut2_4[21] , \nOut2_4[20] , \nOut2_4[19] , 
        \nOut2_4[18] , \nOut2_4[17] , \nOut2_4[16] , \nOut2_4[15] , 
        \nOut2_4[14] , \nOut2_4[13] , \nOut2_4[12] , \nOut2_4[11] , 
        \nOut2_4[10] , \nOut2_4[9] , \nOut2_4[8] , \nOut2_4[7] , \nOut2_4[6] , 
        \nOut2_4[5] , \nOut2_4[4] , \nOut2_4[3] , \nOut2_4[2] , \nOut2_4[1] , 
        \nOut2_4[0] }), .NORTH_EDGE({\nOut2_3[31] , \nOut2_3[30] , 
        \nOut2_3[29] , \nOut2_3[28] , \nOut2_3[27] , \nOut2_3[26] , 
        \nOut2_3[25] , \nOut2_3[24] , \nOut2_3[23] , \nOut2_3[22] , 
        \nOut2_3[21] , \nOut2_3[20] , \nOut2_3[19] , \nOut2_3[18] , 
        \nOut2_3[17] , \nOut2_3[16] , \nOut2_3[15] , \nOut2_3[14] , 
        \nOut2_3[13] , \nOut2_3[12] , \nOut2_3[11] , \nOut2_3[10] , 
        \nOut2_3[9] , \nOut2_3[8] , \nOut2_3[7] , \nOut2_3[6] , \nOut2_3[5] , 
        \nOut2_3[4] , \nOut2_3[3] , \nOut2_3[2] , \nOut2_3[1] , \nOut2_3[0] }), 
        .SOUTH_EDGE({\nOut2_5[31] , \nOut2_5[30] , \nOut2_5[29] , 
        \nOut2_5[28] , \nOut2_5[27] , \nOut2_5[26] , \nOut2_5[25] , 
        \nOut2_5[24] , \nOut2_5[23] , \nOut2_5[22] , \nOut2_5[21] , 
        \nOut2_5[20] , \nOut2_5[19] , \nOut2_5[18] , \nOut2_5[17] , 
        \nOut2_5[16] , \nOut2_5[15] , \nOut2_5[14] , \nOut2_5[13] , 
        \nOut2_5[12] , \nOut2_5[11] , \nOut2_5[10] , \nOut2_5[9] , 
        \nOut2_5[8] , \nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , \nOut2_5[4] , 
        \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_4[0] ), .NW_EDGE(\nOut1_3[0] ), .SW_EDGE(
        \nOut1_5[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_18 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut19[31] , \nScanOut19[30] , \nScanOut19[29] , 
        \nScanOut19[28] , \nScanOut19[27] , \nScanOut19[26] , \nScanOut19[25] , 
        \nScanOut19[24] , \nScanOut19[23] , \nScanOut19[22] , \nScanOut19[21] , 
        \nScanOut19[20] , \nScanOut19[19] , \nScanOut19[18] , \nScanOut19[17] , 
        \nScanOut19[16] , \nScanOut19[15] , \nScanOut19[14] , \nScanOut19[13] , 
        \nScanOut19[12] , \nScanOut19[11] , \nScanOut19[10] , \nScanOut19[9] , 
        \nScanOut19[8] , \nScanOut19[7] , \nScanOut19[6] , \nScanOut19[5] , 
        \nScanOut19[4] , \nScanOut19[3] , \nScanOut19[2] , \nScanOut19[1] , 
        \nScanOut19[0] }), .ScanOut({\nScanOut18[31] , \nScanOut18[30] , 
        \nScanOut18[29] , \nScanOut18[28] , \nScanOut18[27] , \nScanOut18[26] , 
        \nScanOut18[25] , \nScanOut18[24] , \nScanOut18[23] , \nScanOut18[22] , 
        \nScanOut18[21] , \nScanOut18[20] , \nScanOut18[19] , \nScanOut18[18] , 
        \nScanOut18[17] , \nScanOut18[16] , \nScanOut18[15] , \nScanOut18[14] , 
        \nScanOut18[13] , \nScanOut18[12] , \nScanOut18[11] , \nScanOut18[10] , 
        \nScanOut18[9] , \nScanOut18[8] , \nScanOut18[7] , \nScanOut18[6] , 
        \nScanOut18[5] , \nScanOut18[4] , \nScanOut18[3] , \nScanOut18[2] , 
        \nScanOut18[1] , \nScanOut18[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_2[31] , 
        \nOut1_2[30] , \nOut1_2[29] , \nOut1_2[28] , \nOut1_2[27] , 
        \nOut1_2[26] , \nOut1_2[25] , \nOut1_2[24] , \nOut1_2[23] , 
        \nOut1_2[22] , \nOut1_2[21] , \nOut1_2[20] , \nOut1_2[19] , 
        \nOut1_2[18] , \nOut1_2[17] , \nOut1_2[16] , \nOut1_2[15] , 
        \nOut1_2[14] , \nOut1_2[13] , \nOut1_2[12] , \nOut1_2[11] , 
        \nOut1_2[10] , \nOut1_2[9] , \nOut1_2[8] , \nOut1_2[7] , \nOut1_2[6] , 
        \nOut1_2[5] , \nOut1_2[4] , \nOut1_2[3] , \nOut1_2[2] , \nOut1_2[1] , 
        \nOut1_2[0] }), .NORTH_EDGE({\nOut1_1[31] , \nOut1_1[30] , 
        \nOut1_1[29] , \nOut1_1[28] , \nOut1_1[27] , \nOut1_1[26] , 
        \nOut1_1[25] , \nOut1_1[24] , \nOut1_1[23] , \nOut1_1[22] , 
        \nOut1_1[21] , \nOut1_1[20] , \nOut1_1[19] , \nOut1_1[18] , 
        \nOut1_1[17] , \nOut1_1[16] , \nOut1_1[15] , \nOut1_1[14] , 
        \nOut1_1[13] , \nOut1_1[12] , \nOut1_1[11] , \nOut1_1[10] , 
        \nOut1_1[9] , \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , 
        \nOut1_1[4] , \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), 
        .SOUTH_EDGE({\nOut1_3[31] , \nOut1_3[30] , \nOut1_3[29] , 
        \nOut1_3[28] , \nOut1_3[27] , \nOut1_3[26] , \nOut1_3[25] , 
        \nOut1_3[24] , \nOut1_3[23] , \nOut1_3[22] , \nOut1_3[21] , 
        \nOut1_3[20] , \nOut1_3[19] , \nOut1_3[18] , \nOut1_3[17] , 
        \nOut1_3[16] , \nOut1_3[15] , \nOut1_3[14] , \nOut1_3[13] , 
        \nOut1_3[12] , \nOut1_3[11] , \nOut1_3[10] , \nOut1_3[9] , 
        \nOut1_3[8] , \nOut1_3[7] , \nOut1_3[6] , \nOut1_3[5] , \nOut1_3[4] , 
        \nOut1_3[3] , \nOut1_3[2] , \nOut1_3[1] , \nOut1_3[0] }), .EAST_EDGE(
        \nOut2_2[31] ), .WEST_EDGE(\nOut0_2[0] ), .NW_EDGE(\nOut0_1[0] ), 
        .SW_EDGE(\nOut0_3[0] ), .NE_EDGE(\nOut2_1[31] ), .SE_EDGE(
        \nOut2_3[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_43 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut44[31] , \nScanOut44[30] , \nScanOut44[29] , 
        \nScanOut44[28] , \nScanOut44[27] , \nScanOut44[26] , \nScanOut44[25] , 
        \nScanOut44[24] , \nScanOut44[23] , \nScanOut44[22] , \nScanOut44[21] , 
        \nScanOut44[20] , \nScanOut44[19] , \nScanOut44[18] , \nScanOut44[17] , 
        \nScanOut44[16] , \nScanOut44[15] , \nScanOut44[14] , \nScanOut44[13] , 
        \nScanOut44[12] , \nScanOut44[11] , \nScanOut44[10] , \nScanOut44[9] , 
        \nScanOut44[8] , \nScanOut44[7] , \nScanOut44[6] , \nScanOut44[5] , 
        \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , \nScanOut44[1] , 
        \nScanOut44[0] }), .ScanOut({\nScanOut43[31] , \nScanOut43[30] , 
        \nScanOut43[29] , \nScanOut43[28] , \nScanOut43[27] , \nScanOut43[26] , 
        \nScanOut43[25] , \nScanOut43[24] , \nScanOut43[23] , \nScanOut43[22] , 
        \nScanOut43[21] , \nScanOut43[20] , \nScanOut43[19] , \nScanOut43[18] , 
        \nScanOut43[17] , \nScanOut43[16] , \nScanOut43[15] , \nScanOut43[14] , 
        \nScanOut43[13] , \nScanOut43[12] , \nScanOut43[11] , \nScanOut43[10] , 
        \nScanOut43[9] , \nScanOut43[8] , \nScanOut43[7] , \nScanOut43[6] , 
        \nScanOut43[5] , \nScanOut43[4] , \nScanOut43[3] , \nScanOut43[2] , 
        \nScanOut43[1] , \nScanOut43[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_11[31] , 
        \nOut2_11[30] , \nOut2_11[29] , \nOut2_11[28] , \nOut2_11[27] , 
        \nOut2_11[26] , \nOut2_11[25] , \nOut2_11[24] , \nOut2_11[23] , 
        \nOut2_11[22] , \nOut2_11[21] , \nOut2_11[20] , \nOut2_11[19] , 
        \nOut2_11[18] , \nOut2_11[17] , \nOut2_11[16] , \nOut2_11[15] , 
        \nOut2_11[14] , \nOut2_11[13] , \nOut2_11[12] , \nOut2_11[11] , 
        \nOut2_11[10] , \nOut2_11[9] , \nOut2_11[8] , \nOut2_11[7] , 
        \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , \nOut2_11[3] , 
        \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), .NORTH_EDGE({
        \nOut2_10[31] , \nOut2_10[30] , \nOut2_10[29] , \nOut2_10[28] , 
        \nOut2_10[27] , \nOut2_10[26] , \nOut2_10[25] , \nOut2_10[24] , 
        \nOut2_10[23] , \nOut2_10[22] , \nOut2_10[21] , \nOut2_10[20] , 
        \nOut2_10[19] , \nOut2_10[18] , \nOut2_10[17] , \nOut2_10[16] , 
        \nOut2_10[15] , \nOut2_10[14] , \nOut2_10[13] , \nOut2_10[12] , 
        \nOut2_10[11] , \nOut2_10[10] , \nOut2_10[9] , \nOut2_10[8] , 
        \nOut2_10[7] , \nOut2_10[6] , \nOut2_10[5] , \nOut2_10[4] , 
        \nOut2_10[3] , \nOut2_10[2] , \nOut2_10[1] , \nOut2_10[0] }), 
        .SOUTH_EDGE({\nOut2_12[31] , \nOut2_12[30] , \nOut2_12[29] , 
        \nOut2_12[28] , \nOut2_12[27] , \nOut2_12[26] , \nOut2_12[25] , 
        \nOut2_12[24] , \nOut2_12[23] , \nOut2_12[22] , \nOut2_12[21] , 
        \nOut2_12[20] , \nOut2_12[19] , \nOut2_12[18] , \nOut2_12[17] , 
        \nOut2_12[16] , \nOut2_12[15] , \nOut2_12[14] , \nOut2_12[13] , 
        \nOut2_12[12] , \nOut2_12[11] , \nOut2_12[10] , \nOut2_12[9] , 
        \nOut2_12[8] , \nOut2_12[7] , \nOut2_12[6] , \nOut2_12[5] , 
        \nOut2_12[4] , \nOut2_12[3] , \nOut2_12[2] , \nOut2_12[1] , 
        \nOut2_12[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_11[0] ), 
        .NW_EDGE(\nOut1_10[0] ), .SW_EDGE(\nOut1_12[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_23 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut24[31] , \nScanOut24[30] , \nScanOut24[29] , 
        \nScanOut24[28] , \nScanOut24[27] , \nScanOut24[26] , \nScanOut24[25] , 
        \nScanOut24[24] , \nScanOut24[23] , \nScanOut24[22] , \nScanOut24[21] , 
        \nScanOut24[20] , \nScanOut24[19] , \nScanOut24[18] , \nScanOut24[17] , 
        \nScanOut24[16] , \nScanOut24[15] , \nScanOut24[14] , \nScanOut24[13] , 
        \nScanOut24[12] , \nScanOut24[11] , \nScanOut24[10] , \nScanOut24[9] , 
        \nScanOut24[8] , \nScanOut24[7] , \nScanOut24[6] , \nScanOut24[5] , 
        \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , \nScanOut24[1] , 
        \nScanOut24[0] }), .ScanOut({\nScanOut23[31] , \nScanOut23[30] , 
        \nScanOut23[29] , \nScanOut23[28] , \nScanOut23[27] , \nScanOut23[26] , 
        \nScanOut23[25] , \nScanOut23[24] , \nScanOut23[23] , \nScanOut23[22] , 
        \nScanOut23[21] , \nScanOut23[20] , \nScanOut23[19] , \nScanOut23[18] , 
        \nScanOut23[17] , \nScanOut23[16] , \nScanOut23[15] , \nScanOut23[14] , 
        \nScanOut23[13] , \nScanOut23[12] , \nScanOut23[11] , \nScanOut23[10] , 
        \nScanOut23[9] , \nScanOut23[8] , \nScanOut23[7] , \nScanOut23[6] , 
        \nScanOut23[5] , \nScanOut23[4] , \nScanOut23[3] , \nScanOut23[2] , 
        \nScanOut23[1] , \nScanOut23[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_7[31] , 
        \nOut1_7[30] , \nOut1_7[29] , \nOut1_7[28] , \nOut1_7[27] , 
        \nOut1_7[26] , \nOut1_7[25] , \nOut1_7[24] , \nOut1_7[23] , 
        \nOut1_7[22] , \nOut1_7[21] , \nOut1_7[20] , \nOut1_7[19] , 
        \nOut1_7[18] , \nOut1_7[17] , \nOut1_7[16] , \nOut1_7[15] , 
        \nOut1_7[14] , \nOut1_7[13] , \nOut1_7[12] , \nOut1_7[11] , 
        \nOut1_7[10] , \nOut1_7[9] , \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , 
        \nOut1_7[5] , \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , 
        \nOut1_7[0] }), .NORTH_EDGE({\nOut1_6[31] , \nOut1_6[30] , 
        \nOut1_6[29] , \nOut1_6[28] , \nOut1_6[27] , \nOut1_6[26] , 
        \nOut1_6[25] , \nOut1_6[24] , \nOut1_6[23] , \nOut1_6[22] , 
        \nOut1_6[21] , \nOut1_6[20] , \nOut1_6[19] , \nOut1_6[18] , 
        \nOut1_6[17] , \nOut1_6[16] , \nOut1_6[15] , \nOut1_6[14] , 
        \nOut1_6[13] , \nOut1_6[12] , \nOut1_6[11] , \nOut1_6[10] , 
        \nOut1_6[9] , \nOut1_6[8] , \nOut1_6[7] , \nOut1_6[6] , \nOut1_6[5] , 
        \nOut1_6[4] , \nOut1_6[3] , \nOut1_6[2] , \nOut1_6[1] , \nOut1_6[0] }), 
        .SOUTH_EDGE({\nOut1_8[31] , \nOut1_8[30] , \nOut1_8[29] , 
        \nOut1_8[28] , \nOut1_8[27] , \nOut1_8[26] , \nOut1_8[25] , 
        \nOut1_8[24] , \nOut1_8[23] , \nOut1_8[22] , \nOut1_8[21] , 
        \nOut1_8[20] , \nOut1_8[19] , \nOut1_8[18] , \nOut1_8[17] , 
        \nOut1_8[16] , \nOut1_8[15] , \nOut1_8[14] , \nOut1_8[13] , 
        \nOut1_8[12] , \nOut1_8[11] , \nOut1_8[10] , \nOut1_8[9] , 
        \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , \nOut1_8[5] , \nOut1_8[4] , 
        \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , \nOut1_8[0] }), .EAST_EDGE(
        \nOut2_7[31] ), .WEST_EDGE(\nOut0_7[0] ), .NW_EDGE(\nOut0_6[0] ), 
        .SW_EDGE(\nOut0_8[0] ), .NE_EDGE(\nOut2_6[31] ), .SE_EDGE(
        \nOut2_8[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_24 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut25[31] , \nScanOut25[30] , \nScanOut25[29] , 
        \nScanOut25[28] , \nScanOut25[27] , \nScanOut25[26] , \nScanOut25[25] , 
        \nScanOut25[24] , \nScanOut25[23] , \nScanOut25[22] , \nScanOut25[21] , 
        \nScanOut25[20] , \nScanOut25[19] , \nScanOut25[18] , \nScanOut25[17] , 
        \nScanOut25[16] , \nScanOut25[15] , \nScanOut25[14] , \nScanOut25[13] , 
        \nScanOut25[12] , \nScanOut25[11] , \nScanOut25[10] , \nScanOut25[9] , 
        \nScanOut25[8] , \nScanOut25[7] , \nScanOut25[6] , \nScanOut25[5] , 
        \nScanOut25[4] , \nScanOut25[3] , \nScanOut25[2] , \nScanOut25[1] , 
        \nScanOut25[0] }), .ScanOut({\nScanOut24[31] , \nScanOut24[30] , 
        \nScanOut24[29] , \nScanOut24[28] , \nScanOut24[27] , \nScanOut24[26] , 
        \nScanOut24[25] , \nScanOut24[24] , \nScanOut24[23] , \nScanOut24[22] , 
        \nScanOut24[21] , \nScanOut24[20] , \nScanOut24[19] , \nScanOut24[18] , 
        \nScanOut24[17] , \nScanOut24[16] , \nScanOut24[15] , \nScanOut24[14] , 
        \nScanOut24[13] , \nScanOut24[12] , \nScanOut24[11] , \nScanOut24[10] , 
        \nScanOut24[9] , \nScanOut24[8] , \nScanOut24[7] , \nScanOut24[6] , 
        \nScanOut24[5] , \nScanOut24[4] , \nScanOut24[3] , \nScanOut24[2] , 
        \nScanOut24[1] , \nScanOut24[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_8[31] , 
        \nOut1_8[30] , \nOut1_8[29] , \nOut1_8[28] , \nOut1_8[27] , 
        \nOut1_8[26] , \nOut1_8[25] , \nOut1_8[24] , \nOut1_8[23] , 
        \nOut1_8[22] , \nOut1_8[21] , \nOut1_8[20] , \nOut1_8[19] , 
        \nOut1_8[18] , \nOut1_8[17] , \nOut1_8[16] , \nOut1_8[15] , 
        \nOut1_8[14] , \nOut1_8[13] , \nOut1_8[12] , \nOut1_8[11] , 
        \nOut1_8[10] , \nOut1_8[9] , \nOut1_8[8] , \nOut1_8[7] , \nOut1_8[6] , 
        \nOut1_8[5] , \nOut1_8[4] , \nOut1_8[3] , \nOut1_8[2] , \nOut1_8[1] , 
        \nOut1_8[0] }), .NORTH_EDGE({\nOut1_7[31] , \nOut1_7[30] , 
        \nOut1_7[29] , \nOut1_7[28] , \nOut1_7[27] , \nOut1_7[26] , 
        \nOut1_7[25] , \nOut1_7[24] , \nOut1_7[23] , \nOut1_7[22] , 
        \nOut1_7[21] , \nOut1_7[20] , \nOut1_7[19] , \nOut1_7[18] , 
        \nOut1_7[17] , \nOut1_7[16] , \nOut1_7[15] , \nOut1_7[14] , 
        \nOut1_7[13] , \nOut1_7[12] , \nOut1_7[11] , \nOut1_7[10] , 
        \nOut1_7[9] , \nOut1_7[8] , \nOut1_7[7] , \nOut1_7[6] , \nOut1_7[5] , 
        \nOut1_7[4] , \nOut1_7[3] , \nOut1_7[2] , \nOut1_7[1] , \nOut1_7[0] }), 
        .SOUTH_EDGE({\nOut1_9[31] , \nOut1_9[30] , \nOut1_9[29] , 
        \nOut1_9[28] , \nOut1_9[27] , \nOut1_9[26] , \nOut1_9[25] , 
        \nOut1_9[24] , \nOut1_9[23] , \nOut1_9[22] , \nOut1_9[21] , 
        \nOut1_9[20] , \nOut1_9[19] , \nOut1_9[18] , \nOut1_9[17] , 
        \nOut1_9[16] , \nOut1_9[15] , \nOut1_9[14] , \nOut1_9[13] , 
        \nOut1_9[12] , \nOut1_9[11] , \nOut1_9[10] , \nOut1_9[9] , 
        \nOut1_9[8] , \nOut1_9[7] , \nOut1_9[6] , \nOut1_9[5] , \nOut1_9[4] , 
        \nOut1_9[3] , \nOut1_9[2] , \nOut1_9[1] , \nOut1_9[0] }), .EAST_EDGE(
        \nOut2_8[31] ), .WEST_EDGE(\nOut0_8[0] ), .NW_EDGE(\nOut0_7[0] ), 
        .SW_EDGE(\nOut0_9[0] ), .NE_EDGE(\nOut2_7[31] ), .SE_EDGE(
        \nOut2_9[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_8 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut9[31] , \nScanOut9[30] , \nScanOut9[29] , 
        \nScanOut9[28] , \nScanOut9[27] , \nScanOut9[26] , \nScanOut9[25] , 
        \nScanOut9[24] , \nScanOut9[23] , \nScanOut9[22] , \nScanOut9[21] , 
        \nScanOut9[20] , \nScanOut9[19] , \nScanOut9[18] , \nScanOut9[17] , 
        \nScanOut9[16] , \nScanOut9[15] , \nScanOut9[14] , \nScanOut9[13] , 
        \nScanOut9[12] , \nScanOut9[11] , \nScanOut9[10] , \nScanOut9[9] , 
        \nScanOut9[8] , \nScanOut9[7] , \nScanOut9[6] , \nScanOut9[5] , 
        \nScanOut9[4] , \nScanOut9[3] , \nScanOut9[2] , \nScanOut9[1] , 
        \nScanOut9[0] }), .ScanOut({\nScanOut8[31] , \nScanOut8[30] , 
        \nScanOut8[29] , \nScanOut8[28] , \nScanOut8[27] , \nScanOut8[26] , 
        \nScanOut8[25] , \nScanOut8[24] , \nScanOut8[23] , \nScanOut8[22] , 
        \nScanOut8[21] , \nScanOut8[20] , \nScanOut8[19] , \nScanOut8[18] , 
        \nScanOut8[17] , \nScanOut8[16] , \nScanOut8[15] , \nScanOut8[14] , 
        \nScanOut8[13] , \nScanOut8[12] , \nScanOut8[11] , \nScanOut8[10] , 
        \nScanOut8[9] , \nScanOut8[8] , \nScanOut8[7] , \nScanOut8[6] , 
        \nScanOut8[5] , \nScanOut8[4] , \nScanOut8[3] , \nScanOut8[2] , 
        \nScanOut8[1] , \nScanOut8[0] }), .ScanEnable(\nScanEnable[0] ), .Id(
        1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut0_8[31] , 
        \nOut0_8[30] , \nOut0_8[29] , \nOut0_8[28] , \nOut0_8[27] , 
        \nOut0_8[26] , \nOut0_8[25] , \nOut0_8[24] , \nOut0_8[23] , 
        \nOut0_8[22] , \nOut0_8[21] , \nOut0_8[20] , \nOut0_8[19] , 
        \nOut0_8[18] , \nOut0_8[17] , \nOut0_8[16] , \nOut0_8[15] , 
        \nOut0_8[14] , \nOut0_8[13] , \nOut0_8[12] , \nOut0_8[11] , 
        \nOut0_8[10] , \nOut0_8[9] , \nOut0_8[8] , \nOut0_8[7] , \nOut0_8[6] , 
        \nOut0_8[5] , \nOut0_8[4] , \nOut0_8[3] , \nOut0_8[2] , \nOut0_8[1] , 
        \nOut0_8[0] }), .NORTH_EDGE({\nOut0_7[31] , \nOut0_7[30] , 
        \nOut0_7[29] , \nOut0_7[28] , \nOut0_7[27] , \nOut0_7[26] , 
        \nOut0_7[25] , \nOut0_7[24] , \nOut0_7[23] , \nOut0_7[22] , 
        \nOut0_7[21] , \nOut0_7[20] , \nOut0_7[19] , \nOut0_7[18] , 
        \nOut0_7[17] , \nOut0_7[16] , \nOut0_7[15] , \nOut0_7[14] , 
        \nOut0_7[13] , \nOut0_7[12] , \nOut0_7[11] , \nOut0_7[10] , 
        \nOut0_7[9] , \nOut0_7[8] , \nOut0_7[7] , \nOut0_7[6] , \nOut0_7[5] , 
        \nOut0_7[4] , \nOut0_7[3] , \nOut0_7[2] , \nOut0_7[1] , \nOut0_7[0] }), 
        .SOUTH_EDGE({\nOut0_9[31] , \nOut0_9[30] , \nOut0_9[29] , 
        \nOut0_9[28] , \nOut0_9[27] , \nOut0_9[26] , \nOut0_9[25] , 
        \nOut0_9[24] , \nOut0_9[23] , \nOut0_9[22] , \nOut0_9[21] , 
        \nOut0_9[20] , \nOut0_9[19] , \nOut0_9[18] , \nOut0_9[17] , 
        \nOut0_9[16] , \nOut0_9[15] , \nOut0_9[14] , \nOut0_9[13] , 
        \nOut0_9[12] , \nOut0_9[11] , \nOut0_9[10] , \nOut0_9[9] , 
        \nOut0_9[8] , \nOut0_9[7] , \nOut0_9[6] , \nOut0_9[5] , \nOut0_9[4] , 
        \nOut0_9[3] , \nOut0_9[2] , \nOut0_9[1] , \nOut0_9[0] }), .EAST_EDGE(
        \nOut1_8[31] ), .WEST_EDGE(1'b0), .NW_EDGE(1'b0), .SW_EDGE(1'b0), 
        .NE_EDGE(\nOut1_7[31] ), .SE_EDGE(\nOut1_9[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_38 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut39[31] , \nScanOut39[30] , \nScanOut39[29] , 
        \nScanOut39[28] , \nScanOut39[27] , \nScanOut39[26] , \nScanOut39[25] , 
        \nScanOut39[24] , \nScanOut39[23] , \nScanOut39[22] , \nScanOut39[21] , 
        \nScanOut39[20] , \nScanOut39[19] , \nScanOut39[18] , \nScanOut39[17] , 
        \nScanOut39[16] , \nScanOut39[15] , \nScanOut39[14] , \nScanOut39[13] , 
        \nScanOut39[12] , \nScanOut39[11] , \nScanOut39[10] , \nScanOut39[9] , 
        \nScanOut39[8] , \nScanOut39[7] , \nScanOut39[6] , \nScanOut39[5] , 
        \nScanOut39[4] , \nScanOut39[3] , \nScanOut39[2] , \nScanOut39[1] , 
        \nScanOut39[0] }), .ScanOut({\nScanOut38[31] , \nScanOut38[30] , 
        \nScanOut38[29] , \nScanOut38[28] , \nScanOut38[27] , \nScanOut38[26] , 
        \nScanOut38[25] , \nScanOut38[24] , \nScanOut38[23] , \nScanOut38[22] , 
        \nScanOut38[21] , \nScanOut38[20] , \nScanOut38[19] , \nScanOut38[18] , 
        \nScanOut38[17] , \nScanOut38[16] , \nScanOut38[15] , \nScanOut38[14] , 
        \nScanOut38[13] , \nScanOut38[12] , \nScanOut38[11] , \nScanOut38[10] , 
        \nScanOut38[9] , \nScanOut38[8] , \nScanOut38[7] , \nScanOut38[6] , 
        \nScanOut38[5] , \nScanOut38[4] , \nScanOut38[3] , \nScanOut38[2] , 
        \nScanOut38[1] , \nScanOut38[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_6[31] , 
        \nOut2_6[30] , \nOut2_6[29] , \nOut2_6[28] , \nOut2_6[27] , 
        \nOut2_6[26] , \nOut2_6[25] , \nOut2_6[24] , \nOut2_6[23] , 
        \nOut2_6[22] , \nOut2_6[21] , \nOut2_6[20] , \nOut2_6[19] , 
        \nOut2_6[18] , \nOut2_6[17] , \nOut2_6[16] , \nOut2_6[15] , 
        \nOut2_6[14] , \nOut2_6[13] , \nOut2_6[12] , \nOut2_6[11] , 
        \nOut2_6[10] , \nOut2_6[9] , \nOut2_6[8] , \nOut2_6[7] , \nOut2_6[6] , 
        \nOut2_6[5] , \nOut2_6[4] , \nOut2_6[3] , \nOut2_6[2] , \nOut2_6[1] , 
        \nOut2_6[0] }), .NORTH_EDGE({\nOut2_5[31] , \nOut2_5[30] , 
        \nOut2_5[29] , \nOut2_5[28] , \nOut2_5[27] , \nOut2_5[26] , 
        \nOut2_5[25] , \nOut2_5[24] , \nOut2_5[23] , \nOut2_5[22] , 
        \nOut2_5[21] , \nOut2_5[20] , \nOut2_5[19] , \nOut2_5[18] , 
        \nOut2_5[17] , \nOut2_5[16] , \nOut2_5[15] , \nOut2_5[14] , 
        \nOut2_5[13] , \nOut2_5[12] , \nOut2_5[11] , \nOut2_5[10] , 
        \nOut2_5[9] , \nOut2_5[8] , \nOut2_5[7] , \nOut2_5[6] , \nOut2_5[5] , 
        \nOut2_5[4] , \nOut2_5[3] , \nOut2_5[2] , \nOut2_5[1] , \nOut2_5[0] }), 
        .SOUTH_EDGE({\nOut2_7[31] , \nOut2_7[30] , \nOut2_7[29] , 
        \nOut2_7[28] , \nOut2_7[27] , \nOut2_7[26] , \nOut2_7[25] , 
        \nOut2_7[24] , \nOut2_7[23] , \nOut2_7[22] , \nOut2_7[21] , 
        \nOut2_7[20] , \nOut2_7[19] , \nOut2_7[18] , \nOut2_7[17] , 
        \nOut2_7[16] , \nOut2_7[15] , \nOut2_7[14] , \nOut2_7[13] , 
        \nOut2_7[12] , \nOut2_7[11] , \nOut2_7[10] , \nOut2_7[9] , 
        \nOut2_7[8] , \nOut2_7[7] , \nOut2_7[6] , \nOut2_7[5] , \nOut2_7[4] , 
        \nOut2_7[3] , \nOut2_7[2] , \nOut2_7[1] , \nOut2_7[0] }), .EAST_EDGE(
        1'b0), .WEST_EDGE(\nOut1_6[0] ), .NW_EDGE(\nOut1_5[0] ), .SW_EDGE(
        \nOut1_7[0] ), .NE_EDGE(1'b0), .SE_EDGE(1'b0) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_44 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut45[31] , \nScanOut45[30] , \nScanOut45[29] , 
        \nScanOut45[28] , \nScanOut45[27] , \nScanOut45[26] , \nScanOut45[25] , 
        \nScanOut45[24] , \nScanOut45[23] , \nScanOut45[22] , \nScanOut45[21] , 
        \nScanOut45[20] , \nScanOut45[19] , \nScanOut45[18] , \nScanOut45[17] , 
        \nScanOut45[16] , \nScanOut45[15] , \nScanOut45[14] , \nScanOut45[13] , 
        \nScanOut45[12] , \nScanOut45[11] , \nScanOut45[10] , \nScanOut45[9] , 
        \nScanOut45[8] , \nScanOut45[7] , \nScanOut45[6] , \nScanOut45[5] , 
        \nScanOut45[4] , \nScanOut45[3] , \nScanOut45[2] , \nScanOut45[1] , 
        \nScanOut45[0] }), .ScanOut({\nScanOut44[31] , \nScanOut44[30] , 
        \nScanOut44[29] , \nScanOut44[28] , \nScanOut44[27] , \nScanOut44[26] , 
        \nScanOut44[25] , \nScanOut44[24] , \nScanOut44[23] , \nScanOut44[22] , 
        \nScanOut44[21] , \nScanOut44[20] , \nScanOut44[19] , \nScanOut44[18] , 
        \nScanOut44[17] , \nScanOut44[16] , \nScanOut44[15] , \nScanOut44[14] , 
        \nScanOut44[13] , \nScanOut44[12] , \nScanOut44[11] , \nScanOut44[10] , 
        \nScanOut44[9] , \nScanOut44[8] , \nScanOut44[7] , \nScanOut44[6] , 
        \nScanOut44[5] , \nScanOut44[4] , \nScanOut44[3] , \nScanOut44[2] , 
        \nScanOut44[1] , \nScanOut44[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut2_12[31] , 
        \nOut2_12[30] , \nOut2_12[29] , \nOut2_12[28] , \nOut2_12[27] , 
        \nOut2_12[26] , \nOut2_12[25] , \nOut2_12[24] , \nOut2_12[23] , 
        \nOut2_12[22] , \nOut2_12[21] , \nOut2_12[20] , \nOut2_12[19] , 
        \nOut2_12[18] , \nOut2_12[17] , \nOut2_12[16] , \nOut2_12[15] , 
        \nOut2_12[14] , \nOut2_12[13] , \nOut2_12[12] , \nOut2_12[11] , 
        \nOut2_12[10] , \nOut2_12[9] , \nOut2_12[8] , \nOut2_12[7] , 
        \nOut2_12[6] , \nOut2_12[5] , \nOut2_12[4] , \nOut2_12[3] , 
        \nOut2_12[2] , \nOut2_12[1] , \nOut2_12[0] }), .NORTH_EDGE({
        \nOut2_11[31] , \nOut2_11[30] , \nOut2_11[29] , \nOut2_11[28] , 
        \nOut2_11[27] , \nOut2_11[26] , \nOut2_11[25] , \nOut2_11[24] , 
        \nOut2_11[23] , \nOut2_11[22] , \nOut2_11[21] , \nOut2_11[20] , 
        \nOut2_11[19] , \nOut2_11[18] , \nOut2_11[17] , \nOut2_11[16] , 
        \nOut2_11[15] , \nOut2_11[14] , \nOut2_11[13] , \nOut2_11[12] , 
        \nOut2_11[11] , \nOut2_11[10] , \nOut2_11[9] , \nOut2_11[8] , 
        \nOut2_11[7] , \nOut2_11[6] , \nOut2_11[5] , \nOut2_11[4] , 
        \nOut2_11[3] , \nOut2_11[2] , \nOut2_11[1] , \nOut2_11[0] }), 
        .SOUTH_EDGE({\nOut2_13[31] , \nOut2_13[30] , \nOut2_13[29] , 
        \nOut2_13[28] , \nOut2_13[27] , \nOut2_13[26] , \nOut2_13[25] , 
        \nOut2_13[24] , \nOut2_13[23] , \nOut2_13[22] , \nOut2_13[21] , 
        \nOut2_13[20] , \nOut2_13[19] , \nOut2_13[18] , \nOut2_13[17] , 
        \nOut2_13[16] , \nOut2_13[15] , \nOut2_13[14] , \nOut2_13[13] , 
        \nOut2_13[12] , \nOut2_13[11] , \nOut2_13[10] , \nOut2_13[9] , 
        \nOut2_13[8] , \nOut2_13[7] , \nOut2_13[6] , \nOut2_13[5] , 
        \nOut2_13[4] , \nOut2_13[3] , \nOut2_13[2] , \nOut2_13[1] , 
        \nOut2_13[0] }), .EAST_EDGE(1'b0), .WEST_EDGE(\nOut1_12[0] ), 
        .NW_EDGE(\nOut1_11[0] ), .SW_EDGE(\nOut1_13[0] ), .NE_EDGE(1'b0), 
        .SE_EDGE(1'b0) );
    Life_Control_WIDTH32_CWIDTH7_IDWIDTH1_SCAN1 U_Life_Control ( .Clk(Clk), 
        .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), 
        .DataOut(DataOut), .ScanIn({\nScanOut0[31] , \nScanOut0[30] , 
        \nScanOut0[29] , \nScanOut0[28] , \nScanOut0[27] , \nScanOut0[26] , 
        \nScanOut0[25] , \nScanOut0[24] , \nScanOut0[23] , \nScanOut0[22] , 
        \nScanOut0[21] , \nScanOut0[20] , \nScanOut0[19] , \nScanOut0[18] , 
        \nScanOut0[17] , \nScanOut0[16] , \nScanOut0[15] , \nScanOut0[14] , 
        \nScanOut0[13] , \nScanOut0[12] , \nScanOut0[11] , \nScanOut0[10] , 
        \nScanOut0[9] , \nScanOut0[8] , \nScanOut0[7] , \nScanOut0[6] , 
        \nScanOut0[5] , \nScanOut0[4] , \nScanOut0[3] , \nScanOut0[2] , 
        \nScanOut0[1] , \nScanOut0[0] }), .ScanOut({\nScanOut48[31] , 
        \nScanOut48[30] , \nScanOut48[29] , \nScanOut48[28] , \nScanOut48[27] , 
        \nScanOut48[26] , \nScanOut48[25] , \nScanOut48[24] , \nScanOut48[23] , 
        \nScanOut48[22] , \nScanOut48[21] , \nScanOut48[20] , \nScanOut48[19] , 
        \nScanOut48[18] , \nScanOut48[17] , \nScanOut48[16] , \nScanOut48[15] , 
        \nScanOut48[14] , \nScanOut48[13] , \nScanOut48[12] , \nScanOut48[11] , 
        \nScanOut48[10] , \nScanOut48[9] , \nScanOut48[8] , \nScanOut48[7] , 
        \nScanOut48[6] , \nScanOut48[5] , \nScanOut48[4] , \nScanOut48[3] , 
        \nScanOut48[2] , \nScanOut48[1] , \nScanOut48[0] }), .ScanEnable(
        \nScanEnable[0] ), .Id(1'b1), .ScanId(1'b0), .Enable(\nEnable[0] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_16 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut17[31] , \nScanOut17[30] , \nScanOut17[29] , 
        \nScanOut17[28] , \nScanOut17[27] , \nScanOut17[26] , \nScanOut17[25] , 
        \nScanOut17[24] , \nScanOut17[23] , \nScanOut17[22] , \nScanOut17[21] , 
        \nScanOut17[20] , \nScanOut17[19] , \nScanOut17[18] , \nScanOut17[17] , 
        \nScanOut17[16] , \nScanOut17[15] , \nScanOut17[14] , \nScanOut17[13] , 
        \nScanOut17[12] , \nScanOut17[11] , \nScanOut17[10] , \nScanOut17[9] , 
        \nScanOut17[8] , \nScanOut17[7] , \nScanOut17[6] , \nScanOut17[5] , 
        \nScanOut17[4] , \nScanOut17[3] , \nScanOut17[2] , \nScanOut17[1] , 
        \nScanOut17[0] }), .ScanOut({\nScanOut16[31] , \nScanOut16[30] , 
        \nScanOut16[29] , \nScanOut16[28] , \nScanOut16[27] , \nScanOut16[26] , 
        \nScanOut16[25] , \nScanOut16[24] , \nScanOut16[23] , \nScanOut16[22] , 
        \nScanOut16[21] , \nScanOut16[20] , \nScanOut16[19] , \nScanOut16[18] , 
        \nScanOut16[17] , \nScanOut16[16] , \nScanOut16[15] , \nScanOut16[14] , 
        \nScanOut16[13] , \nScanOut16[12] , \nScanOut16[11] , \nScanOut16[10] , 
        \nScanOut16[9] , \nScanOut16[8] , \nScanOut16[7] , \nScanOut16[6] , 
        \nScanOut16[5] , \nScanOut16[4] , \nScanOut16[3] , \nScanOut16[2] , 
        \nScanOut16[1] , \nScanOut16[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_0[31] , 
        \nOut1_0[30] , \nOut1_0[29] , \nOut1_0[28] , \nOut1_0[27] , 
        \nOut1_0[26] , \nOut1_0[25] , \nOut1_0[24] , \nOut1_0[23] , 
        \nOut1_0[22] , \nOut1_0[21] , \nOut1_0[20] , \nOut1_0[19] , 
        \nOut1_0[18] , \nOut1_0[17] , \nOut1_0[16] , \nOut1_0[15] , 
        \nOut1_0[14] , \nOut1_0[13] , \nOut1_0[12] , \nOut1_0[11] , 
        \nOut1_0[10] , \nOut1_0[9] , \nOut1_0[8] , \nOut1_0[7] , \nOut1_0[6] , 
        \nOut1_0[5] , \nOut1_0[4] , \nOut1_0[3] , \nOut1_0[2] , \nOut1_0[1] , 
        \nOut1_0[0] }), .NORTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SOUTH_EDGE({\nOut1_1[31] , \nOut1_1[30] , \nOut1_1[29] , 
        \nOut1_1[28] , \nOut1_1[27] , \nOut1_1[26] , \nOut1_1[25] , 
        \nOut1_1[24] , \nOut1_1[23] , \nOut1_1[22] , \nOut1_1[21] , 
        \nOut1_1[20] , \nOut1_1[19] , \nOut1_1[18] , \nOut1_1[17] , 
        \nOut1_1[16] , \nOut1_1[15] , \nOut1_1[14] , \nOut1_1[13] , 
        \nOut1_1[12] , \nOut1_1[11] , \nOut1_1[10] , \nOut1_1[9] , 
        \nOut1_1[8] , \nOut1_1[7] , \nOut1_1[6] , \nOut1_1[5] , \nOut1_1[4] , 
        \nOut1_1[3] , \nOut1_1[2] , \nOut1_1[1] , \nOut1_1[0] }), .EAST_EDGE(
        \nOut2_0[31] ), .WEST_EDGE(\nOut0_0[0] ), .NW_EDGE(1'b0), .SW_EDGE(
        \nOut0_1[0] ), .NE_EDGE(1'b0), .SE_EDGE(\nOut2_1[31] ) );
    Life_Block_IDWIDTH1_SCAN1 U_Life_Block_31 ( .Clk(Clk), .Reset(Reset), .RD(
        RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), 
        .ScanIn({\nScanOut32[31] , \nScanOut32[30] , \nScanOut32[29] , 
        \nScanOut32[28] , \nScanOut32[27] , \nScanOut32[26] , \nScanOut32[25] , 
        \nScanOut32[24] , \nScanOut32[23] , \nScanOut32[22] , \nScanOut32[21] , 
        \nScanOut32[20] , \nScanOut32[19] , \nScanOut32[18] , \nScanOut32[17] , 
        \nScanOut32[16] , \nScanOut32[15] , \nScanOut32[14] , \nScanOut32[13] , 
        \nScanOut32[12] , \nScanOut32[11] , \nScanOut32[10] , \nScanOut32[9] , 
        \nScanOut32[8] , \nScanOut32[7] , \nScanOut32[6] , \nScanOut32[5] , 
        \nScanOut32[4] , \nScanOut32[3] , \nScanOut32[2] , \nScanOut32[1] , 
        \nScanOut32[0] }), .ScanOut({\nScanOut31[31] , \nScanOut31[30] , 
        \nScanOut31[29] , \nScanOut31[28] , \nScanOut31[27] , \nScanOut31[26] , 
        \nScanOut31[25] , \nScanOut31[24] , \nScanOut31[23] , \nScanOut31[22] , 
        \nScanOut31[21] , \nScanOut31[20] , \nScanOut31[19] , \nScanOut31[18] , 
        \nScanOut31[17] , \nScanOut31[16] , \nScanOut31[15] , \nScanOut31[14] , 
        \nScanOut31[13] , \nScanOut31[12] , \nScanOut31[11] , \nScanOut31[10] , 
        \nScanOut31[9] , \nScanOut31[8] , \nScanOut31[7] , \nScanOut31[6] , 
        \nScanOut31[5] , \nScanOut31[4] , \nScanOut31[3] , \nScanOut31[2] , 
        \nScanOut31[1] , \nScanOut31[0] }), .ScanEnable(\nScanEnable[0] ), 
        .Id(1'b0), .Enable(\nEnable[0] ), .BLOCK_VALUE({\nOut1_15[31] , 
        \nOut1_15[30] , \nOut1_15[29] , \nOut1_15[28] , \nOut1_15[27] , 
        \nOut1_15[26] , \nOut1_15[25] , \nOut1_15[24] , \nOut1_15[23] , 
        \nOut1_15[22] , \nOut1_15[21] , \nOut1_15[20] , \nOut1_15[19] , 
        \nOut1_15[18] , \nOut1_15[17] , \nOut1_15[16] , \nOut1_15[15] , 
        \nOut1_15[14] , \nOut1_15[13] , \nOut1_15[12] , \nOut1_15[11] , 
        \nOut1_15[10] , \nOut1_15[9] , \nOut1_15[8] , \nOut1_15[7] , 
        \nOut1_15[6] , \nOut1_15[5] , \nOut1_15[4] , \nOut1_15[3] , 
        \nOut1_15[2] , \nOut1_15[1] , \nOut1_15[0] }), .NORTH_EDGE({
        \nOut1_14[31] , \nOut1_14[30] , \nOut1_14[29] , \nOut1_14[28] , 
        \nOut1_14[27] , \nOut1_14[26] , \nOut1_14[25] , \nOut1_14[24] , 
        \nOut1_14[23] , \nOut1_14[22] , \nOut1_14[21] , \nOut1_14[20] , 
        \nOut1_14[19] , \nOut1_14[18] , \nOut1_14[17] , \nOut1_14[16] , 
        \nOut1_14[15] , \nOut1_14[14] , \nOut1_14[13] , \nOut1_14[12] , 
        \nOut1_14[11] , \nOut1_14[10] , \nOut1_14[9] , \nOut1_14[8] , 
        \nOut1_14[7] , \nOut1_14[6] , \nOut1_14[5] , \nOut1_14[4] , 
        \nOut1_14[3] , \nOut1_14[2] , \nOut1_14[1] , \nOut1_14[0] }), 
        .SOUTH_EDGE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .EAST_EDGE(\nOut2_15[31] ), .WEST_EDGE(\nOut0_15[0] ), .NW_EDGE(
        \nOut0_14[0] ), .SW_EDGE(1'b0), .NE_EDGE(\nOut2_14[31] ), .SE_EDGE(
        1'b0) );
endmodule

